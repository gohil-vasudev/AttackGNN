module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n1024_, new_n1125_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n1145_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1150_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n1070_, new_n176_, new_n1109_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n1142_, new_n654_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n861_, new_n1095_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g0000 ( new_n138_, N1 );
not g0001 ( new_n139_, N73 );
nor g0002 ( new_n140_, new_n139_, N77 );
not g0003 ( new_n141_, N77 );
nor g0004 ( new_n142_, new_n141_, N73 );
nor g0005 ( new_n143_, new_n140_, new_n142_ );
nand g0006 ( new_n144_, N65, N69 );
not g0007 ( new_n145_, new_n144_ );
nor g0008 ( new_n146_, N65, N69 );
nor g0009 ( new_n147_, new_n145_, new_n146_ );
nor g0010 ( new_n148_, new_n143_, new_n147_ );
nand g0011 ( new_n149_, new_n143_, new_n147_ );
not g0012 ( new_n150_, new_n149_ );
nor g0013 ( new_n151_, new_n150_, new_n148_ );
not g0014 ( new_n152_, N89 );
nor g0015 ( new_n153_, new_n152_, N93 );
not g0016 ( new_n154_, N93 );
nor g0017 ( new_n155_, new_n154_, N89 );
nor g0018 ( new_n156_, new_n153_, new_n155_ );
nand g0019 ( new_n157_, N81, N85 );
not g0020 ( new_n158_, new_n157_ );
nor g0021 ( new_n159_, N81, N85 );
nor g0022 ( new_n160_, new_n158_, new_n159_ );
nor g0023 ( new_n161_, new_n156_, new_n160_ );
nand g0024 ( new_n162_, new_n156_, new_n160_ );
not g0025 ( new_n163_, new_n162_ );
nor g0026 ( new_n164_, new_n163_, new_n161_ );
not g0027 ( new_n165_, new_n164_ );
nor g0028 ( new_n166_, new_n165_, new_n151_ );
not g0029 ( new_n167_, new_n151_ );
nor g0030 ( new_n168_, new_n167_, new_n164_ );
nor g0031 ( new_n169_, new_n166_, new_n168_ );
not g0032 ( new_n170_, new_n169_ );
nand g0033 ( new_n171_, N129, N137 );
nand g0034 ( new_n172_, new_n170_, new_n171_ );
not g0035 ( new_n173_, new_n172_ );
nor g0036 ( new_n174_, new_n170_, new_n171_ );
nor g0037 ( new_n175_, new_n173_, new_n174_ );
not g0038 ( new_n176_, N33 );
nor g0039 ( new_n177_, new_n176_, N49 );
not g0040 ( new_n178_, N49 );
nor g0041 ( new_n179_, new_n178_, N33 );
nor g0042 ( new_n180_, new_n177_, new_n179_ );
nand g0043 ( new_n181_, N1, N17 );
not g0044 ( new_n182_, new_n181_ );
nor g0045 ( new_n183_, N1, N17 );
nor g0046 ( new_n184_, new_n182_, new_n183_ );
nor g0047 ( new_n185_, new_n180_, new_n184_ );
nand g0048 ( new_n186_, new_n180_, new_n184_ );
not g0049 ( new_n187_, new_n186_ );
nor g0050 ( new_n188_, new_n187_, new_n185_ );
nor g0051 ( new_n189_, new_n175_, new_n188_ );
nand g0052 ( new_n190_, new_n175_, new_n188_ );
not g0053 ( new_n191_, new_n190_ );
nor g0054 ( new_n192_, new_n191_, new_n189_ );
not g0055 ( new_n193_, new_n192_ );
not g0056 ( new_n194_, N105 );
nor g0057 ( new_n195_, new_n194_, N109 );
not g0058 ( new_n196_, N109 );
nor g0059 ( new_n197_, new_n196_, N105 );
nor g0060 ( new_n198_, new_n195_, new_n197_ );
nand g0061 ( new_n199_, N97, N101 );
not g0062 ( new_n200_, new_n199_ );
nor g0063 ( new_n201_, N97, N101 );
nor g0064 ( new_n202_, new_n200_, new_n201_ );
nor g0065 ( new_n203_, new_n198_, new_n202_ );
nand g0066 ( new_n204_, new_n198_, new_n202_ );
not g0067 ( new_n205_, new_n204_ );
nor g0068 ( new_n206_, new_n205_, new_n203_ );
not g0069 ( new_n207_, new_n206_ );
nor g0070 ( new_n208_, new_n207_, new_n151_ );
nor g0071 ( new_n209_, new_n167_, new_n206_ );
nor g0072 ( new_n210_, new_n208_, new_n209_ );
not g0073 ( new_n211_, new_n210_ );
nand g0074 ( new_n212_, N131, N137 );
nand g0075 ( new_n213_, new_n211_, new_n212_ );
not g0076 ( new_n214_, new_n213_ );
nor g0077 ( new_n215_, new_n211_, new_n212_ );
nor g0078 ( new_n216_, new_n214_, new_n215_ );
not g0079 ( new_n217_, N41 );
nor g0080 ( new_n218_, new_n217_, N57 );
not g0081 ( new_n219_, N57 );
nor g0082 ( new_n220_, new_n219_, N41 );
nor g0083 ( new_n221_, new_n218_, new_n220_ );
nand g0084 ( new_n222_, N9, N25 );
not g0085 ( new_n223_, new_n222_ );
nor g0086 ( new_n224_, N9, N25 );
nor g0087 ( new_n225_, new_n223_, new_n224_ );
nor g0088 ( new_n226_, new_n221_, new_n225_ );
nand g0089 ( new_n227_, new_n221_, new_n225_ );
not g0090 ( new_n228_, new_n227_ );
nor g0091 ( new_n229_, new_n228_, new_n226_ );
nor g0092 ( new_n230_, new_n216_, new_n229_ );
nand g0093 ( new_n231_, new_n216_, new_n229_ );
not g0094 ( new_n232_, new_n231_ );
nor g0095 ( new_n233_, new_n232_, new_n230_ );
nand g0096 ( new_n234_, new_n233_, keyIn_0_24 );
nor g0097 ( new_n235_, new_n234_, new_n193_ );
nand g0098 ( new_n236_, new_n234_, new_n193_ );
not g0099 ( new_n237_, N121 );
nor g0100 ( new_n238_, new_n237_, N125 );
not g0101 ( new_n239_, N125 );
nor g0102 ( new_n240_, new_n239_, N121 );
nor g0103 ( new_n241_, new_n238_, new_n240_ );
nand g0104 ( new_n242_, N113, N117 );
not g0105 ( new_n243_, new_n242_ );
nor g0106 ( new_n244_, N113, N117 );
nor g0107 ( new_n245_, new_n243_, new_n244_ );
nor g0108 ( new_n246_, new_n241_, new_n245_ );
nand g0109 ( new_n247_, new_n241_, new_n245_ );
not g0110 ( new_n248_, new_n247_ );
nor g0111 ( new_n249_, new_n248_, new_n246_ );
not g0112 ( new_n250_, new_n249_ );
nor g0113 ( new_n251_, new_n250_, new_n206_ );
nor g0114 ( new_n252_, new_n207_, new_n249_ );
nor g0115 ( new_n253_, new_n251_, new_n252_ );
not g0116 ( new_n254_, new_n253_ );
nand g0117 ( new_n255_, N130, N137 );
nand g0118 ( new_n256_, new_n254_, new_n255_ );
not g0119 ( new_n257_, new_n256_ );
nor g0120 ( new_n258_, new_n254_, new_n255_ );
nor g0121 ( new_n259_, new_n257_, new_n258_ );
not g0122 ( new_n260_, N37 );
nor g0123 ( new_n261_, new_n260_, N53 );
not g0124 ( new_n262_, N53 );
nor g0125 ( new_n263_, new_n262_, N37 );
nor g0126 ( new_n264_, new_n261_, new_n263_ );
nand g0127 ( new_n265_, N5, N21 );
not g0128 ( new_n266_, new_n265_ );
nor g0129 ( new_n267_, N5, N21 );
nor g0130 ( new_n268_, new_n266_, new_n267_ );
nor g0131 ( new_n269_, new_n264_, new_n268_ );
nand g0132 ( new_n270_, new_n264_, new_n268_ );
not g0133 ( new_n271_, new_n270_ );
nor g0134 ( new_n272_, new_n271_, new_n269_ );
nor g0135 ( new_n273_, new_n259_, new_n272_ );
nand g0136 ( new_n274_, new_n259_, new_n272_ );
not g0137 ( new_n275_, new_n274_ );
nor g0138 ( new_n276_, new_n275_, new_n273_ );
not g0139 ( new_n277_, new_n276_ );
nand g0140 ( new_n278_, new_n236_, new_n277_ );
nor g0141 ( new_n279_, new_n278_, new_n235_ );
not g0142 ( new_n280_, new_n233_ );
nand g0143 ( new_n281_, new_n193_, new_n280_ );
nor g0144 ( new_n282_, new_n281_, new_n277_ );
nor g0145 ( new_n283_, new_n279_, new_n282_ );
nor g0146 ( new_n284_, new_n250_, new_n164_ );
nor g0147 ( new_n285_, new_n165_, new_n249_ );
nor g0148 ( new_n286_, new_n284_, new_n285_ );
not g0149 ( new_n287_, new_n286_ );
nand g0150 ( new_n288_, N132, N137 );
nand g0151 ( new_n289_, new_n287_, new_n288_ );
not g0152 ( new_n290_, new_n289_ );
nor g0153 ( new_n291_, new_n287_, new_n288_ );
nor g0154 ( new_n292_, new_n290_, new_n291_ );
not g0155 ( new_n293_, keyIn_0_15 );
not g0156 ( new_n294_, N45 );
nor g0157 ( new_n295_, new_n294_, N61 );
not g0158 ( new_n296_, N61 );
nor g0159 ( new_n297_, new_n296_, N45 );
nor g0160 ( new_n298_, new_n295_, new_n297_ );
nand g0161 ( new_n299_, N13, N29 );
not g0162 ( new_n300_, new_n299_ );
nor g0163 ( new_n301_, N13, N29 );
nor g0164 ( new_n302_, new_n300_, new_n301_ );
nor g0165 ( new_n303_, new_n298_, new_n302_ );
nand g0166 ( new_n304_, new_n298_, new_n302_ );
not g0167 ( new_n305_, new_n304_ );
nor g0168 ( new_n306_, new_n305_, new_n303_ );
nor g0169 ( new_n307_, new_n306_, new_n293_ );
nand g0170 ( new_n308_, new_n306_, new_n293_ );
not g0171 ( new_n309_, new_n308_ );
nor g0172 ( new_n310_, new_n309_, new_n307_ );
nor g0173 ( new_n311_, new_n292_, new_n310_ );
nand g0174 ( new_n312_, new_n292_, new_n310_ );
not g0175 ( new_n313_, new_n312_ );
nor g0176 ( new_n314_, new_n313_, new_n311_ );
nor g0177 ( new_n315_, new_n283_, new_n314_ );
not g0178 ( new_n316_, new_n314_ );
nor g0179 ( new_n317_, new_n316_, new_n276_ );
not g0180 ( new_n318_, new_n317_ );
nor g0181 ( new_n319_, new_n318_, new_n281_ );
nor g0182 ( new_n320_, new_n315_, new_n319_ );
not g0183 ( new_n321_, keyIn_0_3 );
nand g0184 ( new_n322_, N25, N29 );
not g0185 ( new_n323_, new_n322_ );
nor g0186 ( new_n324_, N25, N29 );
nor g0187 ( new_n325_, new_n323_, new_n324_ );
nand g0188 ( new_n326_, new_n325_, new_n321_ );
not g0189 ( new_n327_, new_n324_ );
nand g0190 ( new_n328_, new_n327_, new_n322_ );
nand g0191 ( new_n329_, new_n328_, keyIn_0_3 );
nand g0192 ( new_n330_, new_n329_, new_n326_ );
nand g0193 ( new_n331_, N17, N21 );
not g0194 ( new_n332_, N17 );
not g0195 ( new_n333_, N21 );
nand g0196 ( new_n334_, new_n332_, new_n333_ );
nand g0197 ( new_n335_, new_n334_, new_n331_ );
nand g0198 ( new_n336_, new_n335_, keyIn_0_2 );
not g0199 ( new_n337_, keyIn_0_2 );
not g0200 ( new_n338_, new_n331_ );
nor g0201 ( new_n339_, N17, N21 );
nor g0202 ( new_n340_, new_n338_, new_n339_ );
nand g0203 ( new_n341_, new_n340_, new_n337_ );
nand g0204 ( new_n342_, new_n341_, new_n336_ );
nor g0205 ( new_n343_, new_n330_, new_n342_ );
not g0206 ( new_n344_, keyIn_0_13 );
nand g0207 ( new_n345_, new_n330_, new_n342_ );
nand g0208 ( new_n346_, new_n345_, new_n344_ );
nor g0209 ( new_n347_, new_n346_, new_n343_ );
not g0210 ( new_n348_, new_n347_ );
not g0211 ( new_n349_, new_n330_ );
not g0212 ( new_n350_, new_n342_ );
nand g0213 ( new_n351_, new_n349_, new_n350_ );
nand g0214 ( new_n352_, new_n351_, new_n345_ );
nand g0215 ( new_n353_, new_n352_, keyIn_0_13 );
nand g0216 ( new_n354_, new_n348_, new_n353_ );
nand g0217 ( new_n355_, N57, N61 );
not g0218 ( new_n356_, new_n355_ );
nor g0219 ( new_n357_, N57, N61 );
nor g0220 ( new_n358_, new_n356_, new_n357_ );
nand g0221 ( new_n359_, N49, N53 );
not g0222 ( new_n360_, new_n359_ );
nor g0223 ( new_n361_, N49, N53 );
nor g0224 ( new_n362_, new_n360_, new_n361_ );
nor g0225 ( new_n363_, new_n358_, new_n362_ );
nand g0226 ( new_n364_, new_n358_, new_n362_ );
not g0227 ( new_n365_, new_n364_ );
nor g0228 ( new_n366_, new_n365_, new_n363_ );
not g0229 ( new_n367_, new_n366_ );
nand g0230 ( new_n368_, new_n354_, new_n367_ );
not g0231 ( new_n369_, new_n368_ );
nor g0232 ( new_n370_, new_n354_, new_n367_ );
nor g0233 ( new_n371_, new_n369_, new_n370_ );
nand g0234 ( new_n372_, N136, N137 );
not g0235 ( new_n373_, new_n372_ );
nor g0236 ( new_n374_, new_n371_, new_n373_ );
nand g0237 ( new_n375_, new_n371_, new_n373_ );
not g0238 ( new_n376_, new_n375_ );
nor g0239 ( new_n377_, new_n376_, new_n374_ );
nand g0240 ( new_n378_, N109, N125 );
not g0241 ( new_n379_, new_n378_ );
nor g0242 ( new_n380_, N109, N125 );
nor g0243 ( new_n381_, new_n379_, new_n380_ );
nand g0244 ( new_n382_, N77, N93 );
not g0245 ( new_n383_, new_n382_ );
nor g0246 ( new_n384_, N77, N93 );
nor g0247 ( new_n385_, new_n383_, new_n384_ );
nor g0248 ( new_n386_, new_n381_, new_n385_ );
nand g0249 ( new_n387_, new_n381_, new_n385_ );
not g0250 ( new_n388_, new_n387_ );
nor g0251 ( new_n389_, new_n388_, new_n386_ );
nor g0252 ( new_n390_, new_n377_, new_n389_ );
nand g0253 ( new_n391_, new_n377_, new_n389_ );
not g0254 ( new_n392_, new_n391_ );
nor g0255 ( new_n393_, new_n392_, new_n390_ );
not g0256 ( new_n394_, keyIn_0_17 );
nor g0257 ( new_n395_, new_n139_, N89 );
nor g0258 ( new_n396_, new_n152_, N73 );
nor g0259 ( new_n397_, new_n395_, new_n396_ );
not g0260 ( new_n398_, new_n397_ );
nand g0261 ( new_n399_, new_n398_, keyIn_0_10 );
not g0262 ( new_n400_, new_n399_ );
nor g0263 ( new_n401_, new_n398_, keyIn_0_10 );
nor g0264 ( new_n402_, new_n400_, new_n401_ );
nor g0265 ( new_n403_, new_n194_, N121 );
nor g0266 ( new_n404_, new_n237_, N105 );
nor g0267 ( new_n405_, new_n403_, new_n404_ );
not g0268 ( new_n406_, new_n405_ );
nand g0269 ( new_n407_, new_n406_, keyIn_0_11 );
not g0270 ( new_n408_, new_n407_ );
nor g0271 ( new_n409_, new_n406_, keyIn_0_11 );
nor g0272 ( new_n410_, new_n408_, new_n409_ );
nor g0273 ( new_n411_, new_n402_, new_n410_ );
nand g0274 ( new_n412_, new_n402_, new_n410_ );
not g0275 ( new_n413_, new_n412_ );
nor g0276 ( new_n414_, new_n413_, new_n411_ );
not g0277 ( new_n415_, new_n414_ );
nand g0278 ( new_n416_, new_n415_, new_n394_ );
not g0279 ( new_n417_, new_n416_ );
nor g0280 ( new_n418_, new_n415_, new_n394_ );
nor g0281 ( new_n419_, new_n417_, new_n418_ );
not g0282 ( new_n420_, new_n419_ );
not g0283 ( new_n421_, keyIn_0_7 );
nand g0284 ( new_n422_, N135, N137 );
nand g0285 ( new_n423_, new_n422_, new_n421_ );
not g0286 ( new_n424_, new_n423_ );
nor g0287 ( new_n425_, new_n422_, new_n421_ );
nor g0288 ( new_n426_, new_n424_, new_n425_ );
not g0289 ( new_n427_, new_n426_ );
not g0290 ( new_n428_, keyIn_0_5 );
nand g0291 ( new_n429_, new_n294_, N41 );
nand g0292 ( new_n430_, new_n217_, N45 );
nand g0293 ( new_n431_, new_n429_, new_n430_ );
nor g0294 ( new_n432_, new_n431_, new_n428_ );
nand g0295 ( new_n433_, new_n431_, new_n428_ );
not g0296 ( new_n434_, new_n433_ );
nor g0297 ( new_n435_, new_n434_, new_n432_ );
not g0298 ( new_n436_, keyIn_0_4 );
nand g0299 ( new_n437_, N33, N37 );
not g0300 ( new_n438_, new_n437_ );
nor g0301 ( new_n439_, N33, N37 );
nor g0302 ( new_n440_, new_n438_, new_n439_ );
nor g0303 ( new_n441_, new_n440_, new_n436_ );
nand g0304 ( new_n442_, new_n176_, new_n260_ );
nand g0305 ( new_n443_, new_n442_, new_n437_ );
nor g0306 ( new_n444_, new_n443_, keyIn_0_4 );
nor g0307 ( new_n445_, new_n441_, new_n444_ );
nor g0308 ( new_n446_, new_n435_, new_n445_ );
not g0309 ( new_n447_, new_n431_ );
nand g0310 ( new_n448_, new_n447_, keyIn_0_5 );
nand g0311 ( new_n449_, new_n448_, new_n433_ );
nand g0312 ( new_n450_, new_n443_, keyIn_0_4 );
nand g0313 ( new_n451_, new_n440_, new_n436_ );
nand g0314 ( new_n452_, new_n451_, new_n450_ );
nor g0315 ( new_n453_, new_n449_, new_n452_ );
nor g0316 ( new_n454_, new_n446_, new_n453_ );
nor g0317 ( new_n455_, new_n454_, keyIn_0_14 );
nand g0318 ( new_n456_, new_n449_, new_n452_ );
nand g0319 ( new_n457_, new_n456_, keyIn_0_14 );
nor g0320 ( new_n458_, new_n457_, new_n453_ );
nor g0321 ( new_n459_, new_n455_, new_n458_ );
nand g0322 ( new_n460_, N1, N5 );
not g0323 ( new_n461_, new_n460_ );
nor g0324 ( new_n462_, N1, N5 );
nor g0325 ( new_n463_, new_n461_, new_n462_ );
nor g0326 ( new_n464_, new_n463_, keyIn_0_0 );
not g0327 ( new_n465_, keyIn_0_0 );
not g0328 ( new_n466_, N5 );
nand g0329 ( new_n467_, new_n138_, new_n466_ );
nand g0330 ( new_n468_, new_n467_, new_n460_ );
nor g0331 ( new_n469_, new_n468_, new_n465_ );
nor g0332 ( new_n470_, new_n464_, new_n469_ );
not g0333 ( new_n471_, keyIn_0_1 );
nand g0334 ( new_n472_, N9, N13 );
not g0335 ( new_n473_, new_n472_ );
nor g0336 ( new_n474_, N9, N13 );
nor g0337 ( new_n475_, new_n473_, new_n474_ );
nor g0338 ( new_n476_, new_n475_, new_n471_ );
not g0339 ( new_n477_, N9 );
not g0340 ( new_n478_, N13 );
nand g0341 ( new_n479_, new_n477_, new_n478_ );
nand g0342 ( new_n480_, new_n479_, new_n472_ );
nor g0343 ( new_n481_, new_n480_, keyIn_0_1 );
nor g0344 ( new_n482_, new_n476_, new_n481_ );
nand g0345 ( new_n483_, new_n470_, new_n482_ );
nand g0346 ( new_n484_, new_n468_, new_n465_ );
nand g0347 ( new_n485_, new_n463_, keyIn_0_0 );
nand g0348 ( new_n486_, new_n485_, new_n484_ );
nand g0349 ( new_n487_, new_n480_, keyIn_0_1 );
nand g0350 ( new_n488_, new_n475_, new_n471_ );
nand g0351 ( new_n489_, new_n488_, new_n487_ );
nand g0352 ( new_n490_, new_n486_, new_n489_ );
nand g0353 ( new_n491_, new_n483_, new_n490_ );
nand g0354 ( new_n492_, new_n491_, keyIn_0_12 );
nor g0355 ( new_n493_, new_n486_, new_n489_ );
nor g0356 ( new_n494_, new_n493_, keyIn_0_12 );
nand g0357 ( new_n495_, new_n494_, new_n490_ );
nand g0358 ( new_n496_, new_n495_, new_n492_ );
not g0359 ( new_n497_, new_n496_ );
nand g0360 ( new_n498_, new_n459_, new_n497_ );
not g0361 ( new_n499_, keyIn_0_14 );
nand g0362 ( new_n500_, new_n435_, new_n445_ );
nand g0363 ( new_n501_, new_n500_, new_n456_ );
nand g0364 ( new_n502_, new_n501_, new_n499_ );
not g0365 ( new_n503_, new_n458_ );
nand g0366 ( new_n504_, new_n503_, new_n502_ );
nand g0367 ( new_n505_, new_n504_, new_n496_ );
nand g0368 ( new_n506_, new_n498_, new_n505_ );
nand g0369 ( new_n507_, new_n506_, keyIn_0_19 );
not g0370 ( new_n508_, keyIn_0_19 );
not g0371 ( new_n509_, keyIn_0_12 );
not g0372 ( new_n510_, new_n490_ );
nor g0373 ( new_n511_, new_n510_, new_n493_ );
nand g0374 ( new_n512_, new_n511_, new_n509_ );
nand g0375 ( new_n513_, new_n512_, new_n492_ );
nand g0376 ( new_n514_, new_n459_, new_n513_ );
nand g0377 ( new_n515_, new_n454_, keyIn_0_14 );
nand g0378 ( new_n516_, new_n515_, new_n502_ );
nand g0379 ( new_n517_, new_n497_, new_n516_ );
nand g0380 ( new_n518_, new_n514_, new_n517_ );
nand g0381 ( new_n519_, new_n518_, new_n508_ );
nand g0382 ( new_n520_, new_n507_, new_n519_ );
nand g0383 ( new_n521_, new_n520_, new_n427_ );
not g0384 ( new_n522_, new_n520_ );
nand g0385 ( new_n523_, new_n522_, new_n426_ );
nand g0386 ( new_n524_, new_n523_, new_n521_ );
nand g0387 ( new_n525_, new_n524_, keyIn_0_21 );
not g0388 ( new_n526_, keyIn_0_21 );
nor g0389 ( new_n527_, new_n520_, new_n427_ );
not g0390 ( new_n528_, new_n519_ );
nor g0391 ( new_n529_, new_n518_, new_n508_ );
nor g0392 ( new_n530_, new_n528_, new_n529_ );
nor g0393 ( new_n531_, new_n530_, new_n426_ );
nor g0394 ( new_n532_, new_n531_, new_n527_ );
nand g0395 ( new_n533_, new_n532_, new_n526_ );
nand g0396 ( new_n534_, new_n533_, new_n525_ );
nand g0397 ( new_n535_, new_n534_, new_n420_ );
not g0398 ( new_n536_, new_n492_ );
nor g0399 ( new_n537_, new_n491_, keyIn_0_12 );
nor g0400 ( new_n538_, new_n536_, new_n537_ );
nor g0401 ( new_n539_, new_n538_, new_n504_ );
nor g0402 ( new_n540_, new_n501_, new_n499_ );
nor g0403 ( new_n541_, new_n455_, new_n540_ );
nor g0404 ( new_n542_, new_n541_, new_n496_ );
nor g0405 ( new_n543_, new_n539_, new_n542_ );
nand g0406 ( new_n544_, new_n543_, keyIn_0_19 );
nand g0407 ( new_n545_, new_n544_, new_n519_ );
nand g0408 ( new_n546_, new_n545_, new_n427_ );
nand g0409 ( new_n547_, new_n523_, new_n546_ );
nand g0410 ( new_n548_, new_n547_, keyIn_0_21 );
nor g0411 ( new_n549_, new_n547_, keyIn_0_21 );
nor g0412 ( new_n550_, new_n549_, new_n420_ );
nand g0413 ( new_n551_, new_n550_, new_n548_ );
nand g0414 ( new_n552_, new_n535_, new_n551_ );
nand g0415 ( new_n553_, new_n552_, keyIn_0_23 );
not g0416 ( new_n554_, keyIn_0_23 );
not g0417 ( new_n555_, new_n521_ );
nor g0418 ( new_n556_, new_n555_, new_n527_ );
nor g0419 ( new_n557_, new_n556_, new_n526_ );
nor g0420 ( new_n558_, new_n557_, new_n549_ );
nor g0421 ( new_n559_, new_n558_, new_n419_ );
not g0422 ( new_n560_, new_n548_ );
nand g0423 ( new_n561_, new_n533_, new_n419_ );
nor g0424 ( new_n562_, new_n561_, new_n560_ );
nor g0425 ( new_n563_, new_n559_, new_n562_ );
nand g0426 ( new_n564_, new_n563_, new_n554_ );
nand g0427 ( new_n565_, new_n564_, new_n553_ );
nand g0428 ( new_n566_, new_n565_, new_n393_ );
nor g0429 ( new_n567_, new_n566_, new_n320_ );
not g0430 ( new_n568_, new_n567_ );
not g0431 ( new_n569_, keyIn_0_22 );
not g0432 ( new_n570_, keyIn_0_16 );
not g0433 ( new_n571_, N65 );
nor g0434 ( new_n572_, new_n571_, N81 );
not g0435 ( new_n573_, N81 );
nor g0436 ( new_n574_, new_n573_, N65 );
nor g0437 ( new_n575_, new_n572_, new_n574_ );
not g0438 ( new_n576_, new_n575_ );
nand g0439 ( new_n577_, new_n576_, keyIn_0_8 );
not g0440 ( new_n578_, new_n577_ );
nor g0441 ( new_n579_, new_n576_, keyIn_0_8 );
nor g0442 ( new_n580_, new_n578_, new_n579_ );
not g0443 ( new_n581_, keyIn_0_9 );
nand g0444 ( new_n582_, N97, N113 );
not g0445 ( new_n583_, new_n582_ );
nor g0446 ( new_n584_, N97, N113 );
nor g0447 ( new_n585_, new_n583_, new_n584_ );
nor g0448 ( new_n586_, new_n585_, new_n581_ );
nand g0449 ( new_n587_, new_n585_, new_n581_ );
not g0450 ( new_n588_, new_n587_ );
nor g0451 ( new_n589_, new_n588_, new_n586_ );
nor g0452 ( new_n590_, new_n580_, new_n589_ );
nand g0453 ( new_n591_, new_n580_, new_n589_ );
not g0454 ( new_n592_, new_n591_ );
nor g0455 ( new_n593_, new_n592_, new_n590_ );
nor g0456 ( new_n594_, new_n593_, new_n570_ );
nand g0457 ( new_n595_, new_n593_, new_n570_ );
not g0458 ( new_n596_, new_n595_ );
nor g0459 ( new_n597_, new_n596_, new_n594_ );
not g0460 ( new_n598_, keyIn_0_20 );
not g0461 ( new_n599_, keyIn_0_6 );
nand g0462 ( new_n600_, N133, N137 );
nand g0463 ( new_n601_, new_n600_, new_n599_ );
not g0464 ( new_n602_, new_n601_ );
nor g0465 ( new_n603_, new_n600_, new_n599_ );
nor g0466 ( new_n604_, new_n602_, new_n603_ );
not g0467 ( new_n605_, new_n604_ );
not g0468 ( new_n606_, keyIn_0_18 );
nand g0469 ( new_n607_, new_n513_, new_n354_ );
not g0470 ( new_n608_, new_n345_ );
nor g0471 ( new_n609_, new_n608_, new_n343_ );
nor g0472 ( new_n610_, new_n609_, new_n344_ );
nor g0473 ( new_n611_, new_n610_, new_n347_ );
nand g0474 ( new_n612_, new_n611_, new_n538_ );
nand g0475 ( new_n613_, new_n612_, new_n607_ );
nand g0476 ( new_n614_, new_n613_, new_n606_ );
nand g0477 ( new_n615_, new_n497_, new_n354_ );
nor g0478 ( new_n616_, new_n352_, keyIn_0_13 );
nor g0479 ( new_n617_, new_n610_, new_n616_ );
nand g0480 ( new_n618_, new_n617_, new_n513_ );
nand g0481 ( new_n619_, new_n618_, new_n615_ );
nand g0482 ( new_n620_, new_n619_, keyIn_0_18 );
nand g0483 ( new_n621_, new_n614_, new_n620_ );
nand g0484 ( new_n622_, new_n621_, new_n605_ );
not g0485 ( new_n623_, new_n622_ );
nor g0486 ( new_n624_, new_n621_, new_n605_ );
nor g0487 ( new_n625_, new_n623_, new_n624_ );
nor g0488 ( new_n626_, new_n625_, new_n598_ );
not g0489 ( new_n627_, new_n621_ );
nand g0490 ( new_n628_, new_n627_, new_n604_ );
not g0491 ( new_n629_, new_n619_ );
nand g0492 ( new_n630_, new_n629_, new_n606_ );
nand g0493 ( new_n631_, new_n630_, new_n620_ );
nand g0494 ( new_n632_, new_n631_, new_n605_ );
nand g0495 ( new_n633_, new_n628_, new_n632_ );
nor g0496 ( new_n634_, new_n633_, keyIn_0_20 );
nor g0497 ( new_n635_, new_n626_, new_n634_ );
nand g0498 ( new_n636_, new_n635_, new_n597_ );
not g0499 ( new_n637_, new_n597_ );
not g0500 ( new_n638_, new_n620_ );
nor g0501 ( new_n639_, new_n619_, keyIn_0_18 );
nor g0502 ( new_n640_, new_n638_, new_n639_ );
nor g0503 ( new_n641_, new_n640_, new_n604_ );
nor g0504 ( new_n642_, new_n641_, new_n624_ );
nand g0505 ( new_n643_, new_n642_, new_n598_ );
nand g0506 ( new_n644_, new_n633_, keyIn_0_20 );
nand g0507 ( new_n645_, new_n643_, new_n644_ );
nand g0508 ( new_n646_, new_n645_, new_n637_ );
nand g0509 ( new_n647_, new_n636_, new_n646_ );
nor g0510 ( new_n648_, new_n647_, new_n569_ );
nand g0511 ( new_n649_, new_n647_, new_n569_ );
not g0512 ( new_n650_, new_n649_ );
nor g0513 ( new_n651_, new_n650_, new_n648_ );
nor g0514 ( new_n652_, new_n541_, new_n366_ );
nor g0515 ( new_n653_, new_n516_, new_n367_ );
nor g0516 ( new_n654_, new_n652_, new_n653_ );
nand g0517 ( new_n655_, N134, N137 );
not g0518 ( new_n656_, new_n655_ );
nor g0519 ( new_n657_, new_n654_, new_n656_ );
nand g0520 ( new_n658_, new_n654_, new_n656_ );
not g0521 ( new_n659_, new_n658_ );
nor g0522 ( new_n660_, new_n659_, new_n657_ );
not g0523 ( new_n661_, N101 );
nor g0524 ( new_n662_, new_n661_, N117 );
not g0525 ( new_n663_, N117 );
nor g0526 ( new_n664_, new_n663_, N101 );
nor g0527 ( new_n665_, new_n662_, new_n664_ );
nand g0528 ( new_n666_, N69, N85 );
not g0529 ( new_n667_, new_n666_ );
nor g0530 ( new_n668_, N69, N85 );
nor g0531 ( new_n669_, new_n667_, new_n668_ );
nor g0532 ( new_n670_, new_n665_, new_n669_ );
nand g0533 ( new_n671_, new_n665_, new_n669_ );
not g0534 ( new_n672_, new_n671_ );
nor g0535 ( new_n673_, new_n672_, new_n670_ );
nor g0536 ( new_n674_, new_n660_, new_n673_ );
nand g0537 ( new_n675_, new_n660_, new_n673_ );
not g0538 ( new_n676_, new_n675_ );
nor g0539 ( new_n677_, new_n676_, new_n674_ );
not g0540 ( new_n678_, new_n677_ );
nand g0541 ( new_n679_, new_n651_, new_n678_ );
nor g0542 ( new_n680_, new_n568_, new_n679_ );
not g0543 ( new_n681_, new_n680_ );
nor g0544 ( new_n682_, new_n681_, new_n193_ );
nand g0545 ( new_n683_, new_n682_, new_n138_ );
not g0546 ( new_n684_, new_n682_ );
nand g0547 ( new_n685_, new_n684_, N1 );
nand g0548 ( N724, new_n685_, new_n683_ );
nor g0549 ( new_n687_, new_n681_, new_n277_ );
nand g0550 ( new_n688_, new_n687_, new_n466_ );
not g0551 ( new_n689_, new_n687_ );
nand g0552 ( new_n690_, new_n689_, N5 );
nand g0553 ( N725, new_n690_, new_n688_ );
nor g0554 ( new_n692_, new_n681_, new_n280_ );
nand g0555 ( new_n693_, new_n692_, new_n477_ );
not g0556 ( new_n694_, new_n692_ );
nand g0557 ( new_n695_, new_n694_, N9 );
nand g0558 ( N726, new_n695_, new_n693_ );
nor g0559 ( new_n697_, new_n681_, new_n316_ );
nand g0560 ( new_n698_, new_n697_, new_n478_ );
not g0561 ( new_n699_, new_n697_ );
nand g0562 ( new_n700_, new_n699_, N13 );
nand g0563 ( N727, new_n700_, new_n698_ );
not g0564 ( new_n702_, new_n320_ );
not g0565 ( new_n703_, new_n393_ );
nand g0566 ( new_n704_, new_n702_, new_n703_ );
nor g0567 ( new_n705_, new_n704_, new_n565_ );
not g0568 ( new_n706_, new_n705_ );
nor g0569 ( new_n707_, new_n706_, new_n679_ );
not g0570 ( new_n708_, new_n707_ );
nor g0571 ( new_n709_, new_n708_, new_n193_ );
nand g0572 ( new_n710_, new_n709_, new_n332_ );
not g0573 ( new_n711_, new_n709_ );
nand g0574 ( new_n712_, new_n711_, N17 );
nand g0575 ( N728, new_n712_, new_n710_ );
nor g0576 ( new_n714_, new_n708_, new_n277_ );
nand g0577 ( new_n715_, new_n714_, new_n333_ );
not g0578 ( new_n716_, new_n714_ );
nand g0579 ( new_n717_, new_n716_, N21 );
nand g0580 ( N729, new_n717_, new_n715_ );
not g0581 ( new_n719_, N25 );
nor g0582 ( new_n720_, new_n708_, new_n280_ );
nand g0583 ( new_n721_, new_n720_, new_n719_ );
not g0584 ( new_n722_, new_n720_ );
nand g0585 ( new_n723_, new_n722_, N25 );
nand g0586 ( N730, new_n723_, new_n721_ );
not g0587 ( new_n725_, N29 );
nor g0588 ( new_n726_, new_n708_, new_n316_ );
nand g0589 ( new_n727_, new_n726_, new_n725_ );
not g0590 ( new_n728_, new_n726_ );
nand g0591 ( new_n729_, new_n728_, N29 );
nand g0592 ( N731, new_n729_, new_n727_ );
nor g0593 ( new_n731_, new_n651_, new_n678_ );
not g0594 ( new_n732_, new_n731_ );
nor g0595 ( new_n733_, new_n568_, new_n732_ );
not g0596 ( new_n734_, new_n733_ );
nor g0597 ( new_n735_, new_n734_, new_n193_ );
not g0598 ( new_n736_, new_n735_ );
nand g0599 ( new_n737_, new_n736_, N33 );
nand g0600 ( new_n738_, new_n735_, new_n176_ );
nand g0601 ( N732, new_n737_, new_n738_ );
nor g0602 ( new_n740_, new_n734_, new_n277_ );
not g0603 ( new_n741_, new_n740_ );
nand g0604 ( new_n742_, new_n741_, N37 );
nand g0605 ( new_n743_, new_n740_, new_n260_ );
nand g0606 ( N733, new_n742_, new_n743_ );
nor g0607 ( new_n745_, new_n734_, new_n280_ );
not g0608 ( new_n746_, new_n745_ );
nand g0609 ( new_n747_, new_n746_, N41 );
nand g0610 ( new_n748_, new_n745_, new_n217_ );
nand g0611 ( N734, new_n747_, new_n748_ );
nor g0612 ( new_n750_, new_n734_, new_n316_ );
not g0613 ( new_n751_, new_n750_ );
nand g0614 ( new_n752_, new_n751_, N45 );
nand g0615 ( new_n753_, new_n750_, new_n294_ );
nand g0616 ( N735, new_n752_, new_n753_ );
nor g0617 ( new_n755_, new_n706_, new_n732_ );
not g0618 ( new_n756_, new_n755_ );
nor g0619 ( new_n757_, new_n756_, new_n193_ );
not g0620 ( new_n758_, new_n757_ );
nand g0621 ( new_n759_, new_n758_, N49 );
nand g0622 ( new_n760_, new_n757_, new_n178_ );
nand g0623 ( N736, new_n759_, new_n760_ );
nor g0624 ( new_n762_, new_n756_, new_n277_ );
not g0625 ( new_n763_, new_n762_ );
nand g0626 ( new_n764_, new_n763_, N53 );
nand g0627 ( new_n765_, new_n762_, new_n262_ );
nand g0628 ( N737, new_n764_, new_n765_ );
nor g0629 ( new_n767_, new_n756_, new_n280_ );
not g0630 ( new_n768_, new_n767_ );
nand g0631 ( new_n769_, new_n768_, N57 );
nand g0632 ( new_n770_, new_n767_, new_n219_ );
nand g0633 ( N738, new_n769_, new_n770_ );
nor g0634 ( new_n772_, new_n756_, new_n316_ );
not g0635 ( new_n773_, new_n772_ );
nand g0636 ( new_n774_, new_n773_, N61 );
nand g0637 ( new_n775_, new_n772_, new_n296_ );
nand g0638 ( N739, new_n774_, new_n775_ );
not g0639 ( new_n777_, keyIn_0_52 );
not g0640 ( new_n778_, keyIn_0_40 );
nor g0641 ( new_n779_, new_n635_, new_n597_ );
nand g0642 ( new_n780_, new_n636_, keyIn_0_22 );
nor g0643 ( new_n781_, new_n780_, new_n779_ );
nor g0644 ( new_n782_, new_n650_, new_n781_ );
not g0645 ( new_n783_, keyIn_0_37 );
not g0646 ( new_n784_, keyIn_0_31 );
not g0647 ( new_n785_, new_n553_ );
nor g0648 ( new_n786_, new_n552_, keyIn_0_23 );
nor g0649 ( new_n787_, new_n785_, new_n786_ );
nor g0650 ( new_n788_, new_n787_, new_n784_ );
nor g0651 ( new_n789_, new_n565_, keyIn_0_31 );
nor g0652 ( new_n790_, new_n788_, new_n789_ );
nor g0653 ( new_n791_, new_n679_, new_n703_ );
nand g0654 ( new_n792_, new_n790_, new_n791_ );
nand g0655 ( new_n793_, new_n792_, keyIn_0_35 );
not g0656 ( new_n794_, new_n793_ );
nand g0657 ( new_n795_, new_n565_, keyIn_0_31 );
nand g0658 ( new_n796_, new_n787_, new_n784_ );
nand g0659 ( new_n797_, new_n796_, new_n795_ );
not g0660 ( new_n798_, keyIn_0_35 );
nand g0661 ( new_n799_, new_n393_, new_n798_ );
nor g0662 ( new_n800_, new_n799_, new_n677_ );
nand g0663 ( new_n801_, new_n782_, new_n800_ );
nor g0664 ( new_n802_, new_n797_, new_n801_ );
nor g0665 ( new_n803_, new_n794_, new_n802_ );
not g0666 ( new_n804_, keyIn_0_36 );
not g0667 ( new_n805_, keyIn_0_33 );
nor g0668 ( new_n806_, new_n566_, new_n677_ );
nor g0669 ( new_n807_, new_n651_, keyIn_0_28 );
not g0670 ( new_n808_, keyIn_0_28 );
not g0671 ( new_n809_, new_n781_ );
nand g0672 ( new_n810_, new_n809_, new_n649_ );
nor g0673 ( new_n811_, new_n810_, new_n808_ );
nor g0674 ( new_n812_, new_n807_, new_n811_ );
nand g0675 ( new_n813_, new_n812_, new_n806_ );
nand g0676 ( new_n814_, new_n813_, new_n805_ );
nor g0677 ( new_n815_, new_n787_, new_n703_ );
nand g0678 ( new_n816_, new_n815_, new_n678_ );
not g0679 ( new_n817_, new_n647_ );
nand g0680 ( new_n818_, new_n817_, keyIn_0_22 );
nand g0681 ( new_n819_, new_n818_, new_n649_ );
nand g0682 ( new_n820_, new_n819_, new_n808_ );
nand g0683 ( new_n821_, new_n782_, keyIn_0_28 );
nand g0684 ( new_n822_, new_n821_, new_n820_ );
nor g0685 ( new_n823_, new_n816_, new_n822_ );
nand g0686 ( new_n824_, new_n823_, keyIn_0_33 );
nand g0687 ( new_n825_, new_n814_, new_n824_ );
nand g0688 ( new_n826_, new_n825_, new_n804_ );
nor g0689 ( new_n827_, new_n826_, new_n803_ );
not g0690 ( new_n828_, keyIn_0_34 );
nand g0691 ( new_n829_, new_n819_, keyIn_0_29 );
not g0692 ( new_n830_, new_n829_ );
nor g0693 ( new_n831_, new_n819_, keyIn_0_29 );
nor g0694 ( new_n832_, new_n830_, new_n831_ );
not g0695 ( new_n833_, keyIn_0_30 );
nor g0696 ( new_n834_, new_n787_, new_n833_ );
not g0697 ( new_n835_, new_n834_ );
nor g0698 ( new_n836_, new_n565_, keyIn_0_30 );
nor g0699 ( new_n837_, new_n678_, new_n703_ );
not g0700 ( new_n838_, new_n837_ );
nor g0701 ( new_n839_, new_n836_, new_n838_ );
nand g0702 ( new_n840_, new_n839_, new_n835_ );
nor g0703 ( new_n841_, new_n840_, new_n832_ );
nor g0704 ( new_n842_, new_n841_, new_n828_ );
not g0705 ( new_n843_, new_n831_ );
nand g0706 ( new_n844_, new_n843_, new_n829_ );
nand g0707 ( new_n845_, new_n787_, new_n833_ );
nand g0708 ( new_n846_, new_n845_, new_n837_ );
nor g0709 ( new_n847_, new_n846_, new_n834_ );
nand g0710 ( new_n848_, new_n847_, new_n844_ );
nor g0711 ( new_n849_, new_n848_, keyIn_0_34 );
nor g0712 ( new_n850_, new_n842_, new_n849_ );
not g0713 ( new_n851_, keyIn_0_32 );
not g0714 ( new_n852_, keyIn_0_27 );
nor g0715 ( new_n853_, new_n787_, new_n852_ );
nor g0716 ( new_n854_, new_n565_, keyIn_0_27 );
nor g0717 ( new_n855_, new_n853_, new_n854_ );
nand g0718 ( new_n856_, new_n810_, keyIn_0_25 );
nor g0719 ( new_n857_, new_n810_, keyIn_0_25 );
nor g0720 ( new_n858_, new_n677_, keyIn_0_26 );
nand g0721 ( new_n859_, new_n677_, keyIn_0_26 );
nand g0722 ( new_n860_, new_n859_, new_n703_ );
nor g0723 ( new_n861_, new_n860_, new_n858_ );
not g0724 ( new_n862_, new_n861_ );
nor g0725 ( new_n863_, new_n857_, new_n862_ );
nand g0726 ( new_n864_, new_n863_, new_n856_ );
nor g0727 ( new_n865_, new_n864_, new_n855_ );
not g0728 ( new_n866_, new_n865_ );
nand g0729 ( new_n867_, new_n866_, new_n851_ );
nand g0730 ( new_n868_, new_n865_, keyIn_0_32 );
nand g0731 ( new_n869_, new_n867_, new_n868_ );
nor g0732 ( new_n870_, new_n869_, new_n850_ );
nand g0733 ( new_n871_, new_n870_, new_n827_ );
nor g0734 ( new_n872_, new_n865_, keyIn_0_32 );
not g0735 ( new_n873_, new_n868_ );
nor g0736 ( new_n874_, new_n873_, new_n872_ );
nor g0737 ( new_n875_, new_n819_, new_n677_ );
nand g0738 ( new_n876_, new_n875_, new_n393_ );
nor g0739 ( new_n877_, new_n876_, new_n797_ );
nand g0740 ( new_n878_, new_n877_, new_n798_ );
nand g0741 ( new_n879_, new_n793_, new_n878_ );
nand g0742 ( new_n880_, new_n825_, new_n879_ );
nor g0743 ( new_n881_, new_n850_, new_n880_ );
nand g0744 ( new_n882_, new_n881_, new_n874_ );
nand g0745 ( new_n883_, new_n882_, keyIn_0_36 );
nand g0746 ( new_n884_, new_n883_, new_n871_ );
nand g0747 ( new_n885_, new_n277_, new_n192_ );
nand g0748 ( new_n886_, new_n316_, new_n233_ );
nor g0749 ( new_n887_, new_n885_, new_n886_ );
nand g0750 ( new_n888_, new_n884_, new_n887_ );
nand g0751 ( new_n889_, new_n888_, new_n783_ );
not g0752 ( new_n890_, new_n889_ );
nor g0753 ( new_n891_, new_n888_, new_n783_ );
nor g0754 ( new_n892_, new_n890_, new_n891_ );
nand g0755 ( new_n893_, new_n892_, new_n782_ );
nand g0756 ( new_n894_, new_n893_, new_n778_ );
not g0757 ( new_n895_, new_n888_ );
nand g0758 ( new_n896_, new_n895_, keyIn_0_37 );
nand g0759 ( new_n897_, new_n896_, new_n889_ );
nor g0760 ( new_n898_, new_n897_, new_n810_ );
nand g0761 ( new_n899_, new_n898_, keyIn_0_40 );
nand g0762 ( new_n900_, new_n894_, new_n899_ );
nand g0763 ( new_n901_, new_n900_, new_n571_ );
nand g0764 ( new_n902_, new_n889_, new_n651_ );
nor g0765 ( new_n903_, new_n902_, new_n891_ );
nor g0766 ( new_n904_, new_n903_, keyIn_0_40 );
not g0767 ( new_n905_, new_n904_ );
nand g0768 ( new_n906_, new_n905_, new_n899_ );
not g0769 ( new_n907_, new_n906_ );
nand g0770 ( new_n908_, new_n907_, N65 );
nand g0771 ( new_n909_, new_n908_, new_n901_ );
nand g0772 ( new_n910_, new_n909_, new_n777_ );
nand g0773 ( new_n911_, new_n906_, new_n571_ );
nor g0774 ( new_n912_, new_n906_, new_n571_ );
nor g0775 ( new_n913_, new_n912_, new_n777_ );
nand g0776 ( new_n914_, new_n913_, new_n911_ );
nand g0777 ( N740, new_n910_, new_n914_ );
not g0778 ( new_n916_, keyIn_0_53 );
not g0779 ( new_n917_, N69 );
nor g0780 ( new_n918_, new_n897_, new_n678_ );
nand g0781 ( new_n919_, new_n918_, keyIn_0_41 );
not g0782 ( new_n920_, keyIn_0_41 );
nand g0783 ( new_n921_, new_n892_, new_n677_ );
nand g0784 ( new_n922_, new_n921_, new_n920_ );
nand g0785 ( new_n923_, new_n919_, new_n922_ );
nand g0786 ( new_n924_, new_n923_, new_n917_ );
not g0787 ( new_n925_, new_n923_ );
nand g0788 ( new_n926_, new_n925_, N69 );
nand g0789 ( new_n927_, new_n926_, new_n924_ );
nand g0790 ( new_n928_, new_n927_, new_n916_ );
not g0791 ( new_n929_, new_n924_ );
nor g0792 ( new_n930_, new_n923_, new_n917_ );
nor g0793 ( new_n931_, new_n929_, new_n930_ );
nand g0794 ( new_n932_, new_n931_, keyIn_0_53 );
nand g0795 ( N741, new_n932_, new_n928_ );
not g0796 ( new_n934_, keyIn_0_54 );
not g0797 ( new_n935_, keyIn_0_42 );
nor g0798 ( new_n936_, new_n897_, new_n787_ );
nand g0799 ( new_n937_, new_n936_, new_n935_ );
nand g0800 ( new_n938_, new_n892_, new_n565_ );
nand g0801 ( new_n939_, new_n938_, keyIn_0_42 );
nand g0802 ( new_n940_, new_n937_, new_n939_ );
nand g0803 ( new_n941_, new_n940_, new_n139_ );
not g0804 ( new_n942_, new_n941_ );
nor g0805 ( new_n943_, new_n940_, new_n139_ );
nor g0806 ( new_n944_, new_n942_, new_n943_ );
nand g0807 ( new_n945_, new_n944_, new_n934_ );
not g0808 ( new_n946_, new_n940_ );
nand g0809 ( new_n947_, new_n946_, N73 );
nand g0810 ( new_n948_, new_n947_, new_n941_ );
nand g0811 ( new_n949_, new_n948_, keyIn_0_54 );
nand g0812 ( N742, new_n945_, new_n949_ );
not g0813 ( new_n951_, keyIn_0_55 );
not g0814 ( new_n952_, keyIn_0_43 );
nor g0815 ( new_n953_, new_n897_, new_n393_ );
nand g0816 ( new_n954_, new_n953_, new_n952_ );
nand g0817 ( new_n955_, new_n892_, new_n703_ );
nand g0818 ( new_n956_, new_n955_, keyIn_0_43 );
nand g0819 ( new_n957_, new_n954_, new_n956_ );
nand g0820 ( new_n958_, new_n957_, N77 );
not g0821 ( new_n959_, new_n957_ );
nand g0822 ( new_n960_, new_n959_, new_n141_ );
nand g0823 ( new_n961_, new_n960_, new_n958_ );
nand g0824 ( new_n962_, new_n961_, new_n951_ );
not g0825 ( new_n963_, new_n958_ );
nor g0826 ( new_n964_, new_n957_, N77 );
nor g0827 ( new_n965_, new_n963_, new_n964_ );
nand g0828 ( new_n966_, new_n965_, keyIn_0_55 );
nand g0829 ( N743, new_n966_, new_n962_ );
not g0830 ( new_n968_, keyIn_0_44 );
nand g0831 ( new_n969_, new_n280_, new_n314_ );
nor g0832 ( new_n970_, new_n885_, new_n969_ );
nand g0833 ( new_n971_, new_n884_, new_n970_ );
nor g0834 ( new_n972_, new_n971_, keyIn_0_38 );
nand g0835 ( new_n973_, new_n971_, keyIn_0_38 );
nand g0836 ( new_n974_, new_n973_, new_n782_ );
nor g0837 ( new_n975_, new_n974_, new_n972_ );
nand g0838 ( new_n976_, new_n975_, new_n968_ );
not g0839 ( new_n977_, new_n976_ );
nor g0840 ( new_n978_, new_n975_, new_n968_ );
nor g0841 ( new_n979_, new_n977_, new_n978_ );
nor g0842 ( new_n980_, new_n979_, N81 );
not g0843 ( new_n981_, new_n978_ );
nand g0844 ( new_n982_, new_n981_, new_n976_ );
nor g0845 ( new_n983_, new_n982_, new_n573_ );
nor g0846 ( new_n984_, new_n980_, new_n983_ );
nand g0847 ( new_n985_, new_n984_, keyIn_0_56 );
not g0848 ( new_n986_, keyIn_0_56 );
nand g0849 ( new_n987_, new_n982_, new_n573_ );
nand g0850 ( new_n988_, new_n979_, N81 );
nand g0851 ( new_n989_, new_n988_, new_n987_ );
nand g0852 ( new_n990_, new_n989_, new_n986_ );
nand g0853 ( N744, new_n985_, new_n990_ );
not g0854 ( new_n992_, keyIn_0_57 );
not g0855 ( new_n993_, keyIn_0_45 );
nand g0856 ( new_n994_, new_n973_, new_n677_ );
nor g0857 ( new_n995_, new_n994_, new_n972_ );
nand g0858 ( new_n996_, new_n995_, new_n993_ );
not g0859 ( new_n997_, new_n996_ );
nor g0860 ( new_n998_, new_n995_, new_n993_ );
nor g0861 ( new_n999_, new_n997_, new_n998_ );
nor g0862 ( new_n1000_, new_n999_, N85 );
not g0863 ( new_n1001_, N85 );
not g0864 ( new_n1002_, new_n998_ );
nand g0865 ( new_n1003_, new_n1002_, new_n996_ );
nor g0866 ( new_n1004_, new_n1003_, new_n1001_ );
nor g0867 ( new_n1005_, new_n1000_, new_n1004_ );
nand g0868 ( new_n1006_, new_n1005_, new_n992_ );
nand g0869 ( new_n1007_, new_n1003_, new_n1001_ );
nand g0870 ( new_n1008_, new_n999_, N85 );
nand g0871 ( new_n1009_, new_n1008_, new_n1007_ );
nand g0872 ( new_n1010_, new_n1009_, keyIn_0_57 );
nand g0873 ( N745, new_n1006_, new_n1010_ );
nand g0874 ( new_n1012_, new_n973_, new_n565_ );
nor g0875 ( new_n1013_, new_n1012_, new_n972_ );
nand g0876 ( new_n1014_, new_n1013_, keyIn_0_46 );
nor g0877 ( new_n1015_, new_n1013_, keyIn_0_46 );
not g0878 ( new_n1016_, new_n1015_ );
nand g0879 ( new_n1017_, new_n1016_, new_n1014_ );
nand g0880 ( new_n1018_, new_n1017_, new_n152_ );
not g0881 ( new_n1019_, new_n1014_ );
nor g0882 ( new_n1020_, new_n1019_, new_n1015_ );
nand g0883 ( new_n1021_, new_n1020_, N89 );
nand g0884 ( new_n1022_, new_n1021_, new_n1018_ );
nand g0885 ( new_n1023_, new_n1022_, keyIn_0_58 );
not g0886 ( new_n1024_, keyIn_0_58 );
nor g0887 ( new_n1025_, new_n1020_, N89 );
nor g0888 ( new_n1026_, new_n1017_, new_n152_ );
nor g0889 ( new_n1027_, new_n1025_, new_n1026_ );
nand g0890 ( new_n1028_, new_n1027_, new_n1024_ );
nand g0891 ( N746, new_n1028_, new_n1023_ );
not g0892 ( new_n1030_, keyIn_0_59 );
nand g0893 ( new_n1031_, new_n973_, new_n703_ );
nor g0894 ( new_n1032_, new_n1031_, new_n972_ );
nand g0895 ( new_n1033_, new_n1032_, keyIn_0_47 );
nor g0896 ( new_n1034_, new_n1032_, keyIn_0_47 );
not g0897 ( new_n1035_, new_n1034_ );
nand g0898 ( new_n1036_, new_n1035_, new_n1033_ );
nand g0899 ( new_n1037_, new_n1036_, new_n154_ );
not g0900 ( new_n1038_, new_n1033_ );
nor g0901 ( new_n1039_, new_n1038_, new_n1034_ );
nand g0902 ( new_n1040_, new_n1039_, N93 );
nand g0903 ( new_n1041_, new_n1040_, new_n1037_ );
nand g0904 ( new_n1042_, new_n1041_, new_n1030_ );
nor g0905 ( new_n1043_, new_n1039_, N93 );
nor g0906 ( new_n1044_, new_n1036_, new_n154_ );
nor g0907 ( new_n1045_, new_n1043_, new_n1044_ );
nand g0908 ( new_n1046_, new_n1045_, keyIn_0_59 );
nand g0909 ( N747, new_n1046_, new_n1042_ );
not g0910 ( new_n1048_, N97 );
not g0911 ( new_n1049_, keyIn_0_39 );
nand g0912 ( new_n1050_, new_n193_, new_n276_ );
nor g0913 ( new_n1051_, new_n886_, new_n1050_ );
nand g0914 ( new_n1052_, new_n884_, new_n1051_ );
nor g0915 ( new_n1053_, new_n1052_, new_n1049_ );
nand g0916 ( new_n1054_, new_n1052_, new_n1049_ );
nand g0917 ( new_n1055_, new_n1054_, new_n782_ );
nor g0918 ( new_n1056_, new_n1055_, new_n1053_ );
nand g0919 ( new_n1057_, new_n1056_, keyIn_0_48 );
nor g0920 ( new_n1058_, new_n1056_, keyIn_0_48 );
not g0921 ( new_n1059_, new_n1058_ );
nand g0922 ( new_n1060_, new_n1059_, new_n1057_ );
nand g0923 ( new_n1061_, new_n1060_, new_n1048_ );
not g0924 ( new_n1062_, new_n1057_ );
nor g0925 ( new_n1063_, new_n1062_, new_n1058_ );
nand g0926 ( new_n1064_, new_n1063_, N97 );
nand g0927 ( new_n1065_, new_n1064_, new_n1061_ );
nand g0928 ( new_n1066_, new_n1065_, keyIn_0_60 );
not g0929 ( new_n1067_, keyIn_0_60 );
nor g0930 ( new_n1068_, new_n1063_, N97 );
nor g0931 ( new_n1069_, new_n1060_, new_n1048_ );
nor g0932 ( new_n1070_, new_n1068_, new_n1069_ );
nand g0933 ( new_n1071_, new_n1070_, new_n1067_ );
nand g0934 ( N748, new_n1071_, new_n1066_ );
not g0935 ( new_n1073_, keyIn_0_49 );
nand g0936 ( new_n1074_, new_n1054_, new_n677_ );
nor g0937 ( new_n1075_, new_n1074_, new_n1053_ );
nand g0938 ( new_n1076_, new_n1075_, new_n1073_ );
nor g0939 ( new_n1077_, new_n1075_, new_n1073_ );
not g0940 ( new_n1078_, new_n1077_ );
nand g0941 ( new_n1079_, new_n1078_, new_n1076_ );
nand g0942 ( new_n1080_, new_n1079_, N101 );
not g0943 ( new_n1081_, new_n1076_ );
nor g0944 ( new_n1082_, new_n1081_, new_n1077_ );
nand g0945 ( new_n1083_, new_n1082_, new_n661_ );
nand g0946 ( new_n1084_, new_n1083_, new_n1080_ );
nand g0947 ( new_n1085_, new_n1084_, keyIn_0_61 );
not g0948 ( new_n1086_, keyIn_0_61 );
nor g0949 ( new_n1087_, new_n1082_, new_n661_ );
nor g0950 ( new_n1088_, new_n1079_, N101 );
nor g0951 ( new_n1089_, new_n1087_, new_n1088_ );
nand g0952 ( new_n1090_, new_n1089_, new_n1086_ );
nand g0953 ( N749, new_n1090_, new_n1085_ );
not g0954 ( new_n1092_, keyIn_0_50 );
nand g0955 ( new_n1093_, new_n1054_, new_n565_ );
nor g0956 ( new_n1094_, new_n1093_, new_n1053_ );
nand g0957 ( new_n1095_, new_n1094_, new_n1092_ );
not g0958 ( new_n1096_, new_n1095_ );
nor g0959 ( new_n1097_, new_n1094_, new_n1092_ );
nor g0960 ( new_n1098_, new_n1096_, new_n1097_ );
nor g0961 ( new_n1099_, new_n1098_, N105 );
not g0962 ( new_n1100_, new_n1097_ );
nand g0963 ( new_n1101_, new_n1100_, new_n1095_ );
nor g0964 ( new_n1102_, new_n1101_, new_n194_ );
nor g0965 ( new_n1103_, new_n1099_, new_n1102_ );
nand g0966 ( new_n1104_, new_n1103_, keyIn_0_62 );
not g0967 ( new_n1105_, keyIn_0_62 );
nand g0968 ( new_n1106_, new_n1101_, new_n194_ );
nand g0969 ( new_n1107_, new_n1098_, N105 );
nand g0970 ( new_n1108_, new_n1107_, new_n1106_ );
nand g0971 ( new_n1109_, new_n1108_, new_n1105_ );
nand g0972 ( N750, new_n1104_, new_n1109_ );
not g0973 ( new_n1111_, keyIn_0_51 );
nand g0974 ( new_n1112_, new_n1054_, new_n703_ );
nor g0975 ( new_n1113_, new_n1112_, new_n1053_ );
nand g0976 ( new_n1114_, new_n1113_, new_n1111_ );
not g0977 ( new_n1115_, new_n1114_ );
nor g0978 ( new_n1116_, new_n1113_, new_n1111_ );
nor g0979 ( new_n1117_, new_n1115_, new_n1116_ );
nor g0980 ( new_n1118_, new_n1117_, N109 );
not g0981 ( new_n1119_, new_n1116_ );
nand g0982 ( new_n1120_, new_n1119_, new_n1114_ );
nor g0983 ( new_n1121_, new_n1120_, new_n196_ );
nor g0984 ( new_n1122_, new_n1118_, new_n1121_ );
nand g0985 ( new_n1123_, new_n1122_, keyIn_0_63 );
not g0986 ( new_n1124_, keyIn_0_63 );
nand g0987 ( new_n1125_, new_n1120_, new_n196_ );
nand g0988 ( new_n1126_, new_n1117_, N109 );
nand g0989 ( new_n1127_, new_n1126_, new_n1125_ );
nand g0990 ( new_n1128_, new_n1127_, new_n1124_ );
nand g0991 ( N751, new_n1123_, new_n1128_ );
not g0992 ( new_n1130_, N113 );
nand g0993 ( new_n1131_, new_n282_, new_n314_ );
nor g0994 ( new_n1132_, new_n810_, new_n1131_ );
nand g0995 ( new_n1133_, new_n884_, new_n1132_ );
not g0996 ( new_n1134_, new_n1133_ );
nand g0997 ( new_n1135_, new_n1134_, new_n1130_ );
nand g0998 ( new_n1136_, new_n1133_, N113 );
nand g0999 ( N752, new_n1135_, new_n1136_ );
nor g1000 ( new_n1138_, new_n1131_, new_n678_ );
nand g1001 ( new_n1139_, new_n884_, new_n1138_ );
not g1002 ( new_n1140_, new_n1139_ );
nand g1003 ( new_n1141_, new_n1140_, new_n663_ );
nand g1004 ( new_n1142_, new_n1139_, N117 );
nand g1005 ( N753, new_n1141_, new_n1142_ );
nor g1006 ( new_n1144_, new_n787_, new_n1131_ );
nand g1007 ( new_n1145_, new_n884_, new_n1144_ );
not g1008 ( new_n1146_, new_n1145_ );
nand g1009 ( new_n1147_, new_n1146_, new_n237_ );
nand g1010 ( new_n1148_, new_n1145_, N121 );
nand g1011 ( N754, new_n1147_, new_n1148_ );
nor g1012 ( new_n1150_, new_n1131_, new_n393_ );
nand g1013 ( new_n1151_, new_n884_, new_n1150_ );
not g1014 ( new_n1152_, new_n1151_ );
nand g1015 ( new_n1153_, new_n1152_, new_n239_ );
nand g1016 ( new_n1154_, new_n1151_, N125 );
nand g1017 ( N755, new_n1153_, new_n1154_ );
endmodule