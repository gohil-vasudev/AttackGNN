module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124;

  INV_X2 U2001 ( .A(n2010), .ZN(n1969) );
  NOR2_X1 U2002 ( .A1(n1969), .A2(n1970), .ZN(Result_9_) );
  XOR2_X1 U2003 ( .A(n1971), .B(n1972), .Z(n1970) );
  NAND2_X1 U2004 ( .A1(n1973), .A2(n1974), .ZN(n1972) );
  NOR2_X1 U2005 ( .A1(n1969), .A2(n1975), .ZN(Result_8_) );
  XOR2_X1 U2006 ( .A(n1976), .B(n1977), .Z(n1975) );
  NAND2_X1 U2007 ( .A1(n1978), .A2(n1979), .ZN(n1977) );
  NOR2_X1 U2008 ( .A1(n1969), .A2(n1980), .ZN(Result_7_) );
  XOR2_X1 U2009 ( .A(n1981), .B(n1982), .Z(n1980) );
  NAND2_X1 U2010 ( .A1(n1983), .A2(n1984), .ZN(n1982) );
  NOR2_X1 U2011 ( .A1(n1969), .A2(n1985), .ZN(Result_6_) );
  XOR2_X1 U2012 ( .A(n1986), .B(n1987), .Z(n1985) );
  NAND2_X1 U2013 ( .A1(n1988), .A2(n1989), .ZN(n1987) );
  NOR2_X1 U2014 ( .A1(n1969), .A2(n1990), .ZN(Result_5_) );
  XOR2_X1 U2015 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND2_X1 U2016 ( .A1(n1993), .A2(n1994), .ZN(n1992) );
  NOR2_X1 U2017 ( .A1(n1969), .A2(n1995), .ZN(Result_4_) );
  XOR2_X1 U2018 ( .A(n1996), .B(n1997), .Z(n1995) );
  NAND2_X1 U2019 ( .A1(n1998), .A2(n1999), .ZN(n1997) );
  NOR2_X1 U2020 ( .A1(n1969), .A2(n2000), .ZN(Result_3_) );
  XOR2_X1 U2021 ( .A(n2001), .B(n2002), .Z(n2000) );
  NAND2_X1 U2022 ( .A1(n2003), .A2(n2004), .ZN(n2002) );
  NAND2_X1 U2023 ( .A1(n2005), .A2(n2006), .ZN(Result_31_) );
  NAND2_X1 U2024 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
  NOR2_X1 U2025 ( .A1(n2009), .A2(n2010), .ZN(n2007) );
  NAND2_X1 U2026 ( .A1(n2011), .A2(b_15_), .ZN(n2005) );
  XOR2_X1 U2027 ( .A(n2009), .B(n2010), .Z(n2011) );
  NAND2_X1 U2028 ( .A1(n2012), .A2(n2013), .ZN(Result_30_) );
  NAND2_X1 U2029 ( .A1(n2014), .A2(n2010), .ZN(n2013) );
  NAND2_X1 U2030 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
  NAND2_X1 U2031 ( .A1(b_14_), .A2(n2017), .ZN(n2016) );
  NAND2_X1 U2032 ( .A1(n2018), .A2(n2019), .ZN(n2017) );
  NAND2_X1 U2033 ( .A1(a_15_), .A2(n2008), .ZN(n2019) );
  NAND2_X1 U2034 ( .A1(b_15_), .A2(n2020), .ZN(n2015) );
  NAND2_X1 U2035 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
  NAND2_X1 U2036 ( .A1(a_14_), .A2(n2023), .ZN(n2022) );
  NAND2_X1 U2037 ( .A1(n2024), .A2(n1969), .ZN(n2012) );
  XOR2_X1 U2038 ( .A(n2025), .B(n2026), .Z(n2024) );
  XOR2_X1 U2039 ( .A(b_14_), .B(a_14_), .Z(n2026) );
  NOR2_X1 U2040 ( .A1(n2008), .A2(n2009), .ZN(n2025) );
  NOR2_X1 U2041 ( .A1(n1969), .A2(n2027), .ZN(Result_2_) );
  XOR2_X1 U2042 ( .A(n2028), .B(n2029), .Z(n2027) );
  NAND2_X1 U2043 ( .A1(n2030), .A2(n2031), .ZN(n2029) );
  NAND2_X1 U2044 ( .A1(n2032), .A2(n2033), .ZN(Result_29_) );
  NAND2_X1 U2045 ( .A1(n1969), .A2(n2034), .ZN(n2033) );
  NAND2_X1 U2046 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  NAND2_X1 U2047 ( .A1(n2037), .A2(n2038), .ZN(n2036) );
  NOR2_X1 U2048 ( .A1(n2039), .A2(n2040), .ZN(n2035) );
  NOR2_X1 U2049 ( .A1(b_13_), .A2(n2041), .ZN(n2040) );
  XOR2_X1 U2050 ( .A(n2042), .B(n2038), .Z(n2041) );
  NOR2_X1 U2051 ( .A1(n2043), .A2(n2044), .ZN(n2039) );
  OR2_X1 U2052 ( .A1(n2038), .A2(a_13_), .ZN(n2044) );
  NAND2_X1 U2053 ( .A1(n2045), .A2(n2010), .ZN(n2032) );
  XOR2_X1 U2054 ( .A(n2046), .B(n2047), .Z(n2045) );
  NOR2_X1 U2055 ( .A1(n2008), .A2(n2042), .ZN(n2047) );
  XOR2_X1 U2056 ( .A(n2048), .B(n2049), .Z(n2046) );
  NAND2_X1 U2057 ( .A1(n2050), .A2(n2051), .ZN(Result_28_) );
  NAND2_X1 U2058 ( .A1(n2052), .A2(n2010), .ZN(n2051) );
  XNOR2_X1 U2059 ( .A(n2053), .B(n2054), .ZN(n2052) );
  XOR2_X1 U2060 ( .A(n2055), .B(n2056), .Z(n2054) );
  NAND2_X1 U2061 ( .A1(a_12_), .A2(b_15_), .ZN(n2056) );
  NAND2_X1 U2062 ( .A1(n2057), .A2(n1969), .ZN(n2050) );
  XOR2_X1 U2063 ( .A(n2058), .B(n2059), .Z(n2057) );
  AND2_X1 U2064 ( .A1(n2060), .A2(n2061), .ZN(n2059) );
  NAND2_X1 U2065 ( .A1(n2062), .A2(n2063), .ZN(Result_27_) );
  NAND2_X1 U2066 ( .A1(n1969), .A2(n2064), .ZN(n2063) );
  NAND2_X1 U2067 ( .A1(n2065), .A2(n2066), .ZN(n2064) );
  NAND2_X1 U2068 ( .A1(n2067), .A2(n2068), .ZN(n2066) );
  NOR2_X1 U2069 ( .A1(n2069), .A2(n2070), .ZN(n2065) );
  NOR2_X1 U2070 ( .A1(b_11_), .A2(n2071), .ZN(n2070) );
  XOR2_X1 U2071 ( .A(n2072), .B(n2068), .Z(n2071) );
  NOR2_X1 U2072 ( .A1(n2073), .A2(n2074), .ZN(n2069) );
  OR2_X1 U2073 ( .A1(n2068), .A2(a_11_), .ZN(n2074) );
  NAND2_X1 U2074 ( .A1(n2075), .A2(n2010), .ZN(n2062) );
  XNOR2_X1 U2075 ( .A(n2076), .B(n2077), .ZN(n2075) );
  NAND2_X1 U2076 ( .A1(n2078), .A2(n2079), .ZN(n2076) );
  NAND2_X1 U2077 ( .A1(n2080), .A2(n2081), .ZN(Result_26_) );
  NAND2_X1 U2078 ( .A1(n2082), .A2(n2010), .ZN(n2081) );
  XOR2_X1 U2079 ( .A(n2083), .B(n2084), .Z(n2082) );
  XNOR2_X1 U2080 ( .A(n2085), .B(n2086), .ZN(n2083) );
  NAND2_X1 U2081 ( .A1(a_10_), .A2(b_15_), .ZN(n2085) );
  NAND2_X1 U2082 ( .A1(n2087), .A2(n1969), .ZN(n2080) );
  XOR2_X1 U2083 ( .A(n2088), .B(n2089), .Z(n2087) );
  AND2_X1 U2084 ( .A1(n2090), .A2(n2091), .ZN(n2089) );
  NAND2_X1 U2085 ( .A1(n2092), .A2(n2093), .ZN(Result_25_) );
  NAND2_X1 U2086 ( .A1(n1969), .A2(n2094), .ZN(n2093) );
  NAND2_X1 U2087 ( .A1(n2095), .A2(n2096), .ZN(n2094) );
  NAND2_X1 U2088 ( .A1(n2097), .A2(n2098), .ZN(n2096) );
  NOR2_X1 U2089 ( .A1(n2099), .A2(n2100), .ZN(n2095) );
  NOR2_X1 U2090 ( .A1(b_9_), .A2(n2101), .ZN(n2100) );
  XOR2_X1 U2091 ( .A(n2102), .B(n2098), .Z(n2101) );
  NOR2_X1 U2092 ( .A1(n2103), .A2(n2104), .ZN(n2099) );
  OR2_X1 U2093 ( .A1(n2098), .A2(a_9_), .ZN(n2104) );
  NAND2_X1 U2094 ( .A1(n2105), .A2(n2010), .ZN(n2092) );
  XNOR2_X1 U2095 ( .A(n2106), .B(n2107), .ZN(n2105) );
  NAND2_X1 U2096 ( .A1(n2108), .A2(n2109), .ZN(n2106) );
  NAND2_X1 U2097 ( .A1(n2110), .A2(n2111), .ZN(Result_24_) );
  NAND2_X1 U2098 ( .A1(n2112), .A2(n2010), .ZN(n2111) );
  XOR2_X1 U2099 ( .A(n2113), .B(n2114), .Z(n2112) );
  XNOR2_X1 U2100 ( .A(n2115), .B(n2116), .ZN(n2114) );
  NAND2_X1 U2101 ( .A1(a_8_), .A2(b_15_), .ZN(n2115) );
  NAND2_X1 U2102 ( .A1(n2117), .A2(n1969), .ZN(n2110) );
  XOR2_X1 U2103 ( .A(n2118), .B(n2119), .Z(n2117) );
  AND2_X1 U2104 ( .A1(n2120), .A2(n2121), .ZN(n2119) );
  NAND2_X1 U2105 ( .A1(n2122), .A2(n2123), .ZN(Result_23_) );
  NAND2_X1 U2106 ( .A1(n1969), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2107 ( .A1(n2125), .A2(n2126), .ZN(n2124) );
  NAND2_X1 U2108 ( .A1(n2127), .A2(n2128), .ZN(n2126) );
  NOR2_X1 U2109 ( .A1(n2129), .A2(n2130), .ZN(n2125) );
  NOR2_X1 U2110 ( .A1(b_7_), .A2(n2131), .ZN(n2130) );
  XOR2_X1 U2111 ( .A(n2132), .B(n2128), .Z(n2131) );
  NOR2_X1 U2112 ( .A1(n2133), .A2(n2134), .ZN(n2129) );
  OR2_X1 U2113 ( .A1(n2128), .A2(a_7_), .ZN(n2134) );
  NAND2_X1 U2114 ( .A1(n2135), .A2(n2010), .ZN(n2122) );
  XNOR2_X1 U2115 ( .A(n2136), .B(n2137), .ZN(n2135) );
  NAND2_X1 U2116 ( .A1(n2138), .A2(n2139), .ZN(n2136) );
  NAND2_X1 U2117 ( .A1(n2140), .A2(n2141), .ZN(Result_22_) );
  NAND2_X1 U2118 ( .A1(n2142), .A2(n2010), .ZN(n2141) );
  XNOR2_X1 U2119 ( .A(n2143), .B(n2144), .ZN(n2142) );
  XOR2_X1 U2120 ( .A(n2145), .B(n2146), .Z(n2144) );
  NAND2_X1 U2121 ( .A1(a_6_), .A2(b_15_), .ZN(n2146) );
  NAND2_X1 U2122 ( .A1(n2147), .A2(n1969), .ZN(n2140) );
  XOR2_X1 U2123 ( .A(n2148), .B(n2149), .Z(n2147) );
  AND2_X1 U2124 ( .A1(n2150), .A2(n2151), .ZN(n2149) );
  NAND2_X1 U2125 ( .A1(n2152), .A2(n2153), .ZN(Result_21_) );
  NAND2_X1 U2126 ( .A1(n1969), .A2(n2154), .ZN(n2153) );
  NAND2_X1 U2127 ( .A1(n2155), .A2(n2156), .ZN(n2154) );
  NAND2_X1 U2128 ( .A1(n2157), .A2(n2158), .ZN(n2156) );
  NOR2_X1 U2129 ( .A1(n2159), .A2(n2160), .ZN(n2155) );
  NOR2_X1 U2130 ( .A1(b_5_), .A2(n2161), .ZN(n2160) );
  XOR2_X1 U2131 ( .A(n2162), .B(n2158), .Z(n2161) );
  NOR2_X1 U2132 ( .A1(n2163), .A2(n2164), .ZN(n2159) );
  OR2_X1 U2133 ( .A1(n2158), .A2(a_5_), .ZN(n2164) );
  NAND2_X1 U2134 ( .A1(n2165), .A2(n2010), .ZN(n2152) );
  XNOR2_X1 U2135 ( .A(n2166), .B(n2167), .ZN(n2165) );
  NAND2_X1 U2136 ( .A1(n2168), .A2(n2169), .ZN(n2166) );
  NAND2_X1 U2137 ( .A1(n2170), .A2(n2171), .ZN(Result_20_) );
  NAND2_X1 U2138 ( .A1(n2172), .A2(n2010), .ZN(n2171) );
  XNOR2_X1 U2139 ( .A(n2173), .B(n2174), .ZN(n2172) );
  XOR2_X1 U2140 ( .A(n2175), .B(n2176), .Z(n2174) );
  NAND2_X1 U2141 ( .A1(a_4_), .A2(b_15_), .ZN(n2176) );
  NAND2_X1 U2142 ( .A1(n2177), .A2(n1969), .ZN(n2170) );
  XOR2_X1 U2143 ( .A(n2178), .B(n2179), .Z(n2177) );
  AND2_X1 U2144 ( .A1(n2180), .A2(n2181), .ZN(n2179) );
  NOR2_X1 U2145 ( .A1(n1969), .A2(n2182), .ZN(Result_1_) );
  XOR2_X1 U2146 ( .A(n2183), .B(n2184), .Z(n2182) );
  NAND2_X1 U2147 ( .A1(n2185), .A2(n2186), .ZN(n2184) );
  NAND2_X1 U2148 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
  NAND2_X1 U2149 ( .A1(n2189), .A2(n2190), .ZN(Result_19_) );
  NAND2_X1 U2150 ( .A1(n1969), .A2(n2191), .ZN(n2190) );
  NAND2_X1 U2151 ( .A1(n2192), .A2(n2193), .ZN(n2191) );
  NAND2_X1 U2152 ( .A1(n2194), .A2(n2195), .ZN(n2193) );
  NOR2_X1 U2153 ( .A1(n2196), .A2(n2197), .ZN(n2192) );
  NOR2_X1 U2154 ( .A1(b_3_), .A2(n2198), .ZN(n2197) );
  XOR2_X1 U2155 ( .A(n2199), .B(n2195), .Z(n2198) );
  NOR2_X1 U2156 ( .A1(n2200), .A2(n2201), .ZN(n2196) );
  OR2_X1 U2157 ( .A1(n2195), .A2(a_3_), .ZN(n2201) );
  NAND2_X1 U2158 ( .A1(n2202), .A2(n2010), .ZN(n2189) );
  XNOR2_X1 U2159 ( .A(n2203), .B(n2204), .ZN(n2202) );
  XOR2_X1 U2160 ( .A(n2205), .B(n2206), .Z(n2204) );
  NAND2_X1 U2161 ( .A1(a_3_), .A2(b_15_), .ZN(n2206) );
  NAND2_X1 U2162 ( .A1(n2207), .A2(n2208), .ZN(Result_18_) );
  NAND2_X1 U2163 ( .A1(n2209), .A2(n2010), .ZN(n2208) );
  XNOR2_X1 U2164 ( .A(n2210), .B(n2211), .ZN(n2209) );
  XOR2_X1 U2165 ( .A(n2212), .B(n2213), .Z(n2211) );
  NAND2_X1 U2166 ( .A1(a_2_), .A2(b_15_), .ZN(n2213) );
  NAND2_X1 U2167 ( .A1(n2214), .A2(n1969), .ZN(n2207) );
  XOR2_X1 U2168 ( .A(n2215), .B(n2216), .Z(n2214) );
  AND2_X1 U2169 ( .A1(n2217), .A2(n2218), .ZN(n2216) );
  NAND2_X1 U2170 ( .A1(n2219), .A2(n2220), .ZN(Result_17_) );
  NAND2_X1 U2171 ( .A1(n2221), .A2(n2010), .ZN(n2220) );
  XNOR2_X1 U2172 ( .A(n2222), .B(n2223), .ZN(n2221) );
  XOR2_X1 U2173 ( .A(n2224), .B(n2225), .Z(n2223) );
  NAND2_X1 U2174 ( .A1(b_15_), .A2(a_1_), .ZN(n2225) );
  NAND2_X1 U2175 ( .A1(n2226), .A2(n1969), .ZN(n2219) );
  NAND2_X1 U2176 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
  NAND2_X1 U2177 ( .A1(n2229), .A2(n2230), .ZN(n2228) );
  OR2_X1 U2178 ( .A1(n2231), .A2(n2232), .ZN(n2229) );
  NAND2_X1 U2179 ( .A1(n2233), .A2(n2234), .ZN(n2227) );
  INV_X1 U2180 ( .A(n2230), .ZN(n2234) );
  XOR2_X1 U2181 ( .A(b_1_), .B(a_1_), .Z(n2233) );
  NAND2_X1 U2182 ( .A1(n2235), .A2(n2236), .ZN(Result_16_) );
  NAND2_X1 U2183 ( .A1(n2237), .A2(n2010), .ZN(n2236) );
  XOR2_X1 U2184 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR2_X1 U2185 ( .A(n2240), .B(n2241), .Z(n2239) );
  NAND2_X1 U2186 ( .A1(n2242), .A2(n1969), .ZN(n2235) );
  XNOR2_X1 U2187 ( .A(n2243), .B(n2244), .ZN(n2242) );
  NOR2_X1 U2188 ( .A1(n2232), .A2(n2245), .ZN(n2243) );
  NOR2_X1 U2189 ( .A1(n2231), .A2(n2230), .ZN(n2245) );
  NAND2_X1 U2190 ( .A1(n2218), .A2(n2246), .ZN(n2230) );
  NAND2_X1 U2191 ( .A1(n2217), .A2(n2215), .ZN(n2246) );
  NAND2_X1 U2192 ( .A1(n2247), .A2(n2248), .ZN(n2215) );
  NAND2_X1 U2193 ( .A1(n2249), .A2(n2195), .ZN(n2248) );
  NAND2_X1 U2194 ( .A1(n2181), .A2(n2250), .ZN(n2195) );
  NAND2_X1 U2195 ( .A1(n2180), .A2(n2178), .ZN(n2250) );
  NAND2_X1 U2196 ( .A1(n2251), .A2(n2252), .ZN(n2178) );
  NAND2_X1 U2197 ( .A1(n2253), .A2(n2158), .ZN(n2252) );
  NAND2_X1 U2198 ( .A1(n2151), .A2(n2254), .ZN(n2158) );
  NAND2_X1 U2199 ( .A1(n2150), .A2(n2148), .ZN(n2254) );
  NAND2_X1 U2200 ( .A1(n2255), .A2(n2256), .ZN(n2148) );
  NAND2_X1 U2201 ( .A1(n2257), .A2(n2128), .ZN(n2256) );
  NAND2_X1 U2202 ( .A1(n2121), .A2(n2258), .ZN(n2128) );
  NAND2_X1 U2203 ( .A1(n2120), .A2(n2118), .ZN(n2258) );
  NAND2_X1 U2204 ( .A1(n2259), .A2(n2260), .ZN(n2118) );
  NAND2_X1 U2205 ( .A1(n2261), .A2(n2098), .ZN(n2260) );
  NAND2_X1 U2206 ( .A1(n2091), .A2(n2262), .ZN(n2098) );
  NAND2_X1 U2207 ( .A1(n2090), .A2(n2088), .ZN(n2262) );
  NAND2_X1 U2208 ( .A1(n2263), .A2(n2264), .ZN(n2088) );
  NAND2_X1 U2209 ( .A1(n2265), .A2(n2068), .ZN(n2264) );
  NAND2_X1 U2210 ( .A1(n2061), .A2(n2266), .ZN(n2068) );
  NAND2_X1 U2211 ( .A1(n2060), .A2(n2058), .ZN(n2266) );
  NAND2_X1 U2212 ( .A1(n2267), .A2(n2268), .ZN(n2058) );
  NAND2_X1 U2213 ( .A1(n2269), .A2(n2038), .ZN(n2268) );
  NAND2_X1 U2214 ( .A1(n2270), .A2(n2271), .ZN(n2038) );
  NAND2_X1 U2215 ( .A1(a_14_), .A2(b_14_), .ZN(n2271) );
  NOR2_X1 U2216 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
  NOR2_X1 U2217 ( .A1(n2008), .A2(n2274), .ZN(n2273) );
  NOR2_X1 U2218 ( .A1(n2009), .A2(n2275), .ZN(n2272) );
  NAND2_X1 U2219 ( .A1(n2043), .A2(n2042), .ZN(n2269) );
  NAND2_X1 U2220 ( .A1(n2276), .A2(n2277), .ZN(n2060) );
  NAND2_X1 U2221 ( .A1(n2073), .A2(n2072), .ZN(n2265) );
  NAND2_X1 U2222 ( .A1(n2278), .A2(n2279), .ZN(n2090) );
  NAND2_X1 U2223 ( .A1(n2103), .A2(n2102), .ZN(n2261) );
  NAND2_X1 U2224 ( .A1(n2280), .A2(n2281), .ZN(n2120) );
  NAND2_X1 U2225 ( .A1(n2133), .A2(n2132), .ZN(n2257) );
  NAND2_X1 U2226 ( .A1(n2282), .A2(n2283), .ZN(n2150) );
  NAND2_X1 U2227 ( .A1(n2163), .A2(n2162), .ZN(n2253) );
  NAND2_X1 U2228 ( .A1(n2284), .A2(n2285), .ZN(n2180) );
  NAND2_X1 U2229 ( .A1(n2200), .A2(n2199), .ZN(n2249) );
  NAND2_X1 U2230 ( .A1(n2286), .A2(n2287), .ZN(n2217) );
  INV_X1 U2231 ( .A(n2288), .ZN(n2231) );
  NOR2_X1 U2232 ( .A1(b_1_), .A2(a_1_), .ZN(n2232) );
  NOR2_X1 U2233 ( .A1(n1969), .A2(n2289), .ZN(Result_15_) );
  XNOR2_X1 U2234 ( .A(n2290), .B(n2291), .ZN(n2289) );
  NOR2_X1 U2235 ( .A1(n2292), .A2(n2293), .ZN(Result_14_) );
  NAND2_X1 U2236 ( .A1(n2294), .A2(n2010), .ZN(n2293) );
  NOR2_X1 U2237 ( .A1(n2295), .A2(n2296), .ZN(n2292) );
  XOR2_X1 U2238 ( .A(n2297), .B(n2298), .Z(n2296) );
  NOR2_X1 U2239 ( .A1(n2290), .A2(n2291), .ZN(n2295) );
  NOR2_X1 U2240 ( .A1(n1969), .A2(n2299), .ZN(Result_13_) );
  NAND2_X1 U2241 ( .A1(n2300), .A2(n2301), .ZN(n2299) );
  NAND2_X1 U2242 ( .A1(n2302), .A2(n2294), .ZN(n2301) );
  NAND2_X1 U2243 ( .A1(n2303), .A2(n2304), .ZN(n2302) );
  NAND2_X1 U2244 ( .A1(n2305), .A2(n2306), .ZN(n2303) );
  NAND2_X1 U2245 ( .A1(n2307), .A2(n2304), .ZN(n2300) );
  NAND2_X1 U2246 ( .A1(n2308), .A2(n2309), .ZN(n2304) );
  INV_X1 U2247 ( .A(n2294), .ZN(n2307) );
  NOR2_X1 U2248 ( .A1(n1969), .A2(n2310), .ZN(Result_12_) );
  XNOR2_X1 U2249 ( .A(n2311), .B(n2312), .ZN(n2310) );
  NOR2_X1 U2250 ( .A1(n1969), .A2(n2313), .ZN(Result_11_) );
  XNOR2_X1 U2251 ( .A(n2314), .B(n2315), .ZN(n2313) );
  NOR2_X1 U2252 ( .A1(n2316), .A2(n2317), .ZN(n2315) );
  NOR2_X1 U2253 ( .A1(n2318), .A2(n2319), .ZN(n2317) );
  INV_X1 U2254 ( .A(n2320), .ZN(n2316) );
  NOR2_X1 U2255 ( .A1(n1969), .A2(n2321), .ZN(Result_10_) );
  XNOR2_X1 U2256 ( .A(n2322), .B(n2323), .ZN(n2321) );
  NOR2_X1 U2257 ( .A1(n2324), .A2(n2325), .ZN(n2323) );
  NOR2_X1 U2258 ( .A1(n2326), .A2(n2327), .ZN(n2325) );
  NOR2_X1 U2259 ( .A1(n1969), .A2(n2328), .ZN(Result_0_) );
  NOR2_X1 U2260 ( .A1(n2329), .A2(n2330), .ZN(n2328) );
  NAND2_X1 U2261 ( .A1(n2188), .A2(n2331), .ZN(n2330) );
  INV_X1 U2262 ( .A(n2187), .ZN(n2331) );
  NOR2_X1 U2263 ( .A1(n2332), .A2(n2333), .ZN(n2187) );
  AND2_X1 U2264 ( .A1(n2183), .A2(n2185), .ZN(n2329) );
  NAND2_X1 U2265 ( .A1(n2332), .A2(n2334), .ZN(n2185) );
  NAND2_X1 U2266 ( .A1(b_0_), .A2(n2188), .ZN(n2334) );
  NAND2_X1 U2267 ( .A1(n2335), .A2(n2336), .ZN(n2188) );
  NAND2_X1 U2268 ( .A1(n2030), .A2(n2337), .ZN(n2183) );
  NAND2_X1 U2269 ( .A1(n2031), .A2(n2028), .ZN(n2337) );
  NAND2_X1 U2270 ( .A1(n2003), .A2(n2338), .ZN(n2028) );
  NAND2_X1 U2271 ( .A1(n2004), .A2(n2001), .ZN(n2338) );
  NAND2_X1 U2272 ( .A1(n1998), .A2(n2339), .ZN(n2001) );
  NAND2_X1 U2273 ( .A1(n1999), .A2(n1996), .ZN(n2339) );
  NAND2_X1 U2274 ( .A1(n1993), .A2(n2340), .ZN(n1996) );
  NAND2_X1 U2275 ( .A1(n1994), .A2(n1991), .ZN(n2340) );
  NAND2_X1 U2276 ( .A1(n1988), .A2(n2341), .ZN(n1991) );
  NAND2_X1 U2277 ( .A1(n1989), .A2(n1986), .ZN(n2341) );
  NAND2_X1 U2278 ( .A1(n1983), .A2(n2342), .ZN(n1986) );
  NAND2_X1 U2279 ( .A1(n1984), .A2(n1981), .ZN(n2342) );
  NAND2_X1 U2280 ( .A1(n1978), .A2(n2343), .ZN(n1981) );
  NAND2_X1 U2281 ( .A1(n1979), .A2(n1976), .ZN(n2343) );
  NAND2_X1 U2282 ( .A1(n1973), .A2(n2344), .ZN(n1976) );
  NAND2_X1 U2283 ( .A1(n1974), .A2(n1971), .ZN(n2344) );
  NAND2_X1 U2284 ( .A1(n2345), .A2(n2346), .ZN(n1971) );
  NAND2_X1 U2285 ( .A1(n2347), .A2(n2348), .ZN(n2346) );
  NAND2_X1 U2286 ( .A1(n2322), .A2(n2349), .ZN(n2345) );
  INV_X1 U2287 ( .A(n2324), .ZN(n2349) );
  NOR2_X1 U2288 ( .A1(n2348), .A2(n2347), .ZN(n2324) );
  INV_X1 U2289 ( .A(n2326), .ZN(n2348) );
  XNOR2_X1 U2290 ( .A(n2350), .B(n2351), .ZN(n2326) );
  NAND2_X1 U2291 ( .A1(n2352), .A2(n2320), .ZN(n2322) );
  NAND2_X1 U2292 ( .A1(n2319), .A2(n2318), .ZN(n2320) );
  AND2_X1 U2293 ( .A1(n2353), .A2(n2354), .ZN(n2318) );
  NAND2_X1 U2294 ( .A1(n2314), .A2(n2319), .ZN(n2352) );
  AND2_X1 U2295 ( .A1(n2327), .A2(n2355), .ZN(n2319) );
  NAND2_X1 U2296 ( .A1(n2356), .A2(n2357), .ZN(n2355) );
  INV_X1 U2297 ( .A(n2347), .ZN(n2327) );
  NOR2_X1 U2298 ( .A1(n2357), .A2(n2356), .ZN(n2347) );
  XOR2_X1 U2299 ( .A(n2358), .B(n2359), .Z(n2356) );
  NAND2_X1 U2300 ( .A1(n2360), .A2(n2361), .ZN(n2358) );
  NAND2_X1 U2301 ( .A1(n2362), .A2(n2363), .ZN(n2357) );
  NAND2_X1 U2302 ( .A1(n2364), .A2(n2365), .ZN(n2363) );
  NAND2_X1 U2303 ( .A1(n2366), .A2(n2367), .ZN(n2365) );
  OR2_X1 U2304 ( .A1(n2367), .A2(n2366), .ZN(n2362) );
  NOR2_X1 U2305 ( .A1(n2312), .A2(n2311), .ZN(n2314) );
  AND2_X1 U2306 ( .A1(n2368), .A2(n2369), .ZN(n2311) );
  NAND2_X1 U2307 ( .A1(n2306), .A2(n2370), .ZN(n2368) );
  NAND2_X1 U2308 ( .A1(n2294), .A2(n2308), .ZN(n2370) );
  NAND2_X1 U2309 ( .A1(n2371), .A2(n2372), .ZN(n2294) );
  NOR2_X1 U2310 ( .A1(n2290), .A2(n2305), .ZN(n2372) );
  INV_X1 U2311 ( .A(n2308), .ZN(n2305) );
  NAND2_X1 U2312 ( .A1(n2298), .A2(n2297), .ZN(n2308) );
  AND2_X1 U2313 ( .A1(n2373), .A2(n2374), .ZN(n2290) );
  NAND2_X1 U2314 ( .A1(n2241), .A2(n2375), .ZN(n2374) );
  NAND2_X1 U2315 ( .A1(n2240), .A2(n2238), .ZN(n2375) );
  NOR2_X1 U2316 ( .A1(n2376), .A2(n2008), .ZN(n2241) );
  OR2_X1 U2317 ( .A1(n2238), .A2(n2240), .ZN(n2373) );
  AND2_X1 U2318 ( .A1(n2377), .A2(n2378), .ZN(n2240) );
  NAND2_X1 U2319 ( .A1(n2379), .A2(b_15_), .ZN(n2378) );
  NOR2_X1 U2320 ( .A1(n2380), .A2(n2381), .ZN(n2379) );
  NOR2_X1 U2321 ( .A1(n2222), .A2(n2224), .ZN(n2380) );
  NAND2_X1 U2322 ( .A1(n2222), .A2(n2224), .ZN(n2377) );
  NAND2_X1 U2323 ( .A1(n2382), .A2(n2383), .ZN(n2224) );
  NAND2_X1 U2324 ( .A1(n2384), .A2(a_2_), .ZN(n2383) );
  NOR2_X1 U2325 ( .A1(n2385), .A2(n2008), .ZN(n2384) );
  NOR2_X1 U2326 ( .A1(n2210), .A2(n2212), .ZN(n2385) );
  NAND2_X1 U2327 ( .A1(n2210), .A2(n2212), .ZN(n2382) );
  NAND2_X1 U2328 ( .A1(n2386), .A2(n2387), .ZN(n2212) );
  NAND2_X1 U2329 ( .A1(n2388), .A2(a_3_), .ZN(n2387) );
  NOR2_X1 U2330 ( .A1(n2389), .A2(n2008), .ZN(n2388) );
  NOR2_X1 U2331 ( .A1(n2203), .A2(n2205), .ZN(n2389) );
  NAND2_X1 U2332 ( .A1(n2203), .A2(n2205), .ZN(n2386) );
  NAND2_X1 U2333 ( .A1(n2390), .A2(n2391), .ZN(n2205) );
  NAND2_X1 U2334 ( .A1(n2392), .A2(a_4_), .ZN(n2391) );
  NOR2_X1 U2335 ( .A1(n2393), .A2(n2008), .ZN(n2392) );
  NOR2_X1 U2336 ( .A1(n2173), .A2(n2175), .ZN(n2393) );
  NAND2_X1 U2337 ( .A1(n2173), .A2(n2175), .ZN(n2390) );
  NAND2_X1 U2338 ( .A1(n2168), .A2(n2394), .ZN(n2175) );
  NAND2_X1 U2339 ( .A1(n2167), .A2(n2169), .ZN(n2394) );
  NAND2_X1 U2340 ( .A1(n2395), .A2(n2396), .ZN(n2169) );
  NAND2_X1 U2341 ( .A1(a_5_), .A2(b_15_), .ZN(n2396) );
  INV_X1 U2342 ( .A(n2397), .ZN(n2395) );
  XOR2_X1 U2343 ( .A(n2398), .B(n2399), .Z(n2167) );
  XOR2_X1 U2344 ( .A(n2400), .B(n2401), .Z(n2398) );
  NOR2_X1 U2345 ( .A1(n2023), .A2(n2283), .ZN(n2401) );
  NAND2_X1 U2346 ( .A1(a_5_), .A2(n2397), .ZN(n2168) );
  NAND2_X1 U2347 ( .A1(n2402), .A2(n2403), .ZN(n2397) );
  NAND2_X1 U2348 ( .A1(n2404), .A2(a_6_), .ZN(n2403) );
  NOR2_X1 U2349 ( .A1(n2405), .A2(n2008), .ZN(n2404) );
  NOR2_X1 U2350 ( .A1(n2143), .A2(n2145), .ZN(n2405) );
  NAND2_X1 U2351 ( .A1(n2143), .A2(n2145), .ZN(n2402) );
  NAND2_X1 U2352 ( .A1(n2138), .A2(n2406), .ZN(n2145) );
  NAND2_X1 U2353 ( .A1(n2137), .A2(n2139), .ZN(n2406) );
  NAND2_X1 U2354 ( .A1(n2407), .A2(n2408), .ZN(n2139) );
  NAND2_X1 U2355 ( .A1(a_7_), .A2(b_15_), .ZN(n2408) );
  INV_X1 U2356 ( .A(n2409), .ZN(n2407) );
  XOR2_X1 U2357 ( .A(n2410), .B(n2411), .Z(n2137) );
  XOR2_X1 U2358 ( .A(n2412), .B(n2413), .Z(n2410) );
  NOR2_X1 U2359 ( .A1(n2023), .A2(n2281), .ZN(n2413) );
  NAND2_X1 U2360 ( .A1(a_7_), .A2(n2409), .ZN(n2138) );
  NAND2_X1 U2361 ( .A1(n2414), .A2(n2415), .ZN(n2409) );
  NAND2_X1 U2362 ( .A1(n2416), .A2(a_8_), .ZN(n2415) );
  NOR2_X1 U2363 ( .A1(n2417), .A2(n2008), .ZN(n2416) );
  NOR2_X1 U2364 ( .A1(n2113), .A2(n2116), .ZN(n2417) );
  NAND2_X1 U2365 ( .A1(n2113), .A2(n2116), .ZN(n2414) );
  NAND2_X1 U2366 ( .A1(n2108), .A2(n2418), .ZN(n2116) );
  NAND2_X1 U2367 ( .A1(n2107), .A2(n2109), .ZN(n2418) );
  NAND2_X1 U2368 ( .A1(n2419), .A2(n2420), .ZN(n2109) );
  NAND2_X1 U2369 ( .A1(a_9_), .A2(b_15_), .ZN(n2420) );
  INV_X1 U2370 ( .A(n2421), .ZN(n2419) );
  XNOR2_X1 U2371 ( .A(n2422), .B(n2423), .ZN(n2107) );
  NAND2_X1 U2372 ( .A1(n2424), .A2(n2425), .ZN(n2422) );
  NAND2_X1 U2373 ( .A1(a_9_), .A2(n2421), .ZN(n2108) );
  NAND2_X1 U2374 ( .A1(n2426), .A2(n2427), .ZN(n2421) );
  NAND2_X1 U2375 ( .A1(n2428), .A2(a_10_), .ZN(n2427) );
  NOR2_X1 U2376 ( .A1(n2429), .A2(n2008), .ZN(n2428) );
  NOR2_X1 U2377 ( .A1(n2084), .A2(n2086), .ZN(n2429) );
  NAND2_X1 U2378 ( .A1(n2084), .A2(n2086), .ZN(n2426) );
  NAND2_X1 U2379 ( .A1(n2078), .A2(n2430), .ZN(n2086) );
  NAND2_X1 U2380 ( .A1(n2077), .A2(n2079), .ZN(n2430) );
  NAND2_X1 U2381 ( .A1(n2431), .A2(n2432), .ZN(n2079) );
  NAND2_X1 U2382 ( .A1(a_11_), .A2(b_15_), .ZN(n2432) );
  INV_X1 U2383 ( .A(n2433), .ZN(n2431) );
  XOR2_X1 U2384 ( .A(n2434), .B(n2435), .Z(n2077) );
  XNOR2_X1 U2385 ( .A(n2436), .B(n2437), .ZN(n2434) );
  NAND2_X1 U2386 ( .A1(a_12_), .A2(b_14_), .ZN(n2436) );
  NAND2_X1 U2387 ( .A1(a_11_), .A2(n2433), .ZN(n2078) );
  NAND2_X1 U2388 ( .A1(n2438), .A2(n2439), .ZN(n2433) );
  NAND2_X1 U2389 ( .A1(n2440), .A2(a_12_), .ZN(n2439) );
  NOR2_X1 U2390 ( .A1(n2441), .A2(n2008), .ZN(n2440) );
  NOR2_X1 U2391 ( .A1(n2053), .A2(n2055), .ZN(n2441) );
  NAND2_X1 U2392 ( .A1(n2053), .A2(n2055), .ZN(n2438) );
  NAND2_X1 U2393 ( .A1(n2442), .A2(n2443), .ZN(n2055) );
  NAND2_X1 U2394 ( .A1(n2444), .A2(a_13_), .ZN(n2443) );
  NOR2_X1 U2395 ( .A1(n2445), .A2(n2008), .ZN(n2444) );
  INV_X1 U2396 ( .A(b_15_), .ZN(n2008) );
  NOR2_X1 U2397 ( .A1(n2049), .A2(n2048), .ZN(n2445) );
  NAND2_X1 U2398 ( .A1(n2049), .A2(n2048), .ZN(n2442) );
  NAND2_X1 U2399 ( .A1(n2446), .A2(n2447), .ZN(n2048) );
  NAND2_X1 U2400 ( .A1(b_13_), .A2(n2448), .ZN(n2447) );
  NAND2_X1 U2401 ( .A1(n2018), .A2(n2449), .ZN(n2448) );
  NAND2_X1 U2402 ( .A1(a_15_), .A2(n2023), .ZN(n2449) );
  NAND2_X1 U2403 ( .A1(b_14_), .A2(n2450), .ZN(n2446) );
  NAND2_X1 U2404 ( .A1(n2021), .A2(n2451), .ZN(n2450) );
  NAND2_X1 U2405 ( .A1(a_14_), .A2(n2043), .ZN(n2451) );
  NOR2_X1 U2406 ( .A1(n2275), .A2(n2274), .ZN(n2049) );
  XOR2_X1 U2407 ( .A(n2452), .B(n2453), .Z(n2053) );
  XOR2_X1 U2408 ( .A(n2454), .B(n2455), .Z(n2452) );
  XNOR2_X1 U2409 ( .A(n2456), .B(n2457), .ZN(n2084) );
  NAND2_X1 U2410 ( .A1(n2458), .A2(n2459), .ZN(n2456) );
  XNOR2_X1 U2411 ( .A(n2460), .B(n2461), .ZN(n2113) );
  XNOR2_X1 U2412 ( .A(n2462), .B(n2463), .ZN(n2461) );
  XOR2_X1 U2413 ( .A(n2464), .B(n2465), .Z(n2143) );
  XOR2_X1 U2414 ( .A(n2466), .B(n2467), .Z(n2464) );
  XNOR2_X1 U2415 ( .A(n2468), .B(n2469), .ZN(n2173) );
  XNOR2_X1 U2416 ( .A(n2470), .B(n2471), .ZN(n2469) );
  XOR2_X1 U2417 ( .A(n2472), .B(n2473), .Z(n2203) );
  XNOR2_X1 U2418 ( .A(n2474), .B(n2475), .ZN(n2472) );
  NAND2_X1 U2419 ( .A1(a_4_), .A2(b_14_), .ZN(n2474) );
  XNOR2_X1 U2420 ( .A(n2476), .B(n2477), .ZN(n2210) );
  XNOR2_X1 U2421 ( .A(n2478), .B(n2479), .ZN(n2477) );
  XOR2_X1 U2422 ( .A(n2480), .B(n2481), .Z(n2222) );
  XNOR2_X1 U2423 ( .A(n2482), .B(n2483), .ZN(n2480) );
  NAND2_X1 U2424 ( .A1(a_2_), .A2(b_14_), .ZN(n2482) );
  XOR2_X1 U2425 ( .A(n2484), .B(n2485), .Z(n2238) );
  XOR2_X1 U2426 ( .A(n2486), .B(n2487), .Z(n2485) );
  NAND2_X1 U2427 ( .A1(b_14_), .A2(a_1_), .ZN(n2487) );
  NOR2_X1 U2428 ( .A1(n2488), .A2(n2291), .ZN(n2371) );
  XOR2_X1 U2429 ( .A(n2489), .B(n2490), .Z(n2291) );
  XNOR2_X1 U2430 ( .A(n2491), .B(n2492), .ZN(n2490) );
  NOR2_X1 U2431 ( .A1(n2298), .A2(n2297), .ZN(n2488) );
  NAND2_X1 U2432 ( .A1(n2493), .A2(n2494), .ZN(n2297) );
  NAND2_X1 U2433 ( .A1(n2492), .A2(n2495), .ZN(n2494) );
  OR2_X1 U2434 ( .A1(n2491), .A2(n2489), .ZN(n2495) );
  NOR2_X1 U2435 ( .A1(n2376), .A2(n2023), .ZN(n2492) );
  NAND2_X1 U2436 ( .A1(n2489), .A2(n2491), .ZN(n2493) );
  NAND2_X1 U2437 ( .A1(n2496), .A2(n2497), .ZN(n2491) );
  NAND2_X1 U2438 ( .A1(n2498), .A2(b_14_), .ZN(n2497) );
  NOR2_X1 U2439 ( .A1(n2499), .A2(n2381), .ZN(n2498) );
  NOR2_X1 U2440 ( .A1(n2484), .A2(n2486), .ZN(n2499) );
  NAND2_X1 U2441 ( .A1(n2484), .A2(n2486), .ZN(n2496) );
  NAND2_X1 U2442 ( .A1(n2500), .A2(n2501), .ZN(n2486) );
  NAND2_X1 U2443 ( .A1(n2502), .A2(a_2_), .ZN(n2501) );
  NOR2_X1 U2444 ( .A1(n2503), .A2(n2023), .ZN(n2502) );
  NOR2_X1 U2445 ( .A1(n2481), .A2(n2483), .ZN(n2503) );
  NAND2_X1 U2446 ( .A1(n2481), .A2(n2483), .ZN(n2500) );
  NAND2_X1 U2447 ( .A1(n2504), .A2(n2505), .ZN(n2483) );
  NAND2_X1 U2448 ( .A1(n2479), .A2(n2506), .ZN(n2505) );
  OR2_X1 U2449 ( .A1(n2478), .A2(n2476), .ZN(n2506) );
  NOR2_X1 U2450 ( .A1(n2199), .A2(n2023), .ZN(n2479) );
  NAND2_X1 U2451 ( .A1(n2476), .A2(n2478), .ZN(n2504) );
  NAND2_X1 U2452 ( .A1(n2507), .A2(n2508), .ZN(n2478) );
  NAND2_X1 U2453 ( .A1(n2509), .A2(a_4_), .ZN(n2508) );
  NOR2_X1 U2454 ( .A1(n2510), .A2(n2023), .ZN(n2509) );
  NOR2_X1 U2455 ( .A1(n2473), .A2(n2475), .ZN(n2510) );
  NAND2_X1 U2456 ( .A1(n2473), .A2(n2475), .ZN(n2507) );
  NAND2_X1 U2457 ( .A1(n2511), .A2(n2512), .ZN(n2475) );
  NAND2_X1 U2458 ( .A1(n2471), .A2(n2513), .ZN(n2512) );
  OR2_X1 U2459 ( .A1(n2470), .A2(n2468), .ZN(n2513) );
  NOR2_X1 U2460 ( .A1(n2162), .A2(n2023), .ZN(n2471) );
  NAND2_X1 U2461 ( .A1(n2468), .A2(n2470), .ZN(n2511) );
  NAND2_X1 U2462 ( .A1(n2514), .A2(n2515), .ZN(n2470) );
  NAND2_X1 U2463 ( .A1(n2516), .A2(a_6_), .ZN(n2515) );
  NOR2_X1 U2464 ( .A1(n2517), .A2(n2023), .ZN(n2516) );
  NOR2_X1 U2465 ( .A1(n2399), .A2(n2400), .ZN(n2517) );
  NAND2_X1 U2466 ( .A1(n2399), .A2(n2400), .ZN(n2514) );
  NAND2_X1 U2467 ( .A1(n2518), .A2(n2519), .ZN(n2400) );
  NAND2_X1 U2468 ( .A1(n2467), .A2(n2520), .ZN(n2519) );
  OR2_X1 U2469 ( .A1(n2466), .A2(n2465), .ZN(n2520) );
  NOR2_X1 U2470 ( .A1(n2132), .A2(n2023), .ZN(n2467) );
  NAND2_X1 U2471 ( .A1(n2465), .A2(n2466), .ZN(n2518) );
  NAND2_X1 U2472 ( .A1(n2521), .A2(n2522), .ZN(n2466) );
  NAND2_X1 U2473 ( .A1(n2523), .A2(a_8_), .ZN(n2522) );
  NOR2_X1 U2474 ( .A1(n2524), .A2(n2023), .ZN(n2523) );
  NOR2_X1 U2475 ( .A1(n2411), .A2(n2412), .ZN(n2524) );
  NAND2_X1 U2476 ( .A1(n2411), .A2(n2412), .ZN(n2521) );
  NAND2_X1 U2477 ( .A1(n2525), .A2(n2526), .ZN(n2412) );
  NAND2_X1 U2478 ( .A1(n2463), .A2(n2527), .ZN(n2526) );
  OR2_X1 U2479 ( .A1(n2462), .A2(n2460), .ZN(n2527) );
  NOR2_X1 U2480 ( .A1(n2102), .A2(n2023), .ZN(n2463) );
  NAND2_X1 U2481 ( .A1(n2460), .A2(n2462), .ZN(n2525) );
  NAND2_X1 U2482 ( .A1(n2424), .A2(n2528), .ZN(n2462) );
  NAND2_X1 U2483 ( .A1(n2423), .A2(n2425), .ZN(n2528) );
  NAND2_X1 U2484 ( .A1(n2529), .A2(n2530), .ZN(n2425) );
  NAND2_X1 U2485 ( .A1(a_10_), .A2(b_14_), .ZN(n2530) );
  INV_X1 U2486 ( .A(n2531), .ZN(n2529) );
  XNOR2_X1 U2487 ( .A(n2532), .B(n2533), .ZN(n2423) );
  NAND2_X1 U2488 ( .A1(n2534), .A2(n2535), .ZN(n2532) );
  NAND2_X1 U2489 ( .A1(a_10_), .A2(n2531), .ZN(n2424) );
  NAND2_X1 U2490 ( .A1(n2458), .A2(n2536), .ZN(n2531) );
  NAND2_X1 U2491 ( .A1(n2457), .A2(n2459), .ZN(n2536) );
  NAND2_X1 U2492 ( .A1(n2537), .A2(n2538), .ZN(n2459) );
  NAND2_X1 U2493 ( .A1(a_11_), .A2(b_14_), .ZN(n2538) );
  INV_X1 U2494 ( .A(n2539), .ZN(n2537) );
  XOR2_X1 U2495 ( .A(n2540), .B(n2541), .Z(n2457) );
  XNOR2_X1 U2496 ( .A(n2542), .B(n2543), .ZN(n2540) );
  NAND2_X1 U2497 ( .A1(a_12_), .A2(b_13_), .ZN(n2542) );
  NAND2_X1 U2498 ( .A1(a_11_), .A2(n2539), .ZN(n2458) );
  NAND2_X1 U2499 ( .A1(n2544), .A2(n2545), .ZN(n2539) );
  NAND2_X1 U2500 ( .A1(n2546), .A2(a_12_), .ZN(n2545) );
  NOR2_X1 U2501 ( .A1(n2547), .A2(n2023), .ZN(n2546) );
  NOR2_X1 U2502 ( .A1(n2435), .A2(n2437), .ZN(n2547) );
  NAND2_X1 U2503 ( .A1(n2435), .A2(n2437), .ZN(n2544) );
  NAND2_X1 U2504 ( .A1(n2548), .A2(n2549), .ZN(n2437) );
  NAND2_X1 U2505 ( .A1(n2453), .A2(n2550), .ZN(n2549) );
  OR2_X1 U2506 ( .A1(n2454), .A2(n2455), .ZN(n2550) );
  NOR2_X1 U2507 ( .A1(n2042), .A2(n2023), .ZN(n2453) );
  NAND2_X1 U2508 ( .A1(n2455), .A2(n2454), .ZN(n2548) );
  NAND2_X1 U2509 ( .A1(n2551), .A2(n2552), .ZN(n2454) );
  NAND2_X1 U2510 ( .A1(b_12_), .A2(n2553), .ZN(n2552) );
  NAND2_X1 U2511 ( .A1(n2018), .A2(n2554), .ZN(n2553) );
  NAND2_X1 U2512 ( .A1(a_15_), .A2(n2043), .ZN(n2554) );
  NAND2_X1 U2513 ( .A1(b_13_), .A2(n2555), .ZN(n2551) );
  NAND2_X1 U2514 ( .A1(n2021), .A2(n2556), .ZN(n2555) );
  NAND2_X1 U2515 ( .A1(a_14_), .A2(n2276), .ZN(n2556) );
  AND2_X1 U2516 ( .A1(n2557), .A2(n2558), .ZN(n2455) );
  NOR2_X1 U2517 ( .A1(n2023), .A2(n2043), .ZN(n2557) );
  XNOR2_X1 U2518 ( .A(n2559), .B(n2267), .ZN(n2435) );
  XOR2_X1 U2519 ( .A(n2560), .B(n2561), .Z(n2559) );
  XNOR2_X1 U2520 ( .A(n2562), .B(n2563), .ZN(n2460) );
  NAND2_X1 U2521 ( .A1(n2564), .A2(n2565), .ZN(n2562) );
  XNOR2_X1 U2522 ( .A(n2566), .B(n2567), .ZN(n2411) );
  XNOR2_X1 U2523 ( .A(n2568), .B(n2569), .ZN(n2566) );
  XNOR2_X1 U2524 ( .A(n2570), .B(n2571), .ZN(n2465) );
  XOR2_X1 U2525 ( .A(n2572), .B(n2573), .Z(n2571) );
  NAND2_X1 U2526 ( .A1(a_8_), .A2(b_13_), .ZN(n2573) );
  XNOR2_X1 U2527 ( .A(n2574), .B(n2575), .ZN(n2399) );
  XNOR2_X1 U2528 ( .A(n2576), .B(n2577), .ZN(n2575) );
  XNOR2_X1 U2529 ( .A(n2578), .B(n2579), .ZN(n2468) );
  XOR2_X1 U2530 ( .A(n2580), .B(n2581), .Z(n2579) );
  NAND2_X1 U2531 ( .A1(a_6_), .A2(b_13_), .ZN(n2581) );
  XNOR2_X1 U2532 ( .A(n2582), .B(n2583), .ZN(n2473) );
  XNOR2_X1 U2533 ( .A(n2584), .B(n2585), .ZN(n2583) );
  XOR2_X1 U2534 ( .A(n2586), .B(n2587), .Z(n2476) );
  XNOR2_X1 U2535 ( .A(n2588), .B(n2589), .ZN(n2586) );
  NAND2_X1 U2536 ( .A1(a_4_), .A2(b_13_), .ZN(n2588) );
  XNOR2_X1 U2537 ( .A(n2590), .B(n2591), .ZN(n2481) );
  XNOR2_X1 U2538 ( .A(n2592), .B(n2593), .ZN(n2591) );
  XNOR2_X1 U2539 ( .A(n2594), .B(n2595), .ZN(n2484) );
  XOR2_X1 U2540 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND2_X1 U2541 ( .A1(a_2_), .A2(b_13_), .ZN(n2597) );
  XOR2_X1 U2542 ( .A(n2598), .B(n2599), .Z(n2489) );
  XOR2_X1 U2543 ( .A(n2600), .B(n2601), .Z(n2598) );
  NOR2_X1 U2544 ( .A1(n2381), .A2(n2043), .ZN(n2601) );
  XNOR2_X1 U2545 ( .A(n2602), .B(n2603), .ZN(n2298) );
  XOR2_X1 U2546 ( .A(n2604), .B(n2605), .Z(n2602) );
  INV_X1 U2547 ( .A(n2309), .ZN(n2306) );
  NAND2_X1 U2548 ( .A1(n2606), .A2(n2369), .ZN(n2309) );
  NAND2_X1 U2549 ( .A1(n2607), .A2(n2608), .ZN(n2369) );
  OR2_X1 U2550 ( .A1(n2608), .A2(n2607), .ZN(n2606) );
  AND2_X1 U2551 ( .A1(n2609), .A2(n2610), .ZN(n2607) );
  NAND2_X1 U2552 ( .A1(n2603), .A2(n2611), .ZN(n2610) );
  NAND2_X1 U2553 ( .A1(n2605), .A2(n2604), .ZN(n2611) );
  XOR2_X1 U2554 ( .A(n2612), .B(n2613), .Z(n2603) );
  XNOR2_X1 U2555 ( .A(n2614), .B(n2615), .ZN(n2612) );
  OR2_X1 U2556 ( .A1(n2604), .A2(n2605), .ZN(n2609) );
  NOR2_X1 U2557 ( .A1(n2376), .A2(n2043), .ZN(n2605) );
  NAND2_X1 U2558 ( .A1(n2616), .A2(n2617), .ZN(n2604) );
  NAND2_X1 U2559 ( .A1(n2618), .A2(b_13_), .ZN(n2617) );
  NOR2_X1 U2560 ( .A1(n2619), .A2(n2381), .ZN(n2618) );
  NOR2_X1 U2561 ( .A1(n2599), .A2(n2600), .ZN(n2619) );
  NAND2_X1 U2562 ( .A1(n2599), .A2(n2600), .ZN(n2616) );
  NAND2_X1 U2563 ( .A1(n2620), .A2(n2621), .ZN(n2600) );
  NAND2_X1 U2564 ( .A1(n2622), .A2(a_2_), .ZN(n2621) );
  NOR2_X1 U2565 ( .A1(n2623), .A2(n2043), .ZN(n2622) );
  NOR2_X1 U2566 ( .A1(n2594), .A2(n2596), .ZN(n2623) );
  NAND2_X1 U2567 ( .A1(n2594), .A2(n2596), .ZN(n2620) );
  NAND2_X1 U2568 ( .A1(n2624), .A2(n2625), .ZN(n2596) );
  NAND2_X1 U2569 ( .A1(n2593), .A2(n2626), .ZN(n2625) );
  OR2_X1 U2570 ( .A1(n2592), .A2(n2590), .ZN(n2626) );
  NOR2_X1 U2571 ( .A1(n2199), .A2(n2043), .ZN(n2593) );
  NAND2_X1 U2572 ( .A1(n2590), .A2(n2592), .ZN(n2624) );
  NAND2_X1 U2573 ( .A1(n2627), .A2(n2628), .ZN(n2592) );
  NAND2_X1 U2574 ( .A1(n2629), .A2(a_4_), .ZN(n2628) );
  NOR2_X1 U2575 ( .A1(n2630), .A2(n2043), .ZN(n2629) );
  NOR2_X1 U2576 ( .A1(n2587), .A2(n2589), .ZN(n2630) );
  NAND2_X1 U2577 ( .A1(n2587), .A2(n2589), .ZN(n2627) );
  NAND2_X1 U2578 ( .A1(n2631), .A2(n2632), .ZN(n2589) );
  NAND2_X1 U2579 ( .A1(n2585), .A2(n2633), .ZN(n2632) );
  OR2_X1 U2580 ( .A1(n2584), .A2(n2582), .ZN(n2633) );
  NOR2_X1 U2581 ( .A1(n2162), .A2(n2043), .ZN(n2585) );
  NAND2_X1 U2582 ( .A1(n2582), .A2(n2584), .ZN(n2631) );
  NAND2_X1 U2583 ( .A1(n2634), .A2(n2635), .ZN(n2584) );
  NAND2_X1 U2584 ( .A1(n2636), .A2(a_6_), .ZN(n2635) );
  NOR2_X1 U2585 ( .A1(n2637), .A2(n2043), .ZN(n2636) );
  NOR2_X1 U2586 ( .A1(n2578), .A2(n2580), .ZN(n2637) );
  NAND2_X1 U2587 ( .A1(n2578), .A2(n2580), .ZN(n2634) );
  NAND2_X1 U2588 ( .A1(n2638), .A2(n2639), .ZN(n2580) );
  NAND2_X1 U2589 ( .A1(n2577), .A2(n2640), .ZN(n2639) );
  OR2_X1 U2590 ( .A1(n2576), .A2(n2574), .ZN(n2640) );
  NOR2_X1 U2591 ( .A1(n2132), .A2(n2043), .ZN(n2577) );
  NAND2_X1 U2592 ( .A1(n2574), .A2(n2576), .ZN(n2638) );
  NAND2_X1 U2593 ( .A1(n2641), .A2(n2642), .ZN(n2576) );
  NAND2_X1 U2594 ( .A1(n2643), .A2(a_8_), .ZN(n2642) );
  NOR2_X1 U2595 ( .A1(n2644), .A2(n2043), .ZN(n2643) );
  NOR2_X1 U2596 ( .A1(n2570), .A2(n2572), .ZN(n2644) );
  NAND2_X1 U2597 ( .A1(n2570), .A2(n2572), .ZN(n2641) );
  NAND2_X1 U2598 ( .A1(n2645), .A2(n2646), .ZN(n2572) );
  NAND2_X1 U2599 ( .A1(n2569), .A2(n2647), .ZN(n2646) );
  NAND2_X1 U2600 ( .A1(n2568), .A2(n2567), .ZN(n2647) );
  NOR2_X1 U2601 ( .A1(n2102), .A2(n2043), .ZN(n2569) );
  OR2_X1 U2602 ( .A1(n2567), .A2(n2568), .ZN(n2645) );
  AND2_X1 U2603 ( .A1(n2564), .A2(n2648), .ZN(n2568) );
  NAND2_X1 U2604 ( .A1(n2563), .A2(n2565), .ZN(n2648) );
  NAND2_X1 U2605 ( .A1(n2649), .A2(n2650), .ZN(n2565) );
  NAND2_X1 U2606 ( .A1(a_10_), .A2(b_13_), .ZN(n2650) );
  INV_X1 U2607 ( .A(n2651), .ZN(n2649) );
  XNOR2_X1 U2608 ( .A(n2652), .B(n2653), .ZN(n2563) );
  NAND2_X1 U2609 ( .A1(n2654), .A2(n2655), .ZN(n2652) );
  NAND2_X1 U2610 ( .A1(a_10_), .A2(n2651), .ZN(n2564) );
  NAND2_X1 U2611 ( .A1(n2534), .A2(n2656), .ZN(n2651) );
  NAND2_X1 U2612 ( .A1(n2533), .A2(n2535), .ZN(n2656) );
  NAND2_X1 U2613 ( .A1(n2657), .A2(n2658), .ZN(n2535) );
  NAND2_X1 U2614 ( .A1(a_11_), .A2(b_13_), .ZN(n2658) );
  INV_X1 U2615 ( .A(n2659), .ZN(n2657) );
  XOR2_X1 U2616 ( .A(n2660), .B(n2661), .Z(n2533) );
  XOR2_X1 U2617 ( .A(n2061), .B(n2662), .Z(n2660) );
  NAND2_X1 U2618 ( .A1(a_11_), .A2(n2659), .ZN(n2534) );
  NAND2_X1 U2619 ( .A1(n2663), .A2(n2664), .ZN(n2659) );
  NAND2_X1 U2620 ( .A1(n2665), .A2(a_12_), .ZN(n2664) );
  NOR2_X1 U2621 ( .A1(n2666), .A2(n2043), .ZN(n2665) );
  NOR2_X1 U2622 ( .A1(n2541), .A2(n2543), .ZN(n2666) );
  NAND2_X1 U2623 ( .A1(n2541), .A2(n2543), .ZN(n2663) );
  NAND2_X1 U2624 ( .A1(n2667), .A2(n2668), .ZN(n2543) );
  NAND2_X1 U2625 ( .A1(n2037), .A2(n2669), .ZN(n2668) );
  OR2_X1 U2626 ( .A1(n2560), .A2(n2561), .ZN(n2669) );
  INV_X1 U2627 ( .A(n2267), .ZN(n2037) );
  NAND2_X1 U2628 ( .A1(a_13_), .A2(b_13_), .ZN(n2267) );
  NAND2_X1 U2629 ( .A1(n2561), .A2(n2560), .ZN(n2667) );
  NAND2_X1 U2630 ( .A1(n2670), .A2(n2671), .ZN(n2560) );
  NAND2_X1 U2631 ( .A1(b_11_), .A2(n2672), .ZN(n2671) );
  NAND2_X1 U2632 ( .A1(n2018), .A2(n2673), .ZN(n2672) );
  NAND2_X1 U2633 ( .A1(a_15_), .A2(n2276), .ZN(n2673) );
  NAND2_X1 U2634 ( .A1(b_12_), .A2(n2674), .ZN(n2670) );
  NAND2_X1 U2635 ( .A1(n2021), .A2(n2675), .ZN(n2674) );
  NAND2_X1 U2636 ( .A1(a_14_), .A2(n2073), .ZN(n2675) );
  AND2_X1 U2637 ( .A1(n2676), .A2(n2558), .ZN(n2561) );
  NOR2_X1 U2638 ( .A1(n2043), .A2(n2276), .ZN(n2676) );
  XOR2_X1 U2639 ( .A(n2677), .B(n2678), .Z(n2541) );
  XOR2_X1 U2640 ( .A(n2679), .B(n2680), .Z(n2677) );
  XOR2_X1 U2641 ( .A(n2681), .B(n2682), .Z(n2567) );
  NAND2_X1 U2642 ( .A1(n2683), .A2(n2684), .ZN(n2681) );
  XNOR2_X1 U2643 ( .A(n2685), .B(n2686), .ZN(n2570) );
  XNOR2_X1 U2644 ( .A(n2687), .B(n2688), .ZN(n2686) );
  XOR2_X1 U2645 ( .A(n2689), .B(n2690), .Z(n2574) );
  XOR2_X1 U2646 ( .A(n2691), .B(n2692), .Z(n2689) );
  NOR2_X1 U2647 ( .A1(n2276), .A2(n2281), .ZN(n2692) );
  XNOR2_X1 U2648 ( .A(n2693), .B(n2694), .ZN(n2578) );
  XNOR2_X1 U2649 ( .A(n2695), .B(n2696), .ZN(n2694) );
  XOR2_X1 U2650 ( .A(n2697), .B(n2698), .Z(n2582) );
  XOR2_X1 U2651 ( .A(n2699), .B(n2700), .Z(n2697) );
  NOR2_X1 U2652 ( .A1(n2276), .A2(n2283), .ZN(n2700) );
  XNOR2_X1 U2653 ( .A(n2701), .B(n2702), .ZN(n2587) );
  XNOR2_X1 U2654 ( .A(n2703), .B(n2704), .ZN(n2702) );
  XOR2_X1 U2655 ( .A(n2705), .B(n2706), .Z(n2590) );
  XNOR2_X1 U2656 ( .A(n2707), .B(n2708), .ZN(n2705) );
  NAND2_X1 U2657 ( .A1(a_4_), .A2(b_12_), .ZN(n2707) );
  XNOR2_X1 U2658 ( .A(n2709), .B(n2710), .ZN(n2594) );
  XOR2_X1 U2659 ( .A(n2711), .B(n2712), .Z(n2710) );
  NAND2_X1 U2660 ( .A1(a_3_), .A2(b_12_), .ZN(n2712) );
  XOR2_X1 U2661 ( .A(n2713), .B(n2714), .Z(n2599) );
  XOR2_X1 U2662 ( .A(n2715), .B(n2716), .Z(n2713) );
  XOR2_X1 U2663 ( .A(n2717), .B(n2718), .Z(n2608) );
  XOR2_X1 U2664 ( .A(n2719), .B(n2720), .Z(n2717) );
  NOR2_X1 U2665 ( .A1(n2276), .A2(n2376), .ZN(n2720) );
  XNOR2_X1 U2666 ( .A(n2354), .B(n2353), .ZN(n2312) );
  XNOR2_X1 U2667 ( .A(n2721), .B(n2364), .ZN(n2353) );
  XOR2_X1 U2668 ( .A(n2722), .B(n2723), .Z(n2364) );
  XNOR2_X1 U2669 ( .A(n2724), .B(n2725), .ZN(n2723) );
  XOR2_X1 U2670 ( .A(n2367), .B(n2366), .Z(n2721) );
  NOR2_X1 U2671 ( .A1(n2376), .A2(n2073), .ZN(n2366) );
  NAND2_X1 U2672 ( .A1(n2726), .A2(n2727), .ZN(n2367) );
  NAND2_X1 U2673 ( .A1(n2728), .A2(b_11_), .ZN(n2727) );
  NOR2_X1 U2674 ( .A1(n2729), .A2(n2381), .ZN(n2728) );
  NOR2_X1 U2675 ( .A1(n2730), .A2(n2731), .ZN(n2729) );
  NAND2_X1 U2676 ( .A1(n2730), .A2(n2731), .ZN(n2726) );
  NAND2_X1 U2677 ( .A1(n2732), .A2(n2733), .ZN(n2354) );
  NAND2_X1 U2678 ( .A1(n2734), .A2(a_0_), .ZN(n2733) );
  NOR2_X1 U2679 ( .A1(n2735), .A2(n2276), .ZN(n2734) );
  NOR2_X1 U2680 ( .A1(n2718), .A2(n2719), .ZN(n2735) );
  NAND2_X1 U2681 ( .A1(n2718), .A2(n2719), .ZN(n2732) );
  NAND2_X1 U2682 ( .A1(n2736), .A2(n2737), .ZN(n2719) );
  NAND2_X1 U2683 ( .A1(n2615), .A2(n2738), .ZN(n2737) );
  NAND2_X1 U2684 ( .A1(n2614), .A2(n2613), .ZN(n2738) );
  NOR2_X1 U2685 ( .A1(n2276), .A2(n2381), .ZN(n2615) );
  OR2_X1 U2686 ( .A1(n2613), .A2(n2614), .ZN(n2736) );
  AND2_X1 U2687 ( .A1(n2739), .A2(n2740), .ZN(n2614) );
  NAND2_X1 U2688 ( .A1(n2716), .A2(n2741), .ZN(n2740) );
  OR2_X1 U2689 ( .A1(n2715), .A2(n2714), .ZN(n2741) );
  NOR2_X1 U2690 ( .A1(n2287), .A2(n2276), .ZN(n2716) );
  NAND2_X1 U2691 ( .A1(n2714), .A2(n2715), .ZN(n2739) );
  NAND2_X1 U2692 ( .A1(n2742), .A2(n2743), .ZN(n2715) );
  NAND2_X1 U2693 ( .A1(n2744), .A2(a_3_), .ZN(n2743) );
  NOR2_X1 U2694 ( .A1(n2745), .A2(n2276), .ZN(n2744) );
  NOR2_X1 U2695 ( .A1(n2709), .A2(n2711), .ZN(n2745) );
  NAND2_X1 U2696 ( .A1(n2709), .A2(n2711), .ZN(n2742) );
  NAND2_X1 U2697 ( .A1(n2746), .A2(n2747), .ZN(n2711) );
  NAND2_X1 U2698 ( .A1(n2748), .A2(a_4_), .ZN(n2747) );
  NOR2_X1 U2699 ( .A1(n2749), .A2(n2276), .ZN(n2748) );
  NOR2_X1 U2700 ( .A1(n2706), .A2(n2708), .ZN(n2749) );
  NAND2_X1 U2701 ( .A1(n2706), .A2(n2708), .ZN(n2746) );
  NAND2_X1 U2702 ( .A1(n2750), .A2(n2751), .ZN(n2708) );
  NAND2_X1 U2703 ( .A1(n2704), .A2(n2752), .ZN(n2751) );
  OR2_X1 U2704 ( .A1(n2703), .A2(n2701), .ZN(n2752) );
  NOR2_X1 U2705 ( .A1(n2162), .A2(n2276), .ZN(n2704) );
  NAND2_X1 U2706 ( .A1(n2701), .A2(n2703), .ZN(n2750) );
  NAND2_X1 U2707 ( .A1(n2753), .A2(n2754), .ZN(n2703) );
  NAND2_X1 U2708 ( .A1(n2755), .A2(a_6_), .ZN(n2754) );
  NOR2_X1 U2709 ( .A1(n2756), .A2(n2276), .ZN(n2755) );
  NOR2_X1 U2710 ( .A1(n2698), .A2(n2699), .ZN(n2756) );
  NAND2_X1 U2711 ( .A1(n2698), .A2(n2699), .ZN(n2753) );
  NAND2_X1 U2712 ( .A1(n2757), .A2(n2758), .ZN(n2699) );
  NAND2_X1 U2713 ( .A1(n2696), .A2(n2759), .ZN(n2758) );
  OR2_X1 U2714 ( .A1(n2695), .A2(n2693), .ZN(n2759) );
  NOR2_X1 U2715 ( .A1(n2132), .A2(n2276), .ZN(n2696) );
  NAND2_X1 U2716 ( .A1(n2693), .A2(n2695), .ZN(n2757) );
  NAND2_X1 U2717 ( .A1(n2760), .A2(n2761), .ZN(n2695) );
  NAND2_X1 U2718 ( .A1(n2762), .A2(a_8_), .ZN(n2761) );
  NOR2_X1 U2719 ( .A1(n2763), .A2(n2276), .ZN(n2762) );
  NOR2_X1 U2720 ( .A1(n2690), .A2(n2691), .ZN(n2763) );
  NAND2_X1 U2721 ( .A1(n2690), .A2(n2691), .ZN(n2760) );
  NAND2_X1 U2722 ( .A1(n2764), .A2(n2765), .ZN(n2691) );
  NAND2_X1 U2723 ( .A1(n2688), .A2(n2766), .ZN(n2765) );
  OR2_X1 U2724 ( .A1(n2687), .A2(n2685), .ZN(n2766) );
  NOR2_X1 U2725 ( .A1(n2102), .A2(n2276), .ZN(n2688) );
  NAND2_X1 U2726 ( .A1(n2685), .A2(n2687), .ZN(n2764) );
  NAND2_X1 U2727 ( .A1(n2683), .A2(n2767), .ZN(n2687) );
  NAND2_X1 U2728 ( .A1(n2682), .A2(n2684), .ZN(n2767) );
  NAND2_X1 U2729 ( .A1(n2768), .A2(n2769), .ZN(n2684) );
  NAND2_X1 U2730 ( .A1(a_10_), .A2(b_12_), .ZN(n2769) );
  INV_X1 U2731 ( .A(n2770), .ZN(n2768) );
  XNOR2_X1 U2732 ( .A(n2771), .B(n2772), .ZN(n2682) );
  XOR2_X1 U2733 ( .A(n2263), .B(n2773), .Z(n2772) );
  NAND2_X1 U2734 ( .A1(a_10_), .A2(n2770), .ZN(n2683) );
  NAND2_X1 U2735 ( .A1(n2654), .A2(n2774), .ZN(n2770) );
  NAND2_X1 U2736 ( .A1(n2653), .A2(n2655), .ZN(n2774) );
  NAND2_X1 U2737 ( .A1(n2775), .A2(n2776), .ZN(n2655) );
  NAND2_X1 U2738 ( .A1(a_11_), .A2(b_12_), .ZN(n2776) );
  INV_X1 U2739 ( .A(n2777), .ZN(n2775) );
  XOR2_X1 U2740 ( .A(n2778), .B(n2779), .Z(n2653) );
  XNOR2_X1 U2741 ( .A(n2780), .B(n2781), .ZN(n2778) );
  NAND2_X1 U2742 ( .A1(b_11_), .A2(a_12_), .ZN(n2780) );
  NAND2_X1 U2743 ( .A1(a_11_), .A2(n2777), .ZN(n2654) );
  NAND2_X1 U2744 ( .A1(n2782), .A2(n2783), .ZN(n2777) );
  NAND2_X1 U2745 ( .A1(n2661), .A2(n2784), .ZN(n2783) );
  NAND2_X1 U2746 ( .A1(n2662), .A2(n2061), .ZN(n2784) );
  INV_X1 U2747 ( .A(n2785), .ZN(n2662) );
  XOR2_X1 U2748 ( .A(n2786), .B(n2787), .Z(n2661) );
  XOR2_X1 U2749 ( .A(n2788), .B(n2789), .Z(n2786) );
  NAND2_X1 U2750 ( .A1(n2790), .A2(n2785), .ZN(n2782) );
  NAND2_X1 U2751 ( .A1(n2791), .A2(n2792), .ZN(n2785) );
  NAND2_X1 U2752 ( .A1(n2678), .A2(n2793), .ZN(n2792) );
  OR2_X1 U2753 ( .A1(n2679), .A2(n2680), .ZN(n2793) );
  NOR2_X1 U2754 ( .A1(n2276), .A2(n2042), .ZN(n2678) );
  NAND2_X1 U2755 ( .A1(n2680), .A2(n2679), .ZN(n2791) );
  NAND2_X1 U2756 ( .A1(n2794), .A2(n2795), .ZN(n2679) );
  NAND2_X1 U2757 ( .A1(b_10_), .A2(n2796), .ZN(n2795) );
  NAND2_X1 U2758 ( .A1(n2018), .A2(n2797), .ZN(n2796) );
  NAND2_X1 U2759 ( .A1(a_15_), .A2(n2073), .ZN(n2797) );
  NAND2_X1 U2760 ( .A1(b_11_), .A2(n2798), .ZN(n2794) );
  NAND2_X1 U2761 ( .A1(n2021), .A2(n2799), .ZN(n2798) );
  NAND2_X1 U2762 ( .A1(a_14_), .A2(n2278), .ZN(n2799) );
  AND2_X1 U2763 ( .A1(n2800), .A2(n2558), .ZN(n2680) );
  NOR2_X1 U2764 ( .A1(n2073), .A2(n2276), .ZN(n2800) );
  INV_X1 U2765 ( .A(n2061), .ZN(n2790) );
  NAND2_X1 U2766 ( .A1(b_12_), .A2(a_12_), .ZN(n2061) );
  XNOR2_X1 U2767 ( .A(n2801), .B(n2802), .ZN(n2685) );
  NAND2_X1 U2768 ( .A1(n2803), .A2(n2804), .ZN(n2801) );
  XNOR2_X1 U2769 ( .A(n2805), .B(n2806), .ZN(n2690) );
  XNOR2_X1 U2770 ( .A(n2807), .B(n2808), .ZN(n2806) );
  XOR2_X1 U2771 ( .A(n2809), .B(n2810), .Z(n2693) );
  XOR2_X1 U2772 ( .A(n2811), .B(n2812), .Z(n2809) );
  NOR2_X1 U2773 ( .A1(n2073), .A2(n2281), .ZN(n2812) );
  XNOR2_X1 U2774 ( .A(n2813), .B(n2814), .ZN(n2698) );
  XNOR2_X1 U2775 ( .A(n2815), .B(n2816), .ZN(n2814) );
  XOR2_X1 U2776 ( .A(n2817), .B(n2818), .Z(n2701) );
  XOR2_X1 U2777 ( .A(n2819), .B(n2820), .Z(n2817) );
  NOR2_X1 U2778 ( .A1(n2073), .A2(n2283), .ZN(n2820) );
  XNOR2_X1 U2779 ( .A(n2821), .B(n2822), .ZN(n2706) );
  XNOR2_X1 U2780 ( .A(n2823), .B(n2824), .ZN(n2822) );
  XNOR2_X1 U2781 ( .A(n2825), .B(n2826), .ZN(n2709) );
  XNOR2_X1 U2782 ( .A(n2827), .B(n2828), .ZN(n2825) );
  XOR2_X1 U2783 ( .A(n2829), .B(n2830), .Z(n2714) );
  XOR2_X1 U2784 ( .A(n2831), .B(n2832), .Z(n2829) );
  NOR2_X1 U2785 ( .A1(n2073), .A2(n2199), .ZN(n2832) );
  XOR2_X1 U2786 ( .A(n2833), .B(n2834), .Z(n2613) );
  XOR2_X1 U2787 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND2_X1 U2788 ( .A1(a_2_), .A2(b_11_), .ZN(n2836) );
  XNOR2_X1 U2789 ( .A(n2730), .B(n2837), .ZN(n2718) );
  XOR2_X1 U2790 ( .A(n2731), .B(n2838), .Z(n2837) );
  NAND2_X1 U2791 ( .A1(b_11_), .A2(a_1_), .ZN(n2838) );
  NAND2_X1 U2792 ( .A1(n2839), .A2(n2840), .ZN(n2731) );
  NAND2_X1 U2793 ( .A1(n2841), .A2(a_2_), .ZN(n2840) );
  NOR2_X1 U2794 ( .A1(n2842), .A2(n2073), .ZN(n2841) );
  NOR2_X1 U2795 ( .A1(n2833), .A2(n2835), .ZN(n2842) );
  NAND2_X1 U2796 ( .A1(n2833), .A2(n2835), .ZN(n2839) );
  NAND2_X1 U2797 ( .A1(n2843), .A2(n2844), .ZN(n2835) );
  NAND2_X1 U2798 ( .A1(n2845), .A2(a_3_), .ZN(n2844) );
  NOR2_X1 U2799 ( .A1(n2846), .A2(n2073), .ZN(n2845) );
  NOR2_X1 U2800 ( .A1(n2830), .A2(n2831), .ZN(n2846) );
  NAND2_X1 U2801 ( .A1(n2830), .A2(n2831), .ZN(n2843) );
  NAND2_X1 U2802 ( .A1(n2847), .A2(n2848), .ZN(n2831) );
  NAND2_X1 U2803 ( .A1(n2828), .A2(n2849), .ZN(n2848) );
  NAND2_X1 U2804 ( .A1(n2827), .A2(n2826), .ZN(n2849) );
  NOR2_X1 U2805 ( .A1(n2285), .A2(n2073), .ZN(n2828) );
  OR2_X1 U2806 ( .A1(n2826), .A2(n2827), .ZN(n2847) );
  AND2_X1 U2807 ( .A1(n2850), .A2(n2851), .ZN(n2827) );
  NAND2_X1 U2808 ( .A1(n2824), .A2(n2852), .ZN(n2851) );
  OR2_X1 U2809 ( .A1(n2823), .A2(n2821), .ZN(n2852) );
  NOR2_X1 U2810 ( .A1(n2162), .A2(n2073), .ZN(n2824) );
  NAND2_X1 U2811 ( .A1(n2821), .A2(n2823), .ZN(n2850) );
  NAND2_X1 U2812 ( .A1(n2853), .A2(n2854), .ZN(n2823) );
  NAND2_X1 U2813 ( .A1(n2855), .A2(a_6_), .ZN(n2854) );
  NOR2_X1 U2814 ( .A1(n2856), .A2(n2073), .ZN(n2855) );
  NOR2_X1 U2815 ( .A1(n2818), .A2(n2819), .ZN(n2856) );
  NAND2_X1 U2816 ( .A1(n2818), .A2(n2819), .ZN(n2853) );
  NAND2_X1 U2817 ( .A1(n2857), .A2(n2858), .ZN(n2819) );
  NAND2_X1 U2818 ( .A1(n2816), .A2(n2859), .ZN(n2858) );
  OR2_X1 U2819 ( .A1(n2815), .A2(n2813), .ZN(n2859) );
  NOR2_X1 U2820 ( .A1(n2132), .A2(n2073), .ZN(n2816) );
  NAND2_X1 U2821 ( .A1(n2813), .A2(n2815), .ZN(n2857) );
  NAND2_X1 U2822 ( .A1(n2860), .A2(n2861), .ZN(n2815) );
  NAND2_X1 U2823 ( .A1(n2862), .A2(a_8_), .ZN(n2861) );
  NOR2_X1 U2824 ( .A1(n2863), .A2(n2073), .ZN(n2862) );
  NOR2_X1 U2825 ( .A1(n2810), .A2(n2811), .ZN(n2863) );
  NAND2_X1 U2826 ( .A1(n2810), .A2(n2811), .ZN(n2860) );
  NAND2_X1 U2827 ( .A1(n2864), .A2(n2865), .ZN(n2811) );
  NAND2_X1 U2828 ( .A1(n2808), .A2(n2866), .ZN(n2865) );
  OR2_X1 U2829 ( .A1(n2807), .A2(n2805), .ZN(n2866) );
  NOR2_X1 U2830 ( .A1(n2102), .A2(n2073), .ZN(n2808) );
  NAND2_X1 U2831 ( .A1(n2805), .A2(n2807), .ZN(n2864) );
  NAND2_X1 U2832 ( .A1(n2803), .A2(n2867), .ZN(n2807) );
  NAND2_X1 U2833 ( .A1(n2802), .A2(n2804), .ZN(n2867) );
  NAND2_X1 U2834 ( .A1(n2868), .A2(n2869), .ZN(n2804) );
  NAND2_X1 U2835 ( .A1(a_10_), .A2(b_11_), .ZN(n2869) );
  INV_X1 U2836 ( .A(n2870), .ZN(n2868) );
  XNOR2_X1 U2837 ( .A(n2871), .B(n2872), .ZN(n2802) );
  NAND2_X1 U2838 ( .A1(n2873), .A2(n2874), .ZN(n2871) );
  NAND2_X1 U2839 ( .A1(a_10_), .A2(n2870), .ZN(n2803) );
  NAND2_X1 U2840 ( .A1(n2875), .A2(n2876), .ZN(n2870) );
  NAND2_X1 U2841 ( .A1(n2771), .A2(n2877), .ZN(n2876) );
  OR2_X1 U2842 ( .A1(n2773), .A2(n2067), .ZN(n2877) );
  XOR2_X1 U2843 ( .A(n2878), .B(n2879), .Z(n2771) );
  XNOR2_X1 U2844 ( .A(n2880), .B(n2881), .ZN(n2878) );
  NAND2_X1 U2845 ( .A1(b_10_), .A2(a_12_), .ZN(n2880) );
  NAND2_X1 U2846 ( .A1(n2067), .A2(n2773), .ZN(n2875) );
  NAND2_X1 U2847 ( .A1(n2882), .A2(n2883), .ZN(n2773) );
  NAND2_X1 U2848 ( .A1(n2884), .A2(b_11_), .ZN(n2883) );
  NOR2_X1 U2849 ( .A1(n2885), .A2(n2277), .ZN(n2884) );
  NOR2_X1 U2850 ( .A1(n2779), .A2(n2781), .ZN(n2885) );
  NAND2_X1 U2851 ( .A1(n2779), .A2(n2781), .ZN(n2882) );
  NAND2_X1 U2852 ( .A1(n2886), .A2(n2887), .ZN(n2781) );
  NAND2_X1 U2853 ( .A1(n2787), .A2(n2888), .ZN(n2887) );
  OR2_X1 U2854 ( .A1(n2788), .A2(n2789), .ZN(n2888) );
  NOR2_X1 U2855 ( .A1(n2073), .A2(n2042), .ZN(n2787) );
  NAND2_X1 U2856 ( .A1(n2789), .A2(n2788), .ZN(n2886) );
  NAND2_X1 U2857 ( .A1(n2889), .A2(n2890), .ZN(n2788) );
  NAND2_X1 U2858 ( .A1(b_10_), .A2(n2891), .ZN(n2890) );
  NAND2_X1 U2859 ( .A1(n2021), .A2(n2892), .ZN(n2891) );
  NAND2_X1 U2860 ( .A1(a_14_), .A2(n2103), .ZN(n2892) );
  NAND2_X1 U2861 ( .A1(b_9_), .A2(n2893), .ZN(n2889) );
  NAND2_X1 U2862 ( .A1(n2018), .A2(n2894), .ZN(n2893) );
  NAND2_X1 U2863 ( .A1(a_15_), .A2(n2278), .ZN(n2894) );
  AND2_X1 U2864 ( .A1(n2895), .A2(n2558), .ZN(n2789) );
  NOR2_X1 U2865 ( .A1(n2073), .A2(n2278), .ZN(n2895) );
  XOR2_X1 U2866 ( .A(n2896), .B(n2897), .Z(n2779) );
  XOR2_X1 U2867 ( .A(n2898), .B(n2899), .Z(n2896) );
  INV_X1 U2868 ( .A(n2263), .ZN(n2067) );
  NAND2_X1 U2869 ( .A1(a_11_), .A2(b_11_), .ZN(n2263) );
  XOR2_X1 U2870 ( .A(n2900), .B(n2901), .Z(n2805) );
  XOR2_X1 U2871 ( .A(n2091), .B(n2902), .Z(n2900) );
  XNOR2_X1 U2872 ( .A(n2903), .B(n2904), .ZN(n2810) );
  XNOR2_X1 U2873 ( .A(n2905), .B(n2906), .ZN(n2904) );
  XOR2_X1 U2874 ( .A(n2907), .B(n2908), .Z(n2813) );
  XOR2_X1 U2875 ( .A(n2909), .B(n2910), .Z(n2907) );
  NOR2_X1 U2876 ( .A1(n2278), .A2(n2281), .ZN(n2910) );
  XNOR2_X1 U2877 ( .A(n2911), .B(n2912), .ZN(n2818) );
  XNOR2_X1 U2878 ( .A(n2913), .B(n2914), .ZN(n2912) );
  XOR2_X1 U2879 ( .A(n2915), .B(n2916), .Z(n2821) );
  XOR2_X1 U2880 ( .A(n2917), .B(n2918), .Z(n2915) );
  NOR2_X1 U2881 ( .A1(n2278), .A2(n2283), .ZN(n2918) );
  XOR2_X1 U2882 ( .A(n2919), .B(n2920), .Z(n2826) );
  XOR2_X1 U2883 ( .A(n2921), .B(n2922), .Z(n2920) );
  NAND2_X1 U2884 ( .A1(a_5_), .A2(b_10_), .ZN(n2922) );
  XNOR2_X1 U2885 ( .A(n2923), .B(n2924), .ZN(n2830) );
  XNOR2_X1 U2886 ( .A(n2925), .B(n2926), .ZN(n2924) );
  XNOR2_X1 U2887 ( .A(n2927), .B(n2928), .ZN(n2833) );
  XNOR2_X1 U2888 ( .A(n2929), .B(n2930), .ZN(n2927) );
  XOR2_X1 U2889 ( .A(n2931), .B(n2932), .Z(n2730) );
  XOR2_X1 U2890 ( .A(n2933), .B(n2934), .Z(n2931) );
  NOR2_X1 U2891 ( .A1(n2278), .A2(n2287), .ZN(n2934) );
  NAND2_X1 U2892 ( .A1(n2935), .A2(n2936), .ZN(n1974) );
  NAND2_X1 U2893 ( .A1(n2351), .A2(n2350), .ZN(n2936) );
  XOR2_X1 U2894 ( .A(n2937), .B(n2938), .Z(n2935) );
  NAND2_X1 U2895 ( .A1(n2939), .A2(n2940), .ZN(n1973) );
  XOR2_X1 U2896 ( .A(n2941), .B(n2938), .Z(n2940) );
  AND2_X1 U2897 ( .A1(n2350), .A2(n2351), .ZN(n2939) );
  XNOR2_X1 U2898 ( .A(n2942), .B(n2943), .ZN(n2351) );
  XOR2_X1 U2899 ( .A(n2944), .B(n2945), .Z(n2943) );
  NAND2_X1 U2900 ( .A1(a_0_), .A2(b_9_), .ZN(n2945) );
  NAND2_X1 U2901 ( .A1(n2360), .A2(n2946), .ZN(n2350) );
  NAND2_X1 U2902 ( .A1(n2359), .A2(n2361), .ZN(n2946) );
  NAND2_X1 U2903 ( .A1(n2947), .A2(n2948), .ZN(n2361) );
  NAND2_X1 U2904 ( .A1(a_0_), .A2(b_10_), .ZN(n2948) );
  INV_X1 U2905 ( .A(n2949), .ZN(n2947) );
  XNOR2_X1 U2906 ( .A(n2950), .B(n2951), .ZN(n2359) );
  XOR2_X1 U2907 ( .A(n2952), .B(n2953), .Z(n2951) );
  NAND2_X1 U2908 ( .A1(b_9_), .A2(a_1_), .ZN(n2953) );
  NAND2_X1 U2909 ( .A1(a_0_), .A2(n2949), .ZN(n2360) );
  NAND2_X1 U2910 ( .A1(n2954), .A2(n2955), .ZN(n2949) );
  NAND2_X1 U2911 ( .A1(n2725), .A2(n2956), .ZN(n2955) );
  OR2_X1 U2912 ( .A1(n2722), .A2(n2724), .ZN(n2956) );
  NOR2_X1 U2913 ( .A1(n2278), .A2(n2381), .ZN(n2725) );
  NAND2_X1 U2914 ( .A1(n2722), .A2(n2724), .ZN(n2954) );
  NAND2_X1 U2915 ( .A1(n2957), .A2(n2958), .ZN(n2724) );
  NAND2_X1 U2916 ( .A1(n2959), .A2(a_2_), .ZN(n2958) );
  NOR2_X1 U2917 ( .A1(n2960), .A2(n2278), .ZN(n2959) );
  NOR2_X1 U2918 ( .A1(n2932), .A2(n2933), .ZN(n2960) );
  NAND2_X1 U2919 ( .A1(n2932), .A2(n2933), .ZN(n2957) );
  NAND2_X1 U2920 ( .A1(n2961), .A2(n2962), .ZN(n2933) );
  NAND2_X1 U2921 ( .A1(n2929), .A2(n2963), .ZN(n2962) );
  NAND2_X1 U2922 ( .A1(n2930), .A2(n2928), .ZN(n2963) );
  NOR2_X1 U2923 ( .A1(n2199), .A2(n2278), .ZN(n2929) );
  OR2_X1 U2924 ( .A1(n2928), .A2(n2930), .ZN(n2961) );
  AND2_X1 U2925 ( .A1(n2964), .A2(n2965), .ZN(n2930) );
  NAND2_X1 U2926 ( .A1(n2926), .A2(n2966), .ZN(n2965) );
  OR2_X1 U2927 ( .A1(n2923), .A2(n2925), .ZN(n2966) );
  NOR2_X1 U2928 ( .A1(n2285), .A2(n2278), .ZN(n2926) );
  NAND2_X1 U2929 ( .A1(n2923), .A2(n2925), .ZN(n2964) );
  NAND2_X1 U2930 ( .A1(n2967), .A2(n2968), .ZN(n2925) );
  NAND2_X1 U2931 ( .A1(n2969), .A2(a_5_), .ZN(n2968) );
  NOR2_X1 U2932 ( .A1(n2970), .A2(n2278), .ZN(n2969) );
  NOR2_X1 U2933 ( .A1(n2921), .A2(n2919), .ZN(n2970) );
  NAND2_X1 U2934 ( .A1(n2919), .A2(n2921), .ZN(n2967) );
  NAND2_X1 U2935 ( .A1(n2971), .A2(n2972), .ZN(n2921) );
  NAND2_X1 U2936 ( .A1(n2973), .A2(a_6_), .ZN(n2972) );
  NOR2_X1 U2937 ( .A1(n2974), .A2(n2278), .ZN(n2973) );
  NOR2_X1 U2938 ( .A1(n2917), .A2(n2916), .ZN(n2974) );
  NAND2_X1 U2939 ( .A1(n2916), .A2(n2917), .ZN(n2971) );
  NAND2_X1 U2940 ( .A1(n2975), .A2(n2976), .ZN(n2917) );
  NAND2_X1 U2941 ( .A1(n2914), .A2(n2977), .ZN(n2976) );
  OR2_X1 U2942 ( .A1(n2911), .A2(n2913), .ZN(n2977) );
  NOR2_X1 U2943 ( .A1(n2132), .A2(n2278), .ZN(n2914) );
  NAND2_X1 U2944 ( .A1(n2911), .A2(n2913), .ZN(n2975) );
  NAND2_X1 U2945 ( .A1(n2978), .A2(n2979), .ZN(n2913) );
  NAND2_X1 U2946 ( .A1(n2980), .A2(a_8_), .ZN(n2979) );
  NOR2_X1 U2947 ( .A1(n2981), .A2(n2278), .ZN(n2980) );
  NOR2_X1 U2948 ( .A1(n2908), .A2(n2909), .ZN(n2981) );
  NAND2_X1 U2949 ( .A1(n2908), .A2(n2909), .ZN(n2978) );
  NAND2_X1 U2950 ( .A1(n2982), .A2(n2983), .ZN(n2909) );
  NAND2_X1 U2951 ( .A1(n2906), .A2(n2984), .ZN(n2983) );
  OR2_X1 U2952 ( .A1(n2903), .A2(n2905), .ZN(n2984) );
  NOR2_X1 U2953 ( .A1(n2102), .A2(n2278), .ZN(n2906) );
  NAND2_X1 U2954 ( .A1(n2903), .A2(n2905), .ZN(n2982) );
  NAND2_X1 U2955 ( .A1(n2985), .A2(n2986), .ZN(n2905) );
  NAND2_X1 U2956 ( .A1(n2901), .A2(n2987), .ZN(n2986) );
  NAND2_X1 U2957 ( .A1(n2902), .A2(n2091), .ZN(n2987) );
  INV_X1 U2958 ( .A(n2988), .ZN(n2902) );
  XNOR2_X1 U2959 ( .A(n2989), .B(n2990), .ZN(n2901) );
  NAND2_X1 U2960 ( .A1(n2991), .A2(n2992), .ZN(n2989) );
  NAND2_X1 U2961 ( .A1(n2993), .A2(n2988), .ZN(n2985) );
  NAND2_X1 U2962 ( .A1(n2873), .A2(n2994), .ZN(n2988) );
  NAND2_X1 U2963 ( .A1(n2872), .A2(n2874), .ZN(n2994) );
  NAND2_X1 U2964 ( .A1(n2995), .A2(n2996), .ZN(n2874) );
  NAND2_X1 U2965 ( .A1(b_10_), .A2(a_11_), .ZN(n2996) );
  INV_X1 U2966 ( .A(n2997), .ZN(n2995) );
  XOR2_X1 U2967 ( .A(n2998), .B(n2999), .Z(n2872) );
  XNOR2_X1 U2968 ( .A(n3000), .B(n3001), .ZN(n2998) );
  NAND2_X1 U2969 ( .A1(b_9_), .A2(a_12_), .ZN(n3000) );
  NAND2_X1 U2970 ( .A1(a_11_), .A2(n2997), .ZN(n2873) );
  NAND2_X1 U2971 ( .A1(n3002), .A2(n3003), .ZN(n2997) );
  NAND2_X1 U2972 ( .A1(n3004), .A2(b_10_), .ZN(n3003) );
  NOR2_X1 U2973 ( .A1(n3005), .A2(n2277), .ZN(n3004) );
  NOR2_X1 U2974 ( .A1(n2879), .A2(n2881), .ZN(n3005) );
  NAND2_X1 U2975 ( .A1(n2879), .A2(n2881), .ZN(n3002) );
  NAND2_X1 U2976 ( .A1(n3006), .A2(n3007), .ZN(n2881) );
  NAND2_X1 U2977 ( .A1(n2897), .A2(n3008), .ZN(n3007) );
  OR2_X1 U2978 ( .A1(n2898), .A2(n2899), .ZN(n3008) );
  NOR2_X1 U2979 ( .A1(n2278), .A2(n2042), .ZN(n2897) );
  NAND2_X1 U2980 ( .A1(n2899), .A2(n2898), .ZN(n3006) );
  NAND2_X1 U2981 ( .A1(n3009), .A2(n3010), .ZN(n2898) );
  NAND2_X1 U2982 ( .A1(b_8_), .A2(n3011), .ZN(n3010) );
  NAND2_X1 U2983 ( .A1(n2018), .A2(n3012), .ZN(n3011) );
  NAND2_X1 U2984 ( .A1(a_15_), .A2(n2103), .ZN(n3012) );
  NAND2_X1 U2985 ( .A1(b_9_), .A2(n3013), .ZN(n3009) );
  NAND2_X1 U2986 ( .A1(n2021), .A2(n3014), .ZN(n3013) );
  NAND2_X1 U2987 ( .A1(a_14_), .A2(n2280), .ZN(n3014) );
  AND2_X1 U2988 ( .A1(n3015), .A2(n2558), .ZN(n2899) );
  NOR2_X1 U2989 ( .A1(n2278), .A2(n2103), .ZN(n3015) );
  XOR2_X1 U2990 ( .A(n3016), .B(n3017), .Z(n2879) );
  XOR2_X1 U2991 ( .A(n3018), .B(n3019), .Z(n3016) );
  INV_X1 U2992 ( .A(n2091), .ZN(n2993) );
  NAND2_X1 U2993 ( .A1(b_10_), .A2(a_10_), .ZN(n2091) );
  XNOR2_X1 U2994 ( .A(n3020), .B(n3021), .ZN(n2903) );
  NAND2_X1 U2995 ( .A1(n3022), .A2(n3023), .ZN(n3020) );
  XNOR2_X1 U2996 ( .A(n3024), .B(n3025), .ZN(n2908) );
  XOR2_X1 U2997 ( .A(n3026), .B(n2259), .Z(n3025) );
  XOR2_X1 U2998 ( .A(n3027), .B(n3028), .Z(n2911) );
  XOR2_X1 U2999 ( .A(n3029), .B(n3030), .Z(n3027) );
  NOR2_X1 U3000 ( .A1(n2103), .A2(n2281), .ZN(n3030) );
  XNOR2_X1 U3001 ( .A(n3031), .B(n3032), .ZN(n2916) );
  XNOR2_X1 U3002 ( .A(n3033), .B(n3034), .ZN(n3032) );
  XNOR2_X1 U3003 ( .A(n3035), .B(n3036), .ZN(n2919) );
  XNOR2_X1 U3004 ( .A(n3037), .B(n3038), .ZN(n3035) );
  XNOR2_X1 U3005 ( .A(n3039), .B(n3040), .ZN(n2923) );
  XOR2_X1 U3006 ( .A(n3041), .B(n3042), .Z(n3040) );
  NAND2_X1 U3007 ( .A1(a_5_), .A2(b_9_), .ZN(n3042) );
  XOR2_X1 U3008 ( .A(n3043), .B(n3044), .Z(n2928) );
  NAND2_X1 U3009 ( .A1(n3045), .A2(n3046), .ZN(n3043) );
  XNOR2_X1 U3010 ( .A(n3047), .B(n3048), .ZN(n2932) );
  XOR2_X1 U3011 ( .A(n3049), .B(n3050), .Z(n3048) );
  NAND2_X1 U3012 ( .A1(a_3_), .A2(b_9_), .ZN(n3050) );
  XNOR2_X1 U3013 ( .A(n3051), .B(n3052), .ZN(n2722) );
  XOR2_X1 U3014 ( .A(n3053), .B(n3054), .Z(n3052) );
  NAND2_X1 U3015 ( .A1(a_2_), .A2(b_9_), .ZN(n3054) );
  NAND2_X1 U3016 ( .A1(n3055), .A2(n3056), .ZN(n1979) );
  NAND2_X1 U3017 ( .A1(n2938), .A2(n2941), .ZN(n3056) );
  NAND2_X1 U3018 ( .A1(n3057), .A2(n2938), .ZN(n1978) );
  XOR2_X1 U3019 ( .A(n3058), .B(n3059), .Z(n2938) );
  XOR2_X1 U3020 ( .A(n3060), .B(n3061), .Z(n3058) );
  NOR2_X1 U3021 ( .A1(n2937), .A2(n3055), .ZN(n3057) );
  XOR2_X1 U3022 ( .A(n3062), .B(n3063), .Z(n3055) );
  INV_X1 U3023 ( .A(n3064), .ZN(n3063) );
  INV_X1 U3024 ( .A(n2941), .ZN(n2937) );
  NAND2_X1 U3025 ( .A1(n3065), .A2(n3066), .ZN(n2941) );
  NAND2_X1 U3026 ( .A1(n3067), .A2(a_0_), .ZN(n3066) );
  NOR2_X1 U3027 ( .A1(n3068), .A2(n2103), .ZN(n3067) );
  NOR2_X1 U3028 ( .A1(n2942), .A2(n2944), .ZN(n3068) );
  NAND2_X1 U3029 ( .A1(n2942), .A2(n2944), .ZN(n3065) );
  NAND2_X1 U3030 ( .A1(n3069), .A2(n3070), .ZN(n2944) );
  NAND2_X1 U3031 ( .A1(n3071), .A2(b_9_), .ZN(n3070) );
  NOR2_X1 U3032 ( .A1(n3072), .A2(n2381), .ZN(n3071) );
  NOR2_X1 U3033 ( .A1(n2952), .A2(n2950), .ZN(n3072) );
  NAND2_X1 U3034 ( .A1(n2950), .A2(n2952), .ZN(n3069) );
  NAND2_X1 U3035 ( .A1(n3073), .A2(n3074), .ZN(n2952) );
  NAND2_X1 U3036 ( .A1(n3075), .A2(a_2_), .ZN(n3074) );
  NOR2_X1 U3037 ( .A1(n3076), .A2(n2103), .ZN(n3075) );
  NOR2_X1 U3038 ( .A1(n3051), .A2(n3053), .ZN(n3076) );
  NAND2_X1 U3039 ( .A1(n3051), .A2(n3053), .ZN(n3073) );
  NAND2_X1 U3040 ( .A1(n3077), .A2(n3078), .ZN(n3053) );
  NAND2_X1 U3041 ( .A1(n3079), .A2(a_3_), .ZN(n3078) );
  NOR2_X1 U3042 ( .A1(n3080), .A2(n2103), .ZN(n3079) );
  NOR2_X1 U3043 ( .A1(n3049), .A2(n3047), .ZN(n3080) );
  NAND2_X1 U3044 ( .A1(n3047), .A2(n3049), .ZN(n3077) );
  NAND2_X1 U3045 ( .A1(n3045), .A2(n3081), .ZN(n3049) );
  NAND2_X1 U3046 ( .A1(n3044), .A2(n3046), .ZN(n3081) );
  NAND2_X1 U3047 ( .A1(n3082), .A2(n3083), .ZN(n3046) );
  NAND2_X1 U3048 ( .A1(a_4_), .A2(b_9_), .ZN(n3083) );
  INV_X1 U3049 ( .A(n3084), .ZN(n3082) );
  XNOR2_X1 U3050 ( .A(n3085), .B(n3086), .ZN(n3044) );
  XOR2_X1 U3051 ( .A(n3087), .B(n3088), .Z(n3086) );
  NAND2_X1 U3052 ( .A1(a_5_), .A2(b_8_), .ZN(n3088) );
  NAND2_X1 U3053 ( .A1(a_4_), .A2(n3084), .ZN(n3045) );
  NAND2_X1 U3054 ( .A1(n3089), .A2(n3090), .ZN(n3084) );
  NAND2_X1 U3055 ( .A1(n3091), .A2(a_5_), .ZN(n3090) );
  NOR2_X1 U3056 ( .A1(n3092), .A2(n2103), .ZN(n3091) );
  NOR2_X1 U3057 ( .A1(n3039), .A2(n3041), .ZN(n3092) );
  NAND2_X1 U3058 ( .A1(n3039), .A2(n3041), .ZN(n3089) );
  NAND2_X1 U3059 ( .A1(n3093), .A2(n3094), .ZN(n3041) );
  NAND2_X1 U3060 ( .A1(n3038), .A2(n3095), .ZN(n3094) );
  NAND2_X1 U3061 ( .A1(n3037), .A2(n3036), .ZN(n3095) );
  NOR2_X1 U3062 ( .A1(n2283), .A2(n2103), .ZN(n3038) );
  OR2_X1 U3063 ( .A1(n3036), .A2(n3037), .ZN(n3093) );
  AND2_X1 U3064 ( .A1(n3096), .A2(n3097), .ZN(n3037) );
  NAND2_X1 U3065 ( .A1(n3034), .A2(n3098), .ZN(n3097) );
  OR2_X1 U3066 ( .A1(n3033), .A2(n3031), .ZN(n3098) );
  NOR2_X1 U3067 ( .A1(n2132), .A2(n2103), .ZN(n3034) );
  NAND2_X1 U3068 ( .A1(n3031), .A2(n3033), .ZN(n3096) );
  NAND2_X1 U3069 ( .A1(n3099), .A2(n3100), .ZN(n3033) );
  NAND2_X1 U3070 ( .A1(n3101), .A2(a_8_), .ZN(n3100) );
  NOR2_X1 U3071 ( .A1(n3102), .A2(n2103), .ZN(n3101) );
  NOR2_X1 U3072 ( .A1(n3028), .A2(n3029), .ZN(n3102) );
  NAND2_X1 U3073 ( .A1(n3028), .A2(n3029), .ZN(n3099) );
  NAND2_X1 U3074 ( .A1(n3103), .A2(n3104), .ZN(n3029) );
  NAND2_X1 U3075 ( .A1(n2097), .A2(n3105), .ZN(n3104) );
  OR2_X1 U3076 ( .A1(n3024), .A2(n3026), .ZN(n3105) );
  INV_X1 U3077 ( .A(n2259), .ZN(n2097) );
  NAND2_X1 U3078 ( .A1(a_9_), .A2(b_9_), .ZN(n2259) );
  NAND2_X1 U3079 ( .A1(n3024), .A2(n3026), .ZN(n3103) );
  NAND2_X1 U3080 ( .A1(n3022), .A2(n3106), .ZN(n3026) );
  NAND2_X1 U3081 ( .A1(n3021), .A2(n3023), .ZN(n3106) );
  NAND2_X1 U3082 ( .A1(n3107), .A2(n3108), .ZN(n3023) );
  NAND2_X1 U3083 ( .A1(b_9_), .A2(a_10_), .ZN(n3108) );
  INV_X1 U3084 ( .A(n3109), .ZN(n3107) );
  XNOR2_X1 U3085 ( .A(n3110), .B(n3111), .ZN(n3021) );
  NAND2_X1 U3086 ( .A1(n3112), .A2(n3113), .ZN(n3110) );
  NAND2_X1 U3087 ( .A1(a_10_), .A2(n3109), .ZN(n3022) );
  NAND2_X1 U3088 ( .A1(n2991), .A2(n3114), .ZN(n3109) );
  NAND2_X1 U3089 ( .A1(n2990), .A2(n2992), .ZN(n3114) );
  NAND2_X1 U3090 ( .A1(n3115), .A2(n3116), .ZN(n2992) );
  NAND2_X1 U3091 ( .A1(b_9_), .A2(a_11_), .ZN(n3116) );
  INV_X1 U3092 ( .A(n3117), .ZN(n3115) );
  XOR2_X1 U3093 ( .A(n3118), .B(n3119), .Z(n2990) );
  XNOR2_X1 U3094 ( .A(n3120), .B(n3121), .ZN(n3118) );
  NAND2_X1 U3095 ( .A1(b_8_), .A2(a_12_), .ZN(n3120) );
  NAND2_X1 U3096 ( .A1(a_11_), .A2(n3117), .ZN(n2991) );
  NAND2_X1 U3097 ( .A1(n3122), .A2(n3123), .ZN(n3117) );
  NAND2_X1 U3098 ( .A1(n3124), .A2(b_9_), .ZN(n3123) );
  NOR2_X1 U3099 ( .A1(n3125), .A2(n2277), .ZN(n3124) );
  NOR2_X1 U3100 ( .A1(n2999), .A2(n3001), .ZN(n3125) );
  NAND2_X1 U3101 ( .A1(n2999), .A2(n3001), .ZN(n3122) );
  NAND2_X1 U3102 ( .A1(n3126), .A2(n3127), .ZN(n3001) );
  NAND2_X1 U3103 ( .A1(n3017), .A2(n3128), .ZN(n3127) );
  OR2_X1 U3104 ( .A1(n3018), .A2(n3019), .ZN(n3128) );
  NOR2_X1 U3105 ( .A1(n2103), .A2(n2042), .ZN(n3017) );
  NAND2_X1 U3106 ( .A1(n3019), .A2(n3018), .ZN(n3126) );
  NAND2_X1 U3107 ( .A1(n3129), .A2(n3130), .ZN(n3018) );
  NAND2_X1 U3108 ( .A1(b_7_), .A2(n3131), .ZN(n3130) );
  NAND2_X1 U3109 ( .A1(n2018), .A2(n3132), .ZN(n3131) );
  NAND2_X1 U3110 ( .A1(a_15_), .A2(n2280), .ZN(n3132) );
  NAND2_X1 U3111 ( .A1(b_8_), .A2(n3133), .ZN(n3129) );
  NAND2_X1 U3112 ( .A1(n2021), .A2(n3134), .ZN(n3133) );
  NAND2_X1 U3113 ( .A1(a_14_), .A2(n2133), .ZN(n3134) );
  AND2_X1 U3114 ( .A1(n3135), .A2(n2558), .ZN(n3019) );
  NOR2_X1 U3115 ( .A1(n2103), .A2(n2280), .ZN(n3135) );
  INV_X1 U3116 ( .A(b_9_), .ZN(n2103) );
  XNOR2_X1 U3117 ( .A(n3136), .B(n3137), .ZN(n2999) );
  XNOR2_X1 U3118 ( .A(n3138), .B(n3139), .ZN(n3137) );
  XNOR2_X1 U3119 ( .A(n3140), .B(n3141), .ZN(n3024) );
  NAND2_X1 U3120 ( .A1(n3142), .A2(n3143), .ZN(n3140) );
  XNOR2_X1 U3121 ( .A(n3144), .B(n3145), .ZN(n3028) );
  XNOR2_X1 U3122 ( .A(n3146), .B(n3147), .ZN(n3145) );
  XOR2_X1 U3123 ( .A(n3148), .B(n3149), .Z(n3031) );
  XOR2_X1 U3124 ( .A(n3150), .B(n3151), .Z(n3148) );
  XNOR2_X1 U3125 ( .A(n3152), .B(n3153), .ZN(n3036) );
  XOR2_X1 U3126 ( .A(n3154), .B(n3155), .Z(n3152) );
  NOR2_X1 U3127 ( .A1(n2280), .A2(n2132), .ZN(n3155) );
  XNOR2_X1 U3128 ( .A(n3156), .B(n3157), .ZN(n3039) );
  XOR2_X1 U3129 ( .A(n3158), .B(n3159), .Z(n3157) );
  NAND2_X1 U3130 ( .A1(a_6_), .A2(b_8_), .ZN(n3159) );
  XNOR2_X1 U3131 ( .A(n3160), .B(n3161), .ZN(n3047) );
  XOR2_X1 U3132 ( .A(n3162), .B(n3163), .Z(n3161) );
  NAND2_X1 U3133 ( .A1(a_4_), .A2(b_8_), .ZN(n3163) );
  XNOR2_X1 U3134 ( .A(n3164), .B(n3165), .ZN(n3051) );
  XNOR2_X1 U3135 ( .A(n3166), .B(n3167), .ZN(n3165) );
  XOR2_X1 U3136 ( .A(n3168), .B(n3169), .Z(n2950) );
  XOR2_X1 U3137 ( .A(n3170), .B(n3171), .Z(n3168) );
  XOR2_X1 U3138 ( .A(n3172), .B(n3173), .Z(n2942) );
  XOR2_X1 U3139 ( .A(n3174), .B(n3175), .Z(n3172) );
  NAND2_X1 U3140 ( .A1(n3176), .A2(n3177), .ZN(n1984) );
  NAND2_X1 U3141 ( .A1(n3064), .A2(n3062), .ZN(n3177) );
  NAND2_X1 U3142 ( .A1(n3178), .A2(n3064), .ZN(n1983) );
  XNOR2_X1 U3143 ( .A(n3179), .B(n3180), .ZN(n3064) );
  XOR2_X1 U3144 ( .A(n3181), .B(n3182), .Z(n3180) );
  NAND2_X1 U3145 ( .A1(a_0_), .A2(b_7_), .ZN(n3182) );
  NOR2_X1 U3146 ( .A1(n3183), .A2(n3176), .ZN(n3178) );
  XOR2_X1 U3147 ( .A(n3184), .B(n3185), .Z(n3176) );
  INV_X1 U3148 ( .A(n3186), .ZN(n3185) );
  INV_X1 U3149 ( .A(n3062), .ZN(n3183) );
  NAND2_X1 U3150 ( .A1(n3187), .A2(n3188), .ZN(n3062) );
  NAND2_X1 U3151 ( .A1(n3061), .A2(n3189), .ZN(n3188) );
  OR2_X1 U3152 ( .A1(n3059), .A2(n3060), .ZN(n3189) );
  NOR2_X1 U3153 ( .A1(n2376), .A2(n2280), .ZN(n3061) );
  NAND2_X1 U3154 ( .A1(n3059), .A2(n3060), .ZN(n3187) );
  NAND2_X1 U3155 ( .A1(n3190), .A2(n3191), .ZN(n3060) );
  NAND2_X1 U3156 ( .A1(n3175), .A2(n3192), .ZN(n3191) );
  OR2_X1 U3157 ( .A1(n3173), .A2(n3174), .ZN(n3192) );
  NOR2_X1 U3158 ( .A1(n2280), .A2(n2381), .ZN(n3175) );
  NAND2_X1 U3159 ( .A1(n3173), .A2(n3174), .ZN(n3190) );
  NAND2_X1 U3160 ( .A1(n3193), .A2(n3194), .ZN(n3174) );
  NAND2_X1 U3161 ( .A1(n3170), .A2(n3195), .ZN(n3194) );
  OR2_X1 U3162 ( .A1(n3171), .A2(n3169), .ZN(n3195) );
  NOR2_X1 U3163 ( .A1(n2287), .A2(n2280), .ZN(n3170) );
  NAND2_X1 U3164 ( .A1(n3169), .A2(n3171), .ZN(n3193) );
  NAND2_X1 U3165 ( .A1(n3196), .A2(n3197), .ZN(n3171) );
  NAND2_X1 U3166 ( .A1(n3167), .A2(n3198), .ZN(n3197) );
  OR2_X1 U3167 ( .A1(n3164), .A2(n3166), .ZN(n3198) );
  NOR2_X1 U3168 ( .A1(n2199), .A2(n2280), .ZN(n3167) );
  NAND2_X1 U3169 ( .A1(n3164), .A2(n3166), .ZN(n3196) );
  NAND2_X1 U3170 ( .A1(n3199), .A2(n3200), .ZN(n3166) );
  NAND2_X1 U3171 ( .A1(n3201), .A2(a_4_), .ZN(n3200) );
  NOR2_X1 U3172 ( .A1(n3202), .A2(n2280), .ZN(n3201) );
  NOR2_X1 U3173 ( .A1(n3160), .A2(n3162), .ZN(n3202) );
  NAND2_X1 U3174 ( .A1(n3160), .A2(n3162), .ZN(n3199) );
  NAND2_X1 U3175 ( .A1(n3203), .A2(n3204), .ZN(n3162) );
  NAND2_X1 U3176 ( .A1(n3205), .A2(a_5_), .ZN(n3204) );
  NOR2_X1 U3177 ( .A1(n3206), .A2(n2280), .ZN(n3205) );
  NOR2_X1 U3178 ( .A1(n3087), .A2(n3085), .ZN(n3206) );
  NAND2_X1 U3179 ( .A1(n3085), .A2(n3087), .ZN(n3203) );
  NAND2_X1 U3180 ( .A1(n3207), .A2(n3208), .ZN(n3087) );
  NAND2_X1 U3181 ( .A1(n3209), .A2(a_6_), .ZN(n3208) );
  NOR2_X1 U3182 ( .A1(n3210), .A2(n2280), .ZN(n3209) );
  NOR2_X1 U3183 ( .A1(n3158), .A2(n3156), .ZN(n3210) );
  NAND2_X1 U3184 ( .A1(n3156), .A2(n3158), .ZN(n3207) );
  NAND2_X1 U3185 ( .A1(n3211), .A2(n3212), .ZN(n3158) );
  NAND2_X1 U3186 ( .A1(n3213), .A2(a_7_), .ZN(n3212) );
  NOR2_X1 U3187 ( .A1(n3214), .A2(n2280), .ZN(n3213) );
  NOR2_X1 U3188 ( .A1(n3154), .A2(n3153), .ZN(n3214) );
  NAND2_X1 U3189 ( .A1(n3153), .A2(n3154), .ZN(n3211) );
  NAND2_X1 U3190 ( .A1(n3215), .A2(n3216), .ZN(n3154) );
  NAND2_X1 U3191 ( .A1(n3149), .A2(n3217), .ZN(n3216) );
  OR2_X1 U3192 ( .A1(n3150), .A2(n3151), .ZN(n3217) );
  XNOR2_X1 U3193 ( .A(n3218), .B(n3219), .ZN(n3149) );
  XNOR2_X1 U3194 ( .A(n3220), .B(n3221), .ZN(n3219) );
  NAND2_X1 U3195 ( .A1(n3151), .A2(n3150), .ZN(n3215) );
  NAND2_X1 U3196 ( .A1(n3222), .A2(n3223), .ZN(n3150) );
  NAND2_X1 U3197 ( .A1(n3147), .A2(n3224), .ZN(n3223) );
  OR2_X1 U3198 ( .A1(n3144), .A2(n3146), .ZN(n3224) );
  NOR2_X1 U3199 ( .A1(n2280), .A2(n2102), .ZN(n3147) );
  NAND2_X1 U3200 ( .A1(n3144), .A2(n3146), .ZN(n3222) );
  NAND2_X1 U3201 ( .A1(n3142), .A2(n3225), .ZN(n3146) );
  NAND2_X1 U3202 ( .A1(n3141), .A2(n3143), .ZN(n3225) );
  NAND2_X1 U3203 ( .A1(n3226), .A2(n3227), .ZN(n3143) );
  NAND2_X1 U3204 ( .A1(b_8_), .A2(a_10_), .ZN(n3227) );
  INV_X1 U3205 ( .A(n3228), .ZN(n3226) );
  XNOR2_X1 U3206 ( .A(n3229), .B(n3230), .ZN(n3141) );
  NAND2_X1 U3207 ( .A1(n3231), .A2(n3232), .ZN(n3229) );
  NAND2_X1 U3208 ( .A1(a_10_), .A2(n3228), .ZN(n3142) );
  NAND2_X1 U3209 ( .A1(n3112), .A2(n3233), .ZN(n3228) );
  NAND2_X1 U3210 ( .A1(n3111), .A2(n3113), .ZN(n3233) );
  NAND2_X1 U3211 ( .A1(n3234), .A2(n3235), .ZN(n3113) );
  NAND2_X1 U3212 ( .A1(b_8_), .A2(a_11_), .ZN(n3235) );
  INV_X1 U3213 ( .A(n3236), .ZN(n3234) );
  XOR2_X1 U3214 ( .A(n3237), .B(n3238), .Z(n3111) );
  XNOR2_X1 U3215 ( .A(n3239), .B(n3240), .ZN(n3237) );
  NAND2_X1 U3216 ( .A1(b_7_), .A2(a_12_), .ZN(n3239) );
  NAND2_X1 U3217 ( .A1(a_11_), .A2(n3236), .ZN(n3112) );
  NAND2_X1 U3218 ( .A1(n3241), .A2(n3242), .ZN(n3236) );
  NAND2_X1 U3219 ( .A1(n3243), .A2(b_8_), .ZN(n3242) );
  NOR2_X1 U3220 ( .A1(n3244), .A2(n2277), .ZN(n3243) );
  NOR2_X1 U3221 ( .A1(n3119), .A2(n3121), .ZN(n3244) );
  NAND2_X1 U3222 ( .A1(n3119), .A2(n3121), .ZN(n3241) );
  NAND2_X1 U3223 ( .A1(n3245), .A2(n3246), .ZN(n3121) );
  NAND2_X1 U3224 ( .A1(n3136), .A2(n3247), .ZN(n3246) );
  NAND2_X1 U3225 ( .A1(n3139), .A2(n3138), .ZN(n3247) );
  NOR2_X1 U3226 ( .A1(n2280), .A2(n2042), .ZN(n3136) );
  OR2_X1 U3227 ( .A1(n3138), .A2(n3139), .ZN(n3245) );
  AND2_X1 U3228 ( .A1(n3248), .A2(n3249), .ZN(n3139) );
  NAND2_X1 U3229 ( .A1(b_6_), .A2(n3250), .ZN(n3249) );
  NAND2_X1 U3230 ( .A1(n2018), .A2(n3251), .ZN(n3250) );
  NAND2_X1 U3231 ( .A1(a_15_), .A2(n2133), .ZN(n3251) );
  NAND2_X1 U3232 ( .A1(b_7_), .A2(n3252), .ZN(n3248) );
  NAND2_X1 U3233 ( .A1(n2021), .A2(n3253), .ZN(n3252) );
  NAND2_X1 U3234 ( .A1(a_14_), .A2(n2282), .ZN(n3253) );
  NAND2_X1 U3235 ( .A1(n3254), .A2(n2558), .ZN(n3138) );
  NOR2_X1 U3236 ( .A1(n2133), .A2(n2280), .ZN(n3254) );
  XOR2_X1 U3237 ( .A(n3255), .B(n3256), .Z(n3119) );
  XOR2_X1 U3238 ( .A(n3257), .B(n3258), .Z(n3255) );
  XNOR2_X1 U3239 ( .A(n3259), .B(n3260), .ZN(n3144) );
  NAND2_X1 U3240 ( .A1(n3261), .A2(n3262), .ZN(n3259) );
  INV_X1 U3241 ( .A(n2121), .ZN(n3151) );
  NAND2_X1 U3242 ( .A1(b_8_), .A2(a_8_), .ZN(n2121) );
  XNOR2_X1 U3243 ( .A(n3263), .B(n3264), .ZN(n3153) );
  XOR2_X1 U3244 ( .A(n3265), .B(n3266), .Z(n3264) );
  NAND2_X1 U3245 ( .A1(b_7_), .A2(a_8_), .ZN(n3266) );
  XNOR2_X1 U3246 ( .A(n3267), .B(n3268), .ZN(n3156) );
  XOR2_X1 U3247 ( .A(n2255), .B(n3269), .Z(n3268) );
  XOR2_X1 U3248 ( .A(n3270), .B(n3271), .Z(n3085) );
  XOR2_X1 U3249 ( .A(n3272), .B(n3273), .Z(n3270) );
  NOR2_X1 U3250 ( .A1(n2133), .A2(n2283), .ZN(n3273) );
  XNOR2_X1 U3251 ( .A(n3274), .B(n3275), .ZN(n3160) );
  XOR2_X1 U3252 ( .A(n3276), .B(n3277), .Z(n3275) );
  NAND2_X1 U3253 ( .A1(a_5_), .A2(b_7_), .ZN(n3277) );
  XNOR2_X1 U3254 ( .A(n3278), .B(n3279), .ZN(n3164) );
  XOR2_X1 U3255 ( .A(n3280), .B(n3281), .Z(n3279) );
  NAND2_X1 U3256 ( .A1(a_4_), .A2(b_7_), .ZN(n3281) );
  XNOR2_X1 U3257 ( .A(n3282), .B(n3283), .ZN(n3169) );
  XOR2_X1 U3258 ( .A(n3284), .B(n3285), .Z(n3283) );
  NAND2_X1 U3259 ( .A1(a_3_), .A2(b_7_), .ZN(n3285) );
  XNOR2_X1 U3260 ( .A(n3286), .B(n3287), .ZN(n3173) );
  XOR2_X1 U3261 ( .A(n3288), .B(n3289), .Z(n3287) );
  NAND2_X1 U3262 ( .A1(a_2_), .A2(b_7_), .ZN(n3289) );
  XNOR2_X1 U3263 ( .A(n3290), .B(n3291), .ZN(n3059) );
  XOR2_X1 U3264 ( .A(n3292), .B(n3293), .Z(n3291) );
  NAND2_X1 U3265 ( .A1(b_7_), .A2(a_1_), .ZN(n3293) );
  NAND2_X1 U3266 ( .A1(n3294), .A2(n3295), .ZN(n1989) );
  NAND2_X1 U3267 ( .A1(n3186), .A2(n3184), .ZN(n3295) );
  NAND2_X1 U3268 ( .A1(n3296), .A2(n3186), .ZN(n1988) );
  XNOR2_X1 U3269 ( .A(n3297), .B(n3298), .ZN(n3186) );
  XNOR2_X1 U3270 ( .A(n3299), .B(n3300), .ZN(n3298) );
  NOR2_X1 U3271 ( .A1(n3301), .A2(n3294), .ZN(n3296) );
  XNOR2_X1 U3272 ( .A(n3302), .B(n3303), .ZN(n3294) );
  INV_X1 U3273 ( .A(n3184), .ZN(n3301) );
  NAND2_X1 U3274 ( .A1(n3304), .A2(n3305), .ZN(n3184) );
  NAND2_X1 U3275 ( .A1(n3306), .A2(a_0_), .ZN(n3305) );
  NOR2_X1 U3276 ( .A1(n3307), .A2(n2133), .ZN(n3306) );
  NOR2_X1 U3277 ( .A1(n3181), .A2(n3179), .ZN(n3307) );
  NAND2_X1 U3278 ( .A1(n3179), .A2(n3181), .ZN(n3304) );
  NAND2_X1 U3279 ( .A1(n3308), .A2(n3309), .ZN(n3181) );
  NAND2_X1 U3280 ( .A1(n3310), .A2(b_7_), .ZN(n3309) );
  NOR2_X1 U3281 ( .A1(n3311), .A2(n2381), .ZN(n3310) );
  NOR2_X1 U3282 ( .A1(n3290), .A2(n3292), .ZN(n3311) );
  NAND2_X1 U3283 ( .A1(n3290), .A2(n3292), .ZN(n3308) );
  NAND2_X1 U3284 ( .A1(n3312), .A2(n3313), .ZN(n3292) );
  NAND2_X1 U3285 ( .A1(n3314), .A2(a_2_), .ZN(n3313) );
  NOR2_X1 U3286 ( .A1(n3315), .A2(n2133), .ZN(n3314) );
  NOR2_X1 U3287 ( .A1(n3286), .A2(n3288), .ZN(n3315) );
  NAND2_X1 U3288 ( .A1(n3286), .A2(n3288), .ZN(n3312) );
  NAND2_X1 U3289 ( .A1(n3316), .A2(n3317), .ZN(n3288) );
  NAND2_X1 U3290 ( .A1(n3318), .A2(a_3_), .ZN(n3317) );
  NOR2_X1 U3291 ( .A1(n3319), .A2(n2133), .ZN(n3318) );
  NOR2_X1 U3292 ( .A1(n3284), .A2(n3282), .ZN(n3319) );
  NAND2_X1 U3293 ( .A1(n3282), .A2(n3284), .ZN(n3316) );
  NAND2_X1 U3294 ( .A1(n3320), .A2(n3321), .ZN(n3284) );
  NAND2_X1 U3295 ( .A1(n3322), .A2(a_4_), .ZN(n3321) );
  NOR2_X1 U3296 ( .A1(n3323), .A2(n2133), .ZN(n3322) );
  NOR2_X1 U3297 ( .A1(n3278), .A2(n3280), .ZN(n3323) );
  NAND2_X1 U3298 ( .A1(n3278), .A2(n3280), .ZN(n3320) );
  NAND2_X1 U3299 ( .A1(n3324), .A2(n3325), .ZN(n3280) );
  NAND2_X1 U3300 ( .A1(n3326), .A2(a_5_), .ZN(n3325) );
  NOR2_X1 U3301 ( .A1(n3327), .A2(n2133), .ZN(n3326) );
  NOR2_X1 U3302 ( .A1(n3276), .A2(n3274), .ZN(n3327) );
  NAND2_X1 U3303 ( .A1(n3274), .A2(n3276), .ZN(n3324) );
  NAND2_X1 U3304 ( .A1(n3328), .A2(n3329), .ZN(n3276) );
  NAND2_X1 U3305 ( .A1(n3330), .A2(a_6_), .ZN(n3329) );
  NOR2_X1 U3306 ( .A1(n3331), .A2(n2133), .ZN(n3330) );
  NOR2_X1 U3307 ( .A1(n3271), .A2(n3272), .ZN(n3331) );
  NAND2_X1 U3308 ( .A1(n3271), .A2(n3272), .ZN(n3328) );
  NAND2_X1 U3309 ( .A1(n3332), .A2(n3333), .ZN(n3272) );
  NAND2_X1 U3310 ( .A1(n3267), .A2(n3334), .ZN(n3333) );
  OR2_X1 U3311 ( .A1(n3269), .A2(n2127), .ZN(n3334) );
  XOR2_X1 U3312 ( .A(n3335), .B(n3336), .Z(n3267) );
  XOR2_X1 U3313 ( .A(n3337), .B(n3338), .Z(n3335) );
  NAND2_X1 U3314 ( .A1(n2127), .A2(n3269), .ZN(n3332) );
  NAND2_X1 U3315 ( .A1(n3339), .A2(n3340), .ZN(n3269) );
  NAND2_X1 U3316 ( .A1(n3341), .A2(b_7_), .ZN(n3340) );
  NOR2_X1 U3317 ( .A1(n3342), .A2(n2281), .ZN(n3341) );
  NOR2_X1 U3318 ( .A1(n3263), .A2(n3265), .ZN(n3342) );
  NAND2_X1 U3319 ( .A1(n3263), .A2(n3265), .ZN(n3339) );
  NAND2_X1 U3320 ( .A1(n3343), .A2(n3344), .ZN(n3265) );
  NAND2_X1 U3321 ( .A1(n3221), .A2(n3345), .ZN(n3344) );
  OR2_X1 U3322 ( .A1(n3220), .A2(n3218), .ZN(n3345) );
  NOR2_X1 U3323 ( .A1(n2133), .A2(n2102), .ZN(n3221) );
  NAND2_X1 U3324 ( .A1(n3218), .A2(n3220), .ZN(n3343) );
  NAND2_X1 U3325 ( .A1(n3261), .A2(n3346), .ZN(n3220) );
  NAND2_X1 U3326 ( .A1(n3260), .A2(n3262), .ZN(n3346) );
  NAND2_X1 U3327 ( .A1(n3347), .A2(n3348), .ZN(n3262) );
  NAND2_X1 U3328 ( .A1(b_7_), .A2(a_10_), .ZN(n3348) );
  INV_X1 U3329 ( .A(n3349), .ZN(n3347) );
  XNOR2_X1 U3330 ( .A(n3350), .B(n3351), .ZN(n3260) );
  NAND2_X1 U3331 ( .A1(n3352), .A2(n3353), .ZN(n3350) );
  NAND2_X1 U3332 ( .A1(a_10_), .A2(n3349), .ZN(n3261) );
  NAND2_X1 U3333 ( .A1(n3231), .A2(n3354), .ZN(n3349) );
  NAND2_X1 U3334 ( .A1(n3230), .A2(n3232), .ZN(n3354) );
  NAND2_X1 U3335 ( .A1(n3355), .A2(n3356), .ZN(n3232) );
  NAND2_X1 U3336 ( .A1(b_7_), .A2(a_11_), .ZN(n3356) );
  INV_X1 U3337 ( .A(n3357), .ZN(n3355) );
  XOR2_X1 U3338 ( .A(n3358), .B(n3359), .Z(n3230) );
  XNOR2_X1 U3339 ( .A(n3360), .B(n3361), .ZN(n3358) );
  NAND2_X1 U3340 ( .A1(b_6_), .A2(a_12_), .ZN(n3360) );
  NAND2_X1 U3341 ( .A1(a_11_), .A2(n3357), .ZN(n3231) );
  NAND2_X1 U3342 ( .A1(n3362), .A2(n3363), .ZN(n3357) );
  NAND2_X1 U3343 ( .A1(n3364), .A2(b_7_), .ZN(n3363) );
  NOR2_X1 U3344 ( .A1(n3365), .A2(n2277), .ZN(n3364) );
  NOR2_X1 U3345 ( .A1(n3238), .A2(n3240), .ZN(n3365) );
  NAND2_X1 U3346 ( .A1(n3238), .A2(n3240), .ZN(n3362) );
  NAND2_X1 U3347 ( .A1(n3366), .A2(n3367), .ZN(n3240) );
  NAND2_X1 U3348 ( .A1(n3256), .A2(n3368), .ZN(n3367) );
  OR2_X1 U3349 ( .A1(n3257), .A2(n3258), .ZN(n3368) );
  NOR2_X1 U3350 ( .A1(n2133), .A2(n2042), .ZN(n3256) );
  NAND2_X1 U3351 ( .A1(n3258), .A2(n3257), .ZN(n3366) );
  NAND2_X1 U3352 ( .A1(n3369), .A2(n3370), .ZN(n3257) );
  NAND2_X1 U3353 ( .A1(b_5_), .A2(n3371), .ZN(n3370) );
  NAND2_X1 U3354 ( .A1(n2018), .A2(n3372), .ZN(n3371) );
  NAND2_X1 U3355 ( .A1(a_15_), .A2(n2282), .ZN(n3372) );
  NAND2_X1 U3356 ( .A1(b_6_), .A2(n3373), .ZN(n3369) );
  NAND2_X1 U3357 ( .A1(n2021), .A2(n3374), .ZN(n3373) );
  NAND2_X1 U3358 ( .A1(a_14_), .A2(n2163), .ZN(n3374) );
  AND2_X1 U3359 ( .A1(n3375), .A2(n2558), .ZN(n3258) );
  NOR2_X1 U3360 ( .A1(n2133), .A2(n2282), .ZN(n3375) );
  XOR2_X1 U3361 ( .A(n3376), .B(n3377), .Z(n3238) );
  XOR2_X1 U3362 ( .A(n3378), .B(n3379), .Z(n3376) );
  XNOR2_X1 U3363 ( .A(n3380), .B(n3381), .ZN(n3218) );
  NAND2_X1 U3364 ( .A1(n3382), .A2(n3383), .ZN(n3380) );
  XNOR2_X1 U3365 ( .A(n3384), .B(n3385), .ZN(n3263) );
  NAND2_X1 U3366 ( .A1(n3386), .A2(n3387), .ZN(n3384) );
  INV_X1 U3367 ( .A(n2255), .ZN(n2127) );
  NAND2_X1 U3368 ( .A1(a_7_), .A2(b_7_), .ZN(n2255) );
  XNOR2_X1 U3369 ( .A(n3388), .B(n3389), .ZN(n3271) );
  NAND2_X1 U3370 ( .A1(n3390), .A2(n3391), .ZN(n3388) );
  XOR2_X1 U3371 ( .A(n3392), .B(n3393), .Z(n3274) );
  XOR2_X1 U3372 ( .A(n3394), .B(n2151), .Z(n3393) );
  XNOR2_X1 U3373 ( .A(n3395), .B(n3396), .ZN(n3278) );
  NAND2_X1 U3374 ( .A1(n3397), .A2(n3398), .ZN(n3395) );
  XOR2_X1 U3375 ( .A(n3399), .B(n3400), .Z(n3282) );
  XOR2_X1 U3376 ( .A(n3401), .B(n3402), .Z(n3400) );
  XNOR2_X1 U3377 ( .A(n3403), .B(n3404), .ZN(n3286) );
  NAND2_X1 U3378 ( .A1(n3405), .A2(n3406), .ZN(n3403) );
  XOR2_X1 U3379 ( .A(n3407), .B(n3408), .Z(n3290) );
  XOR2_X1 U3380 ( .A(n3409), .B(n3410), .Z(n3407) );
  NOR2_X1 U3381 ( .A1(n2282), .A2(n2287), .ZN(n3410) );
  XNOR2_X1 U3382 ( .A(n3411), .B(n3412), .ZN(n3179) );
  XOR2_X1 U3383 ( .A(n3413), .B(n3414), .Z(n3412) );
  NAND2_X1 U3384 ( .A1(b_6_), .A2(a_1_), .ZN(n3414) );
  NAND2_X1 U3385 ( .A1(n3415), .A2(n3416), .ZN(n1994) );
  OR2_X1 U3386 ( .A1(n3303), .A2(n3302), .ZN(n3416) );
  XOR2_X1 U3387 ( .A(n3417), .B(n3418), .Z(n3415) );
  NAND2_X1 U3388 ( .A1(n3419), .A2(n3420), .ZN(n1993) );
  XOR2_X1 U3389 ( .A(n3417), .B(n3421), .Z(n3420) );
  NOR2_X1 U3390 ( .A1(n3302), .A2(n3303), .ZN(n3419) );
  XOR2_X1 U3391 ( .A(n3422), .B(n3423), .Z(n3303) );
  XOR2_X1 U3392 ( .A(n3424), .B(n3425), .Z(n3423) );
  NAND2_X1 U3393 ( .A1(a_0_), .A2(b_5_), .ZN(n3425) );
  AND2_X1 U3394 ( .A1(n3426), .A2(n3427), .ZN(n3302) );
  NAND2_X1 U3395 ( .A1(n3300), .A2(n3428), .ZN(n3427) );
  OR2_X1 U3396 ( .A1(n3297), .A2(n3299), .ZN(n3428) );
  NOR2_X1 U3397 ( .A1(n2376), .A2(n2282), .ZN(n3300) );
  NAND2_X1 U3398 ( .A1(n3297), .A2(n3299), .ZN(n3426) );
  NAND2_X1 U3399 ( .A1(n3429), .A2(n3430), .ZN(n3299) );
  NAND2_X1 U3400 ( .A1(n3431), .A2(b_6_), .ZN(n3430) );
  NOR2_X1 U3401 ( .A1(n3432), .A2(n2381), .ZN(n3431) );
  NOR2_X1 U3402 ( .A1(n3411), .A2(n3413), .ZN(n3432) );
  NAND2_X1 U3403 ( .A1(n3411), .A2(n3413), .ZN(n3429) );
  NAND2_X1 U3404 ( .A1(n3433), .A2(n3434), .ZN(n3413) );
  NAND2_X1 U3405 ( .A1(n3435), .A2(a_2_), .ZN(n3434) );
  NOR2_X1 U3406 ( .A1(n3436), .A2(n2282), .ZN(n3435) );
  NOR2_X1 U3407 ( .A1(n3409), .A2(n3408), .ZN(n3436) );
  NAND2_X1 U3408 ( .A1(n3408), .A2(n3409), .ZN(n3433) );
  NAND2_X1 U3409 ( .A1(n3405), .A2(n3437), .ZN(n3409) );
  NAND2_X1 U3410 ( .A1(n3404), .A2(n3406), .ZN(n3437) );
  NAND2_X1 U3411 ( .A1(n3438), .A2(n3439), .ZN(n3406) );
  NAND2_X1 U3412 ( .A1(a_3_), .A2(b_6_), .ZN(n3439) );
  INV_X1 U3413 ( .A(n3440), .ZN(n3438) );
  XOR2_X1 U3414 ( .A(n3441), .B(n3442), .Z(n3404) );
  XNOR2_X1 U3415 ( .A(n3443), .B(n3444), .ZN(n3441) );
  NAND2_X1 U3416 ( .A1(a_4_), .A2(b_5_), .ZN(n3443) );
  NAND2_X1 U3417 ( .A1(a_3_), .A2(n3440), .ZN(n3405) );
  NAND2_X1 U3418 ( .A1(n3445), .A2(n3446), .ZN(n3440) );
  NAND2_X1 U3419 ( .A1(n3402), .A2(n3447), .ZN(n3446) );
  NAND2_X1 U3420 ( .A1(n3401), .A2(n3399), .ZN(n3447) );
  NOR2_X1 U3421 ( .A1(n2285), .A2(n2282), .ZN(n3402) );
  OR2_X1 U3422 ( .A1(n3399), .A2(n3401), .ZN(n3445) );
  AND2_X1 U3423 ( .A1(n3397), .A2(n3448), .ZN(n3401) );
  NAND2_X1 U3424 ( .A1(n3396), .A2(n3398), .ZN(n3448) );
  NAND2_X1 U3425 ( .A1(n3449), .A2(n3450), .ZN(n3398) );
  NAND2_X1 U3426 ( .A1(a_5_), .A2(b_6_), .ZN(n3450) );
  XNOR2_X1 U3427 ( .A(n3451), .B(n3452), .ZN(n3396) );
  XOR2_X1 U3428 ( .A(n3453), .B(n3454), .Z(n3452) );
  NAND2_X1 U3429 ( .A1(b_5_), .A2(a_6_), .ZN(n3454) );
  OR2_X1 U3430 ( .A1(n3449), .A2(n2162), .ZN(n3397) );
  NAND2_X1 U3431 ( .A1(n3455), .A2(n3456), .ZN(n3449) );
  NAND2_X1 U3432 ( .A1(n3392), .A2(n3457), .ZN(n3456) );
  NAND2_X1 U3433 ( .A1(n3458), .A2(n3394), .ZN(n3457) );
  XOR2_X1 U3434 ( .A(n3459), .B(n3460), .Z(n3392) );
  XOR2_X1 U3435 ( .A(n3461), .B(n3462), .Z(n3460) );
  NAND2_X1 U3436 ( .A1(b_5_), .A2(a_7_), .ZN(n3462) );
  OR2_X1 U3437 ( .A1(n3394), .A2(n3458), .ZN(n3455) );
  INV_X1 U3438 ( .A(n2151), .ZN(n3458) );
  NAND2_X1 U3439 ( .A1(b_6_), .A2(a_6_), .ZN(n2151) );
  NAND2_X1 U3440 ( .A1(n3390), .A2(n3463), .ZN(n3394) );
  NAND2_X1 U3441 ( .A1(n3389), .A2(n3391), .ZN(n3463) );
  NAND2_X1 U3442 ( .A1(n3464), .A2(n3465), .ZN(n3391) );
  NAND2_X1 U3443 ( .A1(b_6_), .A2(a_7_), .ZN(n3465) );
  INV_X1 U3444 ( .A(n3466), .ZN(n3464) );
  XOR2_X1 U3445 ( .A(n3467), .B(n3468), .Z(n3389) );
  XOR2_X1 U3446 ( .A(n3469), .B(n3470), .Z(n3467) );
  NOR2_X1 U3447 ( .A1(n2281), .A2(n2163), .ZN(n3470) );
  NAND2_X1 U3448 ( .A1(a_7_), .A2(n3466), .ZN(n3390) );
  NAND2_X1 U3449 ( .A1(n3471), .A2(n3472), .ZN(n3466) );
  NAND2_X1 U3450 ( .A1(n3338), .A2(n3473), .ZN(n3472) );
  OR2_X1 U3451 ( .A1(n3336), .A2(n3337), .ZN(n3473) );
  NOR2_X1 U3452 ( .A1(n2282), .A2(n2281), .ZN(n3338) );
  NAND2_X1 U3453 ( .A1(n3336), .A2(n3337), .ZN(n3471) );
  NAND2_X1 U3454 ( .A1(n3386), .A2(n3474), .ZN(n3337) );
  NAND2_X1 U3455 ( .A1(n3385), .A2(n3387), .ZN(n3474) );
  NAND2_X1 U3456 ( .A1(n3475), .A2(n3476), .ZN(n3387) );
  NAND2_X1 U3457 ( .A1(b_6_), .A2(a_9_), .ZN(n3476) );
  INV_X1 U3458 ( .A(n3477), .ZN(n3475) );
  XNOR2_X1 U3459 ( .A(n3478), .B(n3479), .ZN(n3385) );
  XNOR2_X1 U3460 ( .A(n3480), .B(n3481), .ZN(n3478) );
  NAND2_X1 U3461 ( .A1(a_9_), .A2(n3477), .ZN(n3386) );
  NAND2_X1 U3462 ( .A1(n3382), .A2(n3482), .ZN(n3477) );
  NAND2_X1 U3463 ( .A1(n3381), .A2(n3383), .ZN(n3482) );
  NAND2_X1 U3464 ( .A1(n3483), .A2(n3484), .ZN(n3383) );
  NAND2_X1 U3465 ( .A1(b_6_), .A2(a_10_), .ZN(n3484) );
  INV_X1 U3466 ( .A(n3485), .ZN(n3483) );
  XNOR2_X1 U3467 ( .A(n3486), .B(n3487), .ZN(n3381) );
  XNOR2_X1 U3468 ( .A(n3488), .B(n3489), .ZN(n3487) );
  NAND2_X1 U3469 ( .A1(a_10_), .A2(n3485), .ZN(n3382) );
  NAND2_X1 U3470 ( .A1(n3352), .A2(n3490), .ZN(n3485) );
  NAND2_X1 U3471 ( .A1(n3351), .A2(n3353), .ZN(n3490) );
  NAND2_X1 U3472 ( .A1(n3491), .A2(n3492), .ZN(n3353) );
  NAND2_X1 U3473 ( .A1(b_6_), .A2(a_11_), .ZN(n3492) );
  INV_X1 U3474 ( .A(n3493), .ZN(n3491) );
  XOR2_X1 U3475 ( .A(n3494), .B(n3495), .Z(n3351) );
  XNOR2_X1 U3476 ( .A(n3496), .B(n3497), .ZN(n3494) );
  NAND2_X1 U3477 ( .A1(b_5_), .A2(a_12_), .ZN(n3496) );
  NAND2_X1 U3478 ( .A1(a_11_), .A2(n3493), .ZN(n3352) );
  NAND2_X1 U3479 ( .A1(n3498), .A2(n3499), .ZN(n3493) );
  NAND2_X1 U3480 ( .A1(n3500), .A2(b_6_), .ZN(n3499) );
  NOR2_X1 U3481 ( .A1(n3501), .A2(n2277), .ZN(n3500) );
  NOR2_X1 U3482 ( .A1(n3359), .A2(n3361), .ZN(n3501) );
  NAND2_X1 U3483 ( .A1(n3359), .A2(n3361), .ZN(n3498) );
  NAND2_X1 U3484 ( .A1(n3502), .A2(n3503), .ZN(n3361) );
  NAND2_X1 U3485 ( .A1(n3377), .A2(n3504), .ZN(n3503) );
  OR2_X1 U3486 ( .A1(n3378), .A2(n3379), .ZN(n3504) );
  NOR2_X1 U3487 ( .A1(n2282), .A2(n2042), .ZN(n3377) );
  NAND2_X1 U3488 ( .A1(n3379), .A2(n3378), .ZN(n3502) );
  NAND2_X1 U3489 ( .A1(n3505), .A2(n3506), .ZN(n3378) );
  NAND2_X1 U3490 ( .A1(b_4_), .A2(n3507), .ZN(n3506) );
  NAND2_X1 U3491 ( .A1(n2018), .A2(n3508), .ZN(n3507) );
  NAND2_X1 U3492 ( .A1(a_15_), .A2(n2163), .ZN(n3508) );
  NAND2_X1 U3493 ( .A1(b_5_), .A2(n3509), .ZN(n3505) );
  NAND2_X1 U3494 ( .A1(n2021), .A2(n3510), .ZN(n3509) );
  NAND2_X1 U3495 ( .A1(a_14_), .A2(n2284), .ZN(n3510) );
  AND2_X1 U3496 ( .A1(n3511), .A2(n2558), .ZN(n3379) );
  NOR2_X1 U3497 ( .A1(n2163), .A2(n2282), .ZN(n3511) );
  XOR2_X1 U3498 ( .A(n3512), .B(n3513), .Z(n3359) );
  XOR2_X1 U3499 ( .A(n3514), .B(n3515), .Z(n3512) );
  XNOR2_X1 U3500 ( .A(n3516), .B(n3517), .ZN(n3336) );
  NAND2_X1 U3501 ( .A1(n3518), .A2(n3519), .ZN(n3516) );
  XOR2_X1 U3502 ( .A(n3520), .B(n3521), .Z(n3399) );
  XOR2_X1 U3503 ( .A(n2251), .B(n3522), .Z(n3521) );
  XNOR2_X1 U3504 ( .A(n3523), .B(n3524), .ZN(n3408) );
  XOR2_X1 U3505 ( .A(n3525), .B(n3526), .Z(n3524) );
  NAND2_X1 U3506 ( .A1(a_3_), .A2(b_5_), .ZN(n3526) );
  XNOR2_X1 U3507 ( .A(n3527), .B(n3528), .ZN(n3411) );
  XOR2_X1 U3508 ( .A(n3529), .B(n3530), .Z(n3528) );
  NAND2_X1 U3509 ( .A1(a_2_), .A2(b_5_), .ZN(n3530) );
  XNOR2_X1 U3510 ( .A(n3531), .B(n3532), .ZN(n3297) );
  XOR2_X1 U3511 ( .A(n3533), .B(n3534), .Z(n3532) );
  NAND2_X1 U3512 ( .A1(b_5_), .A2(a_1_), .ZN(n3534) );
  NAND2_X1 U3513 ( .A1(n3535), .A2(n3536), .ZN(n1999) );
  NAND2_X1 U3514 ( .A1(n3421), .A2(n3417), .ZN(n3536) );
  XNOR2_X1 U3515 ( .A(n3537), .B(n3538), .ZN(n3535) );
  NAND2_X1 U3516 ( .A1(n3539), .A2(n3540), .ZN(n1998) );
  XOR2_X1 U3517 ( .A(n3537), .B(n3538), .Z(n3540) );
  AND2_X1 U3518 ( .A1(n3417), .A2(n3421), .ZN(n3539) );
  INV_X1 U3519 ( .A(n3418), .ZN(n3421) );
  XNOR2_X1 U3520 ( .A(n3541), .B(n3542), .ZN(n3418) );
  XOR2_X1 U3521 ( .A(n3543), .B(n3544), .Z(n3541) );
  NOR2_X1 U3522 ( .A1(n2284), .A2(n2376), .ZN(n3544) );
  NAND2_X1 U3523 ( .A1(n3545), .A2(n3546), .ZN(n3417) );
  NAND2_X1 U3524 ( .A1(n3547), .A2(a_0_), .ZN(n3546) );
  NOR2_X1 U3525 ( .A1(n3548), .A2(n2163), .ZN(n3547) );
  NOR2_X1 U3526 ( .A1(n3424), .A2(n3422), .ZN(n3548) );
  NAND2_X1 U3527 ( .A1(n3422), .A2(n3424), .ZN(n3545) );
  NAND2_X1 U3528 ( .A1(n3549), .A2(n3550), .ZN(n3424) );
  NAND2_X1 U3529 ( .A1(n3551), .A2(b_5_), .ZN(n3550) );
  NOR2_X1 U3530 ( .A1(n3552), .A2(n2381), .ZN(n3551) );
  NOR2_X1 U3531 ( .A1(n3531), .A2(n3533), .ZN(n3552) );
  NAND2_X1 U3532 ( .A1(n3531), .A2(n3533), .ZN(n3549) );
  NAND2_X1 U3533 ( .A1(n3553), .A2(n3554), .ZN(n3533) );
  NAND2_X1 U3534 ( .A1(n3555), .A2(a_2_), .ZN(n3554) );
  NOR2_X1 U3535 ( .A1(n3556), .A2(n2163), .ZN(n3555) );
  NOR2_X1 U3536 ( .A1(n3529), .A2(n3527), .ZN(n3556) );
  NAND2_X1 U3537 ( .A1(n3527), .A2(n3529), .ZN(n3553) );
  NAND2_X1 U3538 ( .A1(n3557), .A2(n3558), .ZN(n3529) );
  NAND2_X1 U3539 ( .A1(n3559), .A2(a_3_), .ZN(n3558) );
  NOR2_X1 U3540 ( .A1(n3560), .A2(n2163), .ZN(n3559) );
  NOR2_X1 U3541 ( .A1(n3523), .A2(n3525), .ZN(n3560) );
  NAND2_X1 U3542 ( .A1(n3523), .A2(n3525), .ZN(n3557) );
  NAND2_X1 U3543 ( .A1(n3561), .A2(n3562), .ZN(n3525) );
  NAND2_X1 U3544 ( .A1(n3563), .A2(a_4_), .ZN(n3562) );
  NOR2_X1 U3545 ( .A1(n3564), .A2(n2163), .ZN(n3563) );
  NOR2_X1 U3546 ( .A1(n3444), .A2(n3442), .ZN(n3564) );
  NAND2_X1 U3547 ( .A1(n3442), .A2(n3444), .ZN(n3561) );
  NAND2_X1 U3548 ( .A1(n3565), .A2(n3566), .ZN(n3444) );
  NAND2_X1 U3549 ( .A1(n3520), .A2(n3567), .ZN(n3566) );
  OR2_X1 U3550 ( .A1(n3522), .A2(n2157), .ZN(n3567) );
  XNOR2_X1 U3551 ( .A(n3568), .B(n3569), .ZN(n3520) );
  XOR2_X1 U3552 ( .A(n3570), .B(n3571), .Z(n3569) );
  NAND2_X1 U3553 ( .A1(b_4_), .A2(a_6_), .ZN(n3571) );
  NAND2_X1 U3554 ( .A1(n2157), .A2(n3522), .ZN(n3565) );
  NAND2_X1 U3555 ( .A1(n3572), .A2(n3573), .ZN(n3522) );
  NAND2_X1 U3556 ( .A1(n3574), .A2(b_5_), .ZN(n3573) );
  NOR2_X1 U3557 ( .A1(n3575), .A2(n2283), .ZN(n3574) );
  NOR2_X1 U3558 ( .A1(n3453), .A2(n3451), .ZN(n3575) );
  NAND2_X1 U3559 ( .A1(n3451), .A2(n3453), .ZN(n3572) );
  NAND2_X1 U3560 ( .A1(n3576), .A2(n3577), .ZN(n3453) );
  NAND2_X1 U3561 ( .A1(n3578), .A2(b_5_), .ZN(n3577) );
  NOR2_X1 U3562 ( .A1(n3579), .A2(n2132), .ZN(n3578) );
  NOR2_X1 U3563 ( .A1(n3461), .A2(n3459), .ZN(n3579) );
  NAND2_X1 U3564 ( .A1(n3459), .A2(n3461), .ZN(n3576) );
  NAND2_X1 U3565 ( .A1(n3580), .A2(n3581), .ZN(n3461) );
  NAND2_X1 U3566 ( .A1(n3582), .A2(b_5_), .ZN(n3581) );
  NOR2_X1 U3567 ( .A1(n3583), .A2(n2281), .ZN(n3582) );
  NOR2_X1 U3568 ( .A1(n3469), .A2(n3468), .ZN(n3583) );
  NAND2_X1 U3569 ( .A1(n3468), .A2(n3469), .ZN(n3580) );
  NAND2_X1 U3570 ( .A1(n3518), .A2(n3584), .ZN(n3469) );
  NAND2_X1 U3571 ( .A1(n3517), .A2(n3519), .ZN(n3584) );
  NAND2_X1 U3572 ( .A1(n3585), .A2(n3586), .ZN(n3519) );
  NAND2_X1 U3573 ( .A1(b_5_), .A2(a_9_), .ZN(n3586) );
  INV_X1 U3574 ( .A(n3587), .ZN(n3585) );
  XNOR2_X1 U3575 ( .A(n3588), .B(n3589), .ZN(n3517) );
  XNOR2_X1 U3576 ( .A(n3590), .B(n3591), .ZN(n3588) );
  NAND2_X1 U3577 ( .A1(a_9_), .A2(n3587), .ZN(n3518) );
  NAND2_X1 U3578 ( .A1(n3592), .A2(n3593), .ZN(n3587) );
  NAND2_X1 U3579 ( .A1(n3481), .A2(n3594), .ZN(n3593) );
  NAND2_X1 U3580 ( .A1(n3479), .A2(n3480), .ZN(n3594) );
  NOR2_X1 U3581 ( .A1(n2163), .A2(n2279), .ZN(n3481) );
  OR2_X1 U3582 ( .A1(n3479), .A2(n3480), .ZN(n3592) );
  AND2_X1 U3583 ( .A1(n3595), .A2(n3596), .ZN(n3480) );
  NAND2_X1 U3584 ( .A1(n3489), .A2(n3597), .ZN(n3596) );
  OR2_X1 U3585 ( .A1(n3486), .A2(n3488), .ZN(n3597) );
  NOR2_X1 U3586 ( .A1(n2163), .A2(n2072), .ZN(n3489) );
  NAND2_X1 U3587 ( .A1(n3486), .A2(n3488), .ZN(n3595) );
  NAND2_X1 U3588 ( .A1(n3598), .A2(n3599), .ZN(n3488) );
  NAND2_X1 U3589 ( .A1(n3600), .A2(b_5_), .ZN(n3599) );
  NOR2_X1 U3590 ( .A1(n3601), .A2(n2277), .ZN(n3600) );
  NOR2_X1 U3591 ( .A1(n3495), .A2(n3497), .ZN(n3601) );
  NAND2_X1 U3592 ( .A1(n3495), .A2(n3497), .ZN(n3598) );
  NAND2_X1 U3593 ( .A1(n3602), .A2(n3603), .ZN(n3497) );
  NAND2_X1 U3594 ( .A1(n3513), .A2(n3604), .ZN(n3603) );
  OR2_X1 U3595 ( .A1(n3514), .A2(n3515), .ZN(n3604) );
  NOR2_X1 U3596 ( .A1(n2163), .A2(n2042), .ZN(n3513) );
  NAND2_X1 U3597 ( .A1(n3515), .A2(n3514), .ZN(n3602) );
  NAND2_X1 U3598 ( .A1(n3605), .A2(n3606), .ZN(n3514) );
  NAND2_X1 U3599 ( .A1(b_3_), .A2(n3607), .ZN(n3606) );
  NAND2_X1 U3600 ( .A1(n2018), .A2(n3608), .ZN(n3607) );
  NAND2_X1 U3601 ( .A1(a_15_), .A2(n2284), .ZN(n3608) );
  NAND2_X1 U3602 ( .A1(b_4_), .A2(n3609), .ZN(n3605) );
  NAND2_X1 U3603 ( .A1(n2021), .A2(n3610), .ZN(n3609) );
  NAND2_X1 U3604 ( .A1(a_14_), .A2(n2200), .ZN(n3610) );
  AND2_X1 U3605 ( .A1(n3611), .A2(n2558), .ZN(n3515) );
  NOR2_X1 U3606 ( .A1(n2163), .A2(n2284), .ZN(n3611) );
  XNOR2_X1 U3607 ( .A(n3612), .B(n3613), .ZN(n3495) );
  XNOR2_X1 U3608 ( .A(n3614), .B(n3615), .ZN(n3613) );
  XOR2_X1 U3609 ( .A(n3616), .B(n3617), .Z(n3486) );
  XNOR2_X1 U3610 ( .A(n3618), .B(n3619), .ZN(n3616) );
  NAND2_X1 U3611 ( .A1(b_4_), .A2(a_12_), .ZN(n3618) );
  XOR2_X1 U3612 ( .A(n3620), .B(n3621), .Z(n3479) );
  NAND2_X1 U3613 ( .A1(n3622), .A2(n3623), .ZN(n3620) );
  XNOR2_X1 U3614 ( .A(n3624), .B(n3625), .ZN(n3468) );
  NAND2_X1 U3615 ( .A1(n3626), .A2(n3627), .ZN(n3624) );
  XOR2_X1 U3616 ( .A(n3628), .B(n3629), .Z(n3459) );
  XOR2_X1 U3617 ( .A(n3630), .B(n3631), .Z(n3628) );
  NOR2_X1 U3618 ( .A1(n2281), .A2(n2284), .ZN(n3631) );
  XNOR2_X1 U3619 ( .A(n3632), .B(n3633), .ZN(n3451) );
  XOR2_X1 U3620 ( .A(n3634), .B(n3635), .Z(n3633) );
  NAND2_X1 U3621 ( .A1(b_4_), .A2(a_7_), .ZN(n3635) );
  INV_X1 U3622 ( .A(n2251), .ZN(n2157) );
  NAND2_X1 U3623 ( .A1(a_5_), .A2(b_5_), .ZN(n2251) );
  XNOR2_X1 U3624 ( .A(n3636), .B(n3637), .ZN(n3442) );
  XOR2_X1 U3625 ( .A(n3638), .B(n3639), .Z(n3637) );
  NAND2_X1 U3626 ( .A1(b_4_), .A2(a_5_), .ZN(n3639) );
  XNOR2_X1 U3627 ( .A(n3640), .B(n3641), .ZN(n3523) );
  XOR2_X1 U3628 ( .A(n3642), .B(n2181), .Z(n3641) );
  XOR2_X1 U3629 ( .A(n3643), .B(n3644), .Z(n3527) );
  XNOR2_X1 U3630 ( .A(n3645), .B(n3646), .ZN(n3643) );
  NAND2_X1 U3631 ( .A1(a_3_), .A2(b_4_), .ZN(n3645) );
  XOR2_X1 U3632 ( .A(n3647), .B(n3648), .Z(n3531) );
  XNOR2_X1 U3633 ( .A(n3649), .B(n3650), .ZN(n3647) );
  NAND2_X1 U3634 ( .A1(a_2_), .A2(b_4_), .ZN(n3649) );
  XOR2_X1 U3635 ( .A(n3651), .B(n3652), .Z(n3422) );
  XOR2_X1 U3636 ( .A(n3653), .B(n3654), .Z(n3651) );
  NOR2_X1 U3637 ( .A1(n2381), .A2(n2284), .ZN(n3654) );
  NAND2_X1 U3638 ( .A1(n3655), .A2(n3656), .ZN(n2004) );
  NAND2_X1 U3639 ( .A1(n3538), .A2(n3537), .ZN(n3656) );
  XOR2_X1 U3640 ( .A(n3657), .B(n3658), .Z(n3655) );
  NAND2_X1 U3641 ( .A1(n3659), .A2(n3660), .ZN(n2003) );
  XOR2_X1 U3642 ( .A(n3657), .B(n3661), .Z(n3660) );
  AND2_X1 U3643 ( .A1(n3537), .A2(n3538), .ZN(n3659) );
  XOR2_X1 U3644 ( .A(n3662), .B(n3663), .Z(n3538) );
  XOR2_X1 U3645 ( .A(n3664), .B(n3665), .Z(n3662) );
  NOR2_X1 U3646 ( .A1(n2200), .A2(n2376), .ZN(n3665) );
  NAND2_X1 U3647 ( .A1(n3666), .A2(n3667), .ZN(n3537) );
  NAND2_X1 U3648 ( .A1(n3668), .A2(a_0_), .ZN(n3667) );
  NOR2_X1 U3649 ( .A1(n3669), .A2(n2284), .ZN(n3668) );
  NOR2_X1 U3650 ( .A1(n3542), .A2(n3543), .ZN(n3669) );
  NAND2_X1 U3651 ( .A1(n3542), .A2(n3543), .ZN(n3666) );
  NAND2_X1 U3652 ( .A1(n3670), .A2(n3671), .ZN(n3543) );
  NAND2_X1 U3653 ( .A1(n3672), .A2(b_4_), .ZN(n3671) );
  NOR2_X1 U3654 ( .A1(n3673), .A2(n2381), .ZN(n3672) );
  NOR2_X1 U3655 ( .A1(n3652), .A2(n3653), .ZN(n3673) );
  NAND2_X1 U3656 ( .A1(n3652), .A2(n3653), .ZN(n3670) );
  NAND2_X1 U3657 ( .A1(n3674), .A2(n3675), .ZN(n3653) );
  NAND2_X1 U3658 ( .A1(n3676), .A2(a_2_), .ZN(n3675) );
  NOR2_X1 U3659 ( .A1(n3677), .A2(n2284), .ZN(n3676) );
  NOR2_X1 U3660 ( .A1(n3650), .A2(n3648), .ZN(n3677) );
  NAND2_X1 U3661 ( .A1(n3648), .A2(n3650), .ZN(n3674) );
  NAND2_X1 U3662 ( .A1(n3678), .A2(n3679), .ZN(n3650) );
  NAND2_X1 U3663 ( .A1(n3680), .A2(a_3_), .ZN(n3679) );
  NOR2_X1 U3664 ( .A1(n3681), .A2(n2284), .ZN(n3680) );
  NOR2_X1 U3665 ( .A1(n3644), .A2(n3646), .ZN(n3681) );
  NAND2_X1 U3666 ( .A1(n3644), .A2(n3646), .ZN(n3678) );
  NAND2_X1 U3667 ( .A1(n3682), .A2(n3683), .ZN(n3646) );
  NAND2_X1 U3668 ( .A1(n3640), .A2(n3684), .ZN(n3683) );
  OR2_X1 U3669 ( .A1(n3642), .A2(n3685), .ZN(n3684) );
  XOR2_X1 U3670 ( .A(n3686), .B(n3687), .Z(n3640) );
  XOR2_X1 U3671 ( .A(n3688), .B(n3689), .Z(n3686) );
  NOR2_X1 U3672 ( .A1(n2162), .A2(n2200), .ZN(n3689) );
  NAND2_X1 U3673 ( .A1(n3685), .A2(n3642), .ZN(n3682) );
  NAND2_X1 U3674 ( .A1(n3690), .A2(n3691), .ZN(n3642) );
  NAND2_X1 U3675 ( .A1(n3692), .A2(b_4_), .ZN(n3691) );
  NOR2_X1 U3676 ( .A1(n3693), .A2(n2162), .ZN(n3692) );
  NOR2_X1 U3677 ( .A1(n3636), .A2(n3638), .ZN(n3693) );
  NAND2_X1 U3678 ( .A1(n3636), .A2(n3638), .ZN(n3690) );
  NAND2_X1 U3679 ( .A1(n3694), .A2(n3695), .ZN(n3638) );
  NAND2_X1 U3680 ( .A1(n3696), .A2(b_4_), .ZN(n3695) );
  NOR2_X1 U3681 ( .A1(n3697), .A2(n2283), .ZN(n3696) );
  NOR2_X1 U3682 ( .A1(n3568), .A2(n3570), .ZN(n3697) );
  NAND2_X1 U3683 ( .A1(n3568), .A2(n3570), .ZN(n3694) );
  NAND2_X1 U3684 ( .A1(n3698), .A2(n3699), .ZN(n3570) );
  NAND2_X1 U3685 ( .A1(n3700), .A2(b_4_), .ZN(n3699) );
  NOR2_X1 U3686 ( .A1(n3701), .A2(n2132), .ZN(n3700) );
  NOR2_X1 U3687 ( .A1(n3632), .A2(n3634), .ZN(n3701) );
  NAND2_X1 U3688 ( .A1(n3632), .A2(n3634), .ZN(n3698) );
  NAND2_X1 U3689 ( .A1(n3702), .A2(n3703), .ZN(n3634) );
  NAND2_X1 U3690 ( .A1(n3704), .A2(b_4_), .ZN(n3703) );
  NOR2_X1 U3691 ( .A1(n3705), .A2(n2281), .ZN(n3704) );
  NOR2_X1 U3692 ( .A1(n3629), .A2(n3630), .ZN(n3705) );
  NAND2_X1 U3693 ( .A1(n3629), .A2(n3630), .ZN(n3702) );
  NAND2_X1 U3694 ( .A1(n3626), .A2(n3706), .ZN(n3630) );
  NAND2_X1 U3695 ( .A1(n3625), .A2(n3627), .ZN(n3706) );
  NAND2_X1 U3696 ( .A1(n3707), .A2(n3708), .ZN(n3627) );
  NAND2_X1 U3697 ( .A1(b_4_), .A2(a_9_), .ZN(n3708) );
  INV_X1 U3698 ( .A(n3709), .ZN(n3707) );
  XNOR2_X1 U3699 ( .A(n3710), .B(n3711), .ZN(n3625) );
  NAND2_X1 U3700 ( .A1(n3712), .A2(n3713), .ZN(n3710) );
  NAND2_X1 U3701 ( .A1(a_9_), .A2(n3709), .ZN(n3626) );
  NAND2_X1 U3702 ( .A1(n3714), .A2(n3715), .ZN(n3709) );
  NAND2_X1 U3703 ( .A1(n3590), .A2(n3716), .ZN(n3715) );
  NAND2_X1 U3704 ( .A1(n3591), .A2(n3589), .ZN(n3716) );
  NOR2_X1 U3705 ( .A1(n2284), .A2(n2279), .ZN(n3590) );
  OR2_X1 U3706 ( .A1(n3589), .A2(n3591), .ZN(n3714) );
  AND2_X1 U3707 ( .A1(n3622), .A2(n3717), .ZN(n3591) );
  NAND2_X1 U3708 ( .A1(n3621), .A2(n3623), .ZN(n3717) );
  NAND2_X1 U3709 ( .A1(n3718), .A2(n3719), .ZN(n3623) );
  NAND2_X1 U3710 ( .A1(b_4_), .A2(a_11_), .ZN(n3719) );
  INV_X1 U3711 ( .A(n3720), .ZN(n3718) );
  XNOR2_X1 U3712 ( .A(n3721), .B(n3722), .ZN(n3621) );
  XNOR2_X1 U3713 ( .A(n3723), .B(n3724), .ZN(n3722) );
  NAND2_X1 U3714 ( .A1(a_11_), .A2(n3720), .ZN(n3622) );
  NAND2_X1 U3715 ( .A1(n3725), .A2(n3726), .ZN(n3720) );
  NAND2_X1 U3716 ( .A1(n3727), .A2(b_4_), .ZN(n3726) );
  NOR2_X1 U3717 ( .A1(n3728), .A2(n2277), .ZN(n3727) );
  NOR2_X1 U3718 ( .A1(n3617), .A2(n3619), .ZN(n3728) );
  NAND2_X1 U3719 ( .A1(n3617), .A2(n3619), .ZN(n3725) );
  NAND2_X1 U3720 ( .A1(n3729), .A2(n3730), .ZN(n3619) );
  NAND2_X1 U3721 ( .A1(n3612), .A2(n3731), .ZN(n3730) );
  OR2_X1 U3722 ( .A1(n3615), .A2(n3614), .ZN(n3731) );
  NOR2_X1 U3723 ( .A1(n2284), .A2(n2042), .ZN(n3612) );
  NAND2_X1 U3724 ( .A1(n3614), .A2(n3615), .ZN(n3729) );
  NAND2_X1 U3725 ( .A1(n3732), .A2(n3733), .ZN(n3615) );
  NAND2_X1 U3726 ( .A1(b_2_), .A2(n3734), .ZN(n3733) );
  NAND2_X1 U3727 ( .A1(n2018), .A2(n3735), .ZN(n3734) );
  NAND2_X1 U3728 ( .A1(a_15_), .A2(n2200), .ZN(n3735) );
  NAND2_X1 U3729 ( .A1(b_3_), .A2(n3736), .ZN(n3732) );
  NAND2_X1 U3730 ( .A1(n2021), .A2(n3737), .ZN(n3736) );
  NAND2_X1 U3731 ( .A1(a_14_), .A2(n2286), .ZN(n3737) );
  AND2_X1 U3732 ( .A1(n3738), .A2(n2558), .ZN(n3614) );
  NOR2_X1 U3733 ( .A1(n2200), .A2(n2284), .ZN(n3738) );
  XOR2_X1 U3734 ( .A(n3739), .B(n3740), .Z(n3617) );
  NOR2_X1 U3735 ( .A1(n2042), .A2(n2200), .ZN(n3740) );
  XOR2_X1 U3736 ( .A(n3741), .B(n3742), .Z(n3739) );
  XOR2_X1 U3737 ( .A(n3743), .B(n3744), .Z(n3589) );
  NAND2_X1 U3738 ( .A1(n3745), .A2(n3746), .ZN(n3743) );
  XNOR2_X1 U3739 ( .A(n3747), .B(n3748), .ZN(n3629) );
  NAND2_X1 U3740 ( .A1(n3749), .A2(n3750), .ZN(n3747) );
  XNOR2_X1 U3741 ( .A(n3751), .B(n3752), .ZN(n3632) );
  XOR2_X1 U3742 ( .A(n3753), .B(n3754), .Z(n3752) );
  NAND2_X1 U3743 ( .A1(b_3_), .A2(a_8_), .ZN(n3754) );
  XNOR2_X1 U3744 ( .A(n3755), .B(n3756), .ZN(n3568) );
  NAND2_X1 U3745 ( .A1(n3757), .A2(n3758), .ZN(n3755) );
  XOR2_X1 U3746 ( .A(n3759), .B(n3760), .Z(n3636) );
  XNOR2_X1 U3747 ( .A(n3761), .B(n3762), .ZN(n3759) );
  NAND2_X1 U3748 ( .A1(b_3_), .A2(a_6_), .ZN(n3761) );
  INV_X1 U3749 ( .A(n2181), .ZN(n3685) );
  NAND2_X1 U3750 ( .A1(b_4_), .A2(a_4_), .ZN(n2181) );
  XOR2_X1 U3751 ( .A(n3763), .B(n3764), .Z(n3644) );
  XOR2_X1 U3752 ( .A(n3765), .B(n3766), .Z(n3763) );
  NOR2_X1 U3753 ( .A1(n2285), .A2(n2200), .ZN(n3766) );
  XOR2_X1 U3754 ( .A(n3767), .B(n3768), .Z(n3648) );
  XOR2_X1 U3755 ( .A(n3769), .B(n2194), .Z(n3767) );
  XOR2_X1 U3756 ( .A(n3770), .B(n3771), .Z(n3652) );
  XNOR2_X1 U3757 ( .A(n3772), .B(n3773), .ZN(n3770) );
  NAND2_X1 U3758 ( .A1(a_2_), .A2(b_3_), .ZN(n3772) );
  XOR2_X1 U3759 ( .A(n3774), .B(n3775), .Z(n3542) );
  XOR2_X1 U3760 ( .A(n3776), .B(n3777), .Z(n3774) );
  NOR2_X1 U3761 ( .A1(n2381), .A2(n2200), .ZN(n3777) );
  NAND2_X1 U3762 ( .A1(n3778), .A2(n3779), .ZN(n2031) );
  NAND2_X1 U3763 ( .A1(n3661), .A2(n3657), .ZN(n3779) );
  XNOR2_X1 U3764 ( .A(n3780), .B(n3781), .ZN(n3778) );
  NAND2_X1 U3765 ( .A1(n3782), .A2(n3783), .ZN(n2030) );
  AND2_X1 U3766 ( .A1(n2332), .A2(n3657), .ZN(n3783) );
  NAND2_X1 U3767 ( .A1(n3784), .A2(n3785), .ZN(n3657) );
  NAND2_X1 U3768 ( .A1(n3786), .A2(a_0_), .ZN(n3785) );
  NOR2_X1 U3769 ( .A1(n3787), .A2(n2200), .ZN(n3786) );
  NOR2_X1 U3770 ( .A1(n3664), .A2(n3663), .ZN(n3787) );
  NAND2_X1 U3771 ( .A1(n3663), .A2(n3664), .ZN(n3784) );
  NAND2_X1 U3772 ( .A1(n3788), .A2(n3789), .ZN(n3664) );
  NAND2_X1 U3773 ( .A1(n3790), .A2(b_3_), .ZN(n3789) );
  NOR2_X1 U3774 ( .A1(n3791), .A2(n2381), .ZN(n3790) );
  NOR2_X1 U3775 ( .A1(n3776), .A2(n3775), .ZN(n3791) );
  NAND2_X1 U3776 ( .A1(n3775), .A2(n3776), .ZN(n3788) );
  NAND2_X1 U3777 ( .A1(n3792), .A2(n3793), .ZN(n3776) );
  NAND2_X1 U3778 ( .A1(n3794), .A2(a_2_), .ZN(n3793) );
  NOR2_X1 U3779 ( .A1(n3795), .A2(n2200), .ZN(n3794) );
  NOR2_X1 U3780 ( .A1(n3773), .A2(n3771), .ZN(n3795) );
  NAND2_X1 U3781 ( .A1(n3771), .A2(n3773), .ZN(n3792) );
  NAND2_X1 U3782 ( .A1(n3796), .A2(n3797), .ZN(n3773) );
  NAND2_X1 U3783 ( .A1(n3768), .A2(n3798), .ZN(n3797) );
  OR2_X1 U3784 ( .A1(n3769), .A2(n2194), .ZN(n3798) );
  XNOR2_X1 U3785 ( .A(n3799), .B(n3800), .ZN(n3768) );
  NAND2_X1 U3786 ( .A1(n3801), .A2(n3802), .ZN(n3799) );
  NAND2_X1 U3787 ( .A1(n2194), .A2(n3769), .ZN(n3796) );
  NAND2_X1 U3788 ( .A1(n3803), .A2(n3804), .ZN(n3769) );
  NAND2_X1 U3789 ( .A1(n3805), .A2(b_3_), .ZN(n3804) );
  NOR2_X1 U3790 ( .A1(n3806), .A2(n2285), .ZN(n3805) );
  NOR2_X1 U3791 ( .A1(n3765), .A2(n3764), .ZN(n3806) );
  NAND2_X1 U3792 ( .A1(n3764), .A2(n3765), .ZN(n3803) );
  NAND2_X1 U3793 ( .A1(n3807), .A2(n3808), .ZN(n3765) );
  NAND2_X1 U3794 ( .A1(n3809), .A2(b_3_), .ZN(n3808) );
  NOR2_X1 U3795 ( .A1(n3810), .A2(n2162), .ZN(n3809) );
  NOR2_X1 U3796 ( .A1(n3687), .A2(n3688), .ZN(n3810) );
  NAND2_X1 U3797 ( .A1(n3687), .A2(n3688), .ZN(n3807) );
  NAND2_X1 U3798 ( .A1(n3811), .A2(n3812), .ZN(n3688) );
  NAND2_X1 U3799 ( .A1(n3813), .A2(b_3_), .ZN(n3812) );
  NOR2_X1 U3800 ( .A1(n3814), .A2(n2283), .ZN(n3813) );
  NOR2_X1 U3801 ( .A1(n3762), .A2(n3760), .ZN(n3814) );
  NAND2_X1 U3802 ( .A1(n3760), .A2(n3762), .ZN(n3811) );
  NAND2_X1 U3803 ( .A1(n3757), .A2(n3815), .ZN(n3762) );
  NAND2_X1 U3804 ( .A1(n3756), .A2(n3758), .ZN(n3815) );
  NAND2_X1 U3805 ( .A1(n3816), .A2(n3817), .ZN(n3758) );
  NAND2_X1 U3806 ( .A1(b_3_), .A2(a_7_), .ZN(n3817) );
  INV_X1 U3807 ( .A(n3818), .ZN(n3816) );
  XNOR2_X1 U3808 ( .A(n3819), .B(n3820), .ZN(n3756) );
  NAND2_X1 U3809 ( .A1(n3821), .A2(n3822), .ZN(n3819) );
  NAND2_X1 U3810 ( .A1(a_7_), .A2(n3818), .ZN(n3757) );
  NAND2_X1 U3811 ( .A1(n3823), .A2(n3824), .ZN(n3818) );
  NAND2_X1 U3812 ( .A1(n3825), .A2(b_3_), .ZN(n3824) );
  NOR2_X1 U3813 ( .A1(n3826), .A2(n2281), .ZN(n3825) );
  NOR2_X1 U3814 ( .A1(n3753), .A2(n3751), .ZN(n3826) );
  NAND2_X1 U3815 ( .A1(n3751), .A2(n3753), .ZN(n3823) );
  NAND2_X1 U3816 ( .A1(n3749), .A2(n3827), .ZN(n3753) );
  NAND2_X1 U3817 ( .A1(n3748), .A2(n3750), .ZN(n3827) );
  NAND2_X1 U3818 ( .A1(n3828), .A2(n3829), .ZN(n3750) );
  NAND2_X1 U3819 ( .A1(b_3_), .A2(a_9_), .ZN(n3829) );
  INV_X1 U3820 ( .A(n3830), .ZN(n3828) );
  XNOR2_X1 U3821 ( .A(n3831), .B(n3832), .ZN(n3748) );
  NAND2_X1 U3822 ( .A1(n3833), .A2(n3834), .ZN(n3831) );
  NAND2_X1 U3823 ( .A1(a_9_), .A2(n3830), .ZN(n3749) );
  NAND2_X1 U3824 ( .A1(n3712), .A2(n3835), .ZN(n3830) );
  NAND2_X1 U3825 ( .A1(n3711), .A2(n3713), .ZN(n3835) );
  NAND2_X1 U3826 ( .A1(n3836), .A2(n3837), .ZN(n3713) );
  NAND2_X1 U3827 ( .A1(b_3_), .A2(a_10_), .ZN(n3837) );
  INV_X1 U3828 ( .A(n3838), .ZN(n3836) );
  XNOR2_X1 U3829 ( .A(n3839), .B(n3840), .ZN(n3711) );
  XNOR2_X1 U3830 ( .A(n3841), .B(n3842), .ZN(n3839) );
  NAND2_X1 U3831 ( .A1(a_10_), .A2(n3838), .ZN(n3712) );
  NAND2_X1 U3832 ( .A1(n3745), .A2(n3843), .ZN(n3838) );
  NAND2_X1 U3833 ( .A1(n3744), .A2(n3746), .ZN(n3843) );
  NAND2_X1 U3834 ( .A1(n3844), .A2(n3845), .ZN(n3746) );
  NAND2_X1 U3835 ( .A1(b_3_), .A2(a_11_), .ZN(n3845) );
  INV_X1 U3836 ( .A(n3846), .ZN(n3844) );
  XNOR2_X1 U3837 ( .A(n3847), .B(n3848), .ZN(n3744) );
  XNOR2_X1 U3838 ( .A(n3849), .B(n3850), .ZN(n3848) );
  NAND2_X1 U3839 ( .A1(a_11_), .A2(n3846), .ZN(n3745) );
  NAND2_X1 U3840 ( .A1(n3851), .A2(n3852), .ZN(n3846) );
  NAND2_X1 U3841 ( .A1(n3724), .A2(n3853), .ZN(n3852) );
  OR2_X1 U3842 ( .A1(n3723), .A2(n3721), .ZN(n3853) );
  NOR2_X1 U3843 ( .A1(n2200), .A2(n2277), .ZN(n3724) );
  NAND2_X1 U3844 ( .A1(n3721), .A2(n3723), .ZN(n3851) );
  NAND2_X1 U3845 ( .A1(n3854), .A2(n3855), .ZN(n3723) );
  NAND2_X1 U3846 ( .A1(n3856), .A2(b_3_), .ZN(n3855) );
  NOR2_X1 U3847 ( .A1(n3857), .A2(n2042), .ZN(n3856) );
  NOR2_X1 U3848 ( .A1(n3742), .A2(n3741), .ZN(n3857) );
  NAND2_X1 U3849 ( .A1(n3742), .A2(n3741), .ZN(n3854) );
  NAND2_X1 U3850 ( .A1(n3858), .A2(n3859), .ZN(n3741) );
  NAND2_X1 U3851 ( .A1(b_1_), .A2(n3860), .ZN(n3859) );
  NAND2_X1 U3852 ( .A1(n2018), .A2(n3861), .ZN(n3860) );
  NAND2_X1 U3853 ( .A1(a_15_), .A2(n2286), .ZN(n3861) );
  NAND2_X1 U3854 ( .A1(b_2_), .A2(n3862), .ZN(n3858) );
  NAND2_X1 U3855 ( .A1(n2021), .A2(n3863), .ZN(n3862) );
  NAND2_X1 U3856 ( .A1(a_14_), .A2(n3864), .ZN(n3863) );
  AND2_X1 U3857 ( .A1(n3865), .A2(n2558), .ZN(n3742) );
  NOR2_X1 U3858 ( .A1(n2200), .A2(n2286), .ZN(n3865) );
  XOR2_X1 U3859 ( .A(n3866), .B(n3867), .Z(n3721) );
  NOR2_X1 U3860 ( .A1(n2042), .A2(n2286), .ZN(n3867) );
  XOR2_X1 U3861 ( .A(n3868), .B(n3869), .Z(n3866) );
  XOR2_X1 U3862 ( .A(n3870), .B(n3871), .Z(n3751) );
  XOR2_X1 U3863 ( .A(n3872), .B(n3873), .Z(n3870) );
  XNOR2_X1 U3864 ( .A(n3874), .B(n3875), .ZN(n3760) );
  XNOR2_X1 U3865 ( .A(n3876), .B(n3877), .ZN(n3874) );
  XNOR2_X1 U3866 ( .A(n3878), .B(n3879), .ZN(n3687) );
  NAND2_X1 U3867 ( .A1(n3880), .A2(n3881), .ZN(n3878) );
  XNOR2_X1 U3868 ( .A(n3882), .B(n3883), .ZN(n3764) );
  XNOR2_X1 U3869 ( .A(n3884), .B(n3885), .ZN(n3882) );
  INV_X1 U3870 ( .A(n2247), .ZN(n2194) );
  NAND2_X1 U3871 ( .A1(a_3_), .A2(b_3_), .ZN(n2247) );
  XNOR2_X1 U3872 ( .A(n3886), .B(n3887), .ZN(n3771) );
  XNOR2_X1 U3873 ( .A(n3888), .B(n3889), .ZN(n3886) );
  XOR2_X1 U3874 ( .A(n3890), .B(n3891), .Z(n3775) );
  XOR2_X1 U3875 ( .A(n3892), .B(n3893), .Z(n3890) );
  XNOR2_X1 U3876 ( .A(n3894), .B(n3895), .ZN(n3663) );
  XNOR2_X1 U3877 ( .A(n3896), .B(n3897), .ZN(n3894) );
  NAND2_X1 U3878 ( .A1(n3780), .A2(n3781), .ZN(n2332) );
  NOR2_X1 U3879 ( .A1(n3898), .A2(n3658), .ZN(n3782) );
  INV_X1 U3880 ( .A(n3661), .ZN(n3658) );
  XOR2_X1 U3881 ( .A(n3899), .B(n3900), .Z(n3661) );
  XNOR2_X1 U3882 ( .A(n3901), .B(n3902), .ZN(n3899) );
  NOR2_X1 U3883 ( .A1(n2286), .A2(n2376), .ZN(n3902) );
  NOR2_X1 U3884 ( .A1(n3781), .A2(n3780), .ZN(n3898) );
  NAND2_X1 U3885 ( .A1(n3903), .A2(n3904), .ZN(n3780) );
  XNOR2_X1 U3886 ( .A(n2335), .B(n2336), .ZN(n3904) );
  NOR2_X1 U3887 ( .A1(n2381), .A2(n2333), .ZN(n2336) );
  NOR2_X1 U3888 ( .A1(n2376), .A2(n3864), .ZN(n2335) );
  NOR2_X1 U3889 ( .A1(n3905), .A2(n3906), .ZN(n3903) );
  NOR2_X1 U3890 ( .A1(n2288), .A2(n3907), .ZN(n3905) );
  NAND2_X1 U3891 ( .A1(n3901), .A2(n3908), .ZN(n3781) );
  NAND2_X1 U3892 ( .A1(n3900), .A2(b_2_), .ZN(n3908) );
  XNOR2_X1 U3893 ( .A(n3907), .B(n3909), .ZN(n3900) );
  NOR2_X1 U3894 ( .A1(n2288), .A2(n3906), .ZN(n3909) );
  NAND2_X1 U3895 ( .A1(n3910), .A2(n3911), .ZN(n3906) );
  NAND2_X1 U3896 ( .A1(n3912), .A2(n3913), .ZN(n3911) );
  OR2_X1 U3897 ( .A1(n3914), .A2(a_2_), .ZN(n3912) );
  NAND2_X1 U3898 ( .A1(b_1_), .A2(a_1_), .ZN(n2288) );
  NAND2_X1 U3899 ( .A1(a_2_), .A2(b_0_), .ZN(n3907) );
  AND2_X1 U3900 ( .A1(n3915), .A2(n3916), .ZN(n3901) );
  NAND2_X1 U3901 ( .A1(n3897), .A2(n3917), .ZN(n3916) );
  NAND2_X1 U3902 ( .A1(n3896), .A2(n3895), .ZN(n3917) );
  NOR2_X1 U3903 ( .A1(n2286), .A2(n2381), .ZN(n3897) );
  INV_X1 U3904 ( .A(a_1_), .ZN(n2381) );
  OR2_X1 U3905 ( .A1(n3895), .A2(n3896), .ZN(n3915) );
  AND2_X1 U3906 ( .A1(n3918), .A2(n3919), .ZN(n3896) );
  NAND2_X1 U3907 ( .A1(n3891), .A2(n3920), .ZN(n3919) );
  OR2_X1 U3908 ( .A1(n3892), .A2(n3893), .ZN(n3920) );
  XOR2_X1 U3909 ( .A(n3921), .B(n3922), .Z(n3891) );
  XNOR2_X1 U3910 ( .A(n3923), .B(n3924), .ZN(n3922) );
  NAND2_X1 U3911 ( .A1(b_1_), .A2(a_3_), .ZN(n3921) );
  NAND2_X1 U3912 ( .A1(n3893), .A2(n3892), .ZN(n3918) );
  NAND2_X1 U3913 ( .A1(n3925), .A2(n3926), .ZN(n3892) );
  NAND2_X1 U3914 ( .A1(n3889), .A2(n3927), .ZN(n3926) );
  NAND2_X1 U3915 ( .A1(n3888), .A2(n3887), .ZN(n3927) );
  NOR2_X1 U3916 ( .A1(n2286), .A2(n2199), .ZN(n3889) );
  OR2_X1 U3917 ( .A1(n3887), .A2(n3888), .ZN(n3925) );
  AND2_X1 U3918 ( .A1(n3801), .A2(n3928), .ZN(n3888) );
  NAND2_X1 U3919 ( .A1(n3800), .A2(n3802), .ZN(n3928) );
  NAND2_X1 U3920 ( .A1(n3929), .A2(n3930), .ZN(n3802) );
  NAND2_X1 U3921 ( .A1(b_2_), .A2(a_4_), .ZN(n3930) );
  INV_X1 U3922 ( .A(n3931), .ZN(n3929) );
  XOR2_X1 U3923 ( .A(n3932), .B(n3933), .Z(n3800) );
  XNOR2_X1 U3924 ( .A(n3934), .B(n3935), .ZN(n3933) );
  NAND2_X1 U3925 ( .A1(b_1_), .A2(a_5_), .ZN(n3932) );
  NAND2_X1 U3926 ( .A1(a_4_), .A2(n3931), .ZN(n3801) );
  NAND2_X1 U3927 ( .A1(n3936), .A2(n3937), .ZN(n3931) );
  NAND2_X1 U3928 ( .A1(n3885), .A2(n3938), .ZN(n3937) );
  NAND2_X1 U3929 ( .A1(n3884), .A2(n3883), .ZN(n3938) );
  NOR2_X1 U3930 ( .A1(n2286), .A2(n2162), .ZN(n3885) );
  OR2_X1 U3931 ( .A1(n3883), .A2(n3884), .ZN(n3936) );
  AND2_X1 U3932 ( .A1(n3880), .A2(n3939), .ZN(n3884) );
  NAND2_X1 U3933 ( .A1(n3879), .A2(n3881), .ZN(n3939) );
  NAND2_X1 U3934 ( .A1(n3940), .A2(n3941), .ZN(n3881) );
  NAND2_X1 U3935 ( .A1(b_2_), .A2(a_6_), .ZN(n3941) );
  INV_X1 U3936 ( .A(n3942), .ZN(n3940) );
  XOR2_X1 U3937 ( .A(n3943), .B(n3944), .Z(n3879) );
  XNOR2_X1 U3938 ( .A(n3945), .B(n3946), .ZN(n3944) );
  NAND2_X1 U3939 ( .A1(b_1_), .A2(a_7_), .ZN(n3943) );
  NAND2_X1 U3940 ( .A1(a_6_), .A2(n3942), .ZN(n3880) );
  NAND2_X1 U3941 ( .A1(n3947), .A2(n3948), .ZN(n3942) );
  NAND2_X1 U3942 ( .A1(n3877), .A2(n3949), .ZN(n3948) );
  NAND2_X1 U3943 ( .A1(n3876), .A2(n3875), .ZN(n3949) );
  NOR2_X1 U3944 ( .A1(n2286), .A2(n2132), .ZN(n3877) );
  OR2_X1 U3945 ( .A1(n3875), .A2(n3876), .ZN(n3947) );
  AND2_X1 U3946 ( .A1(n3821), .A2(n3950), .ZN(n3876) );
  NAND2_X1 U3947 ( .A1(n3820), .A2(n3822), .ZN(n3950) );
  NAND2_X1 U3948 ( .A1(n3951), .A2(n3952), .ZN(n3822) );
  NAND2_X1 U3949 ( .A1(b_2_), .A2(a_8_), .ZN(n3952) );
  INV_X1 U3950 ( .A(n3953), .ZN(n3951) );
  XOR2_X1 U3951 ( .A(n3954), .B(n3955), .Z(n3820) );
  XNOR2_X1 U3952 ( .A(n3956), .B(n3957), .ZN(n3955) );
  NAND2_X1 U3953 ( .A1(b_1_), .A2(a_9_), .ZN(n3954) );
  NAND2_X1 U3954 ( .A1(a_8_), .A2(n3953), .ZN(n3821) );
  NAND2_X1 U3955 ( .A1(n3958), .A2(n3959), .ZN(n3953) );
  NAND2_X1 U3956 ( .A1(n3872), .A2(n3960), .ZN(n3959) );
  OR2_X1 U3957 ( .A1(n3873), .A2(n3871), .ZN(n3960) );
  NOR2_X1 U3958 ( .A1(n2286), .A2(n2102), .ZN(n3872) );
  NAND2_X1 U3959 ( .A1(n3871), .A2(n3873), .ZN(n3958) );
  NAND2_X1 U3960 ( .A1(n3833), .A2(n3961), .ZN(n3873) );
  NAND2_X1 U3961 ( .A1(n3832), .A2(n3834), .ZN(n3961) );
  NAND2_X1 U3962 ( .A1(n3962), .A2(n3963), .ZN(n3834) );
  NAND2_X1 U3963 ( .A1(b_2_), .A2(a_10_), .ZN(n3963) );
  INV_X1 U3964 ( .A(n3964), .ZN(n3962) );
  XOR2_X1 U3965 ( .A(n3965), .B(n3966), .Z(n3832) );
  XNOR2_X1 U3966 ( .A(n3967), .B(n3968), .ZN(n3966) );
  NAND2_X1 U3967 ( .A1(b_1_), .A2(a_11_), .ZN(n3965) );
  NAND2_X1 U3968 ( .A1(a_10_), .A2(n3964), .ZN(n3833) );
  NAND2_X1 U3969 ( .A1(n3969), .A2(n3970), .ZN(n3964) );
  NAND2_X1 U3970 ( .A1(n3841), .A2(n3971), .ZN(n3970) );
  NAND2_X1 U3971 ( .A1(n3842), .A2(n3840), .ZN(n3971) );
  NOR2_X1 U3972 ( .A1(n2286), .A2(n2072), .ZN(n3841) );
  OR2_X1 U3973 ( .A1(n3840), .A2(n3842), .ZN(n3969) );
  AND2_X1 U3974 ( .A1(n3972), .A2(n3973), .ZN(n3842) );
  NAND2_X1 U3975 ( .A1(n3850), .A2(n3974), .ZN(n3973) );
  OR2_X1 U3976 ( .A1(n3847), .A2(n3849), .ZN(n3974) );
  NOR2_X1 U3977 ( .A1(n2286), .A2(n2277), .ZN(n3850) );
  NAND2_X1 U3978 ( .A1(n3847), .A2(n3849), .ZN(n3972) );
  NAND2_X1 U3979 ( .A1(n3975), .A2(n3976), .ZN(n3849) );
  NAND2_X1 U3980 ( .A1(n3977), .A2(b_2_), .ZN(n3976) );
  NOR2_X1 U3981 ( .A1(n3978), .A2(n2042), .ZN(n3977) );
  NOR2_X1 U3982 ( .A1(n3869), .A2(n3868), .ZN(n3978) );
  NAND2_X1 U3983 ( .A1(n3869), .A2(n3868), .ZN(n3975) );
  NAND2_X1 U3984 ( .A1(n3979), .A2(n3980), .ZN(n3868) );
  NAND2_X1 U3985 ( .A1(b_0_), .A2(n3981), .ZN(n3980) );
  NAND2_X1 U3986 ( .A1(n3982), .A2(n2018), .ZN(n3981) );
  NAND2_X1 U3987 ( .A1(a_15_), .A2(n3983), .ZN(n2018) );
  NAND2_X1 U3988 ( .A1(a_15_), .A2(n3864), .ZN(n3982) );
  NAND2_X1 U3989 ( .A1(b_1_), .A2(n3984), .ZN(n3979) );
  NAND2_X1 U3990 ( .A1(n3985), .A2(n2021), .ZN(n3984) );
  NAND2_X1 U3991 ( .A1(a_14_), .A2(n2009), .ZN(n2021) );
  NAND2_X1 U3992 ( .A1(a_14_), .A2(n2333), .ZN(n3985) );
  AND2_X1 U3993 ( .A1(n3986), .A2(n2558), .ZN(n3869) );
  NOR2_X1 U3994 ( .A1(n3864), .A2(n2286), .ZN(n3986) );
  XNOR2_X1 U3995 ( .A(n3987), .B(n3988), .ZN(n3847) );
  XOR2_X1 U3996 ( .A(n3989), .B(n3990), .Z(n3987) );
  XNOR2_X1 U3997 ( .A(n3991), .B(n3992), .ZN(n3840) );
  NOR2_X1 U3998 ( .A1(n2277), .A2(n3864), .ZN(n3992) );
  XOR2_X1 U3999 ( .A(n3993), .B(n3994), .Z(n3991) );
  XNOR2_X1 U4000 ( .A(n3995), .B(n3996), .ZN(n3871) );
  NAND2_X1 U4001 ( .A1(n3997), .A2(n3998), .ZN(n3995) );
  NAND2_X1 U4002 ( .A1(n3999), .A2(n4000), .ZN(n3998) );
  NAND2_X1 U4003 ( .A1(b_1_), .A2(a_10_), .ZN(n3999) );
  XOR2_X1 U4004 ( .A(n4001), .B(n4002), .Z(n3875) );
  NAND2_X1 U4005 ( .A1(n4003), .A2(n4004), .ZN(n4001) );
  NAND2_X1 U4006 ( .A1(n4005), .A2(n4006), .ZN(n4004) );
  NAND2_X1 U4007 ( .A1(b_1_), .A2(a_8_), .ZN(n4005) );
  XOR2_X1 U4008 ( .A(n4007), .B(n4008), .Z(n3883) );
  NAND2_X1 U4009 ( .A1(n4009), .A2(n4010), .ZN(n4007) );
  NAND2_X1 U4010 ( .A1(n4011), .A2(n4012), .ZN(n4010) );
  NAND2_X1 U4011 ( .A1(b_1_), .A2(a_6_), .ZN(n4011) );
  XOR2_X1 U4012 ( .A(n4013), .B(n4014), .Z(n3887) );
  NAND2_X1 U4013 ( .A1(n4015), .A2(n4016), .ZN(n4013) );
  NAND2_X1 U4014 ( .A1(n4017), .A2(n4018), .ZN(n4016) );
  NAND2_X1 U4015 ( .A1(b_1_), .A2(a_4_), .ZN(n4017) );
  INV_X1 U4016 ( .A(n2218), .ZN(n3893) );
  NAND2_X1 U4017 ( .A1(b_2_), .A2(a_2_), .ZN(n2218) );
  XNOR2_X1 U4018 ( .A(n3913), .B(n4019), .ZN(n3895) );
  NOR2_X1 U4019 ( .A1(n4020), .A2(n4021), .ZN(n4019) );
  INV_X1 U4020 ( .A(n3910), .ZN(n4021) );
  NAND2_X1 U4021 ( .A1(n4022), .A2(n3914), .ZN(n3910) );
  NOR2_X1 U4022 ( .A1(n3914), .A2(n4022), .ZN(n4020) );
  NOR2_X1 U4023 ( .A1(n2287), .A2(n3864), .ZN(n4022) );
  NOR2_X1 U4024 ( .A1(n2199), .A2(n2333), .ZN(n3914) );
  NAND2_X1 U4025 ( .A1(n4023), .A2(n4024), .ZN(n3913) );
  NAND2_X1 U4026 ( .A1(n4025), .A2(b_1_), .ZN(n4024) );
  NOR2_X1 U4027 ( .A1(n4026), .A2(n2199), .ZN(n4025) );
  NOR2_X1 U4028 ( .A1(n3923), .A2(n3924), .ZN(n4026) );
  NAND2_X1 U4029 ( .A1(n3923), .A2(n3924), .ZN(n4023) );
  NAND2_X1 U4030 ( .A1(n4015), .A2(n4027), .ZN(n3924) );
  NAND2_X1 U4031 ( .A1(n4028), .A2(n4014), .ZN(n4027) );
  NAND2_X1 U4032 ( .A1(n4029), .A2(n4030), .ZN(n4014) );
  NAND2_X1 U4033 ( .A1(n4031), .A2(b_1_), .ZN(n4030) );
  NOR2_X1 U4034 ( .A1(n4032), .A2(n2162), .ZN(n4031) );
  NOR2_X1 U4035 ( .A1(n3934), .A2(n3935), .ZN(n4032) );
  NAND2_X1 U4036 ( .A1(n3934), .A2(n3935), .ZN(n4029) );
  NAND2_X1 U4037 ( .A1(n4009), .A2(n4033), .ZN(n3935) );
  NAND2_X1 U4038 ( .A1(n4034), .A2(n4008), .ZN(n4033) );
  NAND2_X1 U4039 ( .A1(n4035), .A2(n4036), .ZN(n4008) );
  NAND2_X1 U4040 ( .A1(n4037), .A2(b_1_), .ZN(n4036) );
  NOR2_X1 U4041 ( .A1(n4038), .A2(n2132), .ZN(n4037) );
  NOR2_X1 U4042 ( .A1(n3945), .A2(n3946), .ZN(n4038) );
  NAND2_X1 U4043 ( .A1(n3945), .A2(n3946), .ZN(n4035) );
  NAND2_X1 U4044 ( .A1(n4003), .A2(n4039), .ZN(n3946) );
  NAND2_X1 U4045 ( .A1(n4040), .A2(n4002), .ZN(n4039) );
  NAND2_X1 U4046 ( .A1(n4041), .A2(n4042), .ZN(n4002) );
  NAND2_X1 U4047 ( .A1(n4043), .A2(b_1_), .ZN(n4042) );
  NOR2_X1 U4048 ( .A1(n4044), .A2(n2102), .ZN(n4043) );
  NOR2_X1 U4049 ( .A1(n3956), .A2(n3957), .ZN(n4044) );
  NAND2_X1 U4050 ( .A1(n3956), .A2(n3957), .ZN(n4041) );
  NAND2_X1 U4051 ( .A1(n3997), .A2(n4045), .ZN(n3957) );
  NAND2_X1 U4052 ( .A1(n4046), .A2(n3996), .ZN(n4045) );
  NAND2_X1 U4053 ( .A1(n4047), .A2(n4048), .ZN(n3996) );
  NAND2_X1 U4054 ( .A1(n4049), .A2(b_1_), .ZN(n4048) );
  NOR2_X1 U4055 ( .A1(n4050), .A2(n2072), .ZN(n4049) );
  NOR2_X1 U4056 ( .A1(n3967), .A2(n3968), .ZN(n4050) );
  NAND2_X1 U4057 ( .A1(n3967), .A2(n3968), .ZN(n4047) );
  NAND2_X1 U4058 ( .A1(n4051), .A2(n4052), .ZN(n3968) );
  NAND2_X1 U4059 ( .A1(n4053), .A2(b_1_), .ZN(n4052) );
  NOR2_X1 U4060 ( .A1(n4054), .A2(n2277), .ZN(n4053) );
  NOR2_X1 U4061 ( .A1(n3993), .A2(n3994), .ZN(n4054) );
  NAND2_X1 U4062 ( .A1(n3993), .A2(n3994), .ZN(n4051) );
  NAND2_X1 U4063 ( .A1(n3990), .A2(n4055), .ZN(n3994) );
  NAND2_X1 U4064 ( .A1(n3988), .A2(n3989), .ZN(n4055) );
  NOR2_X1 U4065 ( .A1(n3864), .A2(n2042), .ZN(n3989) );
  NOR2_X1 U4066 ( .A1(n2333), .A2(n3983), .ZN(n3988) );
  INV_X1 U4067 ( .A(a_14_), .ZN(n3983) );
  NAND2_X1 U4068 ( .A1(n4056), .A2(n2558), .ZN(n3990) );
  NOR2_X1 U4069 ( .A1(n2333), .A2(n3864), .ZN(n4056) );
  NOR2_X1 U4070 ( .A1(n2042), .A2(n2333), .ZN(n3993) );
  NOR2_X1 U4071 ( .A1(n2277), .A2(n2333), .ZN(n3967) );
  NAND2_X1 U4072 ( .A1(n4000), .A2(n2279), .ZN(n4046) );
  NAND2_X1 U4073 ( .A1(n4057), .A2(n4058), .ZN(n3997) );
  INV_X1 U4074 ( .A(n4000), .ZN(n4058) );
  NAND2_X1 U4075 ( .A1(a_11_), .A2(b_0_), .ZN(n4000) );
  NOR2_X1 U4076 ( .A1(n2279), .A2(n3864), .ZN(n4057) );
  NOR2_X1 U4077 ( .A1(n2279), .A2(n2333), .ZN(n3956) );
  INV_X1 U4078 ( .A(a_10_), .ZN(n2279) );
  NAND2_X1 U4079 ( .A1(n4006), .A2(n2281), .ZN(n4040) );
  NAND2_X1 U4080 ( .A1(n4059), .A2(n4060), .ZN(n4003) );
  INV_X1 U4081 ( .A(n4006), .ZN(n4060) );
  NAND2_X1 U4082 ( .A1(a_9_), .A2(b_0_), .ZN(n4006) );
  NOR2_X1 U4083 ( .A1(n2281), .A2(n3864), .ZN(n4059) );
  NOR2_X1 U4084 ( .A1(n2281), .A2(n2333), .ZN(n3945) );
  NAND2_X1 U4085 ( .A1(n4012), .A2(n2283), .ZN(n4034) );
  NAND2_X1 U4086 ( .A1(n4061), .A2(n4062), .ZN(n4009) );
  INV_X1 U4087 ( .A(n4012), .ZN(n4062) );
  NAND2_X1 U4088 ( .A1(a_7_), .A2(b_0_), .ZN(n4012) );
  NOR2_X1 U4089 ( .A1(n2283), .A2(n3864), .ZN(n4061) );
  NOR2_X1 U4090 ( .A1(n2283), .A2(n2333), .ZN(n3934) );
  NAND2_X1 U4091 ( .A1(n4018), .A2(n2285), .ZN(n4028) );
  NAND2_X1 U4092 ( .A1(n4063), .A2(n4064), .ZN(n4015) );
  INV_X1 U4093 ( .A(n4018), .ZN(n4064) );
  NAND2_X1 U4094 ( .A1(a_5_), .A2(b_0_), .ZN(n4018) );
  NOR2_X1 U4095 ( .A1(n2285), .A2(n3864), .ZN(n4063) );
  NOR2_X1 U4096 ( .A1(n2285), .A2(n2333), .ZN(n3923) );
  NAND2_X1 U4097 ( .A1(n4065), .A2(n4066), .ZN(n2010) );
  NAND2_X1 U4098 ( .A1(n4067), .A2(n2244), .ZN(n4066) );
  NAND2_X1 U4099 ( .A1(b_0_), .A2(n2376), .ZN(n2244) );
  INV_X1 U4100 ( .A(a_0_), .ZN(n2376) );
  NAND2_X1 U4101 ( .A1(n4068), .A2(n4069), .ZN(n4067) );
  NAND2_X1 U4102 ( .A1(a_1_), .A2(n3864), .ZN(n4069) );
  NAND2_X1 U4103 ( .A1(n4070), .A2(n4071), .ZN(n4068) );
  NAND2_X1 U4104 ( .A1(b_2_), .A2(n2287), .ZN(n4071) );
  INV_X1 U4105 ( .A(a_2_), .ZN(n2287) );
  NOR2_X1 U4106 ( .A1(n4072), .A2(n4073), .ZN(n4070) );
  NOR2_X1 U4107 ( .A1(a_1_), .A2(n3864), .ZN(n4073) );
  INV_X1 U4108 ( .A(b_1_), .ZN(n3864) );
  NOR2_X1 U4109 ( .A1(n4074), .A2(n4075), .ZN(n4072) );
  NAND2_X1 U4110 ( .A1(n4076), .A2(n4077), .ZN(n4075) );
  NAND2_X1 U4111 ( .A1(n4078), .A2(n4079), .ZN(n4077) );
  NAND2_X1 U4112 ( .A1(b_4_), .A2(n2285), .ZN(n4079) );
  INV_X1 U4113 ( .A(a_4_), .ZN(n2285) );
  NOR2_X1 U4114 ( .A1(n4080), .A2(n4081), .ZN(n4078) );
  NOR2_X1 U4115 ( .A1(a_3_), .A2(n2200), .ZN(n4081) );
  INV_X1 U4116 ( .A(b_3_), .ZN(n2200) );
  NOR2_X1 U4117 ( .A1(n4082), .A2(n4083), .ZN(n4080) );
  NAND2_X1 U4118 ( .A1(n4084), .A2(n4085), .ZN(n4083) );
  NAND2_X1 U4119 ( .A1(n4086), .A2(n4087), .ZN(n4085) );
  NAND2_X1 U4120 ( .A1(b_6_), .A2(n2283), .ZN(n4087) );
  INV_X1 U4121 ( .A(a_6_), .ZN(n2283) );
  NOR2_X1 U4122 ( .A1(n4088), .A2(n4089), .ZN(n4086) );
  NOR2_X1 U4123 ( .A1(a_5_), .A2(n2163), .ZN(n4089) );
  INV_X1 U4124 ( .A(b_5_), .ZN(n2163) );
  NOR2_X1 U4125 ( .A1(n4090), .A2(n4091), .ZN(n4088) );
  NAND2_X1 U4126 ( .A1(n4092), .A2(n4093), .ZN(n4091) );
  NAND2_X1 U4127 ( .A1(n4094), .A2(n4095), .ZN(n4093) );
  NAND2_X1 U4128 ( .A1(b_8_), .A2(n2281), .ZN(n4095) );
  INV_X1 U4129 ( .A(a_8_), .ZN(n2281) );
  NOR2_X1 U4130 ( .A1(n4096), .A2(n4097), .ZN(n4094) );
  NOR2_X1 U4131 ( .A1(a_7_), .A2(n2133), .ZN(n4097) );
  INV_X1 U4132 ( .A(b_7_), .ZN(n2133) );
  NOR2_X1 U4133 ( .A1(n4098), .A2(n4099), .ZN(n4096) );
  NAND2_X1 U4134 ( .A1(n4100), .A2(n4101), .ZN(n4099) );
  NAND2_X1 U4135 ( .A1(n4102), .A2(n4103), .ZN(n4101) );
  NAND2_X1 U4136 ( .A1(b_9_), .A2(n2102), .ZN(n4103) );
  NOR2_X1 U4137 ( .A1(n4104), .A2(n4105), .ZN(n4102) );
  NOR2_X1 U4138 ( .A1(a_10_), .A2(n2278), .ZN(n4105) );
  NOR2_X1 U4139 ( .A1(n4106), .A2(n4107), .ZN(n4104) );
  NAND2_X1 U4140 ( .A1(n4108), .A2(n4109), .ZN(n4107) );
  NAND2_X1 U4141 ( .A1(n4110), .A2(n4111), .ZN(n4109) );
  NAND2_X1 U4142 ( .A1(b_12_), .A2(n2277), .ZN(n4111) );
  INV_X1 U4143 ( .A(a_12_), .ZN(n2277) );
  NOR2_X1 U4144 ( .A1(n4112), .A2(n4113), .ZN(n4110) );
  NOR2_X1 U4145 ( .A1(a_11_), .A2(n2073), .ZN(n4113) );
  INV_X1 U4146 ( .A(b_11_), .ZN(n2073) );
  NOR2_X1 U4147 ( .A1(n4114), .A2(n4115), .ZN(n4112) );
  NAND2_X1 U4148 ( .A1(n4116), .A2(n4117), .ZN(n4115) );
  NAND2_X1 U4149 ( .A1(n4118), .A2(n4119), .ZN(n4117) );
  NOR2_X1 U4150 ( .A1(n4120), .A2(n4121), .ZN(n4119) );
  NOR2_X1 U4151 ( .A1(a_14_), .A2(n4122), .ZN(n4121) );
  NOR2_X1 U4152 ( .A1(b_15_), .A2(n2009), .ZN(n4122) );
  INV_X1 U4153 ( .A(a_15_), .ZN(n2009) );
  INV_X1 U4154 ( .A(n2275), .ZN(n4120) );
  NAND2_X1 U4155 ( .A1(b_15_), .A2(b_14_), .ZN(n2275) );
  NOR2_X1 U4156 ( .A1(n4123), .A2(n4124), .ZN(n4118) );
  NOR2_X1 U4157 ( .A1(a_13_), .A2(n2043), .ZN(n4124) );
  INV_X1 U4158 ( .A(b_13_), .ZN(n2043) );
  NOR2_X1 U4159 ( .A1(n2558), .A2(n2023), .ZN(n4123) );
  INV_X1 U4160 ( .A(b_14_), .ZN(n2023) );
  INV_X1 U4161 ( .A(n2274), .ZN(n2558) );
  NAND2_X1 U4162 ( .A1(a_14_), .A2(a_15_), .ZN(n2274) );
  NAND2_X1 U4163 ( .A1(a_12_), .A2(n2276), .ZN(n4116) );
  INV_X1 U4164 ( .A(b_12_), .ZN(n2276) );
  NOR2_X1 U4165 ( .A1(b_13_), .A2(n2042), .ZN(n4114) );
  INV_X1 U4166 ( .A(a_13_), .ZN(n2042) );
  NAND2_X1 U4167 ( .A1(a_10_), .A2(n2278), .ZN(n4108) );
  INV_X1 U4168 ( .A(b_10_), .ZN(n2278) );
  NOR2_X1 U4169 ( .A1(b_11_), .A2(n2072), .ZN(n4106) );
  INV_X1 U4170 ( .A(a_11_), .ZN(n2072) );
  NAND2_X1 U4171 ( .A1(a_8_), .A2(n2280), .ZN(n4100) );
  INV_X1 U4172 ( .A(b_8_), .ZN(n2280) );
  NOR2_X1 U4173 ( .A1(b_9_), .A2(n2102), .ZN(n4098) );
  INV_X1 U4174 ( .A(a_9_), .ZN(n2102) );
  NAND2_X1 U4175 ( .A1(a_6_), .A2(n2282), .ZN(n4092) );
  INV_X1 U4176 ( .A(b_6_), .ZN(n2282) );
  NOR2_X1 U4177 ( .A1(b_7_), .A2(n2132), .ZN(n4090) );
  INV_X1 U4178 ( .A(a_7_), .ZN(n2132) );
  NAND2_X1 U4179 ( .A1(a_4_), .A2(n2284), .ZN(n4084) );
  INV_X1 U4180 ( .A(b_4_), .ZN(n2284) );
  NOR2_X1 U4181 ( .A1(b_5_), .A2(n2162), .ZN(n4082) );
  INV_X1 U4182 ( .A(a_5_), .ZN(n2162) );
  NAND2_X1 U4183 ( .A1(a_2_), .A2(n2286), .ZN(n4076) );
  INV_X1 U4184 ( .A(b_2_), .ZN(n2286) );
  NOR2_X1 U4185 ( .A1(b_3_), .A2(n2199), .ZN(n4074) );
  INV_X1 U4186 ( .A(a_3_), .ZN(n2199) );
  NAND2_X1 U4187 ( .A1(a_0_), .A2(n2333), .ZN(n4065) );
  INV_X1 U4188 ( .A(b_0_), .ZN(n2333) );
endmodule

