module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n556_, new_n456_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n418_, new_n292_, new_n215_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n314_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n570_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n407_, new_n480_, new_n151_, new_n513_, new_n558_, new_n231_, new_n382_, new_n239_, new_n522_, new_n199_, new_n487_, new_n360_, new_n546_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n440_, new_n531_, new_n252_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n412_, new_n327_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n226_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

nand g000 ( new_n151_, N29, N42, N75 );
xor g001 ( N388, new_n151_, keyIn_0_3 );
nand g002 ( new_n153_, N29, N36, N80 );
not g003 ( N389, new_n153_ );
nand g004 ( new_n155_, N29, N36, N42 );
xnor g005 ( N390, new_n155_, keyIn_0_4 );
nand g006 ( new_n157_, N85, N86 );
not g007 ( N391, new_n157_ );
nand g008 ( new_n159_, N1, N8 );
not g009 ( new_n160_, new_n159_ );
nand g010 ( new_n161_, new_n160_, N13, N17 );
xnor g011 ( N418, new_n161_, keyIn_0_0 );
xor g012 ( new_n163_, new_n155_, keyIn_0_1 );
not g013 ( new_n164_, new_n163_ );
nand g014 ( new_n165_, N1, N26 );
nand g015 ( new_n166_, N13, N17 );
nor g016 ( new_n167_, new_n165_, new_n166_ );
nand g017 ( N419, new_n164_, new_n167_ );
nand g018 ( N420, N59, N75, N80 );
nand g019 ( N421, N36, N59, N80 );
nand g020 ( new_n171_, N36, N42, N59 );
xor g021 ( N422, new_n171_, keyIn_0_5 );
not g022 ( new_n173_, N90 );
nor g023 ( new_n174_, N87, N88 );
nor g024 ( N423, new_n174_, new_n173_ );
nand g025 ( N446, new_n163_, new_n167_ );
nand g026 ( new_n177_, keyIn_0_2, N1, N26, N51 );
not g027 ( new_n178_, keyIn_0_2 );
nand g028 ( new_n179_, N1, N26, N51 );
nand g029 ( new_n180_, new_n179_, new_n178_ );
nand g030 ( new_n181_, new_n180_, new_n177_ );
not g031 ( N447, new_n181_ );
nand g032 ( new_n183_, new_n160_, N13, N55 );
nand g033 ( new_n184_, N29, N68 );
nor g034 ( N448, new_n183_, new_n184_ );
not g035 ( new_n186_, new_n183_ );
nand g036 ( new_n187_, N59, N68 );
not g037 ( new_n188_, new_n187_ );
nand g038 ( new_n189_, new_n186_, N74, new_n188_ );
xor g039 ( N449, new_n189_, keyIn_0_12 );
not g040 ( new_n191_, N89 );
nor g041 ( new_n192_, new_n174_, new_n191_ );
xnor g042 ( N450, new_n192_, keyIn_0_9 );
not g043 ( new_n194_, keyIn_0_19 );
not g044 ( new_n195_, N135 );
nor g045 ( new_n196_, N111, N116 );
xnor g046 ( new_n197_, new_n196_, keyIn_0_6 );
nand g047 ( new_n198_, N111, N116 );
nand g048 ( new_n199_, new_n197_, new_n198_ );
xor g049 ( new_n200_, N121, N126 );
xnor g050 ( new_n201_, new_n199_, new_n200_ );
not g051 ( new_n202_, new_n201_ );
nand g052 ( new_n203_, new_n202_, new_n194_, new_n195_ );
nand g053 ( new_n204_, new_n202_, new_n195_ );
nand g054 ( new_n205_, new_n204_, keyIn_0_19 );
nand g055 ( new_n206_, new_n201_, N135 );
xnor g056 ( new_n207_, N91, N96 );
xnor g057 ( new_n208_, N101, N106 );
xnor g058 ( new_n209_, new_n207_, new_n208_ );
xnor g059 ( new_n210_, new_n209_, N130 );
nand g060 ( new_n211_, new_n205_, new_n203_, new_n206_, new_n210_ );
nand g061 ( new_n212_, new_n211_, keyIn_0_32 );
not g062 ( new_n213_, new_n212_ );
nor g063 ( new_n214_, new_n211_, keyIn_0_32 );
nand g064 ( new_n215_, new_n205_, new_n203_, new_n206_ );
not g065 ( new_n216_, new_n210_ );
nand g066 ( new_n217_, new_n215_, new_n216_ );
not g067 ( new_n218_, new_n217_ );
nor g068 ( N767, new_n213_, new_n218_, new_n214_ );
not g069 ( new_n220_, N207 );
xnor g070 ( new_n221_, N183, N189 );
xnor g071 ( new_n222_, N195, N201 );
xnor g072 ( new_n223_, new_n221_, new_n222_ );
nand g073 ( new_n224_, new_n223_, new_n220_ );
xor g074 ( new_n225_, new_n224_, keyIn_0_26 );
not g075 ( new_n226_, new_n223_ );
nand g076 ( new_n227_, new_n226_, N207 );
nand g077 ( new_n228_, new_n225_, new_n227_ );
not g078 ( new_n229_, keyIn_0_25 );
not g079 ( new_n230_, N130 );
not g080 ( new_n231_, keyIn_0_13 );
not g081 ( new_n232_, N159 );
not g082 ( new_n233_, N165 );
nand g083 ( new_n234_, new_n232_, new_n233_ );
nand g084 ( new_n235_, N159, N165 );
nand g085 ( new_n236_, new_n234_, new_n231_, new_n235_ );
xor g086 ( new_n237_, N171, N177 );
xor g087 ( new_n238_, new_n237_, new_n236_ );
nand g088 ( new_n239_, new_n238_, new_n229_, new_n230_ );
nand g089 ( new_n240_, new_n238_, new_n230_ );
nand g090 ( new_n241_, new_n240_, keyIn_0_25 );
not g091 ( new_n242_, new_n238_ );
nand g092 ( new_n243_, new_n242_, N130 );
nand g093 ( new_n244_, new_n241_, new_n243_, keyIn_0_31, new_n239_ );
xor g094 ( N768, new_n228_, new_n244_ );
not g095 ( new_n246_, keyIn_0_52 );
not g096 ( new_n247_, keyIn_0_24 );
nand g097 ( new_n248_, N17, N42 );
nor g098 ( new_n249_, N17, N42 );
nand g099 ( new_n250_, N59, N156 );
nor g100 ( new_n251_, new_n249_, new_n250_ );
nand g101 ( new_n252_, new_n251_, new_n180_, new_n177_, new_n248_ );
nand g102 ( new_n253_, N42, N59, N75 );
nand g103 ( new_n254_, new_n160_, N17, N51, new_n253_ );
nand g104 ( new_n255_, new_n252_, new_n254_ );
nand g105 ( new_n256_, new_n255_, new_n247_, N126 );
nand g106 ( new_n257_, new_n255_, N126 );
nand g107 ( new_n258_, new_n257_, keyIn_0_24 );
nand g108 ( new_n259_, new_n258_, new_n256_ );
not g109 ( new_n260_, keyIn_0_15 );
nand g110 ( new_n261_, N29, N55, N75, N80 );
not g111 ( new_n262_, new_n261_ );
nand g112 ( new_n263_, new_n262_, new_n180_, new_n177_ );
nand g113 ( new_n264_, new_n263_, new_n260_ );
nand g114 ( new_n265_, new_n262_, new_n180_, keyIn_0_15, new_n177_ );
nand g115 ( new_n266_, new_n264_, new_n265_ );
xor g116 ( new_n267_, keyIn_0_10, N268 );
nand g117 ( new_n268_, new_n266_, new_n267_ );
nand g118 ( new_n269_, new_n180_, N17, new_n177_, new_n250_ );
nand g119 ( new_n270_, new_n269_, N1 );
nand g120 ( new_n271_, new_n270_, N153 );
nand g121 ( new_n272_, new_n259_, new_n268_, new_n271_ );
nand g122 ( new_n273_, new_n272_, keyIn_0_37, N201 );
not g123 ( new_n274_, keyIn_0_37 );
nand g124 ( new_n275_, new_n272_, N201 );
nand g125 ( new_n276_, new_n275_, new_n274_ );
nand g126 ( new_n277_, new_n276_, new_n273_ );
not g127 ( new_n278_, new_n277_ );
not g128 ( new_n279_, keyIn_0_38 );
not g129 ( new_n280_, N201 );
nand g130 ( new_n281_, new_n259_, new_n280_, new_n268_, new_n271_ );
xnor g131 ( new_n282_, new_n281_, new_n279_ );
nand g132 ( new_n283_, new_n278_, new_n282_ );
xnor g133 ( new_n284_, new_n283_, N261 );
nand g134 ( new_n285_, new_n284_, new_n246_ );
not g135 ( new_n286_, new_n284_ );
nand g136 ( new_n287_, new_n286_, keyIn_0_52 );
nand g137 ( new_n288_, new_n287_, N219, new_n285_ );
nand g138 ( new_n289_, N121, N210 );
nand g139 ( new_n290_, new_n288_, new_n289_ );
xnor g140 ( new_n291_, new_n290_, keyIn_0_56 );
nand g141 ( new_n292_, new_n186_, N42, N72, new_n188_ );
not g142 ( new_n293_, new_n292_ );
nand g143 ( new_n294_, new_n293_, keyIn_0_8 );
not g144 ( new_n295_, keyIn_0_8 );
nand g145 ( new_n296_, new_n292_, new_n295_ );
nand g146 ( new_n297_, new_n294_, N73, new_n296_ );
xnor g147 ( new_n298_, new_n297_, keyIn_0_11 );
xnor g148 ( new_n299_, new_n298_, keyIn_0_14 );
xnor g149 ( new_n300_, new_n299_, keyIn_0_16 );
nand g150 ( new_n301_, new_n300_, N201 );
xor g151 ( new_n302_, new_n301_, keyIn_0_28 );
nand g152 ( new_n303_, new_n277_, N237 );
nand g153 ( new_n304_, new_n303_, keyIn_0_50 );
nand g154 ( new_n305_, new_n272_, N246 );
nand g155 ( new_n306_, N255, N267 );
nand g156 ( new_n307_, new_n304_, new_n305_, new_n306_ );
not g157 ( new_n308_, keyIn_0_50 );
nand g158 ( new_n309_, new_n277_, new_n308_, N237 );
nand g159 ( new_n310_, new_n278_, N228, new_n282_ );
nand g160 ( new_n311_, new_n310_, new_n309_ );
nor g161 ( new_n312_, new_n302_, new_n307_, new_n311_ );
nand g162 ( N850, new_n291_, new_n312_ );
not g163 ( new_n314_, keyIn_0_51 );
not g164 ( new_n315_, N189 );
nand g165 ( new_n316_, new_n270_, N146 );
nand g166 ( new_n317_, new_n255_, keyIn_0_23, N116 );
not g167 ( new_n318_, keyIn_0_23 );
nand g168 ( new_n319_, new_n255_, N116 );
nand g169 ( new_n320_, new_n319_, new_n318_ );
nand g170 ( new_n321_, new_n320_, new_n268_, new_n316_, new_n317_ );
xnor g171 ( new_n322_, new_n321_, keyIn_0_30 );
nand g172 ( new_n323_, new_n322_, new_n315_ );
not g173 ( new_n324_, N195 );
nand g174 ( new_n325_, new_n270_, N149 );
nand g175 ( new_n326_, new_n255_, N121 );
nand g176 ( new_n327_, new_n268_, new_n324_, new_n325_, new_n326_ );
nand g177 ( new_n328_, new_n277_, new_n323_, new_n327_ );
nand g178 ( new_n329_, new_n328_, new_n314_ );
nand g179 ( new_n330_, new_n277_, new_n323_, keyIn_0_51, new_n327_ );
nand g180 ( new_n331_, new_n329_, new_n330_ );
not g181 ( new_n332_, keyIn_0_42 );
nand g182 ( new_n333_, new_n282_, N261 );
not g183 ( new_n334_, new_n333_ );
nand g184 ( new_n335_, new_n334_, new_n332_, new_n323_, new_n327_ );
nand g185 ( new_n336_, new_n282_, new_n323_, N261, new_n327_ );
nand g186 ( new_n337_, new_n336_, keyIn_0_42 );
nand g187 ( new_n338_, new_n268_, new_n325_, new_n326_ );
nand g188 ( new_n339_, new_n338_, N195 );
not g189 ( new_n340_, new_n339_ );
nand g190 ( new_n341_, new_n323_, new_n340_ );
not g191 ( new_n342_, new_n322_ );
nand g192 ( new_n343_, new_n342_, N189 );
nand g193 ( new_n344_, new_n341_, new_n343_ );
not g194 ( new_n345_, new_n344_ );
nand g195 ( new_n346_, new_n331_, new_n335_, new_n337_, new_n345_ );
not g196 ( new_n347_, new_n346_ );
not g197 ( new_n348_, keyIn_0_29 );
not g198 ( new_n349_, keyIn_0_22 );
nand g199 ( new_n350_, new_n255_, N111 );
nand g200 ( new_n351_, new_n350_, new_n349_ );
nand g201 ( new_n352_, new_n255_, keyIn_0_22, N111 );
nand g202 ( new_n353_, new_n351_, new_n352_ );
nand g203 ( new_n354_, new_n270_, N143 );
nand g204 ( new_n355_, new_n353_, new_n268_, new_n354_ );
nand g205 ( new_n356_, new_n355_, new_n348_ );
nand g206 ( new_n357_, new_n353_, keyIn_0_29, new_n268_, new_n354_ );
nand g207 ( new_n358_, new_n356_, new_n357_ );
nand g208 ( new_n359_, new_n358_, keyIn_0_36, N183 );
not g209 ( new_n360_, keyIn_0_36 );
nand g210 ( new_n361_, new_n358_, N183 );
nand g211 ( new_n362_, new_n361_, new_n360_ );
nand g212 ( new_n363_, new_n362_, new_n359_ );
not g213 ( new_n364_, N183 );
nand g214 ( new_n365_, new_n356_, new_n364_, new_n357_ );
nand g215 ( new_n366_, new_n363_, new_n365_ );
nor g216 ( new_n367_, new_n347_, new_n366_ );
nand g217 ( new_n368_, new_n367_, keyIn_0_53 );
not g218 ( new_n369_, keyIn_0_53 );
not g219 ( new_n370_, new_n367_ );
nand g220 ( new_n371_, new_n370_, new_n369_ );
nand g221 ( new_n372_, new_n347_, new_n366_ );
nand g222 ( new_n373_, new_n371_, keyIn_0_55, new_n368_, new_n372_ );
not g223 ( new_n374_, keyIn_0_55 );
nand g224 ( new_n375_, new_n371_, new_n368_, new_n372_ );
nand g225 ( new_n376_, new_n375_, new_n374_ );
nand g226 ( new_n377_, new_n376_, N219, new_n373_ );
not g227 ( new_n378_, keyIn_0_47 );
not g228 ( new_n379_, new_n366_ );
nand g229 ( new_n380_, new_n379_, N228 );
nand g230 ( new_n381_, new_n380_, new_n378_ );
nand g231 ( new_n382_, new_n300_, N183 );
xnor g232 ( new_n383_, new_n382_, keyIn_0_27 );
nand g233 ( new_n384_, new_n358_, N246 );
nand g234 ( new_n385_, N106, N210 );
nand g235 ( new_n386_, new_n383_, new_n381_, new_n384_, new_n385_ );
not g236 ( new_n387_, new_n386_ );
not g237 ( new_n388_, keyIn_0_40 );
nand g238 ( new_n389_, new_n362_, new_n388_, new_n359_ );
nand g239 ( new_n390_, new_n363_, keyIn_0_40 );
nand g240 ( new_n391_, new_n390_, N237, new_n389_ );
nand g241 ( new_n392_, new_n379_, keyIn_0_47, N228 );
nand g242 ( N863, new_n377_, new_n387_, new_n391_, new_n392_ );
nor g243 ( new_n394_, new_n334_, new_n277_ );
not g244 ( new_n395_, new_n394_ );
nand g245 ( new_n396_, new_n395_, new_n327_ );
xnor g246 ( new_n397_, new_n339_, keyIn_0_49 );
nand g247 ( new_n398_, new_n396_, new_n397_ );
nand g248 ( new_n399_, new_n343_, new_n323_ );
not g249 ( new_n400_, new_n399_ );
nand g250 ( new_n401_, new_n398_, new_n400_ );
nand g251 ( new_n402_, new_n396_, new_n397_, new_n399_ );
nand g252 ( new_n403_, new_n401_, N219, new_n402_ );
nand g253 ( new_n404_, new_n342_, N189, N237 );
nand g254 ( new_n405_, new_n300_, N189 );
nand g255 ( new_n406_, N111, N210 );
nand g256 ( new_n407_, new_n405_, new_n404_, new_n406_ );
nand g257 ( new_n408_, new_n342_, N246 );
nand g258 ( new_n409_, N255, N259 );
nand g259 ( new_n410_, new_n408_, new_n409_ );
xor g260 ( new_n411_, new_n410_, keyIn_0_41 );
nor g261 ( new_n412_, new_n407_, new_n411_ );
nand g262 ( new_n413_, new_n400_, N228 );
xnor g263 ( new_n414_, new_n413_, keyIn_0_48 );
nand g264 ( N864, new_n403_, new_n412_, new_n414_ );
nand g265 ( new_n416_, new_n395_, new_n327_, new_n339_ );
nand g266 ( new_n417_, new_n339_, new_n327_ );
nand g267 ( new_n418_, new_n394_, new_n417_ );
nand g268 ( new_n419_, new_n416_, N219, new_n418_ );
nand g269 ( new_n420_, new_n300_, N195 );
nand g270 ( new_n421_, new_n339_, N228, new_n327_ );
nand g271 ( new_n422_, new_n340_, N237 );
nand g272 ( new_n423_, new_n338_, N246 );
nand g273 ( new_n424_, N255, N260 );
nand g274 ( new_n425_, N116, N210 );
nand g275 ( new_n426_, new_n422_, new_n423_, new_n424_, new_n425_ );
not g276 ( new_n427_, new_n426_ );
nand g277 ( N865, new_n419_, new_n420_, new_n421_, new_n427_ );
not g278 ( new_n429_, keyIn_0_54 );
nand g279 ( new_n430_, new_n346_, new_n365_ );
nand g280 ( new_n431_, new_n390_, keyIn_0_46, new_n389_ );
not g281 ( new_n432_, keyIn_0_46 );
nand g282 ( new_n433_, new_n390_, new_n389_ );
nand g283 ( new_n434_, new_n433_, new_n432_ );
nand g284 ( new_n435_, new_n430_, new_n429_, new_n431_, new_n434_ );
nand g285 ( new_n436_, new_n430_, new_n431_, new_n434_ );
nand g286 ( new_n437_, new_n436_, keyIn_0_54 );
nand g287 ( new_n438_, new_n437_, new_n435_ );
not g288 ( new_n439_, N177 );
nand g289 ( new_n440_, N29, N75, N80 );
nor g290 ( new_n441_, new_n440_, N268 );
nand g291 ( new_n442_, N447, N17, new_n441_ );
xnor g292 ( new_n443_, new_n442_, keyIn_0_18 );
not g293 ( new_n444_, new_n443_ );
nand g294 ( new_n445_, new_n255_, N106 );
nand g295 ( new_n446_, new_n250_, N55 );
nor g296 ( new_n447_, new_n181_, new_n446_ );
nand g297 ( new_n448_, new_n447_, N153 );
nand g298 ( new_n449_, N138, N152 );
nand g299 ( new_n450_, new_n444_, new_n445_, new_n448_, new_n449_ );
not g300 ( new_n451_, new_n450_ );
nand g301 ( new_n452_, new_n451_, new_n439_ );
nand g302 ( new_n453_, new_n438_, new_n452_ );
nand g303 ( new_n454_, new_n450_, N177 );
nand g304 ( new_n455_, new_n453_, new_n454_ );
not g305 ( new_n456_, N171 );
nand g306 ( new_n457_, new_n447_, N149 );
xnor g307 ( new_n458_, new_n457_, keyIn_0_17 );
nand g308 ( new_n459_, new_n255_, N101 );
nand g309 ( new_n460_, N17, N138 );
nand g310 ( new_n461_, new_n459_, new_n442_, new_n460_ );
nor g311 ( new_n462_, new_n458_, new_n461_ );
nand g312 ( new_n463_, new_n462_, new_n456_ );
nand g313 ( new_n464_, new_n455_, new_n463_ );
not g314 ( new_n465_, new_n462_ );
nand g315 ( new_n466_, new_n465_, N171 );
xnor g316 ( new_n467_, new_n466_, keyIn_0_35 );
nand g317 ( new_n468_, new_n464_, new_n467_ );
nand g318 ( new_n469_, new_n447_, N146 );
nand g319 ( new_n470_, new_n469_, new_n442_, keyIn_0_21 );
not g320 ( new_n471_, keyIn_0_21 );
nand g321 ( new_n472_, new_n469_, new_n442_ );
nand g322 ( new_n473_, new_n472_, new_n471_ );
nand g323 ( new_n474_, new_n255_, N96 );
nand g324 ( new_n475_, N51, N138 );
nand g325 ( new_n476_, new_n473_, new_n470_, new_n474_, new_n475_ );
nor g326 ( new_n477_, new_n476_, N165 );
not g327 ( new_n478_, new_n477_ );
nand g328 ( new_n479_, new_n468_, new_n478_ );
nand g329 ( new_n480_, new_n476_, N165 );
nand g330 ( new_n481_, new_n479_, new_n480_ );
not g331 ( new_n482_, keyIn_0_20 );
nand g332 ( new_n483_, new_n447_, N143 );
nand g333 ( new_n484_, new_n483_, new_n442_, new_n482_ );
nand g334 ( new_n485_, new_n483_, new_n442_ );
nand g335 ( new_n486_, new_n485_, keyIn_0_20 );
nand g336 ( new_n487_, new_n255_, N91 );
nand g337 ( new_n488_, N8, N138 );
nand g338 ( new_n489_, new_n486_, new_n484_, new_n487_, new_n488_ );
nor g339 ( new_n490_, new_n489_, N159 );
xnor g340 ( new_n491_, new_n490_, keyIn_0_33 );
not g341 ( new_n492_, new_n491_ );
nand g342 ( new_n493_, new_n481_, new_n492_ );
nand g343 ( new_n494_, new_n489_, N159 );
xnor g344 ( new_n495_, new_n494_, keyIn_0_43 );
nand g345 ( new_n496_, new_n493_, new_n495_ );
xnor g346 ( N866, new_n496_, keyIn_0_59 );
not g347 ( new_n498_, new_n438_ );
nand g348 ( new_n499_, new_n452_, new_n454_ );
nand g349 ( new_n500_, new_n498_, keyIn_0_57, new_n499_ );
not g350 ( new_n501_, keyIn_0_57 );
nand g351 ( new_n502_, new_n498_, new_n499_ );
nand g352 ( new_n503_, new_n502_, new_n501_ );
not g353 ( new_n504_, new_n499_ );
nand g354 ( new_n505_, new_n438_, new_n504_ );
nand g355 ( new_n506_, new_n503_, N219, new_n500_, new_n505_ );
nand g356 ( new_n507_, new_n300_, N177 );
nand g357 ( new_n508_, new_n504_, N228 );
nand g358 ( new_n509_, new_n450_, N177, N237 );
nand g359 ( new_n510_, new_n450_, N246 );
nand g360 ( new_n511_, N101, N210 );
nand g361 ( new_n512_, new_n509_, new_n510_, new_n511_ );
not g362 ( new_n513_, new_n512_ );
nand g363 ( new_n514_, new_n506_, new_n507_, new_n508_, new_n513_ );
xor g364 ( N874, new_n514_, keyIn_0_62 );
not g365 ( new_n516_, new_n494_ );
nor g366 ( new_n517_, new_n491_, new_n516_ );
nand g367 ( new_n518_, new_n481_, new_n517_ );
not g368 ( new_n519_, new_n517_ );
nand g369 ( new_n520_, new_n479_, new_n480_, new_n519_ );
nand g370 ( new_n521_, new_n518_, N219, new_n520_ );
nand g371 ( new_n522_, new_n300_, N159 );
nand g372 ( new_n523_, new_n489_, N246 );
xor g373 ( new_n524_, new_n523_, keyIn_0_34 );
nand g374 ( new_n525_, new_n522_, new_n524_ );
xor g375 ( new_n526_, new_n525_, keyIn_0_39 );
nand g376 ( new_n527_, new_n517_, N228 );
nand g377 ( new_n528_, new_n516_, N237 );
not g378 ( new_n529_, new_n267_ );
nand g379 ( new_n530_, new_n529_, N210 );
nand g380 ( new_n531_, new_n527_, new_n528_, new_n530_ );
not g381 ( new_n532_, new_n531_ );
nand g382 ( N878, new_n521_, new_n526_, new_n532_ );
not g383 ( new_n534_, keyIn_0_60 );
not g384 ( new_n535_, keyIn_0_58 );
xnor g385 ( new_n536_, new_n467_, keyIn_0_44 );
not g386 ( new_n537_, new_n480_ );
nor g387 ( new_n538_, new_n537_, new_n477_ );
not g388 ( new_n539_, new_n538_ );
nand g389 ( new_n540_, new_n464_, new_n535_, new_n536_, new_n539_ );
nand g390 ( new_n541_, new_n464_, new_n536_, new_n539_ );
nand g391 ( new_n542_, new_n541_, keyIn_0_58 );
nand g392 ( new_n543_, new_n542_, new_n540_ );
nand g393 ( new_n544_, new_n464_, new_n536_ );
nand g394 ( new_n545_, new_n544_, new_n538_ );
nand g395 ( new_n546_, new_n543_, N219, new_n545_ );
nand g396 ( new_n547_, N91, N210 );
xor g397 ( new_n548_, new_n547_, keyIn_0_7 );
nand g398 ( new_n549_, new_n546_, new_n548_ );
nand g399 ( new_n550_, new_n549_, new_n534_ );
nand g400 ( new_n551_, new_n546_, keyIn_0_60, new_n548_ );
nand g401 ( new_n552_, new_n550_, new_n551_ );
nand g402 ( new_n553_, new_n300_, N165 );
nand g403 ( new_n554_, new_n538_, N228 );
nand g404 ( new_n555_, new_n537_, N237 );
nand g405 ( new_n556_, new_n476_, N246 );
nand g406 ( new_n557_, new_n553_, new_n554_, new_n555_, new_n556_ );
not g407 ( new_n558_, new_n557_ );
nand g408 ( N879, new_n552_, new_n558_ );
not g409 ( new_n560_, keyIn_0_63 );
nand g410 ( new_n561_, new_n467_, new_n463_ );
not g411 ( new_n562_, new_n561_ );
nand g412 ( new_n563_, new_n455_, new_n562_ );
nand g413 ( new_n564_, new_n453_, new_n454_, new_n561_ );
nand g414 ( new_n565_, new_n563_, N219, new_n564_ );
nand g415 ( new_n566_, N96, N210 );
nand g416 ( new_n567_, new_n565_, new_n566_ );
xor g417 ( new_n568_, new_n567_, keyIn_0_61 );
not g418 ( new_n569_, new_n467_ );
nand g419 ( new_n570_, new_n569_, N237 );
xor g420 ( new_n571_, new_n570_, keyIn_0_45 );
nand g421 ( new_n572_, new_n300_, N171 );
nand g422 ( new_n573_, new_n562_, N228 );
nand g423 ( new_n574_, new_n465_, N246 );
nand g424 ( new_n575_, new_n572_, new_n573_, new_n574_ );
nor g425 ( new_n576_, new_n571_, new_n575_ );
nand g426 ( new_n577_, new_n568_, new_n560_, new_n576_ );
nand g427 ( new_n578_, new_n568_, new_n576_ );
nand g428 ( new_n579_, new_n578_, keyIn_0_63 );
nand g429 ( N880, new_n579_, new_n577_ );
endmodule