module top ( G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, keyinput0_G223gat, keyinput1_G223gat, keyinput2_G223gat, keyinput3_G223gat, keyinput0_G329gat, keyinput1_G329gat, keyinput2_G329gat, keyinput3_G329gat, keyinput0_G370gat, keyinput1_G370gat, keyinput2_G370gat, keyinput3_G370gat, keyinput0_G421gat, keyinput1_G421gat, keyinput2_G421gat, keyinput3_G421gat, keyinput0_G430gat, keyinput1_G430gat, keyinput2_G430gat, keyinput3_G430gat, keyinput0_G431gat, keyinput1_G431gat, keyinput2_G431gat, keyinput3_G431gat, keyinput0_G432gat, keyinput1_G432gat, keyinput2_G432gat, keyinput3_G432gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat );
input G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, keyinput0_G223gat, keyinput1_G223gat, keyinput2_G223gat, keyinput3_G223gat, keyinput0_G329gat, keyinput1_G329gat, keyinput2_G329gat, keyinput3_G329gat, keyinput0_G370gat, keyinput1_G370gat, keyinput2_G370gat, keyinput3_G370gat, keyinput0_G421gat, keyinput1_G421gat, keyinput2_G421gat, keyinput3_G421gat, keyinput0_G430gat, keyinput1_G430gat, keyinput2_G430gat, keyinput3_G430gat, keyinput0_G431gat, keyinput1_G431gat, keyinput2_G431gat, keyinput3_G431gat, keyinput0_G432gat, keyinput1_G432gat, keyinput2_G432gat, keyinput3_G432gat;
output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
wire new_n1668_, new_n595_, new_n2051_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n1743_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1988_, new_n1433_, new_n2260_, new_n1517_, new_n1472_, new_n1785_, new_n439_, new_n1532_, new_n223_, new_n743_, new_n1962_, new_n1327_, new_n241_, new_n1535_, new_n2041_, new_n641_, new_n339_, new_n1849_, new_n389_, new_n514_, new_n1865_, new_n2431_, new_n1351_, new_n636_, new_n691_, new_n1024_, new_n2291_, new_n911_, new_n679_, new_n937_, new_n1879_, new_n173_, new_n2054_, new_n728_, new_n1071_, new_n2114_, new_n1294_, new_n214_, new_n853_, new_n695_, new_n660_, new_n2038_, new_n1311_, new_n2424_, new_n552_, new_n342_, new_n1662_, new_n706_, new_n2132_, new_n2063_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n1769_, new_n317_, new_n2107_, new_n1188_, new_n2231_, new_n2264_, new_n2244_, new_n504_, new_n1414_, new_n234_, new_n873_, new_n1300_, new_n2135_, new_n1898_, new_n774_, new_n1777_, new_n2176_, new_n1620_, new_n1786_, new_n1946_, new_n1580_, new_n766_, new_n1973_, new_n2387_, new_n2421_, new_n1262_, new_n1212_, new_n2452_, new_n1332_, new_n1447_, new_n2293_, new_n685_, new_n326_, new_n2348_, new_n903_, new_n1595_, new_n2468_, new_n822_, new_n1760_, new_n1018_, new_n1884_, new_n1864_, new_n1054_, new_n1288_, new_n385_, new_n1049_, new_n1330_, new_n2318_, new_n461_, new_n2171_, new_n2369_, new_n1323_, new_n297_, new_n150_, new_n1196_, new_n1366_, new_n137_, new_n2104_, new_n303_, new_n2334_, new_n2251_, new_n325_, new_n1285_, new_n1733_, new_n1842_, new_n1216_, new_n1632_, new_n1889_, new_n1987_, new_n629_, new_n2320_, new_n1214_, new_n883_, new_n1647_, new_n960_, new_n2433_, new_n1377_, new_n1522_, new_n549_, new_n2248_, new_n995_, new_n1035_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n2072_, new_n1678_, new_n568_, new_n1950_, new_n1936_, new_n423_, new_n496_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n85_, new_n912_, new_n1424_, new_n2350_, new_n680_, new_n981_, new_n2102_, new_n2337_, new_n1527_, new_n1275_, new_n1800_, new_n1198_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n2414_, new_n2397_, new_n194_, new_n2012_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n2184_, new_n142_, new_n2155_, new_n657_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n165_, new_n785_, new_n1501_, new_n477_, new_n664_, new_n280_, new_n1041_, new_n1989_, new_n426_, new_n1036_, new_n235_, new_n2142_, new_n1576_, new_n301_, new_n1718_, new_n169_, new_n1333_, new_n1132_, new_n395_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n1740_, new_n473_, new_n1624_, new_n1147_, new_n2217_, new_n1827_, new_n2401_, new_n1468_, new_n969_, new_n2332_, new_n1234_, new_n2343_, new_n1360_, new_n378_, new_n621_, new_n1637_, new_n244_, new_n943_, new_n1798_, new_n1321_, new_n1690_, new_n1209_, new_n1709_, new_n347_, new_n2084_, new_n2100_, new_n700_, new_n1419_, new_n921_, new_n396_, new_n1003_, new_n208_, new_n1671_, new_n1239_, new_n528_, new_n1667_, new_n2331_, new_n2213_, new_n2195_, new_n1218_, new_n1346_, new_n1201_, new_n1282_, new_n1630_, new_n2274_, new_n1349_, new_n2317_, new_n1547_, new_n1994_, new_n1437_, new_n2128_, new_n1598_, new_n1205_, new_n1966_, new_n1154_, new_n2411_, new_n295_, new_n1453_, new_n1850_, new_n2194_, new_n628_, new_n409_, new_n1090_, new_n1489_, new_n553_, new_n1061_, new_n2447_, new_n333_, new_n290_, new_n834_, new_n1991_, new_n1781_, new_n1738_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n276_, new_n688_, new_n1704_, new_n410_, new_n1518_, new_n932_, new_n878_, new_n1981_, new_n509_, new_n1761_, new_n202_, new_n296_, new_n2187_, new_n1358_, new_n724_, new_n1070_, new_n1686_, new_n1416_, new_n156_, new_n261_, new_n672_, new_n1496_, new_n616_, new_n529_, new_n323_, new_n914_, new_n1875_, new_n362_, new_n1600_, new_n1631_, new_n2432_, new_n1771_, new_n460_, new_n1267_, new_n2237_, new_n1705_, new_n2090_, new_n1466_, new_n2370_, new_n1707_, new_n1716_, new_n1516_, new_n380_, new_n861_, new_n1564_, new_n1656_, new_n2149_, new_n1252_, new_n1993_, new_n2288_, new_n2371_, new_n352_, new_n1553_, new_n1593_, new_n944_, new_n1542_, new_n1064_, new_n1949_, new_n2280_, new_n2444_, new_n1480_, new_n1745_, new_n1860_, new_n2436_, new_n273_, new_n224_, new_n586_, new_n963_, new_n993_, new_n1357_, new_n102_, new_n143_, new_n1628_, new_n2441_, new_n403_, new_n868_, new_n1242_, new_n2190_, new_n149_, new_n1612_, new_n1343_, new_n936_, new_n1459_, new_n189_, new_n1438_, new_n106_, new_n1016_, new_n1904_, new_n1144_, new_n2461_, new_n1465_, new_n182_, new_n666_, new_n1290_, new_n2065_, new_n2233_, new_n2277_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n1700_, new_n219_, new_n382_, new_n2232_, new_n239_, new_n718_, new_n1310_, new_n2239_, new_n88_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n2103_, new_n95_, new_n1635_, new_n1509_, new_n1559_, new_n2152_, new_n1789_, new_n2440_, new_n544_, new_n2172_, new_n1941_, new_n2465_, new_n1324_, new_n1293_, new_n1336_, new_n345_, new_n2066_, new_n2427_, new_n499_, new_n131_, new_n533_, new_n2416_, new_n795_, new_n459_, new_n1441_, new_n1728_, new_n2363_, new_n2354_, new_n2458_, new_n1510_, new_n1174_, new_n1655_, new_n80_, new_n613_, new_n1464_, new_n417_, new_n837_, new_n801_, new_n2039_, new_n2336_, new_n631_, new_n453_, new_n2430_, new_n1723_, new_n2126_, new_n519_, new_n148_, new_n2319_, new_n662_, new_n864_, new_n2322_, new_n440_, new_n2218_, new_n1826_, new_n2407_, new_n1765_, new_n974_, new_n1907_, new_n2118_, new_n1565_, new_n751_, new_n2289_, new_n2141_, new_n1038_, new_n372_, new_n1758_, new_n2211_, new_n852_, new_n1474_, new_n1328_, new_n1430_, new_n213_, new_n769_, new_n433_, new_n2096_, new_n1956_, new_n109_, new_n1450_, new_n992_, new_n1098_, new_n1729_, new_n2069_, new_n732_, new_n1832_, new_n689_, new_n933_, new_n1608_, new_n1492_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n1379_, new_n712_, new_n550_, new_n1068_, new_n269_, new_n2106_, new_n512_, new_n2375_, new_n2131_, new_n1673_, new_n1220_, new_n989_, new_n1741_, new_n1421_, new_n644_, new_n1856_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n2366_, new_n913_, new_n594_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n881_, new_n1268_, new_n2052_, new_n1381_, new_n1566_, new_n684_, new_n1274_, new_n1893_, new_n1665_, new_n1787_, new_n905_, new_n1539_, new_n1643_, new_n1958_, new_n962_, new_n2399_, new_n86_, new_n627_, new_n760_, new_n1391_, new_n1986_, new_n2408_, new_n1353_, new_n1033_, new_n2050_, new_n2180_, new_n2273_, new_n1153_, new_n320_, new_n984_, new_n1183_, new_n2133_, new_n2353_, new_n89_, new_n2376_, new_n1316_, new_n2391_, new_n1460_, new_n1878_, new_n1602_, new_n128_, new_n610_, new_n1369_, new_n159_, new_n1694_, new_n2226_, new_n1401_, new_n175_, new_n226_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n2446_, new_n171_, new_n1320_, new_n1861_, new_n434_, new_n200_, new_n2021_, new_n2279_, new_n581_, new_n329_, new_n2301_, new_n686_, new_n1567_, new_n168_, new_n1389_, new_n1400_, new_n757_, new_n793_, new_n406_, new_n1597_, new_n1089_, new_n1192_, new_n135_, new_n2347_, new_n405_, new_n2115_, new_n942_, new_n2382_, new_n614_, new_n895_, new_n976_, new_n1405_, new_n1249_, new_n1354_, new_n847_, new_n250_, new_n288_, new_n798_, new_n1926_, new_n1969_, new_n1948_, new_n753_, new_n2345_, new_n1361_, new_n941_, new_n2073_, new_n827_, new_n1356_, new_n1747_, new_n366_, new_n779_, new_n1025_, new_n365_, new_n1207_, new_n1799_, new_n601_, new_n1057_, new_n1644_, new_n1677_, new_n2266_, new_n812_, new_n266_, new_n542_, new_n548_, new_n1397_, new_n1313_, new_n1120_, new_n819_, new_n451_, new_n489_, new_n804_, new_n602_, new_n114_, new_n1060_, new_n1303_, new_n413_, new_n1906_, new_n1544_, new_n1382_, new_n1896_, new_n442_, new_n677_, new_n642_, new_n211_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n1814_, new_n735_, new_n2146_, new_n2202_, new_n1304_, new_n1537_, new_n1834_, new_n1108_, new_n2246_, new_n862_, new_n1606_, new_n532_, new_n2159_, new_n393_, new_n2110_, new_n1617_, new_n292_, new_n2258_, new_n215_, new_n1319_, new_n626_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n2426_, new_n1238_, new_n2062_, new_n133_, new_n2037_, new_n2250_, new_n1880_, new_n1162_, new_n1730_, new_n2018_, new_n212_, new_n2003_, new_n1278_, new_n902_, new_n2113_, new_n2144_, new_n2309_, new_n201_, new_n1996_, new_n414_, new_n2028_, new_n2364_, new_n2011_, new_n1482_, new_n554_, new_n2303_, new_n230_, new_n1151_, new_n2094_, new_n1302_, new_n2212_, new_n855_, new_n103_, new_n1037_, new_n2154_, new_n759_, new_n167_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n1858_, new_n478_, new_n1307_, new_n73_, new_n2339_, new_n1486_, new_n361_, new_n764_, new_n2349_, new_n2081_, new_n2007_, new_n1955_, new_n1683_, new_n510_, new_n966_, new_n351_, new_n1877_, new_n1292_, new_n2036_, new_n609_, new_n180_, new_n1759_, new_n961_, new_n530_, new_n890_, new_n1006_, new_n1836_, new_n1701_, new_n1905_, new_n811_, new_n1445_, new_n1902_, new_n956_, new_n486_, new_n970_, new_n1618_, new_n768_, new_n1691_, new_n773_, new_n1452_, new_n2121_, new_n1823_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n254_, new_n355_, new_n432_, new_n925_, new_n2463_, new_n2040_, new_n1940_, new_n778_, new_n2267_, new_n452_, new_n1483_, new_n2177_, new_n820_, new_n1386_, new_n508_, new_n1844_, new_n714_, new_n1748_, new_n116_, new_n1007_, new_n1613_, new_n882_, new_n2162_, new_n1557_, new_n1159_, new_n118_, new_n1584_, new_n1337_, new_n77_, new_n1348_, new_n1555_, new_n1636_, new_n1322_, new_n1751_, new_n1133_, new_n2164_, new_n1177_, new_n2197_, new_n646_, new_n538_, new_n1026_, new_n2019_, new_n541_, new_n1388_, new_n1550_, new_n2372_, new_n311_, new_n587_, new_n2010_, new_n2220_, new_n465_, new_n84_, new_n783_, new_n1380_, new_n2016_, new_n263_, new_n2080_, new_n1601_, new_n488_, new_n524_, new_n1725_, new_n1245_, new_n663_, new_n1499_, new_n2392_, new_n1791_, new_n2035_, new_n1908_, new_n1689_, new_n198_, new_n1857_, new_n1393_, new_n1335_, new_n1364_, new_n965_, new_n572_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n945_, new_n1882_, new_n1115_, new_n1846_, new_n1231_, new_n2460_, new_n1055_, new_n2043_, new_n1431_, new_n923_, new_n1674_, new_n469_, new_n1633_, new_n2242_, new_n1607_, new_n2373_, new_n1924_, new_n2368_, new_n2188_, new_n457_, new_n1852_, new_n2170_, new_n1301_, new_n1999_, new_n1128_, new_n1002_, new_n1169_, new_n384_, new_n900_, new_n1722_, new_n1824_, new_n2316_, new_n1788_, new_n113_, new_n1648_, new_n2191_, new_n2418_, new_n775_, new_n454_, new_n1872_, new_n1124_, new_n1000_, new_n2225_, new_n1947_, new_n1273_, new_n1491_, new_n1554_, new_n176_, new_n1923_, new_n2013_, new_n291_, new_n309_, new_n1160_, new_n82_, new_n259_, new_n1536_, new_n2305_, new_n2381_, new_n227_, new_n2393_, new_n690_, new_n416_, new_n744_, new_n1175_, new_n2125_, new_n1136_, new_n1272_, new_n1287_, new_n1462_, new_n619_, new_n2410_, new_n1890_, new_n577_, new_n2179_, new_n376_, new_n1538_, new_n1579_, new_n2147_, new_n2310_, new_n2183_, new_n749_, new_n1091_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n2429_, new_n1776_, new_n1030_, new_n485_, new_n578_, new_n918_, new_n126_, new_n1586_, new_n1805_, new_n2380_, new_n2390_, new_n1572_, new_n665_, new_n800_, new_n1387_, new_n719_, new_n1178_, new_n270_, new_n570_, new_n893_, new_n520_, new_n1347_, new_n145_, new_n253_, new_n825_, new_n2312_, new_n1627_, new_n557_, new_n1642_, new_n1807_, new_n2281_, new_n1742_, new_n507_, new_n741_, new_n1699_, new_n1224_, new_n2008_, new_n748_, new_n2117_, new_n1137_, new_n1286_, new_n107_, new_n813_, new_n830_, new_n1107_, new_n730_, new_n1326_, new_n592_, new_n1820_, new_n231_, new_n1080_, new_n1279_, new_n522_, new_n588_, new_n916_, new_n199_, new_n675_, new_n1155_, new_n1186_, new_n1848_, new_n2448_, new_n225_, new_n2002_, new_n1863_, new_n1246_, new_n2119_, new_n387_, new_n112_, new_n2105_, new_n1951_, new_n121_, new_n949_, new_n2048_, new_n221_, new_n450_, new_n1394_, new_n2379_, new_n1179_, new_n298_, new_n184_, new_n1088_, new_n2394_, new_n2374_, new_n1756_, new_n2163_, new_n569_, new_n555_, new_n1139_, new_n1793_, new_n392_, new_n2404_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n147_, new_n692_, new_n502_, new_n1821_, new_n209_, new_n623_, new_n446_, new_n316_, new_n826_, new_n2079_, new_n1476_, new_n1854_, new_n332_, new_n972_, new_n1634_, new_n2285_, new_n2287_, new_n2413_, new_n2178_, new_n1916_, new_n2046_, new_n733_, new_n1983_, new_n122_, new_n1021_, new_n585_, new_n2076_, new_n2116_, new_n2189_, new_n1976_, new_n2307_, new_n242_, new_n503_, new_n2323_, new_n772_, new_n1244_, new_n307_, new_n1736_, new_n1181_, new_n1093_, new_n1451_, new_n2138_, new_n1097_, new_n1069_, new_n1164_, new_n1779_, new_n1869_, new_n2265_, new_n435_, new_n1891_, new_n1719_, new_n1830_, new_n1885_, new_n687_, new_n1029_, new_n1862_, new_n1654_, new_n1688_, new_n1963_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n129_, new_n1112_, new_n1715_, new_n1156_, new_n1938_, new_n930_, new_n1475_, new_n1604_, new_n412_, new_n607_, new_n1731_, new_n645_, new_n1087_, new_n723_, new_n2326_, new_n2282_, new_n1933_, new_n1577_, new_n574_, new_n1548_, new_n1578_, new_n2204_, new_n2435_, new_n1661_, new_n1615_, new_n957_, new_n1047_, new_n75_, new_n787_, new_n336_, new_n2243_, new_n1399_, new_n1531_, new_n1927_, new_n294_, new_n1589_, new_n1792_, new_n1965_, new_n1173_, new_n704_, new_n2087_, new_n1809_, new_n2315_, new_n2443_, new_n1570_, new_n1811_, new_n2004_, new_n2130_, new_n1502_, new_n1778_, new_n2325_, new_n2469_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n2186_, new_n1243_, new_n1077_, new_n2196_, new_n2067_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1506_, new_n1583_, new_n2085_, new_n1011_, new_n802_, new_n104_, new_n1236_, new_n1829_, new_n2150_, new_n2464_, new_n947_, new_n1813_, new_n982_, new_n1449_, new_n1961_, new_n2346_, new_n279_, new_n455_, new_n1982_, new_n1569_, new_n120_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1918_, new_n2222_, new_n1605_, new_n2097_, new_n1964_, new_n1314_, new_n2292_, new_n1359_, new_n1233_, new_n1839_, new_n2236_, new_n501_, new_n1157_, new_n2086_, new_n1575_, new_n1048_, new_n885_, new_n1808_, new_n283_, new_n390_, new_n1910_, new_n1922_, new_n566_, new_n186_, new_n386_, new_n767_, new_n401_, new_n2454_, new_n2173_, new_n556_, new_n1899_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n2095_, new_n246_, new_n1881_, new_n2127_, new_n667_, new_n367_, new_n2099_, new_n1237_, new_n2026_, new_n1837_, new_n1568_, new_n1479_, new_n2240_, new_n2321_, new_n894_, new_n2199_, new_n526_, new_n908_, new_n1886_, new_n2023_, new_n2192_, new_n678_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n2033_, new_n2045_, new_n2160_, new_n2328_, new_n2169_, new_n2283_, new_n2456_, new_n1415_, new_n1390_, new_n721_, new_n742_, new_n892_, new_n1368_, new_n2384_, new_n472_, new_n1919_, new_n1985_, new_n1768_, new_n2111_, new_n1167_, new_n1530_, new_n2070_, new_n1490_, new_n2313_, new_n2278_, new_n792_, new_n953_, new_n257_, new_n2403_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n192_, new_n1851_, new_n635_, new_n1774_, new_n110_, new_n2108_, new_n648_, new_n2450_, new_n164_, new_n1803_, new_n983_, new_n1406_, new_n1990_, new_n1082_, new_n2238_, new_n606_, new_n796_, new_n655_, new_n630_, new_n1717_, new_n1670_, new_n694_, new_n565_, new_n1979_, new_n1984_, new_n108_, new_n183_, new_n511_, new_n2359_, new_n1714_, new_n2034_, new_n2165_, new_n1640_, new_n1031_, new_n2405_, new_n1281_, new_n2129_, new_n1911_, new_n1005_, new_n999_, new_n321_, new_n1816_, new_n324_, new_n1713_, new_n491_, new_n676_, new_n2300_, new_n2112_, new_n271_, new_n674_, new_n274_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n1753_, new_n420_, new_n876_, new_n1894_, new_n1900_, new_n498_, new_n1217_, new_n2032_, new_n1463_, new_n429_, new_n2109_, new_n2122_, new_n1222_, new_n353_, new_n2470_, new_n734_, new_n1062_, new_n506_, new_n872_, new_n1277_, new_n1428_, new_n1440_, new_n656_, new_n2311_, new_n394_, new_n935_, new_n1972_, new_n139_, new_n1150_, new_n1735_, new_n441_, new_n1752_, new_n600_, new_n1737_, new_n1930_, new_n1657_, new_n1797_, new_n1562_, new_n1939_, new_n1953_, new_n398_, new_n2434_, new_n383_, new_n207_, new_n267_, new_n2161_, new_n1395_, new_n1682_, new_n1795_, new_n1373_, new_n1229_, new_n1422_, new_n187_, new_n1523_, new_n1698_, new_n1679_, new_n334_, new_n331_, new_n835_, new_n1574_, new_n1614_, new_n2261_, new_n1423_, new_n1732_, new_n172_, new_n705_, new_n874_, new_n402_, new_n335_, new_n659_, new_n346_, new_n1954_, new_n1315_, new_n696_, new_n1868_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1952_, new_n1365_, new_n952_, new_n1870_, new_n179_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1385_, new_n2185_, new_n559_, new_n762_, new_n2134_, new_n1193_, new_n2467_, new_n1780_, new_n1187_, new_n1253_, new_n1546_, new_n1256_, new_n166_, new_n1513_, new_n162_, new_n1669_, new_n745_, new_n161_, new_n1114_, new_n1084_, new_n668_, new_n1573_, new_n2200_, new_n369_, new_n1693_, new_n1032_, new_n1545_, new_n901_, new_n1757_, new_n1255_, new_n2205_, new_n155_, new_n985_, new_n2074_, new_n1995_, new_n851_, new_n543_, new_n1943_, new_n1975_, new_n886_, new_n371_, new_n1712_, new_n2058_, new_n2075_, new_n2284_, new_n661_, new_n797_, new_n232_, new_n2145_, new_n76_, new_n2466_, new_n1109_, new_n1269_, new_n1653_, new_n2453_, new_n884_, new_n938_, new_n1592_, new_n809_, new_n1142_, new_n1623_, new_n2439_, new_n604_, new_n1461_, new_n1104_, new_n1703_, new_n1511_, new_n571_, new_n1859_, new_n1504_, new_n758_, new_n1802_, new_n328_, new_n2168_, new_n2015_, new_n2327_, new_n130_, new_n2329_, new_n1794_, new_n268_, new_n2124_, new_n1299_, new_n1477_, new_n1079_, new_n144_, new_n2271_, new_n1804_, new_n931_, new_n575_, new_n1493_, new_n2438_, new_n2451_, new_n562_, new_n1929_, new_n2254_, new_n1638_, new_n1065_, new_n1118_, new_n177_, new_n1645_, new_n493_, new_n547_, new_n1934_, new_n264_, new_n379_, new_n1825_, new_n1481_, new_n1325_, new_n1625_, new_n1191_, new_n1931_, new_n824_, new_n2304_, new_n125_, new_n717_, new_n1455_, new_n475_, new_n2249_, new_n237_, new_n858_, new_n2306_, new_n1384_, new_n1434_, new_n411_, new_n673_, new_n1766_, new_n2025_, new_n2082_, new_n407_, new_n1897_, new_n81_, new_n1833_, new_n1692_, new_n1726_, new_n736_, new_n513_, new_n1903_, new_n558_, new_n313_, new_n1370_, new_n2093_, new_n2042_, new_n2415_, new_n1710_, new_n146_, new_n2047_, new_n2167_, new_n919_, new_n302_, new_n755_, new_n2017_, new_n1040_, new_n615_, new_n2298_, new_n722_, new_n856_, new_n415_, new_n537_, new_n2068_, new_n255_, new_n2437_, new_n1130_, new_n2064_, new_n2256_, new_n2360_, new_n1122_, new_n1185_, new_n1240_, new_n2031_, new_n354_, new_n968_, new_n2001_, new_n105_, new_n2419_, new_n2055_, new_n2215_, new_n1508_, new_n337_, new_n1195_, new_n658_, new_n591_, new_n1458_, new_n2091_, new_n163_, new_n1818_, new_n997_, new_n563_, new_n2209_, new_n910_, new_n1521_, new_n1334_, new_n2044_, new_n531_, new_n1675_, new_n2308_, new_n593_, new_n111_, new_n1543_, new_n252_, new_n1248_, new_n1812_, new_n2259_, new_n1978_, new_n2208_, new_n2206_, new_n1454_, new_n978_, new_n1308_, new_n408_, new_n470_, new_n134_, new_n1660_, new_n871_, new_n265_, new_n584_, new_n815_, new_n2223_, new_n1619_, new_n1425_, new_n1980_, new_n857_, new_n1828_, new_n2207_, new_n2272_, new_n1017_, new_n2203_, new_n2314_, new_n1853_, new_n101_, new_n2140_, new_n1471_, new_n1117_, new_n1594_, new_n836_, new_n1684_, new_n2148_, new_n2378_, new_n327_, new_n681_, new_n561_, new_n1427_, new_n2210_, new_n196_, new_n818_, new_n1815_, new_n1376_, new_n1876_, new_n2092_, new_n1534_, new_n640_, new_n2262_, new_n754_, new_n653_, new_n1659_, new_n377_, new_n1258_, new_n2247_, new_n375_, new_n1841_, new_n1724_, new_n1436_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n1339_, new_n1784_, new_n1970_, new_n780_, new_n245_, new_n643_, new_n1194_, new_n1338_, new_n91_, new_n1230_, new_n1027_, new_n348_, new_n2409_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1259_, new_n2297_, new_n1208_, new_n2299_, new_n185_, new_n2241_, new_n1942_, new_n373_, new_n1235_, new_n540_, new_n1149_, new_n1928_, new_n1066_, new_n422_, new_n1944_, new_n99_, new_n1664_, new_n249_, new_n284_, new_n119_, new_n293_, new_n934_, new_n1651_, new_n2457_, new_n770_, new_n1225_, new_n521_, new_n2123_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n2333_, new_n2083_, new_n1616_, new_n1806_, new_n2352_, new_n958_, new_n699_, new_n236_, new_n74_, new_n955_, new_n1895_, new_n79_, new_n888_, new_n1505_, new_n1340_, new_n1180_, new_n817_, new_n720_, new_n1801_, new_n620_, new_n368_, new_n1410_, new_n738_, new_n2201_, new_n1363_, new_n2198_, new_n1317_, new_n2385_, new_n1232_, new_n859_, new_n197_, new_n1211_, new_n1412_, new_n1176_, new_n1374_, new_n2269_, new_n2417_, new_n842_, new_n1552_, new_n170_, new_n682_, new_n1075_, new_n1790_, new_n2030_, new_n1563_, new_n821_, new_n1937_, new_n669_, new_n220_, new_n1402_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n637_, new_n1603_, new_n1971_, new_n1342_, new_n424_, new_n2422_, new_n2182_, new_n1210_, new_n188_, new_n240_, new_n1843_, new_n1487_, new_n1646_, new_n123_, new_n127_, new_n1418_, new_n1871_, new_n761_, new_n2027_, new_n2428_, new_n2156_, new_n840_, new_n1283_, new_n1913_, new_n1873_, new_n898_, new_n1734_, new_n799_, new_n946_, new_n1764_, new_n344_, new_n287_, new_n1977_, new_n2362_, new_n2166_, new_n1901_, new_n1469_, new_n1749_, new_n1838_, new_n427_, new_n2449_, new_n1739_, new_n418_, new_n746_, new_n1221_, new_n1585_, new_n1587_, new_n1264_, new_n1680_, new_n152_, new_n2005_, new_n157_, new_n716_, new_n153_, new_n701_, new_n1676_, new_n1058_, new_n2365_, new_n364_, new_n832_, new_n1696_, new_n2193_, new_n1968_, new_n1101_, new_n1250_, new_n1681_, new_n315_, new_n124_, new_n1050_, new_n2455_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n2234_, new_n589_, new_n248_, new_n350_, new_n117_, new_n1083_, new_n2295_, new_n1297_, new_n2361_, new_n1959_, new_n1720_, new_n2330_, new_n2358_, new_n1228_, new_n710_, new_n971_, new_n2462_, new_n906_, new_n2151_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n1685_, new_n1721_, new_n1184_, new_n1960_, new_n1426_, new_n517_, new_n2077_, new_n1892_, new_n1992_, new_n318_, new_n622_, new_n1706_, new_n2006_, new_n702_, new_n2014_, new_n2230_, new_n833_, new_n1560_, new_n715_, new_n1371_, new_n443_, new_n1086_, new_n158_, new_n763_, new_n1622_, new_n1138_, new_n466_, new_n262_, new_n1652_, new_n2356_, new_n2137_, new_n1847_, new_n2406_, new_n2057_, new_n218_, new_n1170_, new_n2276_, new_n845_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n2398_, new_n1540_, new_n1611_, new_n2143_, new_n205_, new_n1708_, new_n1533_, new_n141_, new_n1754_, new_n1750_, new_n1767_, new_n2235_, new_n887_, new_n926_, new_n2060_, new_n875_, new_n256_, new_n1226_, new_n1727_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n771_, new_n979_, new_n1819_, new_n1435_, new_n2342_, new_n1280_, new_n1241_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n216_, new_n1782_, new_n917_, new_n2275_, new_n2071_, new_n1822_, new_n1887_, new_n210_, new_n447_, new_n2181_, new_n1967_, new_n140_, new_n790_, new_n1081_, new_n1247_, new_n1411_, new_n2000_, new_n739_, new_n2221_, new_n341_, new_n996_, new_n1318_, new_n2088_, new_n846_, new_n915_, new_n349_, new_n2294_, new_n848_, new_n277_, new_n1921_, new_n1772_, new_n1497_, new_n579_, new_n286_, new_n1711_, new_n1254_, new_n2216_, new_n438_, new_n1344_, new_n939_, new_n632_, new_n671_, new_n83_, new_n1514_, new_n2253_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n1446_, new_n2136_, new_n596_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1866_, new_n1383_, new_n948_, new_n1520_, new_n838_, new_n1609_, new_n2324_, new_n2377_, new_n1755_, new_n233_, new_n391_, new_n96_, new_n178_, new_n1085_, new_n2245_, new_n359_, new_n132_, new_n794_, new_n2098_, new_n1582_, new_n2056_, new_n2009_, new_n1702_, new_n1909_, new_n2153_, new_n1810_, new_n448_, new_n1932_, new_n1329_, new_n1161_, new_n2341_, new_n2383_, new_n2367_, new_n2395_, new_n92_, new_n1914_, new_n924_, new_n1867_, new_n97_, new_n1034_, new_n1957_, new_n1663_, new_n308_, new_n2214_, new_n633_, new_n784_, new_n2396_, new_n1396_, new_n258_, new_n860_, new_n306_, new_n494_, new_n2286_, new_n2219_, new_n1166_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n1920_, new_n1043_, new_n222_, new_n400_, new_n693_, new_n1485_, new_n505_, new_n471_, new_n967_, new_n374_, new_n1135_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n2252_, new_n138_, new_n310_, new_n2389_, new_n2388_, new_n1331_, new_n1094_, new_n1621_, new_n839_, new_n2078_, new_n525_, new_n1695_, new_n2412_, new_n940_, new_n810_, new_n2400_, new_n808_, new_n2101_, new_n1284_, new_n907_, new_n897_, new_n1012_, new_n869_, new_n1775_, new_n1525_, new_n2120_, new_n598_, new_n2255_, new_n1935_, new_n1063_, new_n1001_, new_n1917_, new_n90_, new_n260_, new_n251_, new_n300_, new_n1503_, new_n806_, new_n2229_, new_n605_, new_n1074_, new_n2175_, new_n93_, new_n1551_, new_n2423_, new_n480_, new_n625_, new_n1141_, new_n1650_, new_n807_, new_n151_, new_n726_, new_n1763_, new_n1263_, new_n1123_, new_n2020_, new_n2402_, new_n583_, new_n617_, new_n78_, new_n1467_, new_n1762_, new_n1997_, new_n781_, new_n1014_, new_n428_, new_n1855_, new_n487_, new_n360_, new_n98_, new_n2139_, new_n2302_, new_n1915_, new_n1596_, new_n191_, new_n1261_, new_n2445_, new_n2022_, new_n1488_, new_n2024_, new_n2224_, new_n922_, new_n2029_, new_n87_, new_n476_, new_n987_, new_n1641_, new_n2420_, new_n243_, new_n154_, new_n1148_, new_n1146_, new_n174_, new_n468_, new_n977_, new_n2049_, new_n782_, new_n444_, new_n518_, new_n1845_, new_n2174_, new_n285_, new_n1888_, new_n203_, new_n2089_, new_n590_, new_n2357_, new_n789_, new_n515_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n1835_, new_n2338_, new_n2425_, new_n1076_, new_n1350_, new_n160_, new_n312_, new_n535_, new_n725_, new_n100_, new_n814_, new_n527_, new_n115_, new_n1378_, new_n1945_, new_n190_, new_n1478_, new_n597_, new_n1092_, new_n1783_, new_n1143_, new_n1072_, new_n1190_, new_n2442_, new_n651_, new_n1296_, new_n1883_, new_n1309_, new_n1796_, new_n776_, new_n2053_, new_n370_, new_n1649_, new_n1515_, new_n1746_, new_n638_, new_n523_, new_n909_, new_n1840_, new_n2296_, new_n1571_, new_n2386_, new_n1773_, new_n2351_, new_n1470_, new_n711_, new_n1298_, new_n731_, new_n599_, new_n2257_, new_n1260_, new_n973_, new_n1529_, new_n1541_, new_n1096_, new_n2344_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n2228_, new_n1500_, new_n928_, new_n319_, new_n1008_, new_n2059_, new_n1687_, new_n338_, new_n707_, new_n740_, new_n1134_, new_n1291_, new_n247_, new_n539_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1817_, new_n1672_, new_n2061_, new_n1295_, new_n1432_, new_n2158_, new_n1189_, new_n2268_, new_n2355_, new_n1197_, new_n1912_, new_n1312_, new_n2340_, new_n467_, new_n404_, new_n193_, new_n2270_, new_n1666_, new_n1744_, new_n358_, new_n877_, new_n1697_, new_n545_, new_n611_, new_n1998_, new_n289_, new_n72_, new_n425_, new_n896_, new_n1831_, new_n2459_, new_n1925_, new_n1770_, new_n866_, new_n1556_, new_n994_, new_n1494_, new_n2335_, new_n2157_, new_n964_, new_n1078_, new_n2227_, new_n136_, new_n551_, new_n1408_, new_n618_, new_n1140_, new_n2263_, new_n2290_, new_n464_, new_n1498_, new_n94_, new_n204_, new_n181_, new_n1588_, new_n1974_, new_n573_, new_n765_, new_n1103_;

not g0000 ( new_n72_, keyinput3_G223gat );
not g0001 ( new_n73_, keyinput2_G223gat );
not g0002 ( new_n74_, G99gat );
not g0003 ( new_n75_, G108gat );
or g0004 ( new_n76_, G112gat, G115gat );
and g0005 ( new_n77_, new_n76_, G102gat );
or g0006 ( new_n78_, new_n77_, new_n75_ );
and g0007 ( new_n79_, new_n78_, G105gat );
not g0008 ( new_n80_, G105gat );
not g0009 ( new_n81_, G102gat );
and g0010 ( new_n82_, new_n81_, G108gat );
not g0011 ( new_n83_, new_n82_ );
and g0012 ( new_n84_, new_n83_, new_n80_ );
or g0013 ( new_n85_, new_n79_, new_n84_ );
and g0014 ( new_n86_, new_n85_, new_n74_ );
and g0015 ( new_n87_, G102gat, G112gat );
not g0016 ( new_n88_, new_n87_ );
and g0017 ( new_n89_, new_n88_, G108gat );
not g0018 ( new_n90_, new_n89_ );
and g0019 ( new_n91_, new_n90_, G99gat );
and g0020 ( new_n92_, new_n91_, new_n80_ );
or g0021 ( new_n93_, new_n86_, new_n92_ );
and g0022 ( new_n94_, new_n93_, G89gat );
not g0023 ( new_n95_, G89gat );
and g0024 ( new_n96_, G112gat, G115gat );
or g0025 ( new_n97_, new_n83_, new_n96_ );
and g0026 ( new_n98_, new_n97_, G105gat );
or g0027 ( new_n99_, G102gat, G112gat );
or g0028 ( new_n100_, new_n99_, new_n75_ );
and g0029 ( new_n101_, new_n100_, new_n80_ );
or g0030 ( new_n102_, new_n98_, new_n101_ );
and g0031 ( new_n103_, new_n102_, G99gat );
not g0032 ( new_n104_, new_n99_ );
not g0033 ( new_n105_, G115gat );
and g0034 ( new_n106_, new_n105_, G108gat );
and g0035 ( new_n107_, new_n104_, new_n106_ );
not g0036 ( new_n108_, new_n107_ );
or g0037 ( new_n109_, new_n108_, new_n80_ );
and g0038 ( new_n110_, new_n109_, new_n74_ );
or g0039 ( new_n111_, new_n103_, new_n110_ );
and g0040 ( new_n112_, new_n111_, new_n95_ );
or g0041 ( new_n113_, new_n94_, new_n112_ );
and g0042 ( new_n114_, new_n87_, G115gat );
or g0043 ( new_n115_, new_n114_, new_n75_ );
and g0044 ( new_n116_, new_n115_, G105gat );
and g0045 ( new_n117_, G89gat, G99gat );
and g0046 ( new_n118_, new_n116_, new_n117_ );
or g0047 ( new_n119_, new_n113_, new_n118_ );
and g0048 ( new_n120_, new_n119_, keyinput0_G223gat );
not g0049 ( new_n121_, keyinput0_G223gat );
and g0050 ( new_n122_, new_n91_, new_n121_ );
or g0051 ( new_n123_, new_n120_, new_n122_ );
and g0052 ( new_n124_, new_n123_, keyinput1_G223gat );
not g0053 ( new_n125_, keyinput1_G223gat );
and g0054 ( new_n126_, new_n82_, new_n105_ );
or g0055 ( new_n127_, new_n101_, new_n126_ );
and g0056 ( new_n128_, new_n127_, G99gat );
or g0057 ( new_n129_, new_n107_, new_n80_ );
and g0058 ( new_n130_, new_n129_, new_n74_ );
or g0059 ( new_n131_, new_n128_, new_n130_ );
and g0060 ( new_n132_, new_n131_, new_n121_ );
and g0061 ( new_n133_, new_n129_, keyinput0_G223gat );
or g0062 ( new_n134_, new_n132_, new_n133_ );
and g0063 ( new_n135_, new_n134_, new_n125_ );
or g0064 ( new_n136_, new_n124_, new_n135_ );
and g0065 ( new_n137_, new_n136_, new_n73_ );
and g0066 ( new_n138_, new_n89_, new_n105_ );
or g0067 ( new_n139_, new_n138_, new_n80_ );
or g0068 ( new_n140_, new_n83_, new_n105_ );
and g0069 ( new_n141_, new_n139_, new_n140_ );
and g0070 ( new_n142_, new_n141_, new_n74_ );
or g0071 ( new_n143_, new_n90_, new_n105_ );
and g0072 ( new_n144_, new_n143_, G99gat );
or g0073 ( new_n145_, new_n106_, new_n80_ );
and g0074 ( new_n146_, new_n144_, new_n145_ );
or g0075 ( new_n147_, new_n142_, new_n146_ );
and g0076 ( new_n148_, new_n147_, new_n121_ );
and g0077 ( new_n149_, new_n141_, keyinput0_G223gat );
or g0078 ( new_n150_, new_n148_, new_n149_ );
and g0079 ( new_n151_, new_n150_, new_n125_ );
and g0080 ( new_n152_, new_n83_, new_n74_ );
not g0081 ( new_n153_, G112gat );
and g0082 ( new_n154_, new_n153_, G108gat );
or g0083 ( new_n155_, new_n152_, new_n154_ );
and g0084 ( new_n156_, new_n155_, G89gat );
not g0085 ( new_n157_, new_n100_ );
or g0086 ( new_n158_, new_n157_, new_n74_ );
and g0087 ( new_n159_, new_n158_, new_n95_ );
or g0088 ( new_n160_, new_n156_, new_n159_ );
and g0089 ( new_n161_, new_n160_, keyinput0_G223gat );
not g0090 ( new_n162_, G95gat );
or g0091 ( new_n163_, new_n117_, new_n162_ );
and g0092 ( new_n164_, new_n90_, new_n163_ );
and g0093 ( new_n165_, new_n164_, new_n121_ );
or g0094 ( new_n166_, new_n161_, new_n165_ );
and g0095 ( new_n167_, new_n166_, keyinput1_G223gat );
or g0096 ( new_n168_, new_n151_, new_n167_ );
and g0097 ( new_n169_, new_n168_, keyinput2_G223gat );
or g0098 ( new_n170_, new_n137_, new_n169_ );
and g0099 ( new_n171_, new_n170_, new_n72_ );
and g0100 ( new_n172_, new_n95_, G95gat );
not g0101 ( new_n173_, new_n172_ );
and g0102 ( new_n174_, new_n83_, new_n173_ );
not g0103 ( new_n175_, G76gat );
and g0104 ( new_n176_, new_n175_, G82gat );
not g0105 ( new_n177_, new_n176_ );
and g0106 ( new_n178_, new_n174_, new_n177_ );
not g0107 ( new_n179_, G63gat );
and g0108 ( new_n180_, new_n179_, G69gat );
not g0109 ( new_n181_, new_n180_ );
and g0110 ( new_n182_, new_n178_, new_n181_ );
not g0111 ( new_n183_, G50gat );
and g0112 ( new_n184_, new_n183_, G56gat );
not g0113 ( new_n185_, new_n184_ );
and g0114 ( new_n186_, new_n182_, new_n185_ );
not g0115 ( new_n187_, G37gat );
and g0116 ( new_n188_, new_n187_, G43gat );
not g0117 ( new_n189_, new_n188_ );
and g0118 ( new_n190_, new_n186_, new_n189_ );
not g0119 ( new_n191_, G24gat );
and g0120 ( new_n192_, new_n191_, G30gat );
not g0121 ( new_n193_, new_n192_ );
and g0122 ( new_n194_, new_n190_, new_n193_ );
not g0123 ( new_n195_, G11gat );
and g0124 ( new_n196_, new_n195_, G17gat );
not g0125 ( new_n197_, new_n196_ );
not g0126 ( new_n198_, G4gat );
or g0127 ( new_n199_, new_n198_, G1gat );
and g0128 ( new_n200_, new_n197_, new_n199_ );
and g0129 ( new_n201_, new_n194_, new_n200_ );
not g0130 ( new_n202_, new_n201_ );
and g0131 ( new_n203_, new_n202_, keyinput0_G223gat );
and g0132 ( new_n204_, new_n121_, G108gat );
or g0133 ( new_n205_, new_n203_, new_n204_ );
and g0134 ( new_n206_, new_n205_, keyinput1_G223gat );
or g0135 ( new_n207_, new_n106_, new_n121_ );
not g0136 ( new_n208_, new_n204_ );
and g0137 ( new_n209_, new_n208_, new_n125_ );
and g0138 ( new_n210_, new_n209_, new_n207_ );
or g0139 ( new_n211_, new_n206_, new_n210_ );
and g0140 ( new_n212_, new_n211_, keyinput2_G223gat );
not g0141 ( new_n213_, new_n116_ );
and g0142 ( new_n214_, new_n213_, new_n121_ );
and g0143 ( new_n215_, new_n115_, keyinput0_G223gat );
or g0144 ( new_n216_, new_n214_, new_n215_ );
and g0145 ( new_n217_, new_n216_, keyinput1_G223gat );
and g0146 ( new_n218_, new_n117_, G105gat );
or g0147 ( new_n219_, new_n218_, new_n162_ );
and g0148 ( new_n220_, new_n115_, new_n219_ );
and g0149 ( new_n221_, new_n220_, keyinput0_G223gat );
or g0150 ( new_n222_, new_n221_, new_n122_ );
and g0151 ( new_n223_, new_n222_, new_n125_ );
or g0152 ( new_n224_, new_n217_, new_n223_ );
and g0153 ( new_n225_, new_n224_, new_n73_ );
or g0154 ( new_n226_, new_n212_, new_n225_ );
and g0155 ( new_n227_, new_n226_, keyinput3_G223gat );
or g0156 ( G223gat, new_n171_, new_n227_ );
not g0157 ( new_n229_, G86gat );
and g0158 ( new_n230_, new_n172_, new_n74_ );
not g0159 ( new_n231_, new_n230_ );
and g0160 ( new_n232_, new_n231_, new_n100_ );
not g0161 ( new_n233_, new_n232_ );
or g0162 ( new_n234_, new_n233_, new_n174_ );
and g0163 ( new_n235_, new_n234_, new_n229_ );
and g0164 ( new_n236_, G89gat, G112gat );
not g0165 ( new_n237_, new_n236_ );
or g0166 ( new_n238_, new_n83_, new_n237_ );
and g0167 ( new_n239_, G99gat, G102gat );
not g0168 ( new_n240_, new_n239_ );
or g0169 ( new_n241_, new_n173_, new_n240_ );
and g0170 ( new_n242_, new_n74_, G95gat );
or g0171 ( new_n243_, new_n154_, new_n242_ );
and g0172 ( new_n244_, new_n241_, new_n243_ );
and g0173 ( new_n245_, new_n244_, new_n238_ );
and g0174 ( new_n246_, new_n245_, G86gat );
or g0175 ( new_n247_, new_n235_, new_n246_ );
and g0176 ( new_n248_, new_n247_, G76gat );
or g0177 ( new_n249_, new_n233_, new_n229_ );
and g0178 ( new_n250_, new_n249_, new_n175_ );
or g0179 ( new_n251_, new_n248_, new_n250_ );
and g0180 ( new_n252_, new_n251_, G82gat );
not g0181 ( new_n253_, G82gat );
and g0182 ( new_n254_, new_n245_, new_n253_ );
or g0183 ( new_n255_, new_n252_, new_n254_ );
and g0184 ( new_n256_, new_n255_, G73gat );
not g0185 ( new_n257_, G73gat );
and g0186 ( new_n258_, new_n176_, new_n229_ );
not g0187 ( new_n259_, new_n258_ );
and g0188 ( new_n260_, new_n232_, new_n259_ );
not g0189 ( new_n261_, new_n260_ );
or g0190 ( new_n262_, new_n261_, new_n178_ );
and g0191 ( new_n263_, new_n262_, new_n257_ );
or g0192 ( new_n264_, new_n256_, new_n263_ );
and g0193 ( new_n265_, new_n264_, G63gat );
not g0194 ( new_n266_, G69gat );
or g0195 ( new_n267_, new_n261_, new_n257_ );
and g0196 ( new_n268_, new_n267_, new_n179_ );
or g0197 ( new_n269_, new_n268_, new_n266_ );
or g0198 ( new_n270_, new_n265_, new_n269_ );
or g0199 ( new_n271_, new_n255_, G69gat );
and g0200 ( new_n272_, new_n270_, new_n271_ );
not g0201 ( new_n273_, G56gat );
and g0202 ( new_n274_, G50gat, G60gat );
or g0203 ( new_n275_, new_n274_, new_n273_ );
not g0204 ( new_n276_, new_n275_ );
or g0205 ( new_n277_, new_n272_, new_n276_ );
and g0206 ( new_n278_, new_n268_, G69gat );
and g0207 ( new_n279_, new_n262_, new_n181_ );
or g0208 ( new_n280_, new_n278_, new_n279_ );
or g0209 ( new_n281_, new_n280_, new_n183_ );
not g0210 ( new_n282_, G60gat );
and g0211 ( new_n283_, new_n180_, new_n257_ );
not g0212 ( new_n284_, new_n283_ );
and g0213 ( new_n285_, new_n260_, new_n284_ );
not g0214 ( new_n286_, new_n285_ );
or g0215 ( new_n287_, new_n286_, new_n282_ );
and g0216 ( new_n288_, new_n281_, new_n287_ );
or g0217 ( new_n289_, new_n288_, new_n275_ );
and g0218 ( new_n290_, new_n277_, new_n289_ );
not g0219 ( new_n291_, G43gat );
and g0220 ( new_n292_, G37gat, G47gat );
or g0221 ( new_n293_, new_n292_, new_n291_ );
not g0222 ( new_n294_, new_n293_ );
or g0223 ( new_n295_, new_n290_, new_n294_ );
or g0224 ( new_n296_, new_n280_, new_n184_ );
or g0225 ( new_n297_, new_n287_, new_n185_ );
and g0226 ( new_n298_, new_n296_, new_n297_ );
or g0227 ( new_n299_, new_n298_, new_n187_ );
and g0228 ( new_n300_, new_n184_, new_n282_ );
not g0229 ( new_n301_, new_n300_ );
and g0230 ( new_n302_, new_n285_, new_n301_ );
and g0231 ( new_n303_, new_n302_, G47gat );
not g0232 ( new_n304_, new_n303_ );
and g0233 ( new_n305_, new_n299_, new_n304_ );
or g0234 ( new_n306_, new_n305_, new_n293_ );
and g0235 ( new_n307_, new_n295_, new_n306_ );
not g0236 ( new_n308_, G30gat );
and g0237 ( new_n309_, G24gat, G34gat );
or g0238 ( new_n310_, new_n309_, new_n308_ );
not g0239 ( new_n311_, new_n310_ );
or g0240 ( new_n312_, new_n307_, new_n311_ );
or g0241 ( new_n313_, new_n298_, new_n188_ );
and g0242 ( new_n314_, new_n303_, new_n188_ );
not g0243 ( new_n315_, new_n314_ );
and g0244 ( new_n316_, new_n313_, new_n315_ );
not g0245 ( new_n317_, G34gat );
and g0246 ( new_n318_, new_n317_, G24gat );
not g0247 ( new_n319_, new_n318_ );
or g0248 ( new_n320_, new_n316_, new_n319_ );
not g0249 ( new_n321_, G47gat );
and g0250 ( new_n322_, new_n188_, new_n321_ );
not g0251 ( new_n323_, new_n322_ );
and g0252 ( new_n324_, new_n191_, G34gat );
and g0253 ( new_n325_, new_n323_, new_n324_ );
and g0254 ( new_n326_, new_n302_, new_n325_ );
not g0255 ( new_n327_, new_n326_ );
and g0256 ( new_n328_, new_n320_, new_n327_ );
or g0257 ( new_n329_, new_n328_, new_n308_ );
and g0258 ( new_n330_, G1gat, G8gat );
or g0259 ( new_n331_, new_n330_, new_n198_ );
not g0260 ( new_n332_, G17gat );
and g0261 ( new_n333_, G11gat, G21gat );
or g0262 ( new_n334_, new_n333_, new_n332_ );
and g0263 ( new_n335_, new_n331_, new_n334_ );
and g0264 ( new_n336_, new_n329_, new_n335_ );
and g0265 ( new_n337_, new_n312_, new_n336_ );
not g0266 ( new_n338_, G21gat );
or g0267 ( new_n339_, new_n316_, new_n192_ );
and g0268 ( new_n340_, new_n326_, G30gat );
not g0269 ( new_n341_, new_n340_ );
and g0270 ( new_n342_, new_n339_, new_n341_ );
and g0271 ( new_n343_, new_n342_, new_n338_ );
and g0272 ( new_n344_, new_n192_, new_n317_ );
not g0273 ( new_n345_, new_n344_ );
and g0274 ( new_n346_, new_n323_, new_n345_ );
and g0275 ( new_n347_, new_n302_, new_n346_ );
and g0276 ( new_n348_, new_n347_, G21gat );
not g0277 ( new_n349_, new_n348_ );
and g0278 ( new_n350_, new_n349_, new_n195_ );
or g0279 ( new_n351_, new_n343_, new_n350_ );
and g0280 ( new_n352_, new_n199_, G17gat );
and g0281 ( new_n353_, new_n351_, new_n352_ );
not g0282 ( new_n354_, G8gat );
and g0283 ( new_n355_, new_n354_, G1gat );
and g0284 ( new_n356_, new_n197_, new_n355_ );
and g0285 ( new_n357_, new_n342_, new_n356_ );
not g0286 ( new_n358_, G1gat );
or g0287 ( new_n359_, new_n197_, G21gat );
and g0288 ( new_n360_, new_n359_, G8gat );
and g0289 ( new_n361_, new_n347_, new_n360_ );
not g0290 ( new_n362_, new_n361_ );
and g0291 ( new_n363_, new_n362_, new_n358_ );
or g0292 ( new_n364_, new_n357_, new_n363_ );
and g0293 ( new_n365_, new_n364_, G4gat );
or g0294 ( new_n366_, new_n353_, new_n365_ );
or g0295 ( new_n367_, new_n337_, new_n366_ );
and g0296 ( new_n368_, new_n367_, keyinput3_G329gat );
not g0297 ( new_n369_, keyinput3_G329gat );
and g0298 ( new_n370_, new_n89_, new_n369_ );
or g0299 ( new_n371_, new_n368_, new_n370_ );
and g0300 ( new_n372_, new_n371_, keyinput2_G329gat );
not g0301 ( new_n373_, keyinput2_G329gat );
or g0302 ( new_n374_, new_n80_, G115gat );
and g0303 ( new_n375_, new_n374_, new_n74_ );
or g0304 ( new_n376_, new_n375_, G112gat );
or g0305 ( new_n377_, new_n374_, new_n74_ );
and g0306 ( new_n378_, new_n376_, new_n377_ );
and g0307 ( new_n379_, new_n378_, new_n369_ );
or g0308 ( new_n380_, new_n379_, new_n83_ );
and g0309 ( new_n381_, new_n380_, new_n373_ );
or g0310 ( new_n382_, new_n372_, new_n381_ );
and g0311 ( new_n383_, new_n382_, keyinput1_G329gat );
or g0312 ( new_n384_, new_n172_, new_n176_ );
or g0313 ( new_n385_, new_n180_, new_n187_ );
or g0314 ( new_n386_, new_n385_, new_n184_ );
or g0315 ( new_n387_, new_n386_, new_n384_ );
and g0316 ( new_n388_, new_n387_, new_n369_ );
or g0317 ( new_n389_, new_n388_, new_n373_ );
or g0318 ( new_n390_, new_n384_, new_n369_ );
and g0319 ( new_n391_, new_n389_, new_n390_ );
or g0320 ( new_n392_, new_n391_, new_n82_ );
not g0321 ( new_n393_, keyinput1_G329gat );
and g0322 ( new_n394_, new_n74_, new_n80_ );
not g0323 ( new_n395_, new_n394_ );
and g0324 ( new_n396_, new_n395_, G89gat );
and g0325 ( new_n397_, new_n78_, new_n396_ );
or g0326 ( new_n398_, keyinput2_G329gat, keyinput3_G329gat );
or g0327 ( new_n399_, new_n397_, new_n398_ );
and g0328 ( new_n400_, new_n399_, new_n393_ );
and g0329 ( new_n401_, new_n392_, new_n400_ );
or g0330 ( new_n402_, new_n383_, new_n401_ );
and g0331 ( new_n403_, new_n402_, keyinput0_G329gat );
not g0332 ( new_n404_, keyinput0_G329gat );
and g0333 ( new_n405_, new_n95_, G102gat );
or g0334 ( new_n406_, new_n378_, new_n405_ );
or g0335 ( new_n407_, new_n95_, G102gat );
and g0336 ( new_n408_, new_n406_, new_n407_ );
or g0337 ( new_n409_, new_n408_, new_n75_ );
and g0338 ( new_n410_, new_n409_, new_n369_ );
and g0339 ( new_n411_, new_n213_, keyinput3_G329gat );
or g0340 ( new_n412_, new_n410_, new_n411_ );
and g0341 ( new_n413_, new_n412_, new_n373_ );
and g0342 ( new_n414_, new_n138_, new_n369_ );
and g0343 ( new_n415_, new_n75_, keyinput3_G329gat );
or g0344 ( new_n416_, new_n414_, new_n415_ );
and g0345 ( new_n417_, new_n416_, keyinput2_G329gat );
or g0346 ( new_n418_, new_n413_, new_n417_ );
and g0347 ( new_n419_, new_n418_, keyinput1_G329gat );
and g0348 ( new_n420_, new_n83_, G89gat );
and g0349 ( new_n421_, new_n95_, new_n74_ );
or g0350 ( new_n422_, new_n157_, new_n421_ );
or g0351 ( new_n423_, new_n422_, new_n420_ );
and g0352 ( new_n424_, new_n423_, new_n369_ );
not g0353 ( new_n425_, new_n420_ );
and g0354 ( new_n426_, new_n425_, keyinput3_G329gat );
or g0355 ( new_n427_, new_n424_, new_n426_ );
and g0356 ( new_n428_, new_n427_, keyinput2_G329gat );
and g0357 ( new_n429_, new_n127_, new_n369_ );
and g0358 ( new_n430_, new_n220_, keyinput3_G329gat );
or g0359 ( new_n431_, new_n429_, new_n430_ );
and g0360 ( new_n432_, new_n431_, new_n373_ );
or g0361 ( new_n433_, new_n428_, new_n432_ );
and g0362 ( new_n434_, new_n433_, new_n393_ );
or g0363 ( new_n435_, new_n419_, new_n434_ );
and g0364 ( new_n436_, new_n435_, new_n404_ );
or g0365 ( G329gat, new_n403_, new_n436_ );
and g0366 ( new_n438_, new_n147_, G89gat );
and g0367 ( new_n439_, new_n131_, new_n95_ );
or g0368 ( new_n440_, new_n438_, new_n439_ );
and g0369 ( new_n441_, new_n440_, G95gat );
and g0370 ( new_n442_, new_n106_, new_n162_ );
or g0371 ( new_n443_, new_n441_, new_n442_ );
and g0372 ( new_n444_, new_n443_, G92gat );
not g0373 ( new_n445_, G92gat );
or g0374 ( new_n446_, new_n142_, new_n144_ );
and g0375 ( new_n447_, new_n446_, G89gat );
or g0376 ( new_n448_, new_n447_, new_n439_ );
and g0377 ( new_n449_, new_n448_, G95gat );
and g0378 ( new_n450_, new_n143_, new_n162_ );
or g0379 ( new_n451_, new_n449_, new_n450_ );
and g0380 ( new_n452_, new_n451_, new_n445_ );
or g0381 ( new_n453_, new_n444_, new_n452_ );
and g0382 ( new_n454_, new_n453_, G86gat );
and g0383 ( new_n455_, new_n138_, G99gat );
or g0384 ( new_n456_, new_n142_, new_n455_ );
and g0385 ( new_n457_, new_n456_, G89gat );
or g0386 ( new_n458_, new_n457_, new_n439_ );
and g0387 ( new_n459_, new_n458_, G95gat );
and g0388 ( new_n460_, new_n138_, new_n162_ );
or g0389 ( new_n461_, new_n459_, new_n460_ );
and g0390 ( new_n462_, new_n461_, G92gat );
or g0391 ( new_n463_, new_n131_, new_n173_ );
or g0392 ( new_n464_, new_n140_, new_n172_ );
and g0393 ( new_n465_, new_n463_, new_n464_ );
and g0394 ( new_n466_, new_n465_, new_n445_ );
or g0395 ( new_n467_, new_n462_, new_n466_ );
and g0396 ( new_n468_, new_n467_, new_n229_ );
or g0397 ( new_n469_, new_n454_, new_n468_ );
and g0398 ( new_n470_, new_n469_, G76gat );
or g0399 ( new_n471_, new_n126_, new_n172_ );
and g0400 ( new_n472_, new_n463_, new_n471_ );
and g0401 ( new_n473_, new_n472_, G92gat );
and g0402 ( new_n474_, new_n157_, G115gat );
not g0403 ( new_n475_, new_n474_ );
or g0404 ( new_n476_, new_n475_, new_n230_ );
or g0405 ( new_n477_, new_n129_, new_n231_ );
and g0406 ( new_n478_, new_n476_, new_n477_ );
and g0407 ( new_n479_, new_n478_, new_n445_ );
or g0408 ( new_n480_, new_n473_, new_n479_ );
and g0409 ( new_n481_, new_n480_, G86gat );
and g0410 ( new_n482_, new_n394_, new_n172_ );
or g0411 ( new_n483_, new_n107_, new_n482_ );
or g0412 ( new_n484_, new_n483_, new_n445_ );
and g0413 ( new_n485_, new_n484_, new_n229_ );
or g0414 ( new_n486_, new_n481_, new_n485_ );
and g0415 ( new_n487_, new_n486_, new_n175_ );
or g0416 ( new_n488_, new_n470_, new_n487_ );
and g0417 ( new_n489_, new_n488_, G82gat );
and g0418 ( new_n490_, new_n443_, new_n253_ );
or g0419 ( new_n491_, new_n489_, new_n490_ );
and g0420 ( new_n492_, new_n491_, G79gat );
not g0421 ( new_n493_, G79gat );
and g0422 ( new_n494_, new_n451_, G86gat );
or g0423 ( new_n495_, new_n468_, new_n494_ );
and g0424 ( new_n496_, new_n495_, G76gat );
or g0425 ( new_n497_, new_n496_, new_n487_ );
and g0426 ( new_n498_, new_n497_, G82gat );
and g0427 ( new_n499_, new_n451_, new_n253_ );
or g0428 ( new_n500_, new_n498_, new_n499_ );
and g0429 ( new_n501_, new_n500_, new_n493_ );
or g0430 ( new_n502_, new_n492_, new_n501_ );
and g0431 ( new_n503_, new_n502_, G73gat );
and g0432 ( new_n504_, new_n461_, G86gat );
or g0433 ( new_n505_, new_n468_, new_n504_ );
and g0434 ( new_n506_, new_n505_, G76gat );
or g0435 ( new_n507_, new_n506_, new_n487_ );
and g0436 ( new_n508_, new_n507_, G82gat );
and g0437 ( new_n509_, new_n461_, new_n253_ );
or g0438 ( new_n510_, new_n508_, new_n509_ );
and g0439 ( new_n511_, new_n510_, G79gat );
and g0440 ( new_n512_, new_n487_, G82gat );
and g0441 ( new_n513_, new_n465_, new_n177_ );
or g0442 ( new_n514_, new_n512_, new_n513_ );
and g0443 ( new_n515_, new_n514_, new_n493_ );
or g0444 ( new_n516_, new_n511_, new_n515_ );
and g0445 ( new_n517_, new_n516_, new_n257_ );
or g0446 ( new_n518_, new_n503_, new_n517_ );
and g0447 ( new_n519_, new_n518_, G63gat );
and g0448 ( new_n520_, new_n472_, new_n177_ );
or g0449 ( new_n521_, new_n512_, new_n520_ );
and g0450 ( new_n522_, new_n521_, G79gat );
or g0451 ( new_n523_, new_n478_, new_n258_ );
or g0452 ( new_n524_, new_n484_, new_n259_ );
and g0453 ( new_n525_, new_n523_, new_n524_ );
and g0454 ( new_n526_, new_n525_, new_n493_ );
or g0455 ( new_n527_, new_n522_, new_n526_ );
and g0456 ( new_n528_, new_n527_, G73gat );
not g0457 ( new_n529_, new_n483_ );
and g0458 ( new_n530_, new_n229_, new_n445_ );
and g0459 ( new_n531_, new_n530_, new_n176_ );
not g0460 ( new_n532_, new_n531_ );
and g0461 ( new_n533_, new_n529_, new_n532_ );
not g0462 ( new_n534_, new_n533_ );
or g0463 ( new_n535_, new_n534_, new_n493_ );
and g0464 ( new_n536_, new_n535_, new_n257_ );
or g0465 ( new_n537_, new_n528_, new_n536_ );
and g0466 ( new_n538_, new_n537_, new_n179_ );
or g0467 ( new_n539_, new_n519_, new_n538_ );
and g0468 ( new_n540_, new_n539_, G69gat );
and g0469 ( new_n541_, new_n491_, new_n266_ );
or g0470 ( new_n542_, new_n540_, new_n541_ );
and g0471 ( new_n543_, new_n542_, G66gat );
not g0472 ( new_n544_, G66gat );
and g0473 ( new_n545_, new_n500_, G73gat );
or g0474 ( new_n546_, new_n517_, new_n545_ );
and g0475 ( new_n547_, new_n546_, G63gat );
or g0476 ( new_n548_, new_n547_, new_n538_ );
and g0477 ( new_n549_, new_n548_, G69gat );
and g0478 ( new_n550_, new_n500_, new_n266_ );
or g0479 ( new_n551_, new_n549_, new_n550_ );
and g0480 ( new_n552_, new_n551_, new_n544_ );
or g0481 ( new_n553_, new_n543_, new_n552_ );
and g0482 ( new_n554_, new_n553_, G60gat );
and g0483 ( new_n555_, new_n510_, G73gat );
or g0484 ( new_n556_, new_n517_, new_n555_ );
and g0485 ( new_n557_, new_n556_, G63gat );
or g0486 ( new_n558_, new_n557_, new_n538_ );
and g0487 ( new_n559_, new_n558_, G69gat );
and g0488 ( new_n560_, new_n510_, new_n266_ );
or g0489 ( new_n561_, new_n559_, new_n560_ );
and g0490 ( new_n562_, new_n561_, G66gat );
and g0491 ( new_n563_, new_n538_, G69gat );
and g0492 ( new_n564_, new_n514_, new_n181_ );
or g0493 ( new_n565_, new_n563_, new_n564_ );
and g0494 ( new_n566_, new_n565_, new_n544_ );
or g0495 ( new_n567_, new_n562_, new_n566_ );
and g0496 ( new_n568_, new_n567_, new_n282_ );
or g0497 ( new_n569_, new_n554_, new_n568_ );
and g0498 ( new_n570_, new_n569_, G50gat );
and g0499 ( new_n571_, new_n521_, new_n181_ );
or g0500 ( new_n572_, new_n563_, new_n571_ );
and g0501 ( new_n573_, new_n572_, G66gat );
or g0502 ( new_n574_, new_n525_, new_n283_ );
or g0503 ( new_n575_, new_n535_, new_n284_ );
and g0504 ( new_n576_, new_n574_, new_n575_ );
and g0505 ( new_n577_, new_n576_, new_n544_ );
or g0506 ( new_n578_, new_n573_, new_n577_ );
and g0507 ( new_n579_, new_n578_, G60gat );
and g0508 ( new_n580_, new_n257_, new_n493_ );
and g0509 ( new_n581_, new_n580_, new_n180_ );
or g0510 ( new_n582_, new_n534_, new_n581_ );
or g0511 ( new_n583_, new_n582_, new_n544_ );
and g0512 ( new_n584_, new_n583_, new_n282_ );
or g0513 ( new_n585_, new_n579_, new_n584_ );
and g0514 ( new_n586_, new_n585_, new_n183_ );
or g0515 ( new_n587_, new_n570_, new_n586_ );
and g0516 ( new_n588_, new_n587_, G56gat );
and g0517 ( new_n589_, new_n542_, new_n273_ );
or g0518 ( new_n590_, new_n588_, new_n589_ );
and g0519 ( new_n591_, new_n590_, G53gat );
not g0520 ( new_n592_, G53gat );
and g0521 ( new_n593_, new_n551_, G60gat );
or g0522 ( new_n594_, new_n568_, new_n593_ );
and g0523 ( new_n595_, new_n594_, G50gat );
or g0524 ( new_n596_, new_n595_, new_n586_ );
and g0525 ( new_n597_, new_n596_, G56gat );
and g0526 ( new_n598_, new_n551_, new_n273_ );
or g0527 ( new_n599_, new_n597_, new_n598_ );
and g0528 ( new_n600_, new_n599_, new_n592_ );
or g0529 ( new_n601_, new_n591_, new_n600_ );
and g0530 ( new_n602_, new_n601_, G47gat );
and g0531 ( new_n603_, new_n561_, G60gat );
or g0532 ( new_n604_, new_n568_, new_n603_ );
and g0533 ( new_n605_, new_n604_, G50gat );
or g0534 ( new_n606_, new_n605_, new_n586_ );
and g0535 ( new_n607_, new_n606_, G56gat );
and g0536 ( new_n608_, new_n561_, new_n273_ );
or g0537 ( new_n609_, new_n607_, new_n608_ );
and g0538 ( new_n610_, new_n609_, G53gat );
and g0539 ( new_n611_, new_n586_, G56gat );
and g0540 ( new_n612_, new_n565_, new_n185_ );
or g0541 ( new_n613_, new_n611_, new_n612_ );
and g0542 ( new_n614_, new_n613_, new_n592_ );
or g0543 ( new_n615_, new_n610_, new_n614_ );
and g0544 ( new_n616_, new_n615_, new_n321_ );
or g0545 ( new_n617_, new_n602_, new_n616_ );
and g0546 ( new_n618_, new_n617_, G37gat );
and g0547 ( new_n619_, new_n572_, new_n185_ );
or g0548 ( new_n620_, new_n611_, new_n619_ );
and g0549 ( new_n621_, new_n620_, G53gat );
or g0550 ( new_n622_, new_n576_, new_n300_ );
or g0551 ( new_n623_, new_n583_, new_n301_ );
and g0552 ( new_n624_, new_n622_, new_n623_ );
and g0553 ( new_n625_, new_n624_, new_n592_ );
or g0554 ( new_n626_, new_n621_, new_n625_ );
and g0555 ( new_n627_, new_n626_, G47gat );
not g0556 ( new_n628_, new_n582_ );
and g0557 ( new_n629_, new_n300_, new_n544_ );
not g0558 ( new_n630_, new_n629_ );
and g0559 ( new_n631_, new_n628_, new_n630_ );
and g0560 ( new_n632_, new_n631_, G53gat );
not g0561 ( new_n633_, new_n632_ );
and g0562 ( new_n634_, new_n633_, new_n321_ );
or g0563 ( new_n635_, new_n627_, new_n634_ );
and g0564 ( new_n636_, new_n635_, new_n187_ );
or g0565 ( new_n637_, new_n618_, new_n636_ );
and g0566 ( new_n638_, new_n637_, G43gat );
and g0567 ( new_n639_, new_n590_, new_n291_ );
or g0568 ( new_n640_, new_n638_, new_n639_ );
and g0569 ( new_n641_, new_n640_, G40gat );
not g0570 ( new_n642_, G40gat );
and g0571 ( new_n643_, new_n599_, G47gat );
or g0572 ( new_n644_, new_n616_, new_n643_ );
and g0573 ( new_n645_, new_n644_, G37gat );
or g0574 ( new_n646_, new_n645_, new_n636_ );
and g0575 ( new_n647_, new_n646_, G43gat );
and g0576 ( new_n648_, new_n599_, new_n291_ );
or g0577 ( new_n649_, new_n647_, new_n648_ );
and g0578 ( new_n650_, new_n649_, new_n642_ );
or g0579 ( new_n651_, new_n641_, new_n650_ );
and g0580 ( new_n652_, new_n651_, G34gat );
and g0581 ( new_n653_, new_n609_, G47gat );
or g0582 ( new_n654_, new_n616_, new_n653_ );
and g0583 ( new_n655_, new_n654_, G37gat );
or g0584 ( new_n656_, new_n655_, new_n636_ );
and g0585 ( new_n657_, new_n656_, G43gat );
and g0586 ( new_n658_, new_n609_, new_n291_ );
or g0587 ( new_n659_, new_n657_, new_n658_ );
and g0588 ( new_n660_, new_n659_, G40gat );
and g0589 ( new_n661_, new_n636_, G43gat );
and g0590 ( new_n662_, new_n613_, new_n189_ );
or g0591 ( new_n663_, new_n661_, new_n662_ );
and g0592 ( new_n664_, new_n663_, new_n642_ );
or g0593 ( new_n665_, new_n660_, new_n664_ );
and g0594 ( new_n666_, new_n665_, new_n317_ );
or g0595 ( new_n667_, new_n652_, new_n666_ );
and g0596 ( new_n668_, new_n667_, G24gat );
and g0597 ( new_n669_, new_n620_, new_n189_ );
or g0598 ( new_n670_, new_n661_, new_n669_ );
and g0599 ( new_n671_, new_n670_, G40gat );
or g0600 ( new_n672_, new_n624_, new_n322_ );
and g0601 ( new_n673_, new_n632_, new_n322_ );
not g0602 ( new_n674_, new_n673_ );
and g0603 ( new_n675_, new_n672_, new_n674_ );
and g0604 ( new_n676_, new_n675_, new_n642_ );
or g0605 ( new_n677_, new_n671_, new_n676_ );
and g0606 ( new_n678_, new_n677_, G34gat );
and g0607 ( new_n679_, new_n321_, new_n592_ );
and g0608 ( new_n680_, new_n679_, new_n188_ );
not g0609 ( new_n681_, new_n680_ );
and g0610 ( new_n682_, new_n631_, new_n681_ );
and g0611 ( new_n683_, new_n682_, G40gat );
not g0612 ( new_n684_, new_n683_ );
and g0613 ( new_n685_, new_n684_, new_n317_ );
or g0614 ( new_n686_, new_n678_, new_n685_ );
and g0615 ( new_n687_, new_n686_, new_n191_ );
or g0616 ( new_n688_, new_n668_, new_n687_ );
and g0617 ( new_n689_, new_n688_, G30gat );
and g0618 ( new_n690_, new_n640_, new_n308_ );
or g0619 ( new_n691_, new_n689_, new_n690_ );
and g0620 ( new_n692_, new_n691_, G27gat );
not g0621 ( new_n693_, G27gat );
and g0622 ( new_n694_, new_n649_, G34gat );
or g0623 ( new_n695_, new_n666_, new_n694_ );
and g0624 ( new_n696_, new_n695_, G24gat );
or g0625 ( new_n697_, new_n696_, new_n687_ );
and g0626 ( new_n698_, new_n697_, G30gat );
and g0627 ( new_n699_, new_n649_, new_n308_ );
or g0628 ( new_n700_, new_n698_, new_n699_ );
and g0629 ( new_n701_, new_n700_, new_n693_ );
or g0630 ( new_n702_, new_n692_, new_n701_ );
and g0631 ( new_n703_, new_n702_, G14gat );
not g0632 ( new_n704_, G14gat );
and g0633 ( new_n705_, new_n700_, new_n704_ );
or g0634 ( new_n706_, new_n703_, new_n705_ );
and g0635 ( new_n707_, new_n706_, G21gat );
and g0636 ( new_n708_, new_n659_, G34gat );
or g0637 ( new_n709_, new_n666_, new_n708_ );
and g0638 ( new_n710_, new_n709_, G24gat );
or g0639 ( new_n711_, new_n710_, new_n687_ );
and g0640 ( new_n712_, new_n711_, G30gat );
and g0641 ( new_n713_, new_n659_, new_n308_ );
or g0642 ( new_n714_, new_n712_, new_n713_ );
and g0643 ( new_n715_, new_n714_, G27gat );
and g0644 ( new_n716_, new_n687_, G30gat );
and g0645 ( new_n717_, new_n663_, new_n193_ );
or g0646 ( new_n718_, new_n716_, new_n717_ );
and g0647 ( new_n719_, new_n718_, new_n693_ );
or g0648 ( new_n720_, new_n715_, new_n719_ );
and g0649 ( new_n721_, new_n720_, new_n338_ );
or g0650 ( new_n722_, new_n707_, new_n721_ );
and g0651 ( new_n723_, new_n722_, G8gat );
and g0652 ( new_n724_, new_n720_, G14gat );
and g0653 ( new_n725_, new_n718_, new_n704_ );
or g0654 ( new_n726_, new_n724_, new_n725_ );
and g0655 ( new_n727_, new_n726_, new_n338_ );
and g0656 ( new_n728_, new_n714_, G14gat );
or g0657 ( new_n729_, new_n728_, new_n725_ );
and g0658 ( new_n730_, new_n729_, G21gat );
or g0659 ( new_n731_, new_n727_, new_n730_ );
and g0660 ( new_n732_, new_n731_, new_n354_ );
or g0661 ( new_n733_, new_n723_, new_n732_ );
and g0662 ( new_n734_, new_n733_, G11gat );
and g0663 ( new_n735_, new_n670_, new_n193_ );
or g0664 ( new_n736_, new_n716_, new_n735_ );
and g0665 ( new_n737_, new_n736_, G27gat );
or g0666 ( new_n738_, new_n675_, new_n344_ );
and g0667 ( new_n739_, new_n683_, new_n344_ );
not g0668 ( new_n740_, new_n739_ );
and g0669 ( new_n741_, new_n738_, new_n740_ );
and g0670 ( new_n742_, new_n741_, new_n693_ );
or g0671 ( new_n743_, new_n737_, new_n742_ );
and g0672 ( new_n744_, new_n743_, G21gat );
and g0673 ( new_n745_, new_n317_, new_n642_ );
and g0674 ( new_n746_, new_n745_, new_n192_ );
not g0675 ( new_n747_, new_n746_ );
and g0676 ( new_n748_, new_n682_, new_n747_ );
and g0677 ( new_n749_, new_n748_, G27gat );
not g0678 ( new_n750_, new_n749_ );
and g0679 ( new_n751_, new_n750_, new_n338_ );
or g0680 ( new_n752_, new_n744_, new_n751_ );
and g0681 ( new_n753_, new_n752_, new_n195_ );
or g0682 ( new_n754_, new_n734_, new_n753_ );
and g0683 ( new_n755_, new_n754_, G17gat );
and g0684 ( new_n756_, new_n691_, G14gat );
or g0685 ( new_n757_, new_n756_, new_n705_ );
and g0686 ( new_n758_, new_n757_, G8gat );
and g0687 ( new_n759_, new_n729_, new_n354_ );
or g0688 ( new_n760_, new_n758_, new_n759_ );
and g0689 ( new_n761_, new_n760_, new_n332_ );
or g0690 ( new_n762_, new_n755_, new_n761_ );
and g0691 ( new_n763_, new_n762_, G1gat );
and g0692 ( new_n764_, G21gat, G27gat );
or g0693 ( new_n765_, new_n197_, new_n764_ );
and g0694 ( new_n766_, G8gat, G14gat );
and g0695 ( new_n767_, new_n765_, new_n766_ );
and g0696 ( new_n768_, new_n736_, new_n767_ );
and g0697 ( new_n769_, new_n742_, G8gat );
or g0698 ( new_n770_, new_n769_, new_n751_ );
and g0699 ( new_n771_, new_n770_, new_n196_ );
and g0700 ( new_n772_, new_n359_, new_n704_ );
and g0701 ( new_n773_, new_n741_, new_n772_ );
and g0702 ( new_n774_, new_n748_, G14gat );
not g0703 ( new_n775_, new_n774_ );
and g0704 ( new_n776_, new_n775_, new_n354_ );
or g0705 ( new_n777_, new_n773_, new_n776_ );
or g0706 ( new_n778_, new_n771_, new_n777_ );
or g0707 ( new_n779_, new_n768_, new_n778_ );
and g0708 ( new_n780_, new_n779_, new_n358_ );
or g0709 ( new_n781_, new_n763_, new_n780_ );
and g0710 ( new_n782_, new_n781_, G4gat );
and g0711 ( new_n783_, new_n702_, G21gat );
or g0712 ( new_n784_, new_n783_, new_n721_ );
and g0713 ( new_n785_, new_n784_, G11gat );
or g0714 ( new_n786_, new_n785_, new_n753_ );
and g0715 ( new_n787_, new_n786_, G17gat );
and g0716 ( new_n788_, new_n691_, new_n332_ );
or g0717 ( new_n789_, new_n787_, new_n788_ );
and g0718 ( new_n790_, new_n789_, new_n198_ );
or g0719 ( new_n791_, new_n782_, new_n790_ );
and g0720 ( new_n792_, new_n791_, keyinput0_G370gat );
not g0721 ( new_n793_, keyinput0_G370gat );
and g0722 ( new_n794_, new_n75_, new_n793_ );
or g0723 ( new_n795_, new_n792_, new_n794_ );
and g0724 ( new_n796_, new_n795_, keyinput1_G370gat );
not g0725 ( new_n797_, keyinput1_G370gat );
and g0726 ( new_n798_, new_n425_, new_n793_ );
and g0727 ( new_n799_, new_n82_, keyinput0_G370gat );
or g0728 ( new_n800_, new_n798_, new_n799_ );
and g0729 ( new_n801_, new_n800_, new_n797_ );
or g0730 ( new_n802_, new_n796_, new_n801_ );
and g0731 ( new_n803_, new_n802_, keyinput2_G370gat );
not g0732 ( new_n804_, keyinput2_G370gat );
and g0733 ( new_n805_, new_n118_, new_n793_ );
not g0734 ( new_n806_, new_n178_ );
and g0735 ( new_n807_, new_n806_, keyinput0_G370gat );
or g0736 ( new_n808_, new_n805_, new_n807_ );
and g0737 ( new_n809_, new_n808_, new_n797_ );
and g0738 ( new_n810_, new_n116_, new_n793_ );
not g0739 ( new_n811_, new_n810_ );
not g0740 ( new_n812_, new_n799_ );
and g0741 ( new_n813_, new_n812_, keyinput1_G370gat );
and g0742 ( new_n814_, new_n811_, new_n813_ );
or g0743 ( new_n815_, new_n809_, new_n814_ );
and g0744 ( new_n816_, new_n815_, new_n804_ );
or g0745 ( new_n817_, new_n803_, new_n816_ );
and g0746 ( new_n818_, new_n817_, keyinput3_G370gat );
not g0747 ( new_n819_, keyinput3_G370gat );
and g0748 ( new_n820_, new_n160_, G95gat );
and g0749 ( new_n821_, new_n154_, new_n162_ );
or g0750 ( new_n822_, new_n820_, new_n821_ );
and g0751 ( new_n823_, new_n822_, new_n793_ );
not g0752 ( new_n824_, new_n186_ );
and g0753 ( new_n825_, new_n824_, keyinput0_G370gat );
or g0754 ( new_n826_, new_n823_, new_n825_ );
and g0755 ( new_n827_, new_n826_, new_n797_ );
and g0756 ( new_n828_, new_n89_, new_n793_ );
or g0757 ( new_n829_, new_n828_, new_n799_ );
and g0758 ( new_n830_, new_n829_, keyinput1_G370gat );
or g0759 ( new_n831_, new_n827_, new_n830_ );
and g0760 ( new_n832_, new_n831_, keyinput2_G370gat );
and g0761 ( new_n833_, new_n79_, keyinput0_G370gat );
and g0762 ( new_n834_, new_n100_, new_n793_ );
or g0763 ( new_n835_, new_n833_, new_n834_ );
and g0764 ( new_n836_, new_n835_, new_n797_ );
and g0765 ( new_n837_, new_n80_, new_n793_ );
or g0766 ( new_n838_, new_n108_, new_n837_ );
and g0767 ( new_n839_, new_n838_, keyinput1_G370gat );
or g0768 ( new_n840_, new_n836_, new_n839_ );
and g0769 ( new_n841_, new_n840_, new_n804_ );
or g0770 ( new_n842_, new_n832_, new_n841_ );
and g0771 ( new_n843_, new_n842_, new_n819_ );
or g0772 ( G370gat, new_n818_, new_n843_ );
not g0773 ( new_n845_, new_n347_ );
and g0774 ( new_n846_, new_n845_, G8gat );
or g0775 ( new_n847_, new_n846_, G14gat );
and g0776 ( new_n848_, new_n748_, new_n354_ );
not g0777 ( new_n849_, new_n848_ );
and g0778 ( new_n850_, G60gat, G66gat );
or g0779 ( new_n851_, new_n185_, new_n850_ );
not g0780 ( new_n852_, new_n851_ );
and g0781 ( new_n853_, G99gat, G105gat );
or g0782 ( new_n854_, new_n173_, new_n853_ );
not g0783 ( new_n855_, new_n854_ );
or g0784 ( new_n856_, new_n852_, new_n855_ );
and g0785 ( new_n857_, G73gat, G79gat );
or g0786 ( new_n858_, new_n181_, new_n857_ );
not g0787 ( new_n859_, new_n858_ );
and g0788 ( new_n860_, G47gat, G53gat );
or g0789 ( new_n861_, new_n189_, new_n860_ );
not g0790 ( new_n862_, new_n861_ );
or g0791 ( new_n863_, new_n859_, new_n862_ );
or g0792 ( new_n864_, new_n856_, new_n863_ );
not g0793 ( new_n865_, new_n766_ );
or g0794 ( new_n866_, new_n126_, new_n865_ );
and g0795 ( new_n867_, G86gat, G92gat );
or g0796 ( new_n868_, new_n177_, new_n867_ );
not g0797 ( new_n869_, new_n868_ );
and g0798 ( new_n870_, G34gat, G40gat );
or g0799 ( new_n871_, new_n193_, new_n870_ );
not g0800 ( new_n872_, new_n871_ );
or g0801 ( new_n873_, new_n869_, new_n872_ );
or g0802 ( new_n874_, new_n873_, new_n866_ );
or g0803 ( new_n875_, new_n874_, new_n474_ );
or g0804 ( new_n876_, new_n875_, new_n864_ );
and g0805 ( new_n877_, new_n849_, new_n876_ );
and g0806 ( new_n878_, new_n877_, new_n847_ );
and g0807 ( new_n879_, new_n693_, G14gat );
or g0808 ( new_n880_, new_n879_, G8gat );
and g0809 ( new_n881_, new_n880_, new_n338_ );
and g0810 ( new_n882_, new_n879_, G8gat );
or g0811 ( new_n883_, new_n881_, new_n882_ );
and g0812 ( new_n884_, new_n883_, new_n196_ );
or g0813 ( new_n885_, new_n884_, G1gat );
or g0814 ( new_n886_, new_n878_, new_n885_ );
not g0815 ( new_n887_, new_n194_ );
and g0816 ( new_n888_, new_n887_, new_n704_ );
not g0817 ( new_n889_, new_n679_ );
and g0818 ( new_n890_, new_n889_, G37gat );
or g0819 ( new_n891_, new_n890_, new_n291_ );
or g0820 ( new_n892_, new_n396_, new_n162_ );
and g0821 ( new_n893_, new_n282_, new_n544_ );
not g0822 ( new_n894_, new_n893_ );
and g0823 ( new_n895_, new_n894_, G50gat );
or g0824 ( new_n896_, new_n895_, new_n273_ );
and g0825 ( new_n897_, new_n892_, new_n896_ );
and g0826 ( new_n898_, new_n897_, new_n891_ );
not g0827 ( new_n899_, new_n530_ );
and g0828 ( new_n900_, new_n899_, G76gat );
or g0829 ( new_n901_, new_n900_, new_n253_ );
not g0830 ( new_n902_, new_n580_ );
and g0831 ( new_n903_, new_n902_, G63gat );
or g0832 ( new_n904_, new_n903_, new_n266_ );
and g0833 ( new_n905_, new_n901_, new_n904_ );
or g0834 ( new_n906_, new_n745_, new_n191_ );
and g0835 ( new_n907_, new_n906_, G30gat );
not g0836 ( new_n908_, new_n907_ );
and g0837 ( new_n909_, new_n908_, new_n78_ );
and g0838 ( new_n910_, new_n905_, new_n909_ );
and g0839 ( new_n911_, new_n910_, new_n898_ );
not g0840 ( new_n912_, new_n911_ );
and g0841 ( new_n913_, new_n912_, G14gat );
or g0842 ( new_n914_, new_n888_, new_n913_ );
and g0843 ( new_n915_, new_n914_, new_n354_ );
and g0844 ( new_n916_, new_n867_, G76gat );
or g0845 ( new_n917_, new_n916_, new_n253_ );
and g0846 ( new_n918_, new_n857_, G63gat );
or g0847 ( new_n919_, new_n918_, new_n266_ );
and g0848 ( new_n920_, new_n917_, new_n919_ );
and g0849 ( new_n921_, new_n220_, new_n920_ );
and g0850 ( new_n922_, new_n274_, G66gat );
or g0851 ( new_n923_, new_n922_, new_n273_ );
and g0852 ( new_n924_, new_n309_, G40gat );
or g0853 ( new_n925_, new_n924_, new_n308_ );
and g0854 ( new_n926_, new_n292_, G53gat );
or g0855 ( new_n927_, new_n926_, new_n291_ );
and g0856 ( new_n928_, new_n925_, new_n927_ );
and g0857 ( new_n929_, new_n928_, new_n923_ );
and g0858 ( new_n930_, new_n921_, new_n929_ );
not g0859 ( new_n931_, new_n930_ );
and g0860 ( new_n932_, new_n931_, G14gat );
and g0861 ( new_n933_, G63gat, G73gat );
or g0862 ( new_n934_, new_n933_, new_n266_ );
and g0863 ( new_n935_, G76gat, G86gat );
or g0864 ( new_n936_, new_n935_, new_n253_ );
and g0865 ( new_n937_, new_n934_, new_n936_ );
and g0866 ( new_n938_, new_n164_, new_n937_ );
and g0867 ( new_n939_, new_n275_, new_n293_ );
and g0868 ( new_n940_, new_n939_, new_n310_ );
and g0869 ( new_n941_, new_n938_, new_n940_ );
not g0870 ( new_n942_, new_n941_ );
and g0871 ( new_n943_, new_n942_, new_n704_ );
or g0872 ( new_n944_, new_n932_, new_n943_ );
and g0873 ( new_n945_, new_n944_, G8gat );
or g0874 ( new_n946_, new_n883_, new_n195_ );
and g0875 ( new_n947_, new_n946_, G17gat );
or g0876 ( new_n948_, new_n947_, new_n358_ );
or g0877 ( new_n949_, new_n945_, new_n948_ );
or g0878 ( new_n950_, new_n915_, new_n949_ );
and g0879 ( new_n951_, new_n950_, G4gat );
and g0880 ( new_n952_, new_n886_, new_n951_ );
or g0881 ( new_n953_, G69gat, G82gat );
or g0882 ( new_n954_, G95gat, G108gat );
or g0883 ( new_n955_, new_n953_, new_n954_ );
or g0884 ( new_n956_, G17gat, G30gat );
or g0885 ( new_n957_, G43gat, G56gat );
or g0886 ( new_n958_, new_n956_, new_n957_ );
or g0887 ( new_n959_, new_n955_, new_n958_ );
and g0888 ( new_n960_, new_n959_, new_n198_ );
or g0889 ( new_n961_, new_n952_, new_n960_ );
and g0890 ( new_n962_, new_n961_, keyinput3_G421gat );
not g0891 ( new_n963_, keyinput3_G421gat );
and g0892 ( new_n964_, new_n160_, new_n963_ );
or g0893 ( new_n965_, new_n962_, new_n964_ );
and g0894 ( new_n966_, new_n965_, keyinput2_G421gat );
not g0895 ( new_n967_, keyinput2_G421gat );
and g0896 ( new_n968_, new_n119_, new_n963_ );
and g0897 ( new_n969_, new_n115_, keyinput3_G421gat );
or g0898 ( new_n970_, new_n968_, new_n969_ );
and g0899 ( new_n971_, new_n970_, new_n967_ );
or g0900 ( new_n972_, new_n966_, new_n971_ );
and g0901 ( new_n973_, new_n972_, keyinput1_G421gat );
not g0902 ( new_n974_, keyinput1_G421gat );
and g0903 ( new_n975_, new_n141_, new_n963_ );
and g0904 ( new_n976_, new_n106_, keyinput3_G421gat );
or g0905 ( new_n977_, new_n975_, new_n976_ );
and g0906 ( new_n978_, new_n977_, keyinput2_G421gat );
and g0907 ( new_n979_, new_n220_, keyinput3_G421gat );
and g0908 ( new_n980_, new_n129_, new_n963_ );
or g0909 ( new_n981_, new_n979_, new_n980_ );
and g0910 ( new_n982_, new_n981_, new_n967_ );
or g0911 ( new_n983_, new_n978_, new_n982_ );
and g0912 ( new_n984_, new_n983_, new_n974_ );
or g0913 ( new_n985_, new_n973_, new_n984_ );
and g0914 ( new_n986_, new_n985_, keyinput0_G421gat );
not g0915 ( new_n987_, keyinput0_G421gat );
and g0916 ( new_n988_, new_n147_, new_n963_ );
and g0917 ( new_n989_, new_n75_, keyinput3_G421gat );
or g0918 ( new_n990_, new_n988_, new_n989_ );
and g0919 ( new_n991_, new_n990_, keyinput2_G421gat );
and g0920 ( new_n992_, new_n131_, new_n963_ );
and g0921 ( new_n993_, new_n91_, keyinput3_G421gat );
or g0922 ( new_n994_, new_n992_, new_n993_ );
and g0923 ( new_n995_, new_n994_, new_n967_ );
or g0924 ( new_n996_, new_n991_, new_n995_ );
and g0925 ( new_n997_, new_n996_, new_n974_ );
and g0926 ( new_n998_, new_n213_, keyinput3_G421gat );
and g0927 ( new_n999_, new_n91_, new_n963_ );
or g0928 ( new_n1000_, new_n998_, new_n999_ );
and g0929 ( new_n1001_, new_n1000_, new_n967_ );
or g0930 ( new_n1002_, new_n164_, keyinput3_G421gat );
not g0931 ( new_n1003_, new_n989_ );
and g0932 ( new_n1004_, new_n1003_, keyinput2_G421gat );
and g0933 ( new_n1005_, new_n1002_, new_n1004_ );
or g0934 ( new_n1006_, new_n1001_, new_n1005_ );
and g0935 ( new_n1007_, new_n1006_, keyinput1_G421gat );
or g0936 ( new_n1008_, new_n997_, new_n1007_ );
and g0937 ( new_n1009_, new_n1008_, new_n987_ );
or g0938 ( G421gat, new_n986_, new_n1009_ );
or g0939 ( new_n1011_, new_n628_, new_n544_ );
and g0940 ( new_n1012_, new_n1011_, new_n282_ );
and g0941 ( new_n1013_, new_n285_, new_n544_ );
or g0942 ( new_n1014_, new_n1012_, new_n1013_ );
and g0943 ( new_n1015_, new_n97_, new_n854_ );
and g0944 ( new_n1016_, new_n858_, new_n868_ );
and g0945 ( new_n1017_, new_n1015_, new_n1016_ );
and g0946 ( new_n1018_, new_n1017_, new_n850_ );
or g0947 ( new_n1019_, new_n1014_, new_n1018_ );
and g0948 ( new_n1020_, new_n1019_, new_n183_ );
and g0949 ( new_n1021_, new_n892_, new_n78_ );
and g0950 ( new_n1022_, new_n905_, G66gat );
and g0951 ( new_n1023_, new_n1022_, new_n1021_ );
and g0952 ( new_n1024_, new_n182_, new_n544_ );
or g0953 ( new_n1025_, new_n1023_, new_n1024_ );
and g0954 ( new_n1026_, new_n1025_, new_n282_ );
and g0955 ( new_n1027_, new_n921_, G66gat );
and g0956 ( new_n1028_, new_n938_, new_n544_ );
or g0957 ( new_n1029_, new_n1027_, new_n1028_ );
and g0958 ( new_n1030_, new_n1029_, G60gat );
or g0959 ( new_n1031_, new_n1026_, new_n1030_ );
and g0960 ( new_n1032_, new_n1031_, G50gat );
or g0961 ( new_n1033_, new_n1020_, new_n1032_ );
and g0962 ( new_n1034_, new_n1033_, G56gat );
and g0963 ( new_n1035_, new_n921_, new_n273_ );
or g0964 ( new_n1036_, new_n1034_, new_n1035_ );
and g0965 ( new_n1037_, new_n1036_, G53gat );
and g0966 ( new_n1038_, new_n938_, G60gat );
or g0967 ( new_n1039_, new_n1026_, new_n1038_ );
and g0968 ( new_n1040_, new_n1039_, G50gat );
or g0969 ( new_n1041_, new_n1020_, new_n1040_ );
and g0970 ( new_n1042_, new_n1041_, G56gat );
and g0971 ( new_n1043_, new_n938_, new_n273_ );
or g0972 ( new_n1044_, new_n1042_, new_n1043_ );
and g0973 ( new_n1045_, new_n1044_, new_n592_ );
or g0974 ( new_n1046_, new_n1037_, new_n1045_ );
and g0975 ( new_n1047_, new_n1046_, G47gat );
and g0976 ( new_n1048_, new_n905_, G60gat );
and g0977 ( new_n1049_, new_n1048_, new_n1021_ );
or g0978 ( new_n1050_, new_n1026_, new_n1049_ );
and g0979 ( new_n1051_, new_n1050_, G50gat );
or g0980 ( new_n1052_, new_n1020_, new_n1051_ );
and g0981 ( new_n1053_, new_n1052_, G56gat );
and g0982 ( new_n1054_, new_n905_, new_n273_ );
and g0983 ( new_n1055_, new_n1054_, new_n1021_ );
or g0984 ( new_n1056_, new_n1053_, new_n1055_ );
or g0985 ( new_n1057_, new_n1056_, new_n592_ );
and g0986 ( new_n1058_, new_n1020_, G56gat );
or g0987 ( new_n1059_, new_n1058_, new_n186_ );
or g0988 ( new_n1060_, new_n1059_, G53gat );
and g0989 ( new_n1061_, new_n1060_, new_n321_ );
and g0990 ( new_n1062_, new_n1057_, new_n1061_ );
or g0991 ( new_n1063_, new_n1047_, new_n1062_ );
and g0992 ( new_n1064_, new_n1063_, G37gat );
and g0993 ( new_n1065_, new_n1017_, new_n185_ );
or g0994 ( new_n1066_, new_n1058_, new_n1065_ );
and g0995 ( new_n1067_, new_n1066_, G53gat );
and g0996 ( new_n1068_, new_n1011_, new_n300_ );
or g0997 ( new_n1069_, new_n1068_, new_n302_ );
and g0998 ( new_n1070_, new_n1069_, new_n592_ );
or g0999 ( new_n1071_, new_n1067_, new_n1070_ );
and g1000 ( new_n1072_, new_n1071_, G47gat );
or g1001 ( new_n1073_, new_n628_, new_n629_ );
or g1002 ( new_n1074_, new_n1073_, new_n592_ );
and g1003 ( new_n1075_, new_n1074_, new_n321_ );
or g1004 ( new_n1076_, new_n1072_, new_n1075_ );
and g1005 ( new_n1077_, new_n1076_, new_n187_ );
or g1006 ( new_n1078_, new_n1064_, new_n1077_ );
and g1007 ( new_n1079_, new_n1078_, G43gat );
and g1008 ( new_n1080_, new_n1036_, new_n291_ );
or g1009 ( new_n1081_, new_n1079_, new_n1080_ );
and g1010 ( new_n1082_, new_n1081_, G40gat );
and g1011 ( new_n1083_, new_n1044_, G47gat );
or g1012 ( new_n1084_, new_n1062_, new_n1083_ );
and g1013 ( new_n1085_, new_n1084_, G37gat );
or g1014 ( new_n1086_, new_n1085_, new_n1077_ );
and g1015 ( new_n1087_, new_n1086_, G43gat );
and g1016 ( new_n1088_, new_n1044_, new_n291_ );
or g1017 ( new_n1089_, new_n1087_, new_n1088_ );
and g1018 ( new_n1090_, new_n1089_, new_n642_ );
or g1019 ( new_n1091_, new_n1082_, new_n1090_ );
and g1020 ( new_n1092_, new_n1091_, G34gat );
and g1021 ( new_n1093_, new_n1056_, G47gat );
or g1022 ( new_n1094_, new_n1062_, new_n1093_ );
and g1023 ( new_n1095_, new_n1094_, G37gat );
or g1024 ( new_n1096_, new_n1095_, new_n1077_ );
and g1025 ( new_n1097_, new_n1096_, G43gat );
and g1026 ( new_n1098_, new_n1056_, new_n291_ );
or g1027 ( new_n1099_, new_n1097_, new_n1098_ );
or g1028 ( new_n1100_, new_n1099_, new_n642_ );
and g1029 ( new_n1101_, new_n1077_, G43gat );
and g1030 ( new_n1102_, new_n1059_, new_n189_ );
or g1031 ( new_n1103_, new_n1101_, new_n1102_ );
or g1032 ( new_n1104_, new_n1103_, G40gat );
and g1033 ( new_n1105_, new_n1104_, new_n317_ );
and g1034 ( new_n1106_, new_n1100_, new_n1105_ );
or g1035 ( new_n1107_, new_n1092_, new_n1106_ );
and g1036 ( new_n1108_, new_n1107_, G24gat );
and g1037 ( new_n1109_, new_n1066_, new_n189_ );
or g1038 ( new_n1110_, new_n1101_, new_n1109_ );
and g1039 ( new_n1111_, new_n1110_, G40gat );
or g1040 ( new_n1112_, new_n1069_, new_n322_ );
or g1041 ( new_n1113_, new_n1074_, new_n323_ );
and g1042 ( new_n1114_, new_n1112_, new_n1113_ );
and g1043 ( new_n1115_, new_n1114_, new_n642_ );
or g1044 ( new_n1116_, new_n1111_, new_n1115_ );
and g1045 ( new_n1117_, new_n1116_, G34gat );
or g1046 ( new_n1118_, new_n1073_, new_n680_ );
or g1047 ( new_n1119_, new_n1118_, new_n642_ );
and g1048 ( new_n1120_, new_n1119_, new_n317_ );
or g1049 ( new_n1121_, new_n1117_, new_n1120_ );
and g1050 ( new_n1122_, new_n1121_, new_n191_ );
or g1051 ( new_n1123_, new_n1108_, new_n1122_ );
and g1052 ( new_n1124_, new_n1123_, G30gat );
and g1053 ( new_n1125_, new_n1081_, new_n308_ );
or g1054 ( new_n1126_, new_n1124_, new_n1125_ );
and g1055 ( new_n1127_, new_n1126_, G14gat );
and g1056 ( new_n1128_, new_n1028_, G60gat );
or g1057 ( new_n1129_, new_n1026_, new_n1128_ );
and g1058 ( new_n1130_, new_n1129_, G50gat );
or g1059 ( new_n1131_, new_n1020_, new_n1130_ );
and g1060 ( new_n1132_, new_n1131_, G56gat );
and g1061 ( new_n1133_, new_n1132_, G53gat );
or g1062 ( new_n1134_, new_n1045_, new_n1133_ );
and g1063 ( new_n1135_, new_n1134_, G47gat );
or g1064 ( new_n1136_, new_n1135_, new_n1062_ );
and g1065 ( new_n1137_, new_n1136_, G37gat );
or g1066 ( new_n1138_, new_n1137_, new_n1077_ );
and g1067 ( new_n1139_, new_n1138_, G43gat );
and g1068 ( new_n1140_, new_n1132_, new_n291_ );
or g1069 ( new_n1141_, new_n1139_, new_n1140_ );
and g1070 ( new_n1142_, new_n1141_, G40gat );
or g1071 ( new_n1143_, new_n1142_, new_n1090_ );
and g1072 ( new_n1144_, new_n1143_, G34gat );
or g1073 ( new_n1145_, new_n1144_, new_n1106_ );
and g1074 ( new_n1146_, new_n1145_, G24gat );
or g1075 ( new_n1147_, new_n1146_, new_n1122_ );
and g1076 ( new_n1148_, new_n1147_, G30gat );
and g1077 ( new_n1149_, new_n1141_, new_n308_ );
or g1078 ( new_n1150_, new_n1148_, new_n1149_ );
and g1079 ( new_n1151_, new_n1150_, new_n704_ );
or g1080 ( new_n1152_, new_n1127_, new_n1151_ );
and g1081 ( new_n1153_, new_n1152_, G27gat );
and g1082 ( new_n1154_, new_n1089_, G34gat );
or g1083 ( new_n1155_, new_n1106_, new_n1154_ );
and g1084 ( new_n1156_, new_n1155_, G24gat );
or g1085 ( new_n1157_, new_n1156_, new_n1122_ );
and g1086 ( new_n1158_, new_n1157_, G30gat );
and g1087 ( new_n1159_, new_n1089_, new_n308_ );
or g1088 ( new_n1160_, new_n1158_, new_n1159_ );
and g1089 ( new_n1161_, new_n1160_, new_n693_ );
or g1090 ( new_n1162_, new_n1153_, new_n1161_ );
and g1091 ( new_n1163_, new_n1162_, G21gat );
and g1092 ( new_n1164_, new_n1099_, G34gat );
or g1093 ( new_n1165_, new_n1106_, new_n1164_ );
and g1094 ( new_n1166_, new_n1165_, G24gat );
or g1095 ( new_n1167_, new_n1166_, new_n1122_ );
and g1096 ( new_n1168_, new_n1167_, G30gat );
and g1097 ( new_n1169_, new_n1099_, new_n308_ );
or g1098 ( new_n1170_, new_n1168_, new_n1169_ );
and g1099 ( new_n1171_, new_n1170_, G27gat );
and g1100 ( new_n1172_, new_n1122_, G30gat );
and g1101 ( new_n1173_, new_n1103_, new_n193_ );
or g1102 ( new_n1174_, new_n1172_, new_n1173_ );
and g1103 ( new_n1175_, new_n1174_, new_n693_ );
or g1104 ( new_n1176_, new_n1171_, new_n1175_ );
and g1105 ( new_n1177_, new_n1176_, new_n338_ );
or g1106 ( new_n1178_, new_n1163_, new_n1177_ );
and g1107 ( new_n1179_, new_n1178_, G8gat );
and g1108 ( new_n1180_, new_n1170_, G14gat );
or g1109 ( new_n1181_, new_n1060_, G47gat );
and g1110 ( new_n1182_, new_n282_, G50gat );
and g1111 ( new_n1183_, new_n1024_, new_n1182_ );
or g1112 ( new_n1184_, new_n1020_, new_n1183_ );
and g1113 ( new_n1185_, new_n1184_, G56gat );
or g1114 ( new_n1186_, new_n1185_, new_n679_ );
and g1115 ( new_n1187_, new_n1186_, G37gat );
and g1116 ( new_n1188_, new_n1181_, new_n1187_ );
or g1117 ( new_n1189_, new_n1077_, new_n1188_ );
and g1118 ( new_n1190_, new_n1189_, G43gat );
and g1119 ( new_n1191_, new_n1185_, new_n291_ );
or g1120 ( new_n1192_, new_n1190_, new_n1191_ );
or g1121 ( new_n1193_, new_n1192_, new_n745_ );
or g1122 ( new_n1194_, new_n1104_, G34gat );
and g1123 ( new_n1195_, new_n1194_, G24gat );
and g1124 ( new_n1196_, new_n1195_, new_n1193_ );
or g1125 ( new_n1197_, new_n1122_, new_n1196_ );
and g1126 ( new_n1198_, new_n1197_, G30gat );
and g1127 ( new_n1199_, new_n1192_, new_n308_ );
or g1128 ( new_n1200_, new_n1198_, new_n1199_ );
and g1129 ( new_n1201_, new_n1200_, new_n704_ );
or g1130 ( new_n1202_, new_n1180_, new_n1201_ );
and g1131 ( new_n1203_, new_n1202_, G27gat );
or g1132 ( new_n1204_, new_n1203_, new_n1175_ );
and g1133 ( new_n1205_, new_n1204_, new_n338_ );
and g1134 ( new_n1206_, new_n1025_, new_n1182_ );
or g1135 ( new_n1207_, new_n1020_, new_n1206_ );
and g1136 ( new_n1208_, new_n1207_, G56gat );
and g1137 ( new_n1209_, new_n1208_, G47gat );
or g1138 ( new_n1210_, new_n1062_, new_n1209_ );
and g1139 ( new_n1211_, new_n1210_, G37gat );
or g1140 ( new_n1212_, new_n1211_, new_n1077_ );
and g1141 ( new_n1213_, new_n1212_, G43gat );
and g1142 ( new_n1214_, new_n1208_, new_n291_ );
or g1143 ( new_n1215_, new_n1213_, new_n1214_ );
and g1144 ( new_n1216_, new_n1215_, G34gat );
or g1145 ( new_n1217_, new_n1106_, new_n1216_ );
and g1146 ( new_n1218_, new_n1217_, G24gat );
or g1147 ( new_n1219_, new_n1218_, new_n1122_ );
and g1148 ( new_n1220_, new_n1219_, G30gat );
and g1149 ( new_n1221_, new_n1215_, new_n308_ );
or g1150 ( new_n1222_, new_n1220_, new_n1221_ );
and g1151 ( new_n1223_, new_n1222_, G14gat );
or g1152 ( new_n1224_, new_n1223_, new_n1201_ );
and g1153 ( new_n1225_, new_n1224_, G21gat );
or g1154 ( new_n1226_, new_n1205_, new_n1225_ );
and g1155 ( new_n1227_, new_n1226_, new_n354_ );
or g1156 ( new_n1228_, new_n1179_, new_n1227_ );
and g1157 ( new_n1229_, new_n1228_, G11gat );
and g1158 ( new_n1230_, new_n1110_, new_n193_ );
or g1159 ( new_n1231_, new_n1172_, new_n1230_ );
and g1160 ( new_n1232_, new_n1231_, G27gat );
or g1161 ( new_n1233_, new_n1114_, new_n344_ );
or g1162 ( new_n1234_, new_n1119_, new_n345_ );
and g1163 ( new_n1235_, new_n1234_, new_n693_ );
and g1164 ( new_n1236_, new_n1233_, new_n1235_ );
or g1165 ( new_n1237_, new_n1232_, new_n1236_ );
or g1166 ( new_n1238_, new_n1237_, new_n338_ );
or g1167 ( new_n1239_, new_n746_, new_n693_ );
or g1168 ( new_n1240_, new_n1118_, new_n1239_ );
or g1169 ( new_n1241_, new_n1240_, G21gat );
and g1170 ( new_n1242_, new_n1241_, new_n195_ );
and g1171 ( new_n1243_, new_n1238_, new_n1242_ );
or g1172 ( new_n1244_, new_n1229_, new_n1243_ );
and g1173 ( new_n1245_, new_n1244_, G17gat );
and g1174 ( new_n1246_, new_n1034_, new_n291_ );
or g1175 ( new_n1247_, new_n1079_, new_n1246_ );
and g1176 ( new_n1248_, new_n1247_, new_n308_ );
or g1177 ( new_n1249_, new_n1124_, new_n1248_ );
and g1178 ( new_n1250_, new_n1249_, G14gat );
or g1179 ( new_n1251_, new_n1250_, new_n1151_ );
and g1180 ( new_n1252_, new_n1251_, G8gat );
and g1181 ( new_n1253_, new_n1224_, new_n354_ );
or g1182 ( new_n1254_, new_n1252_, new_n1253_ );
and g1183 ( new_n1255_, new_n1254_, new_n332_ );
or g1184 ( new_n1256_, new_n1245_, new_n1255_ );
and g1185 ( new_n1257_, new_n1256_, G1gat );
and g1186 ( new_n1258_, new_n1237_, G14gat );
and g1187 ( new_n1259_, new_n1014_, new_n184_ );
and g1188 ( new_n1260_, new_n1259_, G53gat );
or g1189 ( new_n1261_, new_n1260_, new_n1070_ );
and g1190 ( new_n1262_, new_n1261_, G47gat );
or g1191 ( new_n1263_, new_n1262_, new_n1075_ );
and g1192 ( new_n1264_, new_n1263_, new_n188_ );
and g1193 ( new_n1265_, new_n1259_, new_n189_ );
or g1194 ( new_n1266_, new_n1264_, new_n1265_ );
and g1195 ( new_n1267_, new_n1266_, G40gat );
or g1196 ( new_n1268_, new_n1267_, new_n1115_ );
and g1197 ( new_n1269_, new_n1268_, G34gat );
or g1198 ( new_n1270_, new_n1120_, new_n193_ );
or g1199 ( new_n1271_, new_n1269_, new_n1270_ );
or g1200 ( new_n1272_, new_n1266_, new_n192_ );
and g1201 ( new_n1273_, new_n1271_, new_n1272_ );
and g1202 ( new_n1274_, new_n1273_, G27gat );
or g1203 ( new_n1275_, new_n1274_, new_n1236_ );
and g1204 ( new_n1276_, new_n1275_, new_n704_ );
or g1205 ( new_n1277_, new_n1276_, new_n338_ );
or g1206 ( new_n1278_, new_n1258_, new_n1277_ );
and g1207 ( new_n1279_, new_n1278_, new_n1241_ );
or g1208 ( new_n1280_, new_n1279_, new_n354_ );
and g1209 ( new_n1281_, new_n1075_, new_n188_ );
and g1210 ( new_n1282_, new_n1068_, new_n323_ );
or g1211 ( new_n1283_, new_n1282_, new_n344_ );
or g1212 ( new_n1284_, new_n1281_, new_n1283_ );
and g1213 ( new_n1285_, new_n1234_, G14gat );
and g1214 ( new_n1286_, new_n1284_, new_n1285_ );
and g1215 ( new_n1287_, new_n630_, new_n681_ );
not g1216 ( new_n1288_, new_n1287_ );
or g1217 ( new_n1289_, new_n1288_, new_n746_ );
and g1218 ( new_n1290_, new_n1289_, new_n704_ );
or g1219 ( new_n1291_, new_n1286_, new_n1290_ );
and g1220 ( new_n1292_, new_n1291_, G21gat );
and g1221 ( new_n1293_, new_n1240_, G14gat );
or g1222 ( new_n1294_, new_n1289_, new_n693_ );
and g1223 ( new_n1295_, new_n1294_, new_n704_ );
or g1224 ( new_n1296_, new_n1293_, new_n1295_ );
and g1225 ( new_n1297_, new_n1296_, new_n338_ );
or g1226 ( new_n1298_, new_n1297_, G8gat );
or g1227 ( new_n1299_, new_n1292_, new_n1298_ );
and g1228 ( new_n1300_, new_n1280_, new_n1299_ );
or g1229 ( new_n1301_, new_n1300_, new_n197_ );
and g1230 ( new_n1302_, new_n1058_, new_n189_ );
or g1231 ( new_n1303_, new_n1101_, new_n1302_ );
and g1232 ( new_n1304_, new_n1303_, new_n193_ );
or g1233 ( new_n1305_, new_n1172_, new_n1304_ );
and g1234 ( new_n1306_, new_n1305_, G14gat );
and g1235 ( new_n1307_, new_n1273_, new_n704_ );
or g1236 ( new_n1308_, new_n1307_, new_n354_ );
or g1237 ( new_n1309_, new_n1306_, new_n1308_ );
or g1238 ( new_n1310_, new_n1291_, G8gat );
and g1239 ( new_n1311_, new_n1309_, new_n1310_ );
or g1240 ( new_n1312_, new_n1311_, new_n196_ );
and g1241 ( new_n1313_, new_n1312_, new_n358_ );
and g1242 ( new_n1314_, new_n1301_, new_n1313_ );
or g1243 ( new_n1315_, new_n1257_, new_n1314_ );
and g1244 ( new_n1316_, new_n1315_, G4gat );
and g1245 ( new_n1317_, new_n1126_, G27gat );
or g1246 ( new_n1318_, new_n1317_, new_n1161_ );
and g1247 ( new_n1319_, new_n1318_, G21gat );
or g1248 ( new_n1320_, new_n1319_, new_n1177_ );
and g1249 ( new_n1321_, new_n1320_, G11gat );
or g1250 ( new_n1322_, new_n1321_, new_n1243_ );
and g1251 ( new_n1323_, new_n1322_, G17gat );
and g1252 ( new_n1324_, new_n1249_, new_n332_ );
or g1253 ( new_n1325_, new_n1323_, new_n1324_ );
and g1254 ( new_n1326_, new_n1325_, new_n198_ );
or g1255 ( new_n1327_, new_n1316_, new_n1326_ );
and g1256 ( new_n1328_, new_n1327_, keyinput0_G430gat );
not g1257 ( new_n1329_, keyinput0_G430gat );
and g1258 ( new_n1330_, new_n75_, new_n1329_ );
or g1259 ( new_n1331_, new_n1328_, new_n1330_ );
and g1260 ( new_n1332_, new_n1331_, keyinput1_G430gat );
not g1261 ( new_n1333_, keyinput1_G430gat );
and g1262 ( new_n1334_, new_n425_, new_n1329_ );
and g1263 ( new_n1335_, new_n82_, keyinput0_G430gat );
or g1264 ( new_n1336_, new_n1334_, new_n1335_ );
and g1265 ( new_n1337_, new_n1336_, new_n1333_ );
or g1266 ( new_n1338_, new_n1332_, new_n1337_ );
and g1267 ( new_n1339_, new_n1338_, keyinput2_G430gat );
not g1268 ( new_n1340_, keyinput2_G430gat );
and g1269 ( new_n1341_, new_n118_, new_n1329_ );
and g1270 ( new_n1342_, new_n806_, keyinput0_G430gat );
or g1271 ( new_n1343_, new_n1341_, new_n1342_ );
and g1272 ( new_n1344_, new_n1343_, new_n1333_ );
and g1273 ( new_n1345_, new_n116_, new_n1329_ );
not g1274 ( new_n1346_, new_n1345_ );
not g1275 ( new_n1347_, new_n1335_ );
and g1276 ( new_n1348_, new_n1347_, keyinput1_G430gat );
and g1277 ( new_n1349_, new_n1346_, new_n1348_ );
or g1278 ( new_n1350_, new_n1344_, new_n1349_ );
and g1279 ( new_n1351_, new_n1350_, new_n1340_ );
or g1280 ( new_n1352_, new_n1339_, new_n1351_ );
and g1281 ( new_n1353_, new_n1352_, keyinput3_G430gat );
not g1282 ( new_n1354_, keyinput3_G430gat );
and g1283 ( new_n1355_, new_n822_, new_n1329_ );
and g1284 ( new_n1356_, new_n824_, keyinput0_G430gat );
or g1285 ( new_n1357_, new_n1355_, new_n1356_ );
and g1286 ( new_n1358_, new_n1357_, new_n1333_ );
and g1287 ( new_n1359_, new_n89_, new_n1329_ );
or g1288 ( new_n1360_, new_n1359_, new_n1335_ );
and g1289 ( new_n1361_, new_n1360_, keyinput1_G430gat );
or g1290 ( new_n1362_, new_n1358_, new_n1361_ );
and g1291 ( new_n1363_, new_n1362_, keyinput2_G430gat );
and g1292 ( new_n1364_, new_n79_, keyinput0_G430gat );
and g1293 ( new_n1365_, new_n100_, new_n1329_ );
or g1294 ( new_n1366_, new_n1364_, new_n1365_ );
and g1295 ( new_n1367_, new_n1366_, new_n1333_ );
and g1296 ( new_n1368_, new_n80_, new_n1329_ );
or g1297 ( new_n1369_, new_n108_, new_n1368_ );
and g1298 ( new_n1370_, new_n1369_, keyinput1_G430gat );
or g1299 ( new_n1371_, new_n1367_, new_n1370_ );
and g1300 ( new_n1372_, new_n1371_, new_n1340_ );
or g1301 ( new_n1373_, new_n1363_, new_n1372_ );
and g1302 ( new_n1374_, new_n1373_, new_n1354_ );
or g1303 ( G430gat, new_n1353_, new_n1374_ );
and g1304 ( new_n1376_, new_n1021_, G92gat );
and g1305 ( new_n1377_, new_n174_, new_n445_ );
or g1306 ( new_n1378_, new_n1376_, new_n1377_ );
and g1307 ( new_n1379_, new_n1378_, new_n229_ );
and g1308 ( new_n1380_, new_n220_, G92gat );
and g1309 ( new_n1381_, new_n164_, new_n445_ );
or g1310 ( new_n1382_, new_n1380_, new_n1381_ );
and g1311 ( new_n1383_, new_n1382_, G86gat );
or g1312 ( new_n1384_, new_n1379_, new_n1383_ );
and g1313 ( new_n1385_, new_n1384_, G76gat );
and g1314 ( new_n1386_, new_n1015_, G92gat );
and g1315 ( new_n1387_, new_n232_, new_n445_ );
or g1316 ( new_n1388_, new_n1386_, new_n1387_ );
and g1317 ( new_n1389_, new_n1388_, G86gat );
or g1318 ( new_n1390_, new_n529_, new_n445_ );
and g1319 ( new_n1391_, new_n1390_, new_n229_ );
or g1320 ( new_n1392_, new_n1389_, new_n1391_ );
and g1321 ( new_n1393_, new_n1392_, new_n175_ );
or g1322 ( new_n1394_, new_n1385_, new_n1393_ );
and g1323 ( new_n1395_, new_n1394_, G82gat );
and g1324 ( new_n1396_, new_n220_, new_n253_ );
or g1325 ( new_n1397_, new_n1395_, new_n1396_ );
and g1326 ( new_n1398_, new_n1397_, G79gat );
and g1327 ( new_n1399_, new_n164_, G86gat );
or g1328 ( new_n1400_, new_n1379_, new_n1399_ );
and g1329 ( new_n1401_, new_n1400_, G76gat );
or g1330 ( new_n1402_, new_n1401_, new_n1393_ );
and g1331 ( new_n1403_, new_n1402_, G82gat );
and g1332 ( new_n1404_, new_n164_, new_n253_ );
or g1333 ( new_n1405_, new_n1403_, new_n1404_ );
and g1334 ( new_n1406_, new_n1405_, new_n493_ );
or g1335 ( new_n1407_, new_n1398_, new_n1406_ );
and g1336 ( new_n1408_, new_n1407_, G73gat );
and g1337 ( new_n1409_, new_n1021_, G86gat );
or g1338 ( new_n1410_, new_n1379_, new_n1409_ );
and g1339 ( new_n1411_, new_n1410_, G76gat );
or g1340 ( new_n1412_, new_n1411_, new_n1393_ );
and g1341 ( new_n1413_, new_n1412_, G82gat );
and g1342 ( new_n1414_, new_n1021_, new_n253_ );
or g1343 ( new_n1415_, new_n1413_, new_n1414_ );
or g1344 ( new_n1416_, new_n1415_, new_n493_ );
and g1345 ( new_n1417_, new_n1393_, G82gat );
or g1346 ( new_n1418_, new_n1417_, new_n178_ );
or g1347 ( new_n1419_, new_n1418_, G79gat );
and g1348 ( new_n1420_, new_n1419_, new_n257_ );
and g1349 ( new_n1421_, new_n1416_, new_n1420_ );
or g1350 ( new_n1422_, new_n1408_, new_n1421_ );
and g1351 ( new_n1423_, new_n1422_, G63gat );
and g1352 ( new_n1424_, new_n1015_, new_n177_ );
or g1353 ( new_n1425_, new_n1417_, new_n1424_ );
and g1354 ( new_n1426_, new_n1425_, G79gat );
and g1355 ( new_n1427_, new_n1391_, new_n176_ );
or g1356 ( new_n1428_, new_n1427_, new_n260_ );
and g1357 ( new_n1429_, new_n1428_, new_n493_ );
or g1358 ( new_n1430_, new_n1426_, new_n1429_ );
and g1359 ( new_n1431_, new_n1430_, G73gat );
or g1360 ( new_n1432_, new_n529_, new_n531_ );
or g1361 ( new_n1433_, new_n1432_, new_n493_ );
and g1362 ( new_n1434_, new_n1433_, new_n257_ );
or g1363 ( new_n1435_, new_n1431_, new_n1434_ );
and g1364 ( new_n1436_, new_n1435_, new_n179_ );
or g1365 ( new_n1437_, new_n1423_, new_n1436_ );
and g1366 ( new_n1438_, new_n1437_, G69gat );
and g1367 ( new_n1439_, new_n1397_, new_n266_ );
or g1368 ( new_n1440_, new_n1438_, new_n1439_ );
and g1369 ( new_n1441_, new_n1440_, G66gat );
and g1370 ( new_n1442_, new_n1379_, G76gat );
or g1371 ( new_n1443_, new_n1393_, new_n1442_ );
and g1372 ( new_n1444_, new_n1443_, G82gat );
and g1373 ( new_n1445_, new_n1444_, G73gat );
or g1374 ( new_n1446_, new_n1421_, new_n1445_ );
and g1375 ( new_n1447_, new_n1446_, G63gat );
or g1376 ( new_n1448_, new_n1447_, new_n1436_ );
and g1377 ( new_n1449_, new_n1448_, G69gat );
and g1378 ( new_n1450_, new_n1444_, new_n266_ );
or g1379 ( new_n1451_, new_n1449_, new_n1450_ );
and g1380 ( new_n1452_, new_n1451_, new_n544_ );
or g1381 ( new_n1453_, new_n1441_, new_n1452_ );
and g1382 ( new_n1454_, new_n1453_, G60gat );
or g1383 ( new_n1455_, new_n1419_, G73gat );
and g1384 ( new_n1456_, new_n229_, G76gat );
and g1385 ( new_n1457_, new_n1377_, new_n1456_ );
or g1386 ( new_n1458_, new_n1393_, new_n1457_ );
and g1387 ( new_n1459_, new_n1458_, G82gat );
or g1388 ( new_n1460_, new_n1459_, new_n580_ );
and g1389 ( new_n1461_, new_n1460_, G63gat );
and g1390 ( new_n1462_, new_n1455_, new_n1461_ );
or g1391 ( new_n1463_, new_n1436_, new_n1462_ );
and g1392 ( new_n1464_, new_n1463_, G69gat );
and g1393 ( new_n1465_, new_n1459_, new_n266_ );
or g1394 ( new_n1466_, new_n1464_, new_n1465_ );
and g1395 ( new_n1467_, new_n1466_, G66gat );
and g1396 ( new_n1468_, new_n1436_, G69gat );
and g1397 ( new_n1469_, new_n1417_, new_n181_ );
or g1398 ( new_n1470_, new_n1468_, new_n1469_ );
and g1399 ( new_n1471_, new_n1470_, new_n544_ );
or g1400 ( new_n1472_, new_n1467_, new_n1471_ );
and g1401 ( new_n1473_, new_n1472_, new_n282_ );
or g1402 ( new_n1474_, new_n1454_, new_n1473_ );
and g1403 ( new_n1475_, new_n1474_, G50gat );
or g1404 ( new_n1476_, new_n1434_, new_n858_ );
or g1405 ( new_n1477_, new_n1429_, new_n1476_ );
or g1406 ( new_n1478_, new_n1391_, new_n1387_ );
and g1407 ( new_n1479_, new_n1478_, new_n176_ );
or g1408 ( new_n1480_, new_n1479_, new_n859_ );
and g1409 ( new_n1481_, new_n1477_, new_n1480_ );
and g1410 ( new_n1482_, new_n1481_, G66gat );
and g1411 ( new_n1483_, new_n1427_, new_n284_ );
and g1412 ( new_n1484_, new_n1433_, new_n283_ );
or g1413 ( new_n1485_, new_n1483_, new_n1484_ );
and g1414 ( new_n1486_, new_n1485_, new_n544_ );
or g1415 ( new_n1487_, new_n1482_, new_n1486_ );
and g1416 ( new_n1488_, new_n1487_, G60gat );
or g1417 ( new_n1489_, new_n531_, new_n581_ );
and g1418 ( new_n1490_, new_n1489_, G66gat );
and g1419 ( new_n1491_, new_n1490_, new_n282_ );
or g1420 ( new_n1492_, new_n1488_, new_n1491_ );
and g1421 ( new_n1493_, new_n1492_, new_n183_ );
or g1422 ( new_n1494_, new_n1475_, new_n1493_ );
and g1423 ( new_n1495_, new_n1494_, G56gat );
and g1424 ( new_n1496_, new_n1440_, new_n273_ );
or g1425 ( new_n1497_, new_n1495_, new_n1496_ );
and g1426 ( new_n1498_, new_n1497_, G53gat );
and g1427 ( new_n1499_, new_n1451_, G60gat );
or g1428 ( new_n1500_, new_n1473_, new_n1499_ );
and g1429 ( new_n1501_, new_n1500_, G50gat );
or g1430 ( new_n1502_, new_n1501_, new_n1493_ );
and g1431 ( new_n1503_, new_n1502_, G56gat );
and g1432 ( new_n1504_, new_n1451_, new_n273_ );
or g1433 ( new_n1505_, new_n1503_, new_n1504_ );
and g1434 ( new_n1506_, new_n1505_, new_n592_ );
or g1435 ( new_n1507_, new_n1498_, new_n1506_ );
and g1436 ( new_n1508_, new_n1507_, G47gat );
and g1437 ( new_n1509_, new_n1471_, new_n282_ );
and g1438 ( new_n1510_, new_n1509_, G50gat );
or g1439 ( new_n1511_, new_n1510_, new_n1493_ );
and g1440 ( new_n1512_, new_n1511_, G56gat );
and g1441 ( new_n1513_, new_n1466_, new_n896_ );
or g1442 ( new_n1514_, new_n1512_, new_n1513_ );
and g1443 ( new_n1515_, new_n1514_, G53gat );
and g1444 ( new_n1516_, new_n1470_, new_n185_ );
and g1445 ( new_n1517_, new_n1493_, G56gat );
or g1446 ( new_n1518_, new_n1516_, new_n1517_ );
and g1447 ( new_n1519_, new_n1518_, new_n592_ );
or g1448 ( new_n1520_, new_n1515_, new_n1519_ );
and g1449 ( new_n1521_, new_n1520_, new_n321_ );
or g1450 ( new_n1522_, new_n1508_, new_n1521_ );
and g1451 ( new_n1523_, new_n1522_, G37gat );
and g1452 ( new_n1524_, new_n1481_, new_n185_ );
or g1453 ( new_n1525_, new_n1517_, new_n1524_ );
and g1454 ( new_n1526_, new_n1525_, G53gat );
and g1455 ( new_n1527_, new_n1485_, new_n301_ );
and g1456 ( new_n1528_, new_n1490_, new_n300_ );
or g1457 ( new_n1529_, new_n1527_, new_n1528_ );
and g1458 ( new_n1530_, new_n1529_, new_n592_ );
or g1459 ( new_n1531_, new_n1526_, new_n1530_ );
and g1460 ( new_n1532_, new_n1531_, G47gat );
and g1461 ( new_n1533_, new_n321_, G53gat );
and g1462 ( new_n1534_, new_n630_, new_n1533_ );
and g1463 ( new_n1535_, new_n1534_, new_n1489_ );
or g1464 ( new_n1536_, new_n1532_, new_n1535_ );
and g1465 ( new_n1537_, new_n1536_, new_n187_ );
or g1466 ( new_n1538_, new_n1523_, new_n1537_ );
and g1467 ( new_n1539_, new_n1538_, G43gat );
and g1468 ( new_n1540_, new_n1497_, new_n291_ );
or g1469 ( new_n1541_, new_n1539_, new_n1540_ );
and g1470 ( new_n1542_, new_n1541_, G40gat );
and g1471 ( new_n1543_, new_n1405_, G73gat );
or g1472 ( new_n1544_, new_n1421_, new_n1543_ );
and g1473 ( new_n1545_, new_n1544_, G63gat );
or g1474 ( new_n1546_, new_n1545_, new_n1436_ );
and g1475 ( new_n1547_, new_n1546_, G69gat );
and g1476 ( new_n1548_, new_n1405_, new_n266_ );
or g1477 ( new_n1549_, new_n1547_, new_n1548_ );
and g1478 ( new_n1550_, new_n1549_, G60gat );
or g1479 ( new_n1551_, new_n1473_, new_n1550_ );
and g1480 ( new_n1552_, new_n1551_, G50gat );
or g1481 ( new_n1553_, new_n1552_, new_n1493_ );
and g1482 ( new_n1554_, new_n1553_, G56gat );
and g1483 ( new_n1555_, new_n1549_, new_n273_ );
or g1484 ( new_n1556_, new_n1554_, new_n1555_ );
and g1485 ( new_n1557_, new_n1556_, G47gat );
or g1486 ( new_n1558_, new_n1557_, new_n1521_ );
and g1487 ( new_n1559_, new_n1558_, G37gat );
or g1488 ( new_n1560_, new_n1559_, new_n1537_ );
and g1489 ( new_n1561_, new_n1560_, G43gat );
and g1490 ( new_n1562_, new_n1556_, new_n291_ );
or g1491 ( new_n1563_, new_n1561_, new_n1562_ );
and g1492 ( new_n1564_, new_n1563_, new_n642_ );
or g1493 ( new_n1565_, new_n1542_, new_n1564_ );
and g1494 ( new_n1566_, new_n1565_, G34gat );
and g1495 ( new_n1567_, new_n1415_, G73gat );
or g1496 ( new_n1568_, new_n1421_, new_n1567_ );
and g1497 ( new_n1569_, new_n1568_, G63gat );
or g1498 ( new_n1570_, new_n1569_, new_n1436_ );
and g1499 ( new_n1571_, new_n1570_, G69gat );
and g1500 ( new_n1572_, new_n1415_, new_n266_ );
or g1501 ( new_n1573_, new_n1571_, new_n1572_ );
and g1502 ( new_n1574_, new_n1573_, new_n894_ );
or g1503 ( new_n1575_, new_n1574_, new_n1509_ );
and g1504 ( new_n1576_, new_n1575_, G50gat );
or g1505 ( new_n1577_, new_n1576_, new_n1493_ );
and g1506 ( new_n1578_, new_n1577_, G56gat );
and g1507 ( new_n1579_, new_n1573_, new_n273_ );
or g1508 ( new_n1580_, new_n1578_, new_n1579_ );
or g1509 ( new_n1581_, new_n1580_, new_n679_ );
or g1510 ( new_n1582_, new_n1518_, new_n889_ );
and g1511 ( new_n1583_, new_n1582_, G37gat );
and g1512 ( new_n1584_, new_n1581_, new_n1583_ );
or g1513 ( new_n1585_, new_n1584_, new_n1537_ );
and g1514 ( new_n1586_, new_n1585_, G43gat );
and g1515 ( new_n1587_, new_n1580_, new_n291_ );
or g1516 ( new_n1588_, new_n1586_, new_n1587_ );
and g1517 ( new_n1589_, new_n1588_, G40gat );
and g1518 ( new_n1590_, new_n1537_, G43gat );
and g1519 ( new_n1591_, new_n1418_, new_n181_ );
or g1520 ( new_n1592_, new_n1468_, new_n1591_ );
and g1521 ( new_n1593_, new_n1592_, new_n185_ );
or g1522 ( new_n1594_, new_n1593_, new_n1517_ );
and g1523 ( new_n1595_, new_n1594_, new_n189_ );
or g1524 ( new_n1596_, new_n1590_, new_n1595_ );
and g1525 ( new_n1597_, new_n1596_, new_n642_ );
or g1526 ( new_n1598_, new_n1589_, new_n1597_ );
and g1527 ( new_n1599_, new_n1598_, new_n317_ );
or g1528 ( new_n1600_, new_n1566_, new_n1599_ );
and g1529 ( new_n1601_, new_n1600_, G24gat );
and g1530 ( new_n1602_, new_n1486_, G60gat );
or g1531 ( new_n1603_, new_n1602_, new_n1491_ );
and g1532 ( new_n1604_, new_n1603_, new_n184_ );
or g1533 ( new_n1605_, new_n1425_, new_n859_ );
and g1534 ( new_n1606_, new_n1477_, new_n851_ );
and g1535 ( new_n1607_, new_n1605_, new_n1606_ );
or g1536 ( new_n1608_, new_n1604_, new_n1607_ );
and g1537 ( new_n1609_, new_n1608_, new_n861_ );
and g1538 ( new_n1610_, new_n1530_, G47gat );
or g1539 ( new_n1611_, new_n1610_, new_n1535_ );
and g1540 ( new_n1612_, new_n1611_, new_n188_ );
or g1541 ( new_n1613_, new_n1609_, new_n1612_ );
and g1542 ( new_n1614_, new_n1613_, G40gat );
and g1543 ( new_n1615_, new_n1428_, new_n284_ );
or g1544 ( new_n1616_, new_n1615_, new_n1484_ );
and g1545 ( new_n1617_, new_n1616_, new_n301_ );
or g1546 ( new_n1618_, new_n1617_, new_n1528_ );
and g1547 ( new_n1619_, new_n1618_, new_n323_ );
and g1548 ( new_n1620_, new_n1535_, new_n188_ );
or g1549 ( new_n1621_, new_n1619_, new_n1620_ );
and g1550 ( new_n1622_, new_n1621_, new_n642_ );
or g1551 ( new_n1623_, new_n1614_, new_n1622_ );
and g1552 ( new_n1624_, new_n1623_, G34gat );
or g1553 ( new_n1625_, new_n1432_, new_n581_ );
and g1554 ( new_n1626_, new_n1625_, new_n1287_ );
or g1555 ( new_n1627_, new_n1626_, new_n642_ );
and g1556 ( new_n1628_, new_n1627_, new_n317_ );
or g1557 ( new_n1629_, new_n1624_, new_n1628_ );
and g1558 ( new_n1630_, new_n1629_, new_n191_ );
or g1559 ( new_n1631_, new_n1601_, new_n1630_ );
and g1560 ( new_n1632_, new_n1631_, G30gat );
and g1561 ( new_n1633_, new_n1541_, new_n308_ );
or g1562 ( new_n1634_, new_n1632_, new_n1633_ );
and g1563 ( new_n1635_, new_n1634_, G14gat );
and g1564 ( new_n1636_, new_n1399_, new_n445_ );
or g1565 ( new_n1637_, new_n1379_, new_n1636_ );
and g1566 ( new_n1638_, new_n1637_, G76gat );
or g1567 ( new_n1639_, new_n1638_, new_n1393_ );
and g1568 ( new_n1640_, new_n1639_, G82gat );
and g1569 ( new_n1641_, new_n1640_, G79gat );
or g1570 ( new_n1642_, new_n1406_, new_n1641_ );
and g1571 ( new_n1643_, new_n1642_, G73gat );
or g1572 ( new_n1644_, new_n1643_, new_n1421_ );
and g1573 ( new_n1645_, new_n1644_, G63gat );
or g1574 ( new_n1646_, new_n1645_, new_n1436_ );
and g1575 ( new_n1647_, new_n1646_, G69gat );
and g1576 ( new_n1648_, new_n1640_, new_n266_ );
or g1577 ( new_n1649_, new_n1647_, new_n1648_ );
and g1578 ( new_n1650_, new_n1649_, G66gat );
or g1579 ( new_n1651_, new_n1650_, new_n1452_ );
and g1580 ( new_n1652_, new_n1651_, G60gat );
or g1581 ( new_n1653_, new_n1652_, new_n1473_ );
and g1582 ( new_n1654_, new_n1653_, G50gat );
or g1583 ( new_n1655_, new_n1654_, new_n1493_ );
and g1584 ( new_n1656_, new_n1655_, G56gat );
and g1585 ( new_n1657_, new_n1649_, new_n273_ );
or g1586 ( new_n1658_, new_n1656_, new_n1657_ );
and g1587 ( new_n1659_, new_n1658_, G53gat );
or g1588 ( new_n1660_, new_n1659_, new_n1506_ );
and g1589 ( new_n1661_, new_n1660_, G47gat );
or g1590 ( new_n1662_, new_n1661_, new_n1521_ );
and g1591 ( new_n1663_, new_n1662_, G37gat );
or g1592 ( new_n1664_, new_n1663_, new_n1537_ );
and g1593 ( new_n1665_, new_n1664_, G43gat );
and g1594 ( new_n1666_, new_n1658_, new_n291_ );
or g1595 ( new_n1667_, new_n1665_, new_n1666_ );
and g1596 ( new_n1668_, new_n1667_, G40gat );
or g1597 ( new_n1669_, new_n1668_, new_n1564_ );
and g1598 ( new_n1670_, new_n1669_, G34gat );
or g1599 ( new_n1671_, new_n1670_, new_n1599_ );
and g1600 ( new_n1672_, new_n1671_, G24gat );
or g1601 ( new_n1673_, new_n1672_, new_n1630_ );
and g1602 ( new_n1674_, new_n1673_, G30gat );
and g1603 ( new_n1675_, new_n1667_, new_n308_ );
or g1604 ( new_n1676_, new_n1674_, new_n1675_ );
and g1605 ( new_n1677_, new_n1676_, new_n704_ );
or g1606 ( new_n1678_, new_n1635_, new_n1677_ );
and g1607 ( new_n1679_, new_n1678_, G27gat );
and g1608 ( new_n1680_, new_n1598_, new_n318_ );
or g1609 ( new_n1681_, new_n1680_, new_n1630_ );
and g1610 ( new_n1682_, new_n1681_, G30gat );
and g1611 ( new_n1683_, new_n1563_, new_n310_ );
or g1612 ( new_n1684_, new_n1682_, new_n1683_ );
and g1613 ( new_n1685_, new_n1684_, new_n693_ );
or g1614 ( new_n1686_, new_n1679_, new_n1685_ );
and g1615 ( new_n1687_, new_n1686_, G21gat );
and g1616 ( new_n1688_, new_n1588_, G34gat );
or g1617 ( new_n1689_, new_n1599_, new_n1688_ );
and g1618 ( new_n1690_, new_n1689_, G24gat );
or g1619 ( new_n1691_, new_n1690_, new_n1630_ );
and g1620 ( new_n1692_, new_n1691_, G30gat );
and g1621 ( new_n1693_, new_n1588_, new_n308_ );
or g1622 ( new_n1694_, new_n1692_, new_n1693_ );
and g1623 ( new_n1695_, new_n1694_, G27gat );
and g1624 ( new_n1696_, new_n1596_, new_n193_ );
and g1625 ( new_n1697_, new_n1630_, G30gat );
or g1626 ( new_n1698_, new_n1696_, new_n1697_ );
and g1627 ( new_n1699_, new_n1698_, new_n693_ );
or g1628 ( new_n1700_, new_n1695_, new_n1699_ );
and g1629 ( new_n1701_, new_n1700_, new_n338_ );
or g1630 ( new_n1702_, new_n1687_, new_n1701_ );
and g1631 ( new_n1703_, new_n1702_, G8gat );
and g1632 ( new_n1704_, new_n1694_, G14gat );
and g1633 ( new_n1705_, new_n1597_, new_n318_ );
or g1634 ( new_n1706_, new_n1705_, new_n1630_ );
and g1635 ( new_n1707_, new_n1706_, G30gat );
and g1636 ( new_n1708_, new_n679_, G37gat );
and g1637 ( new_n1709_, new_n1518_, new_n1708_ );
or g1638 ( new_n1710_, new_n1537_, new_n1709_ );
and g1639 ( new_n1711_, new_n1710_, G43gat );
and g1640 ( new_n1712_, new_n1514_, new_n891_ );
or g1641 ( new_n1713_, new_n1711_, new_n1712_ );
and g1642 ( new_n1714_, new_n1713_, new_n908_ );
or g1643 ( new_n1715_, new_n1707_, new_n1714_ );
and g1644 ( new_n1716_, new_n1715_, new_n704_ );
or g1645 ( new_n1717_, new_n1704_, new_n1716_ );
and g1646 ( new_n1718_, new_n1717_, G27gat );
or g1647 ( new_n1719_, new_n1718_, new_n1699_ );
and g1648 ( new_n1720_, new_n1719_, new_n338_ );
and g1649 ( new_n1721_, new_n1521_, G37gat );
or g1650 ( new_n1722_, new_n1721_, new_n1537_ );
and g1651 ( new_n1723_, new_n1722_, G43gat );
and g1652 ( new_n1724_, new_n1505_, new_n293_ );
or g1653 ( new_n1725_, new_n1723_, new_n1724_ );
and g1654 ( new_n1726_, new_n1725_, new_n310_ );
or g1655 ( new_n1727_, new_n1682_, new_n1726_ );
and g1656 ( new_n1728_, new_n1727_, G14gat );
or g1657 ( new_n1729_, new_n1728_, new_n1716_ );
and g1658 ( new_n1730_, new_n1729_, G21gat );
or g1659 ( new_n1731_, new_n1720_, new_n1730_ );
and g1660 ( new_n1732_, new_n1731_, new_n354_ );
or g1661 ( new_n1733_, new_n1703_, new_n1732_ );
and g1662 ( new_n1734_, new_n1733_, G11gat );
and g1663 ( new_n1735_, new_n1613_, new_n193_ );
or g1664 ( new_n1736_, new_n1697_, new_n1735_ );
and g1665 ( new_n1737_, new_n1736_, G27gat );
or g1666 ( new_n1738_, new_n1621_, new_n344_ );
or g1667 ( new_n1739_, new_n1627_, new_n345_ );
and g1668 ( new_n1740_, new_n1739_, new_n693_ );
and g1669 ( new_n1741_, new_n1738_, new_n1740_ );
or g1670 ( new_n1742_, new_n1737_, new_n1741_ );
and g1671 ( new_n1743_, new_n1742_, G21gat );
or g1672 ( new_n1744_, new_n1626_, new_n1239_ );
and g1673 ( new_n1745_, new_n1744_, new_n338_ );
or g1674 ( new_n1746_, new_n1743_, new_n1745_ );
and g1675 ( new_n1747_, new_n1746_, new_n195_ );
or g1676 ( new_n1748_, new_n1734_, new_n1747_ );
and g1677 ( new_n1749_, new_n1748_, G17gat );
and g1678 ( new_n1750_, new_n1395_, new_n266_ );
or g1679 ( new_n1751_, new_n1438_, new_n1750_ );
and g1680 ( new_n1752_, new_n1751_, new_n273_ );
or g1681 ( new_n1753_, new_n1656_, new_n1752_ );
and g1682 ( new_n1754_, new_n1753_, new_n291_ );
or g1683 ( new_n1755_, new_n1665_, new_n1754_ );
and g1684 ( new_n1756_, new_n1755_, new_n308_ );
or g1685 ( new_n1757_, new_n1632_, new_n1756_ );
and g1686 ( new_n1758_, new_n1757_, G14gat );
or g1687 ( new_n1759_, new_n1758_, new_n1677_ );
and g1688 ( new_n1760_, new_n1759_, G8gat );
and g1689 ( new_n1761_, new_n1729_, new_n354_ );
or g1690 ( new_n1762_, new_n1760_, new_n1761_ );
and g1691 ( new_n1763_, new_n1762_, new_n332_ );
or g1692 ( new_n1764_, new_n1749_, new_n1763_ );
and g1693 ( new_n1765_, new_n1764_, G1gat );
and g1694 ( new_n1766_, new_n1525_, new_n861_ );
or g1695 ( new_n1767_, new_n1766_, new_n1612_ );
and g1696 ( new_n1768_, new_n1767_, G40gat );
or g1697 ( new_n1769_, new_n1768_, new_n1622_ );
and g1698 ( new_n1770_, new_n1769_, G34gat );
or g1699 ( new_n1771_, new_n1628_, new_n193_ );
or g1700 ( new_n1772_, new_n1770_, new_n1771_ );
or g1701 ( new_n1773_, new_n1767_, new_n192_ );
and g1702 ( new_n1774_, new_n1773_, new_n704_ );
and g1703 ( new_n1775_, new_n1772_, new_n1774_ );
and g1704 ( new_n1776_, new_n1736_, G14gat );
or g1705 ( new_n1777_, new_n1775_, new_n1776_ );
and g1706 ( new_n1778_, new_n1777_, G27gat );
or g1707 ( new_n1779_, new_n1778_, new_n1741_ );
and g1708 ( new_n1780_, new_n1779_, G21gat );
or g1709 ( new_n1781_, new_n1780_, new_n1745_ );
and g1710 ( new_n1782_, new_n1781_, G8gat );
and g1711 ( new_n1783_, new_n1529_, new_n323_ );
or g1712 ( new_n1784_, new_n1620_, new_n344_ );
or g1713 ( new_n1785_, new_n1783_, new_n1784_ );
and g1714 ( new_n1786_, new_n1739_, G14gat );
and g1715 ( new_n1787_, new_n1785_, new_n1786_ );
and g1716 ( new_n1788_, new_n1287_, new_n1489_ );
or g1717 ( new_n1789_, new_n1788_, new_n746_ );
and g1718 ( new_n1790_, new_n1789_, new_n704_ );
or g1719 ( new_n1791_, new_n1787_, new_n1790_ );
and g1720 ( new_n1792_, new_n1791_, G21gat );
and g1721 ( new_n1793_, new_n1744_, G14gat );
or g1722 ( new_n1794_, new_n1789_, new_n693_ );
and g1723 ( new_n1795_, new_n1794_, new_n704_ );
or g1724 ( new_n1796_, new_n1793_, new_n1795_ );
and g1725 ( new_n1797_, new_n1796_, new_n338_ );
or g1726 ( new_n1798_, new_n1792_, new_n1797_ );
and g1727 ( new_n1799_, new_n1798_, new_n354_ );
or g1728 ( new_n1800_, new_n1782_, new_n1799_ );
and g1729 ( new_n1801_, new_n1800_, new_n196_ );
and g1730 ( new_n1802_, new_n1518_, new_n189_ );
or g1731 ( new_n1803_, new_n1590_, new_n1802_ );
and g1732 ( new_n1804_, new_n1803_, new_n193_ );
or g1733 ( new_n1805_, new_n1804_, new_n1697_ );
and g1734 ( new_n1806_, new_n1805_, G14gat );
or g1735 ( new_n1807_, new_n1806_, new_n1775_ );
and g1736 ( new_n1808_, new_n1807_, G8gat );
and g1737 ( new_n1809_, new_n1791_, new_n354_ );
or g1738 ( new_n1810_, new_n1808_, new_n1809_ );
and g1739 ( new_n1811_, new_n1810_, new_n197_ );
or g1740 ( new_n1812_, new_n1801_, new_n1811_ );
and g1741 ( new_n1813_, new_n1812_, new_n358_ );
or g1742 ( new_n1814_, new_n1765_, new_n1813_ );
and g1743 ( new_n1815_, new_n1814_, G4gat );
and g1744 ( new_n1816_, new_n1634_, G27gat );
or g1745 ( new_n1817_, new_n1816_, new_n1685_ );
and g1746 ( new_n1818_, new_n1817_, G21gat );
or g1747 ( new_n1819_, new_n1818_, new_n1701_ );
and g1748 ( new_n1820_, new_n1819_, G11gat );
or g1749 ( new_n1821_, new_n1820_, new_n1747_ );
and g1750 ( new_n1822_, new_n1821_, G17gat );
and g1751 ( new_n1823_, new_n1757_, new_n332_ );
or g1752 ( new_n1824_, new_n1822_, new_n1823_ );
and g1753 ( new_n1825_, new_n1824_, new_n198_ );
or g1754 ( new_n1826_, new_n1815_, new_n1825_ );
and g1755 ( new_n1827_, new_n1826_, keyinput0_G431gat );
not g1756 ( new_n1828_, keyinput0_G431gat );
and g1757 ( new_n1829_, new_n75_, new_n1828_ );
or g1758 ( new_n1830_, new_n1827_, new_n1829_ );
and g1759 ( new_n1831_, new_n1830_, keyinput1_G431gat );
not g1760 ( new_n1832_, keyinput1_G431gat );
and g1761 ( new_n1833_, new_n425_, new_n1828_ );
and g1762 ( new_n1834_, new_n82_, keyinput0_G431gat );
or g1763 ( new_n1835_, new_n1833_, new_n1834_ );
and g1764 ( new_n1836_, new_n1835_, new_n1832_ );
or g1765 ( new_n1837_, new_n1831_, new_n1836_ );
and g1766 ( new_n1838_, new_n1837_, keyinput2_G431gat );
not g1767 ( new_n1839_, keyinput2_G431gat );
and g1768 ( new_n1840_, new_n118_, new_n1828_ );
and g1769 ( new_n1841_, new_n806_, keyinput0_G431gat );
or g1770 ( new_n1842_, new_n1840_, new_n1841_ );
and g1771 ( new_n1843_, new_n1842_, new_n1832_ );
and g1772 ( new_n1844_, new_n116_, new_n1828_ );
not g1773 ( new_n1845_, new_n1844_ );
not g1774 ( new_n1846_, new_n1834_ );
and g1775 ( new_n1847_, new_n1846_, keyinput1_G431gat );
and g1776 ( new_n1848_, new_n1845_, new_n1847_ );
or g1777 ( new_n1849_, new_n1843_, new_n1848_ );
and g1778 ( new_n1850_, new_n1849_, new_n1839_ );
or g1779 ( new_n1851_, new_n1838_, new_n1850_ );
and g1780 ( new_n1852_, new_n1851_, keyinput3_G431gat );
not g1781 ( new_n1853_, keyinput3_G431gat );
and g1782 ( new_n1854_, new_n822_, new_n1828_ );
and g1783 ( new_n1855_, new_n824_, keyinput0_G431gat );
or g1784 ( new_n1856_, new_n1854_, new_n1855_ );
and g1785 ( new_n1857_, new_n1856_, new_n1832_ );
and g1786 ( new_n1858_, new_n89_, new_n1828_ );
or g1787 ( new_n1859_, new_n1858_, new_n1834_ );
and g1788 ( new_n1860_, new_n1859_, keyinput1_G431gat );
or g1789 ( new_n1861_, new_n1857_, new_n1860_ );
and g1790 ( new_n1862_, new_n1861_, keyinput2_G431gat );
and g1791 ( new_n1863_, new_n79_, keyinput0_G431gat );
and g1792 ( new_n1864_, new_n100_, new_n1828_ );
or g1793 ( new_n1865_, new_n1863_, new_n1864_ );
and g1794 ( new_n1866_, new_n1865_, new_n1832_ );
and g1795 ( new_n1867_, new_n80_, new_n1828_ );
or g1796 ( new_n1868_, new_n108_, new_n1867_ );
and g1797 ( new_n1869_, new_n1868_, keyinput1_G431gat );
or g1798 ( new_n1870_, new_n1866_, new_n1869_ );
and g1799 ( new_n1871_, new_n1870_, new_n1839_ );
or g1800 ( new_n1872_, new_n1862_, new_n1871_ );
and g1801 ( new_n1873_, new_n1872_, new_n1853_ );
or g1802 ( G431gat, new_n1852_, new_n1873_ );
and g1803 ( new_n1875_, new_n86_, G89gat );
or g1804 ( new_n1876_, new_n112_, new_n1875_ );
and g1805 ( new_n1877_, new_n1876_, G95gat );
and g1806 ( new_n1878_, new_n1877_, new_n445_ );
and g1807 ( new_n1879_, G92gat, G95gat );
and g1808 ( new_n1880_, new_n113_, new_n1879_ );
or g1809 ( new_n1881_, new_n1878_, new_n1880_ );
and g1810 ( new_n1882_, new_n1881_, G86gat );
and g1811 ( new_n1883_, new_n420_, new_n394_ );
or g1812 ( new_n1884_, new_n112_, new_n1883_ );
and g1813 ( new_n1885_, new_n1884_, G95gat );
and g1814 ( new_n1886_, new_n1885_, G92gat );
and g1815 ( new_n1887_, new_n112_, G95gat );
and g1816 ( new_n1888_, new_n1887_, new_n445_ );
or g1817 ( new_n1889_, new_n1886_, new_n1888_ );
and g1818 ( new_n1890_, new_n1889_, new_n229_ );
or g1819 ( new_n1891_, new_n1882_, new_n1890_ );
and g1820 ( new_n1892_, new_n1891_, G76gat );
or g1821 ( new_n1893_, new_n110_, new_n101_ );
and g1822 ( new_n1894_, new_n1893_, new_n172_ );
and g1823 ( new_n1895_, new_n1894_, G92gat );
and g1824 ( new_n1896_, new_n110_, new_n172_ );
and g1825 ( new_n1897_, new_n1896_, new_n445_ );
or g1826 ( new_n1898_, new_n1895_, new_n1897_ );
and g1827 ( new_n1899_, new_n1898_, G86gat );
and g1828 ( new_n1900_, new_n482_, G92gat );
and g1829 ( new_n1901_, new_n1900_, new_n229_ );
or g1830 ( new_n1902_, new_n1899_, new_n1901_ );
and g1831 ( new_n1903_, new_n1902_, new_n175_ );
or g1832 ( new_n1904_, new_n1892_, new_n1903_ );
and g1833 ( new_n1905_, new_n1904_, G82gat );
and g1834 ( new_n1906_, new_n253_, G95gat );
and g1835 ( new_n1907_, new_n113_, new_n1906_ );
or g1836 ( new_n1908_, new_n1905_, new_n1907_ );
and g1837 ( new_n1909_, new_n1908_, G79gat );
or g1838 ( new_n1910_, new_n86_, new_n91_ );
and g1839 ( new_n1911_, new_n1910_, G89gat );
or g1840 ( new_n1912_, new_n1911_, new_n112_ );
and g1841 ( new_n1913_, new_n1912_, G95gat );
and g1842 ( new_n1914_, new_n90_, new_n162_ );
or g1843 ( new_n1915_, new_n1913_, new_n1914_ );
and g1844 ( new_n1916_, new_n1915_, G86gat );
or g1845 ( new_n1917_, new_n1890_, new_n1916_ );
and g1846 ( new_n1918_, new_n1917_, G76gat );
or g1847 ( new_n1919_, new_n1918_, new_n1903_ );
and g1848 ( new_n1920_, new_n1919_, G82gat );
and g1849 ( new_n1921_, new_n1915_, new_n253_ );
or g1850 ( new_n1922_, new_n1920_, new_n1921_ );
and g1851 ( new_n1923_, new_n1922_, new_n493_ );
or g1852 ( new_n1924_, new_n1909_, new_n1923_ );
and g1853 ( new_n1925_, new_n1924_, G73gat );
and g1854 ( new_n1926_, new_n78_, G99gat );
or g1855 ( new_n1927_, new_n86_, new_n1926_ );
and g1856 ( new_n1928_, new_n1927_, G89gat );
or g1857 ( new_n1929_, new_n1928_, new_n112_ );
and g1858 ( new_n1930_, new_n1929_, G95gat );
and g1859 ( new_n1931_, new_n78_, new_n162_ );
or g1860 ( new_n1932_, new_n1930_, new_n1931_ );
or g1861 ( new_n1933_, new_n1932_, new_n530_ );
or g1862 ( new_n1934_, new_n1887_, new_n899_ );
and g1863 ( new_n1935_, new_n1934_, G76gat );
and g1864 ( new_n1936_, new_n1933_, new_n1935_ );
or g1865 ( new_n1937_, new_n1936_, new_n1903_ );
and g1866 ( new_n1938_, new_n1937_, G82gat );
and g1867 ( new_n1939_, new_n1932_, new_n253_ );
or g1868 ( new_n1940_, new_n1938_, new_n1939_ );
and g1869 ( new_n1941_, new_n1940_, G79gat );
and g1870 ( new_n1942_, new_n1903_, G82gat );
and g1871 ( new_n1943_, new_n1887_, new_n177_ );
or g1872 ( new_n1944_, new_n1942_, new_n1943_ );
or g1873 ( new_n1945_, new_n1944_, new_n178_ );
and g1874 ( new_n1946_, new_n1945_, new_n493_ );
or g1875 ( new_n1947_, new_n1941_, new_n1946_ );
and g1876 ( new_n1948_, new_n1947_, new_n257_ );
or g1877 ( new_n1949_, new_n1925_, new_n1948_ );
and g1878 ( new_n1950_, new_n1949_, G63gat );
and g1879 ( new_n1951_, new_n97_, new_n173_ );
or g1880 ( new_n1952_, new_n1887_, new_n1951_ );
and g1881 ( new_n1953_, new_n1952_, new_n868_ );
and g1882 ( new_n1954_, new_n1897_, G86gat );
or g1883 ( new_n1955_, new_n1954_, new_n1901_ );
and g1884 ( new_n1956_, new_n1955_, new_n176_ );
or g1885 ( new_n1957_, new_n1953_, new_n1956_ );
and g1886 ( new_n1958_, new_n1957_, G79gat );
and g1887 ( new_n1959_, new_n230_, new_n374_ );
or g1888 ( new_n1960_, new_n1959_, new_n100_ );
and g1889 ( new_n1961_, new_n1960_, new_n259_ );
or g1890 ( new_n1962_, new_n1961_, new_n1900_ );
and g1891 ( new_n1963_, new_n1962_, new_n493_ );
or g1892 ( new_n1964_, new_n1958_, new_n1963_ );
and g1893 ( new_n1965_, new_n1964_, G73gat );
or g1894 ( new_n1966_, new_n108_, new_n482_ );
and g1895 ( new_n1967_, new_n1966_, new_n532_ );
or g1896 ( new_n1968_, new_n1967_, new_n493_ );
and g1897 ( new_n1969_, new_n1968_, new_n257_ );
or g1898 ( new_n1970_, new_n1965_, new_n1969_ );
and g1899 ( new_n1971_, new_n1970_, new_n179_ );
or g1900 ( new_n1972_, new_n1950_, new_n1971_ );
and g1901 ( new_n1973_, new_n1972_, G69gat );
and g1902 ( new_n1974_, new_n1908_, new_n266_ );
or g1903 ( new_n1975_, new_n1973_, new_n1974_ );
and g1904 ( new_n1976_, new_n1975_, G66gat );
and g1905 ( new_n1977_, new_n1908_, G73gat );
or g1906 ( new_n1978_, new_n1948_, new_n1977_ );
and g1907 ( new_n1979_, new_n1978_, G63gat );
or g1908 ( new_n1980_, new_n1979_, new_n1971_ );
and g1909 ( new_n1981_, new_n1980_, G69gat );
or g1910 ( new_n1982_, new_n1981_, new_n1974_ );
and g1911 ( new_n1983_, new_n1982_, new_n544_ );
or g1912 ( new_n1984_, new_n1976_, new_n1983_ );
and g1913 ( new_n1985_, new_n1984_, G60gat );
and g1914 ( new_n1986_, new_n1877_, G86gat );
or g1915 ( new_n1987_, new_n1890_, new_n1986_ );
and g1916 ( new_n1988_, new_n1987_, G76gat );
or g1917 ( new_n1989_, new_n1988_, new_n1903_ );
and g1918 ( new_n1990_, new_n1989_, G82gat );
and g1919 ( new_n1991_, new_n1877_, new_n253_ );
or g1920 ( new_n1992_, new_n1990_, new_n1991_ );
and g1921 ( new_n1993_, new_n1992_, new_n904_ );
and g1922 ( new_n1994_, new_n1945_, new_n580_ );
and g1923 ( new_n1995_, G63gat, G69gat );
and g1924 ( new_n1996_, new_n1994_, new_n1995_ );
or g1925 ( new_n1997_, new_n1993_, new_n1996_ );
and g1926 ( new_n1998_, new_n1997_, G66gat );
and g1927 ( new_n1999_, new_n1971_, G69gat );
and g1928 ( new_n2000_, new_n1888_, new_n1456_ );
or g1929 ( new_n2001_, new_n1903_, new_n2000_ );
and g1930 ( new_n2002_, new_n2001_, G82gat );
and g1931 ( new_n2003_, new_n1885_, new_n901_ );
or g1932 ( new_n2004_, new_n2002_, new_n2003_ );
and g1933 ( new_n2005_, new_n2004_, new_n181_ );
and g1934 ( new_n2006_, new_n2005_, new_n544_ );
or g1935 ( new_n2007_, new_n1999_, new_n2006_ );
or g1936 ( new_n2008_, new_n1998_, new_n2007_ );
and g1937 ( new_n2009_, new_n2008_, new_n282_ );
or g1938 ( new_n2010_, new_n1985_, new_n2009_ );
and g1939 ( new_n2011_, new_n2010_, G50gat );
and g1940 ( new_n2012_, new_n1944_, new_n858_ );
or g1941 ( new_n2013_, new_n1963_, new_n1969_ );
and g1942 ( new_n2014_, new_n2013_, new_n180_ );
or g1943 ( new_n2015_, new_n2012_, new_n2014_ );
and g1944 ( new_n2016_, new_n2015_, G66gat );
and g1945 ( new_n2017_, new_n1894_, new_n868_ );
or g1946 ( new_n2018_, new_n1956_, new_n2017_ );
or g1947 ( new_n2019_, new_n2018_, new_n283_ );
or g1948 ( new_n2020_, new_n1968_, new_n284_ );
and g1949 ( new_n2021_, new_n2020_, new_n544_ );
and g1950 ( new_n2022_, new_n2019_, new_n2021_ );
or g1951 ( new_n2023_, new_n2016_, new_n2022_ );
and g1952 ( new_n2024_, new_n2023_, G60gat );
and g1953 ( new_n2025_, new_n1896_, new_n259_ );
and g1954 ( new_n2026_, new_n1900_, new_n258_ );
or g1955 ( new_n2027_, new_n2025_, new_n2026_ );
or g1956 ( new_n2028_, new_n2027_, new_n581_ );
and g1957 ( new_n2029_, new_n2028_, G66gat );
and g1958 ( new_n2030_, new_n532_, new_n482_ );
and g1959 ( new_n2031_, new_n2030_, new_n544_ );
or g1960 ( new_n2032_, new_n2029_, new_n2031_ );
and g1961 ( new_n2033_, new_n2032_, new_n282_ );
or g1962 ( new_n2034_, new_n2024_, new_n2033_ );
and g1963 ( new_n2035_, new_n2034_, new_n183_ );
or g1964 ( new_n2036_, new_n2011_, new_n2035_ );
and g1965 ( new_n2037_, new_n2036_, G56gat );
and g1966 ( new_n2038_, new_n1975_, new_n273_ );
or g1967 ( new_n2039_, new_n2037_, new_n2038_ );
and g1968 ( new_n2040_, new_n2039_, G53gat );
not g1969 ( new_n2041_, new_n1182_ );
or g1970 ( new_n2042_, new_n2008_, new_n2041_ );
or g1971 ( new_n2043_, new_n2034_, G50gat );
and g1972 ( new_n2044_, new_n2042_, new_n2043_ );
or g1973 ( new_n2045_, new_n2044_, new_n273_ );
and g1974 ( new_n2046_, new_n1922_, G73gat );
or g1975 ( new_n2047_, new_n1948_, new_n2046_ );
and g1976 ( new_n2048_, new_n2047_, G63gat );
or g1977 ( new_n2049_, new_n1971_, new_n266_ );
or g1978 ( new_n2050_, new_n2048_, new_n2049_ );
or g1979 ( new_n2051_, new_n1922_, G69gat );
and g1980 ( new_n2052_, new_n2050_, new_n2051_ );
or g1981 ( new_n2053_, new_n2052_, new_n276_ );
and g1982 ( new_n2054_, new_n2045_, new_n2053_ );
and g1983 ( new_n2055_, new_n2054_, new_n592_ );
or g1984 ( new_n2056_, new_n2040_, new_n2055_ );
and g1985 ( new_n2057_, new_n2056_, G47gat );
and g1986 ( new_n2058_, new_n1940_, G73gat );
or g1987 ( new_n2059_, new_n1948_, new_n2058_ );
and g1988 ( new_n2060_, new_n2059_, G63gat );
or g1989 ( new_n2061_, new_n2060_, new_n1971_ );
and g1990 ( new_n2062_, new_n2061_, G69gat );
and g1991 ( new_n2063_, new_n1940_, new_n266_ );
or g1992 ( new_n2064_, new_n2062_, new_n2063_ );
or g1993 ( new_n2065_, new_n2064_, new_n893_ );
or g1994 ( new_n2066_, new_n2005_, new_n894_ );
or g1995 ( new_n2067_, new_n1999_, new_n2066_ );
and g1996 ( new_n2068_, new_n2067_, G50gat );
and g1997 ( new_n2069_, new_n2065_, new_n2068_ );
or g1998 ( new_n2070_, new_n2069_, new_n2035_ );
and g1999 ( new_n2071_, new_n2070_, G56gat );
and g2000 ( new_n2072_, new_n2064_, new_n273_ );
or g2001 ( new_n2073_, new_n2071_, new_n2072_ );
and g2002 ( new_n2074_, new_n2073_, G53gat );
and g2003 ( new_n2075_, new_n2035_, G56gat );
and g2004 ( new_n2076_, new_n1945_, new_n181_ );
or g2005 ( new_n2077_, new_n1999_, new_n2076_ );
and g2006 ( new_n2078_, new_n2077_, new_n185_ );
or g2007 ( new_n2079_, new_n2075_, new_n2078_ );
and g2008 ( new_n2080_, new_n2079_, new_n592_ );
or g2009 ( new_n2081_, new_n2074_, new_n2080_ );
and g2010 ( new_n2082_, new_n2081_, new_n321_ );
or g2011 ( new_n2083_, new_n2057_, new_n2082_ );
and g2012 ( new_n2084_, new_n2083_, G37gat );
and g2013 ( new_n2085_, new_n1957_, new_n181_ );
or g2014 ( new_n2086_, new_n1999_, new_n2085_ );
and g2015 ( new_n2087_, new_n2086_, G66gat );
or g2016 ( new_n2088_, new_n2087_, new_n2022_ );
and g2017 ( new_n2089_, new_n2088_, G60gat );
or g2018 ( new_n2090_, new_n2033_, new_n185_ );
or g2019 ( new_n2091_, new_n2089_, new_n2090_ );
or g2020 ( new_n2092_, new_n2086_, new_n184_ );
and g2021 ( new_n2093_, new_n2091_, new_n2092_ );
or g2022 ( new_n2094_, new_n2093_, new_n592_ );
and g2023 ( new_n2095_, new_n2033_, new_n184_ );
or g2024 ( new_n2096_, new_n1962_, new_n283_ );
and g2025 ( new_n2097_, new_n2020_, new_n301_ );
and g2026 ( new_n2098_, new_n2097_, new_n2096_ );
or g2027 ( new_n2099_, new_n2095_, new_n2098_ );
or g2028 ( new_n2100_, new_n2099_, G53gat );
and g2029 ( new_n2101_, new_n2094_, new_n2100_ );
or g2030 ( new_n2102_, new_n2101_, new_n321_ );
or g2031 ( new_n2103_, new_n1967_, new_n581_ );
or g2032 ( new_n2104_, new_n2030_, new_n630_ );
and g2033 ( new_n2105_, new_n2103_, new_n2104_ );
or g2034 ( new_n2106_, new_n2105_, new_n592_ );
or g2035 ( new_n2107_, new_n2106_, G47gat );
and g2036 ( new_n2108_, new_n2102_, new_n2107_ );
and g2037 ( new_n2109_, new_n2108_, new_n187_ );
or g2038 ( new_n2110_, new_n2084_, new_n2109_ );
and g2039 ( new_n2111_, new_n2110_, G43gat );
and g2040 ( new_n2112_, new_n2039_, new_n291_ );
or g2041 ( new_n2113_, new_n2111_, new_n2112_ );
and g2042 ( new_n2114_, new_n2113_, G40gat );
and g2043 ( new_n2115_, new_n1992_, G73gat );
or g2044 ( new_n2116_, new_n1948_, new_n2115_ );
and g2045 ( new_n2117_, new_n2116_, G63gat );
or g2046 ( new_n2118_, new_n2117_, new_n2049_ );
or g2047 ( new_n2119_, new_n1992_, G69gat );
and g2048 ( new_n2120_, new_n2118_, new_n2119_ );
or g2049 ( new_n2121_, new_n2120_, new_n276_ );
and g2050 ( new_n2122_, new_n2045_, new_n2121_ );
and g2051 ( new_n2123_, new_n2122_, G47gat );
or g2052 ( new_n2124_, new_n2082_, new_n2123_ );
and g2053 ( new_n2125_, new_n2124_, G37gat );
or g2054 ( new_n2126_, new_n2125_, new_n2109_ );
and g2055 ( new_n2127_, new_n2126_, G43gat );
and g2056 ( new_n2128_, new_n2122_, new_n291_ );
or g2057 ( new_n2129_, new_n2127_, new_n2128_ );
and g2058 ( new_n2130_, new_n2129_, new_n642_ );
or g2059 ( new_n2131_, new_n2114_, new_n2130_ );
and g2060 ( new_n2132_, new_n2131_, G34gat );
and g2061 ( new_n2133_, new_n2079_, G37gat );
or g2062 ( new_n2134_, new_n2133_, new_n891_ );
or g2063 ( new_n2135_, new_n2109_, new_n2134_ );
not g2064 ( new_n2136_, new_n891_ );
or g2065 ( new_n2137_, new_n2068_, new_n273_ );
or g2066 ( new_n2138_, new_n2035_, new_n2137_ );
not g2067 ( new_n2139_, new_n896_ );
and g2068 ( new_n2140_, new_n2004_, new_n902_ );
or g2069 ( new_n2141_, new_n1994_, new_n2140_ );
and g2070 ( new_n2142_, new_n2141_, G63gat );
or g2071 ( new_n2143_, new_n2142_, new_n2049_ );
or g2072 ( new_n2144_, new_n2004_, G69gat );
and g2073 ( new_n2145_, new_n2143_, new_n2144_ );
or g2074 ( new_n2146_, new_n2145_, new_n2139_ );
and g2075 ( new_n2147_, new_n2138_, new_n2146_ );
or g2076 ( new_n2148_, new_n2147_, new_n2136_ );
and g2077 ( new_n2149_, new_n2135_, new_n2148_ );
and g2078 ( new_n2150_, new_n2149_, G40gat );
or g2079 ( new_n2151_, new_n2108_, new_n189_ );
or g2080 ( new_n2152_, new_n2075_, new_n188_ );
and g2081 ( new_n2153_, new_n1944_, new_n181_ );
or g2082 ( new_n2154_, new_n1999_, new_n2153_ );
and g2083 ( new_n2155_, new_n2154_, new_n185_ );
or g2084 ( new_n2156_, new_n2152_, new_n2155_ );
and g2085 ( new_n2157_, new_n2151_, new_n2156_ );
and g2086 ( new_n2158_, new_n2157_, new_n642_ );
or g2087 ( new_n2159_, new_n2150_, new_n2158_ );
and g2088 ( new_n2160_, new_n2159_, new_n317_ );
or g2089 ( new_n2161_, new_n2132_, new_n2160_ );
and g2090 ( new_n2162_, new_n2161_, G24gat );
and g2091 ( new_n2163_, new_n2018_, new_n858_ );
or g2092 ( new_n2164_, new_n2163_, new_n2014_ );
and g2093 ( new_n2165_, new_n2164_, G66gat );
or g2094 ( new_n2166_, new_n2165_, new_n2022_ );
and g2095 ( new_n2167_, new_n2166_, G60gat );
or g2096 ( new_n2168_, new_n2167_, new_n2033_ );
and g2097 ( new_n2169_, new_n2168_, new_n184_ );
and g2098 ( new_n2170_, new_n2164_, new_n185_ );
or g2099 ( new_n2171_, new_n2170_, new_n862_ );
or g2100 ( new_n2172_, new_n2169_, new_n2171_ );
or g2101 ( new_n2173_, new_n2100_, new_n321_ );
and g2102 ( new_n2174_, new_n2173_, new_n2107_ );
or g2103 ( new_n2175_, new_n2174_, new_n189_ );
and g2104 ( new_n2176_, new_n2172_, new_n2175_ );
and g2105 ( new_n2177_, new_n2176_, G40gat );
or g2106 ( new_n2178_, new_n2032_, new_n301_ );
or g2107 ( new_n2179_, new_n2027_, new_n283_ );
and g2108 ( new_n2180_, new_n2179_, new_n2020_ );
or g2109 ( new_n2181_, new_n2180_, new_n300_ );
and g2110 ( new_n2182_, new_n2181_, new_n323_ );
and g2111 ( new_n2183_, new_n2178_, new_n2182_ );
and g2112 ( new_n2184_, new_n2106_, new_n322_ );
or g2113 ( new_n2185_, new_n2183_, new_n2184_ );
and g2114 ( new_n2186_, new_n2185_, new_n642_ );
or g2115 ( new_n2187_, new_n2177_, new_n2186_ );
and g2116 ( new_n2188_, new_n2187_, G34gat );
and g2117 ( new_n2189_, new_n630_, new_n581_ );
or g2118 ( new_n2190_, new_n2030_, new_n680_ );
or g2119 ( new_n2191_, new_n2190_, new_n2189_ );
and g2120 ( new_n2192_, new_n2191_, G40gat );
and g2121 ( new_n2193_, new_n2192_, new_n317_ );
or g2122 ( new_n2194_, new_n2188_, new_n2193_ );
and g2123 ( new_n2195_, new_n2194_, new_n191_ );
or g2124 ( new_n2196_, new_n2162_, new_n2195_ );
and g2125 ( new_n2197_, new_n2196_, G30gat );
and g2126 ( new_n2198_, new_n2113_, new_n308_ );
or g2127 ( new_n2199_, new_n2197_, new_n2198_ );
and g2128 ( new_n2200_, new_n2199_, new_n704_ );
and g2129 ( new_n2201_, new_n119_, G95gat );
and g2130 ( new_n2202_, new_n115_, new_n162_ );
or g2131 ( new_n2203_, new_n2201_, new_n2202_ );
and g2132 ( new_n2204_, new_n2203_, G92gat );
or g2133 ( new_n2205_, new_n2204_, new_n1878_ );
and g2134 ( new_n2206_, new_n2205_, G86gat );
or g2135 ( new_n2207_, new_n2206_, new_n1890_ );
and g2136 ( new_n2208_, new_n2207_, G76gat );
or g2137 ( new_n2209_, new_n2208_, new_n1903_ );
and g2138 ( new_n2210_, new_n2209_, G82gat );
and g2139 ( new_n2211_, new_n2203_, new_n253_ );
or g2140 ( new_n2212_, new_n2210_, new_n2211_ );
and g2141 ( new_n2213_, new_n2212_, G79gat );
or g2142 ( new_n2214_, new_n2213_, new_n1923_ );
and g2143 ( new_n2215_, new_n2214_, G73gat );
or g2144 ( new_n2216_, new_n2215_, new_n1948_ );
and g2145 ( new_n2217_, new_n2216_, G63gat );
or g2146 ( new_n2218_, new_n2217_, new_n1971_ );
and g2147 ( new_n2219_, new_n2218_, G69gat );
and g2148 ( new_n2220_, new_n2212_, new_n266_ );
or g2149 ( new_n2221_, new_n2219_, new_n2220_ );
and g2150 ( new_n2222_, new_n2221_, G66gat );
or g2151 ( new_n2223_, new_n2222_, new_n1983_ );
and g2152 ( new_n2224_, new_n2223_, G60gat );
or g2153 ( new_n2225_, new_n2224_, new_n2009_ );
and g2154 ( new_n2226_, new_n2225_, G50gat );
or g2155 ( new_n2227_, new_n2226_, new_n2035_ );
and g2156 ( new_n2228_, new_n2227_, G56gat );
and g2157 ( new_n2229_, new_n2221_, new_n273_ );
or g2158 ( new_n2230_, new_n2228_, new_n2229_ );
and g2159 ( new_n2231_, new_n2230_, G53gat );
or g2160 ( new_n2232_, new_n2231_, new_n2055_ );
and g2161 ( new_n2233_, new_n2232_, G47gat );
or g2162 ( new_n2234_, new_n2233_, new_n2082_ );
and g2163 ( new_n2235_, new_n2234_, G37gat );
or g2164 ( new_n2236_, new_n2235_, new_n2109_ );
and g2165 ( new_n2237_, new_n2236_, G43gat );
and g2166 ( new_n2238_, new_n2230_, new_n291_ );
or g2167 ( new_n2239_, new_n2237_, new_n2238_ );
and g2168 ( new_n2240_, new_n2239_, new_n925_ );
and g2169 ( new_n2241_, new_n2130_, G34gat );
or g2170 ( new_n2242_, new_n2241_, new_n2160_ );
and g2171 ( new_n2243_, new_n2242_, G24gat );
or g2172 ( new_n2244_, new_n2243_, new_n2195_ );
and g2173 ( new_n2245_, new_n2244_, G30gat );
or g2174 ( new_n2246_, new_n2240_, new_n2245_ );
and g2175 ( new_n2247_, new_n2246_, G14gat );
or g2176 ( new_n2248_, new_n2200_, new_n2247_ );
and g2177 ( new_n2249_, new_n2248_, G27gat );
and g2178 ( new_n2250_, new_n2082_, G37gat );
or g2179 ( new_n2251_, new_n2250_, new_n2109_ );
and g2180 ( new_n2252_, new_n2251_, G43gat );
and g2181 ( new_n2253_, new_n2054_, new_n293_ );
or g2182 ( new_n2254_, new_n2253_, new_n311_ );
or g2183 ( new_n2255_, new_n2252_, new_n2254_ );
or g2184 ( new_n2256_, new_n2159_, new_n319_ );
or g2185 ( new_n2257_, new_n2194_, G24gat );
and g2186 ( new_n2258_, new_n2256_, new_n2257_ );
or g2187 ( new_n2259_, new_n2258_, new_n308_ );
and g2188 ( new_n2260_, new_n2259_, new_n693_ );
and g2189 ( new_n2261_, new_n2260_, new_n2255_ );
or g2190 ( new_n2262_, new_n2249_, new_n2261_ );
and g2191 ( new_n2263_, new_n2262_, G21gat );
or g2192 ( new_n2264_, new_n319_, G40gat );
or g2193 ( new_n2265_, new_n2157_, new_n2264_ );
and g2194 ( new_n2266_, new_n2265_, new_n2257_ );
or g2195 ( new_n2267_, new_n2266_, new_n308_ );
and g2196 ( new_n2268_, new_n2073_, new_n891_ );
and g2197 ( new_n2269_, new_n2133_, new_n679_ );
or g2198 ( new_n2270_, new_n2109_, new_n2269_ );
and g2199 ( new_n2271_, new_n2270_, G43gat );
or g2200 ( new_n2272_, new_n2271_, new_n907_ );
or g2201 ( new_n2273_, new_n2272_, new_n2268_ );
and g2202 ( new_n2274_, new_n2273_, G27gat );
and g2203 ( new_n2275_, new_n2274_, new_n2267_ );
or g2204 ( new_n2276_, new_n2152_, new_n2078_ );
and g2205 ( new_n2277_, new_n2151_, new_n2276_ );
or g2206 ( new_n2278_, new_n2277_, new_n192_ );
or g2207 ( new_n2279_, new_n2257_, new_n308_ );
and g2208 ( new_n2280_, new_n2279_, new_n693_ );
and g2209 ( new_n2281_, new_n2278_, new_n2280_ );
or g2210 ( new_n2282_, new_n2275_, new_n2281_ );
and g2211 ( new_n2283_, new_n2282_, new_n338_ );
or g2212 ( new_n2284_, new_n2263_, new_n2283_ );
and g2213 ( new_n2285_, new_n2284_, G8gat );
and g2214 ( new_n2286_, new_n2129_, new_n310_ );
and g2215 ( new_n2287_, new_n2159_, new_n318_ );
or g2216 ( new_n2288_, new_n2287_, new_n2195_ );
and g2217 ( new_n2289_, new_n2288_, G30gat );
or g2218 ( new_n2290_, new_n2286_, new_n2289_ );
and g2219 ( new_n2291_, new_n2290_, G14gat );
and g2220 ( new_n2292_, new_n2158_, new_n318_ );
or g2221 ( new_n2293_, new_n2292_, new_n2195_ );
and g2222 ( new_n2294_, new_n2293_, G30gat );
and g2223 ( new_n2295_, new_n2149_, new_n908_ );
or g2224 ( new_n2296_, new_n2294_, new_n2295_ );
and g2225 ( new_n2297_, new_n2296_, new_n704_ );
or g2226 ( new_n2298_, new_n2291_, new_n2297_ );
and g2227 ( new_n2299_, new_n2298_, G21gat );
and g2228 ( new_n2300_, new_n2296_, G27gat );
or g2229 ( new_n2301_, new_n2300_, new_n2281_ );
and g2230 ( new_n2302_, new_n2301_, new_n704_ );
and g2231 ( new_n2303_, new_n2282_, G14gat );
or g2232 ( new_n2304_, new_n2302_, new_n2303_ );
and g2233 ( new_n2305_, new_n2304_, new_n338_ );
or g2234 ( new_n2306_, new_n2299_, new_n2305_ );
and g2235 ( new_n2307_, new_n2306_, new_n354_ );
or g2236 ( new_n2308_, new_n2285_, new_n2307_ );
and g2237 ( new_n2309_, new_n2308_, G11gat );
or g2238 ( new_n2310_, new_n2093_, new_n862_ );
and g2239 ( new_n2311_, new_n2175_, new_n871_ );
and g2240 ( new_n2312_, new_n2310_, new_n2311_ );
and g2241 ( new_n2313_, new_n2186_, G34gat );
or g2242 ( new_n2314_, new_n2313_, new_n2193_ );
and g2243 ( new_n2315_, new_n2314_, new_n192_ );
or g2244 ( new_n2316_, new_n2312_, new_n2315_ );
and g2245 ( new_n2317_, new_n2316_, G27gat );
and g2246 ( new_n2318_, new_n2099_, new_n323_ );
or g2247 ( new_n2319_, new_n2318_, new_n2184_ );
and g2248 ( new_n2320_, new_n2319_, new_n345_ );
and g2249 ( new_n2321_, new_n2192_, new_n344_ );
or g2250 ( new_n2322_, new_n2320_, new_n2321_ );
and g2251 ( new_n2323_, new_n2322_, new_n693_ );
or g2252 ( new_n2324_, new_n2317_, new_n2323_ );
and g2253 ( new_n2325_, new_n2324_, G21gat );
or g2254 ( new_n2326_, new_n2105_, new_n680_ );
and g2255 ( new_n2327_, new_n2326_, new_n747_ );
or g2256 ( new_n2328_, new_n2327_, new_n693_ );
and g2257 ( new_n2329_, new_n2328_, new_n338_ );
or g2258 ( new_n2330_, new_n2325_, new_n2329_ );
and g2259 ( new_n2331_, new_n2330_, new_n195_ );
or g2260 ( new_n2332_, new_n2309_, new_n2331_ );
and g2261 ( new_n2333_, new_n2332_, G17gat );
and g2262 ( new_n2334_, new_n2046_, new_n493_ );
or g2263 ( new_n2335_, new_n2334_, new_n1948_ );
and g2264 ( new_n2336_, new_n2335_, G63gat );
or g2265 ( new_n2337_, new_n2336_, new_n1971_ );
and g2266 ( new_n2338_, new_n2337_, G69gat );
and g2267 ( new_n2339_, new_n2201_, new_n253_ );
or g2268 ( new_n2340_, new_n1905_, new_n2339_ );
and g2269 ( new_n2341_, new_n2340_, new_n919_ );
or g2270 ( new_n2342_, new_n2338_, new_n2341_ );
and g2271 ( new_n2343_, new_n2342_, G66gat );
or g2272 ( new_n2344_, new_n2343_, new_n1983_ );
and g2273 ( new_n2345_, new_n2344_, G60gat );
or g2274 ( new_n2346_, new_n2345_, new_n2009_ );
and g2275 ( new_n2347_, new_n2346_, G50gat );
or g2276 ( new_n2348_, new_n2347_, new_n2035_ );
and g2277 ( new_n2349_, new_n2348_, G56gat );
and g2278 ( new_n2350_, new_n2340_, new_n266_ );
or g2279 ( new_n2351_, new_n2219_, new_n2350_ );
and g2280 ( new_n2352_, new_n2351_, new_n273_ );
or g2281 ( new_n2353_, new_n2349_, new_n2352_ );
and g2282 ( new_n2354_, new_n2353_, new_n291_ );
or g2283 ( new_n2355_, new_n2237_, new_n2354_ );
and g2284 ( new_n2356_, new_n2355_, new_n308_ );
or g2285 ( new_n2357_, new_n2197_, new_n2356_ );
and g2286 ( new_n2358_, new_n2357_, G14gat );
or g2287 ( new_n2359_, new_n2200_, new_n2358_ );
and g2288 ( new_n2360_, new_n2359_, G8gat );
and g2289 ( new_n2361_, new_n2298_, new_n354_ );
or g2290 ( new_n2362_, new_n2360_, new_n2361_ );
and g2291 ( new_n2363_, new_n2362_, new_n332_ );
or g2292 ( new_n2364_, new_n2333_, new_n2363_ );
and g2293 ( new_n2365_, new_n2364_, G1gat );
or g2294 ( new_n2366_, new_n2157_, new_n192_ );
and g2295 ( new_n2367_, new_n2366_, new_n2279_ );
or g2296 ( new_n2368_, new_n2367_, new_n704_ );
and g2297 ( new_n2369_, new_n2176_, new_n871_ );
or g2298 ( new_n2370_, new_n2369_, new_n2315_ );
or g2299 ( new_n2371_, new_n2370_, G14gat );
and g2300 ( new_n2372_, new_n2368_, new_n2371_ );
or g2301 ( new_n2373_, new_n2372_, new_n354_ );
and g2302 ( new_n2374_, new_n2185_, new_n345_ );
or g2303 ( new_n2375_, new_n2374_, new_n2321_ );
and g2304 ( new_n2376_, new_n2375_, G14gat );
and g2305 ( new_n2377_, new_n747_, new_n704_ );
and g2306 ( new_n2378_, new_n2191_, new_n2377_ );
or g2307 ( new_n2379_, new_n2376_, new_n2378_ );
or g2308 ( new_n2380_, new_n2379_, G8gat );
and g2309 ( new_n2381_, new_n2373_, new_n2380_ );
or g2310 ( new_n2382_, new_n2381_, new_n196_ );
and g2311 ( new_n2383_, new_n2324_, G14gat );
and g2312 ( new_n2384_, new_n2370_, G27gat );
or g2313 ( new_n2385_, new_n2384_, new_n2323_ );
and g2314 ( new_n2386_, new_n2385_, new_n704_ );
or g2315 ( new_n2387_, new_n2383_, new_n2386_ );
and g2316 ( new_n2388_, new_n2387_, G21gat );
or g2317 ( new_n2389_, new_n2329_, new_n354_ );
or g2318 ( new_n2390_, new_n2388_, new_n2389_ );
and g2319 ( new_n2391_, new_n2379_, G21gat );
and g2320 ( new_n2392_, new_n2327_, G14gat );
or g2321 ( new_n2393_, new_n2378_, new_n693_ );
or g2322 ( new_n2394_, new_n2392_, new_n2393_ );
and g2323 ( new_n2395_, new_n2394_, new_n338_ );
or g2324 ( new_n2396_, new_n2395_, G8gat );
or g2325 ( new_n2397_, new_n2391_, new_n2396_ );
and g2326 ( new_n2398_, new_n2390_, new_n2397_ );
or g2327 ( new_n2399_, new_n2398_, new_n197_ );
and g2328 ( new_n2400_, new_n2399_, new_n358_ );
and g2329 ( new_n2401_, new_n2382_, new_n2400_ );
or g2330 ( new_n2402_, new_n2365_, new_n2401_ );
and g2331 ( new_n2403_, new_n2402_, G4gat );
and g2332 ( new_n2404_, new_n2246_, G27gat );
or g2333 ( new_n2405_, new_n2404_, new_n2261_ );
and g2334 ( new_n2406_, new_n2405_, G21gat );
or g2335 ( new_n2407_, new_n2406_, new_n2283_ );
and g2336 ( new_n2408_, new_n2407_, G11gat );
or g2337 ( new_n2409_, new_n2408_, new_n2331_ );
and g2338 ( new_n2410_, new_n2409_, G17gat );
and g2339 ( new_n2411_, new_n2357_, new_n332_ );
or g2340 ( new_n2412_, new_n2410_, new_n2411_ );
and g2341 ( new_n2413_, new_n2412_, new_n198_ );
or g2342 ( new_n2414_, new_n2403_, new_n2413_ );
and g2343 ( new_n2415_, new_n2414_, keyinput2_G432gat );
not g2344 ( new_n2416_, keyinput2_G432gat );
and g2345 ( new_n2417_, new_n115_, new_n2416_ );
or g2346 ( new_n2418_, new_n2415_, new_n2417_ );
and g2347 ( new_n2419_, new_n2418_, keyinput3_G432gat );
not g2348 ( new_n2420_, keyinput3_G432gat );
not g2349 ( new_n2421_, new_n190_ );
and g2350 ( new_n2422_, new_n2421_, new_n2416_ );
and g2351 ( new_n2423_, new_n220_, keyinput2_G432gat );
or g2352 ( new_n2424_, new_n2422_, new_n2423_ );
and g2353 ( new_n2425_, new_n2424_, new_n2420_ );
or g2354 ( new_n2426_, new_n2419_, new_n2425_ );
and g2355 ( new_n2427_, new_n2426_, keyinput1_G432gat );
not g2356 ( new_n2428_, keyinput1_G432gat );
and g2357 ( new_n2429_, new_n143_, new_n2416_ );
and g2358 ( new_n2430_, new_n82_, keyinput2_G432gat );
or g2359 ( new_n2431_, new_n2429_, new_n2430_ );
and g2360 ( new_n2432_, new_n2431_, keyinput3_G432gat );
and g2361 ( new_n2433_, new_n857_, new_n2416_ );
and g2362 ( new_n2434_, new_n917_, new_n2433_ );
and g2363 ( new_n2435_, new_n867_, keyinput2_G432gat );
or g2364 ( new_n2436_, new_n2434_, new_n2435_ );
and g2365 ( new_n2437_, new_n220_, new_n2420_ );
and g2366 ( new_n2438_, new_n2436_, new_n2437_ );
or g2367 ( new_n2439_, new_n2432_, new_n2438_ );
and g2368 ( new_n2440_, new_n2439_, new_n2428_ );
or g2369 ( new_n2441_, new_n2427_, new_n2440_ );
and g2370 ( new_n2442_, new_n2441_, keyinput0_G432gat );
not g2371 ( new_n2443_, keyinput0_G432gat );
and g2372 ( new_n2444_, new_n194_, G11gat );
not g2373 ( new_n2445_, new_n2444_ );
and g2374 ( new_n2446_, new_n2445_, new_n2416_ );
and g2375 ( new_n2447_, new_n186_, G37gat );
not g2376 ( new_n2448_, new_n2447_ );
and g2377 ( new_n2449_, new_n2448_, keyinput2_G432gat );
or g2378 ( new_n2450_, new_n2446_, new_n2449_ );
and g2379 ( new_n2451_, new_n2450_, new_n2420_ );
or g2380 ( new_n2452_, new_n179_, keyinput2_G432gat );
or g2381 ( new_n2453_, new_n806_, new_n2452_ );
and g2382 ( new_n2454_, new_n89_, keyinput2_G432gat );
not g2383 ( new_n2455_, new_n2454_ );
and g2384 ( new_n2456_, new_n2455_, keyinput3_G432gat );
and g2385 ( new_n2457_, new_n2453_, new_n2456_ );
or g2386 ( new_n2458_, new_n2451_, new_n2457_ );
and g2387 ( new_n2459_, new_n2458_, new_n2428_ );
and g2388 ( new_n2460_, new_n147_, new_n2416_ );
or g2389 ( new_n2461_, new_n2460_, new_n2454_ );
and g2390 ( new_n2462_, new_n2461_, new_n2420_ );
and g2391 ( new_n2463_, new_n116_, new_n2416_ );
and g2392 ( new_n2464_, G108gat, keyinput2_G432gat );
or g2393 ( new_n2465_, new_n2463_, new_n2464_ );
and g2394 ( new_n2466_, new_n2465_, keyinput3_G432gat );
or g2395 ( new_n2467_, new_n2462_, new_n2466_ );
and g2396 ( new_n2468_, new_n2467_, keyinput1_G432gat );
or g2397 ( new_n2469_, new_n2459_, new_n2468_ );
and g2398 ( new_n2470_, new_n2469_, new_n2443_ );
or g2399 ( G432gat, new_n2442_, new_n2470_ );
endmodule