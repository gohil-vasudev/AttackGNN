module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n698_, new_n425_, new_n226_, new_n697_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N42 );
nand g001 ( new_n152_, N29, N75 );
nor g002 ( new_n153_, new_n152_, new_n151_ );
xnor g003 ( N388, new_n153_, keyIn_0_3 );
not g004 ( new_n155_, N80 );
nand g005 ( new_n156_, N29, N36 );
nor g006 ( N389, new_n156_, new_n155_ );
nor g007 ( new_n158_, new_n156_, new_n151_ );
xor g008 ( N390, new_n158_, keyIn_0_4 );
nand g009 ( new_n160_, N85, N86 );
not g010 ( N391, new_n160_ );
not g011 ( new_n162_, N13 );
nand g012 ( new_n163_, N1, N8 );
nor g013 ( new_n164_, new_n163_, new_n162_ );
nand g014 ( new_n165_, new_n164_, N17 );
xnor g015 ( N418, new_n165_, keyIn_0_0 );
xnor g016 ( new_n167_, new_n158_, keyIn_0_1 );
not g017 ( new_n168_, new_n167_ );
nand g018 ( new_n169_, N1, N26 );
nand g019 ( new_n170_, N13, N17 );
nor g020 ( new_n171_, new_n169_, new_n170_ );
nand g021 ( N419, new_n168_, new_n171_ );
nand g022 ( new_n173_, N59, N75 );
not g023 ( new_n174_, new_n173_ );
nand g024 ( N420, new_n174_, N80 );
nand g025 ( new_n176_, N36, N59 );
not g026 ( new_n177_, new_n176_ );
nand g027 ( N421, new_n177_, N80 );
nor g028 ( new_n179_, new_n176_, new_n151_ );
xnor g029 ( N422, new_n179_, keyIn_0_5 );
not g030 ( new_n181_, N90 );
nor g031 ( new_n182_, N87, N88 );
nor g032 ( N423, new_n182_, new_n181_ );
nand g033 ( N446, new_n167_, new_n171_ );
not g034 ( new_n185_, keyIn_0_2 );
not g035 ( new_n186_, N51 );
nor g036 ( new_n187_, new_n169_, new_n186_ );
xnor g037 ( N447, new_n187_, new_n185_ );
nand g038 ( new_n189_, new_n164_, N55 );
nand g039 ( new_n190_, N29, N68 );
nor g040 ( N448, new_n189_, new_n190_ );
nand g041 ( new_n192_, N59, N68 );
not g042 ( new_n193_, new_n192_ );
nand g043 ( new_n194_, new_n193_, N74 );
nor g044 ( new_n195_, new_n189_, new_n194_ );
xnor g045 ( N449, new_n195_, keyIn_0_12 );
not g046 ( new_n197_, N89 );
nor g047 ( new_n198_, new_n182_, new_n197_ );
xnor g048 ( N450, new_n198_, keyIn_0_9 );
nor g049 ( new_n200_, N111, N116 );
xnor g050 ( new_n201_, new_n200_, keyIn_0_6 );
nand g051 ( new_n202_, N111, N116 );
nand g052 ( new_n203_, new_n201_, new_n202_ );
xor g053 ( new_n204_, N121, N126 );
xnor g054 ( new_n205_, new_n203_, new_n204_ );
nor g055 ( new_n206_, new_n205_, N135 );
not g056 ( new_n207_, new_n206_ );
nor g057 ( new_n208_, new_n207_, keyIn_0_19 );
nand g058 ( new_n209_, new_n207_, keyIn_0_19 );
nand g059 ( new_n210_, new_n205_, N135 );
nand g060 ( new_n211_, new_n209_, new_n210_ );
nor g061 ( new_n212_, new_n211_, new_n208_ );
xnor g062 ( new_n213_, N91, N96 );
xnor g063 ( new_n214_, N101, N106 );
xnor g064 ( new_n215_, new_n213_, new_n214_ );
xnor g065 ( new_n216_, new_n215_, N130 );
nand g066 ( new_n217_, new_n212_, new_n216_ );
nor g067 ( new_n218_, new_n217_, keyIn_0_32 );
nand g068 ( new_n219_, new_n217_, keyIn_0_32 );
not g069 ( new_n220_, new_n212_ );
not g070 ( new_n221_, new_n216_ );
nand g071 ( new_n222_, new_n220_, new_n221_ );
nand g072 ( new_n223_, new_n219_, new_n222_ );
nor g073 ( N767, new_n223_, new_n218_ );
not g074 ( new_n225_, keyIn_0_25 );
nor g075 ( new_n226_, N159, N165 );
not g076 ( new_n227_, keyIn_0_13 );
nand g077 ( new_n228_, N159, N165 );
nand g078 ( new_n229_, new_n228_, new_n227_ );
nor g079 ( new_n230_, new_n229_, new_n226_ );
xnor g080 ( new_n231_, N171, N177 );
xnor g081 ( new_n232_, new_n230_, new_n231_ );
nor g082 ( new_n233_, new_n232_, N130 );
nand g083 ( new_n234_, new_n233_, new_n225_ );
nor g084 ( new_n235_, new_n233_, new_n225_ );
nand g085 ( new_n236_, new_n232_, N130 );
nand g086 ( new_n237_, new_n236_, keyIn_0_31 );
nor g087 ( new_n238_, new_n235_, new_n237_ );
nand g088 ( new_n239_, new_n238_, new_n234_ );
xor g089 ( new_n240_, N183, N189 );
xnor g090 ( new_n241_, N195, N201 );
xnor g091 ( new_n242_, new_n240_, new_n241_ );
nor g092 ( new_n243_, new_n242_, N207 );
not g093 ( new_n244_, new_n243_ );
nor g094 ( new_n245_, new_n244_, keyIn_0_26 );
nand g095 ( new_n246_, new_n244_, keyIn_0_26 );
nand g096 ( new_n247_, new_n242_, N207 );
nand g097 ( new_n248_, new_n246_, new_n247_ );
nor g098 ( new_n249_, new_n248_, new_n245_ );
xnor g099 ( N768, new_n249_, new_n239_ );
not g100 ( new_n251_, keyIn_0_52 );
not g101 ( new_n252_, N261 );
not g102 ( new_n253_, N153 );
not g103 ( new_n254_, N1 );
nand g104 ( new_n255_, N447, N17 );
nand g105 ( new_n256_, N59, N156 );
not g106 ( new_n257_, new_n256_ );
nor g107 ( new_n258_, new_n255_, new_n257_ );
nor g108 ( new_n259_, new_n258_, new_n254_ );
nor g109 ( new_n260_, new_n259_, new_n253_ );
nor g110 ( new_n261_, new_n152_, new_n155_ );
nand g111 ( new_n262_, new_n261_, N55 );
not g112 ( new_n263_, new_n262_ );
nand g113 ( new_n264_, N447, new_n263_ );
nor g114 ( new_n265_, new_n264_, keyIn_0_15 );
nand g115 ( new_n266_, new_n264_, keyIn_0_15 );
xor g116 ( new_n267_, keyIn_0_10, N268 );
nand g117 ( new_n268_, new_n266_, new_n267_ );
nor g118 ( new_n269_, new_n268_, new_n265_ );
nor g119 ( new_n270_, new_n260_, new_n269_ );
nor g120 ( new_n271_, new_n173_, new_n151_ );
nand g121 ( new_n272_, N17, N51 );
nor g122 ( new_n273_, new_n163_, new_n272_ );
not g123 ( new_n274_, new_n273_ );
nor g124 ( new_n275_, new_n274_, new_n271_ );
not g125 ( new_n276_, new_n275_ );
nor g126 ( new_n277_, N17, N42 );
nand g127 ( new_n278_, N17, N42 );
nand g128 ( new_n279_, new_n257_, new_n278_ );
nor g129 ( new_n280_, new_n279_, new_n277_ );
nand g130 ( new_n281_, N447, new_n280_ );
nand g131 ( new_n282_, new_n281_, new_n276_ );
nand g132 ( new_n283_, new_n282_, N126 );
xnor g133 ( new_n284_, new_n283_, keyIn_0_24 );
nand g134 ( new_n285_, new_n270_, new_n284_ );
nand g135 ( new_n286_, new_n285_, N201 );
xor g136 ( new_n287_, new_n286_, keyIn_0_37 );
not g137 ( new_n288_, N201 );
not g138 ( new_n289_, N17 );
xnor g139 ( new_n290_, new_n187_, keyIn_0_2 );
nor g140 ( new_n291_, new_n290_, new_n289_ );
nand g141 ( new_n292_, new_n291_, new_n256_ );
nand g142 ( new_n293_, new_n292_, N1 );
nand g143 ( new_n294_, new_n293_, N153 );
not g144 ( new_n295_, new_n265_ );
not g145 ( new_n296_, new_n268_ );
nand g146 ( new_n297_, new_n296_, new_n295_ );
nand g147 ( new_n298_, new_n297_, new_n294_ );
not g148 ( new_n299_, keyIn_0_24 );
xnor g149 ( new_n300_, new_n283_, new_n299_ );
nor g150 ( new_n301_, new_n298_, new_n300_ );
nand g151 ( new_n302_, new_n301_, new_n288_ );
nand g152 ( new_n303_, new_n302_, keyIn_0_38 );
not g153 ( new_n304_, keyIn_0_38 );
nor g154 ( new_n305_, new_n285_, N201 );
nand g155 ( new_n306_, new_n305_, new_n304_ );
nand g156 ( new_n307_, new_n306_, new_n303_ );
nor g157 ( new_n308_, new_n287_, new_n307_ );
xnor g158 ( new_n309_, new_n308_, new_n252_ );
nor g159 ( new_n310_, new_n309_, new_n251_ );
nand g160 ( new_n311_, new_n309_, new_n251_ );
nand g161 ( new_n312_, new_n311_, N219 );
nor g162 ( new_n313_, new_n312_, new_n310_ );
nand g163 ( new_n314_, N121, N210 );
not g164 ( new_n315_, new_n314_ );
nor g165 ( new_n316_, new_n313_, new_n315_ );
nand g166 ( new_n317_, new_n316_, keyIn_0_56 );
nor g167 ( new_n318_, new_n316_, keyIn_0_56 );
not g168 ( new_n319_, N237 );
not g169 ( new_n320_, new_n287_ );
nor g170 ( new_n321_, new_n320_, new_n319_ );
not g171 ( new_n322_, new_n321_ );
nand g172 ( new_n323_, new_n322_, keyIn_0_50 );
not g173 ( new_n324_, N246 );
nor g174 ( new_n325_, new_n301_, new_n324_ );
nand g175 ( new_n326_, N255, N267 );
not g176 ( new_n327_, new_n326_ );
nor g177 ( new_n328_, new_n325_, new_n327_ );
nand g178 ( new_n329_, new_n323_, new_n328_ );
not g179 ( new_n330_, new_n329_ );
not g180 ( new_n331_, keyIn_0_28 );
nand g181 ( new_n332_, N42, N72 );
not g182 ( new_n333_, new_n332_ );
nand g183 ( new_n334_, new_n193_, new_n333_ );
nor g184 ( new_n335_, new_n189_, new_n334_ );
nand g185 ( new_n336_, new_n335_, keyIn_0_8 );
not g186 ( new_n337_, N73 );
nor g187 ( new_n338_, new_n335_, keyIn_0_8 );
nor g188 ( new_n339_, new_n338_, new_n337_ );
nand g189 ( new_n340_, new_n339_, new_n336_ );
xnor g190 ( new_n341_, new_n340_, keyIn_0_11 );
xnor g191 ( new_n342_, new_n341_, keyIn_0_14 );
xor g192 ( new_n343_, new_n342_, keyIn_0_16 );
nor g193 ( new_n344_, new_n343_, new_n288_ );
not g194 ( new_n345_, new_n344_ );
nand g195 ( new_n346_, new_n345_, new_n331_ );
nand g196 ( new_n347_, new_n308_, N228 );
nand g197 ( new_n348_, new_n346_, new_n347_ );
not g198 ( new_n349_, keyIn_0_50 );
nand g199 ( new_n350_, new_n321_, new_n349_ );
nand g200 ( new_n351_, new_n344_, keyIn_0_28 );
nand g201 ( new_n352_, new_n350_, new_n351_ );
nor g202 ( new_n353_, new_n348_, new_n352_ );
nand g203 ( new_n354_, new_n353_, new_n330_ );
nor g204 ( new_n355_, new_n318_, new_n354_ );
nand g205 ( N850, new_n355_, new_n317_ );
not g206 ( new_n357_, keyIn_0_53 );
not g207 ( new_n358_, keyIn_0_51 );
not g208 ( new_n359_, keyIn_0_30 );
not g209 ( new_n360_, N146 );
nor g210 ( new_n361_, new_n259_, new_n360_ );
nor g211 ( new_n362_, new_n361_, new_n269_ );
nand g212 ( new_n363_, new_n282_, N116 );
xnor g213 ( new_n364_, new_n363_, keyIn_0_23 );
nand g214 ( new_n365_, new_n362_, new_n364_ );
nand g215 ( new_n366_, new_n365_, new_n359_ );
nand g216 ( new_n367_, new_n293_, N146 );
nand g217 ( new_n368_, new_n297_, new_n367_ );
not g218 ( new_n369_, keyIn_0_23 );
xnor g219 ( new_n370_, new_n363_, new_n369_ );
nor g220 ( new_n371_, new_n368_, new_n370_ );
nand g221 ( new_n372_, new_n371_, keyIn_0_30 );
nand g222 ( new_n373_, new_n372_, new_n366_ );
nor g223 ( new_n374_, new_n373_, N189 );
not g224 ( new_n375_, N149 );
nor g225 ( new_n376_, new_n259_, new_n375_ );
not g226 ( new_n377_, new_n376_ );
nand g227 ( new_n378_, new_n282_, N121 );
not g228 ( new_n379_, new_n378_ );
nor g229 ( new_n380_, new_n269_, new_n379_ );
nand g230 ( new_n381_, new_n380_, new_n377_ );
nor g231 ( new_n382_, new_n381_, N195 );
nor g232 ( new_n383_, new_n374_, new_n382_ );
nand g233 ( new_n384_, new_n383_, new_n287_ );
xnor g234 ( new_n385_, new_n384_, new_n358_ );
nor g235 ( new_n386_, new_n307_, new_n252_ );
nand g236 ( new_n387_, new_n383_, new_n386_ );
nor g237 ( new_n388_, new_n387_, keyIn_0_42 );
nand g238 ( new_n389_, new_n387_, keyIn_0_42 );
nand g239 ( new_n390_, new_n381_, N195 );
nor g240 ( new_n391_, new_n374_, new_n390_ );
not g241 ( new_n392_, N189 );
not g242 ( new_n393_, new_n373_ );
nor g243 ( new_n394_, new_n393_, new_n392_ );
nor g244 ( new_n395_, new_n391_, new_n394_ );
nand g245 ( new_n396_, new_n389_, new_n395_ );
nor g246 ( new_n397_, new_n396_, new_n388_ );
nand g247 ( new_n398_, new_n397_, new_n385_ );
not g248 ( new_n399_, keyIn_0_36 );
not g249 ( new_n400_, keyIn_0_22 );
nand g250 ( new_n401_, new_n282_, N111 );
not g251 ( new_n402_, new_n401_ );
nand g252 ( new_n403_, new_n402_, new_n400_ );
nand g253 ( new_n404_, new_n297_, new_n403_ );
nand g254 ( new_n405_, new_n293_, N143 );
nand g255 ( new_n406_, new_n401_, keyIn_0_22 );
nand g256 ( new_n407_, new_n405_, new_n406_ );
nor g257 ( new_n408_, new_n404_, new_n407_ );
nand g258 ( new_n409_, new_n408_, keyIn_0_29 );
not g259 ( new_n410_, keyIn_0_29 );
nor g260 ( new_n411_, new_n401_, keyIn_0_22 );
nor g261 ( new_n412_, new_n269_, new_n411_ );
not g262 ( new_n413_, new_n407_ );
nand g263 ( new_n414_, new_n413_, new_n412_ );
nand g264 ( new_n415_, new_n414_, new_n410_ );
nand g265 ( new_n416_, new_n409_, new_n415_ );
nand g266 ( new_n417_, new_n416_, N183 );
xnor g267 ( new_n418_, new_n417_, new_n399_ );
nor g268 ( new_n419_, new_n416_, N183 );
not g269 ( new_n420_, new_n419_ );
nand g270 ( new_n421_, new_n418_, new_n420_ );
not g271 ( new_n422_, new_n421_ );
nand g272 ( new_n423_, new_n398_, new_n422_ );
nor g273 ( new_n424_, new_n423_, new_n357_ );
nand g274 ( new_n425_, new_n423_, new_n357_ );
not g275 ( new_n426_, new_n398_ );
nand g276 ( new_n427_, new_n426_, new_n421_ );
nand g277 ( new_n428_, new_n425_, new_n427_ );
nor g278 ( new_n429_, new_n428_, new_n424_ );
nand g279 ( new_n430_, new_n429_, keyIn_0_55 );
not g280 ( new_n431_, N219 );
nor g281 ( new_n432_, new_n429_, keyIn_0_55 );
nor g282 ( new_n433_, new_n432_, new_n431_ );
nand g283 ( new_n434_, new_n433_, new_n430_ );
not g284 ( new_n435_, keyIn_0_47 );
not g285 ( new_n436_, N228 );
nor g286 ( new_n437_, new_n421_, new_n436_ );
not g287 ( new_n438_, new_n437_ );
nand g288 ( new_n439_, new_n438_, new_n435_ );
not g289 ( new_n440_, keyIn_0_27 );
not g290 ( new_n441_, new_n343_ );
nand g291 ( new_n442_, new_n441_, N183 );
nor g292 ( new_n443_, new_n442_, new_n440_ );
nand g293 ( new_n444_, new_n442_, new_n440_ );
nand g294 ( new_n445_, new_n416_, N246 );
nand g295 ( new_n446_, N106, N210 );
nand g296 ( new_n447_, new_n445_, new_n446_ );
not g297 ( new_n448_, new_n447_ );
nand g298 ( new_n449_, new_n444_, new_n448_ );
nor g299 ( new_n450_, new_n449_, new_n443_ );
nand g300 ( new_n451_, new_n439_, new_n450_ );
nand g301 ( new_n452_, new_n437_, keyIn_0_47 );
not g302 ( new_n453_, keyIn_0_40 );
xnor g303 ( new_n454_, new_n418_, new_n453_ );
nand g304 ( new_n455_, new_n454_, N237 );
nand g305 ( new_n456_, new_n455_, new_n452_ );
nor g306 ( new_n457_, new_n451_, new_n456_ );
nand g307 ( N863, new_n434_, new_n457_ );
not g308 ( new_n459_, new_n382_ );
not g309 ( new_n460_, new_n386_ );
nand g310 ( new_n461_, new_n460_, new_n320_ );
nand g311 ( new_n462_, new_n461_, new_n459_ );
xnor g312 ( new_n463_, new_n390_, keyIn_0_49 );
nand g313 ( new_n464_, new_n462_, new_n463_ );
nor g314 ( new_n465_, new_n394_, new_n374_ );
nand g315 ( new_n466_, new_n464_, new_n465_ );
nor g316 ( new_n467_, new_n464_, new_n465_ );
nor g317 ( new_n468_, new_n467_, new_n431_ );
nand g318 ( new_n469_, new_n468_, new_n466_ );
not g319 ( new_n470_, keyIn_0_48 );
nand g320 ( new_n471_, new_n465_, N228 );
nand g321 ( new_n472_, new_n471_, new_n470_ );
nor g322 ( new_n473_, new_n343_, new_n392_ );
nand g323 ( new_n474_, new_n394_, N237 );
nand g324 ( new_n475_, N111, N210 );
nand g325 ( new_n476_, new_n474_, new_n475_ );
nor g326 ( new_n477_, new_n476_, new_n473_ );
nand g327 ( new_n478_, new_n477_, new_n472_ );
not g328 ( new_n479_, new_n471_ );
nand g329 ( new_n480_, new_n479_, keyIn_0_48 );
nand g330 ( new_n481_, new_n373_, N246 );
nand g331 ( new_n482_, N255, N259 );
nand g332 ( new_n483_, new_n481_, new_n482_ );
xnor g333 ( new_n484_, new_n483_, keyIn_0_41 );
nand g334 ( new_n485_, new_n480_, new_n484_ );
nor g335 ( new_n486_, new_n485_, new_n478_ );
nand g336 ( N864, new_n469_, new_n486_ );
not g337 ( new_n488_, new_n390_ );
nor g338 ( new_n489_, new_n488_, new_n382_ );
nand g339 ( new_n490_, new_n461_, new_n489_ );
nor g340 ( new_n491_, new_n461_, new_n489_ );
nor g341 ( new_n492_, new_n491_, new_n431_ );
nand g342 ( new_n493_, new_n492_, new_n490_ );
not g343 ( new_n494_, N195 );
nor g344 ( new_n495_, new_n343_, new_n494_ );
nand g345 ( new_n496_, new_n489_, N228 );
nor g346 ( new_n497_, new_n390_, new_n319_ );
nand g347 ( new_n498_, new_n381_, N246 );
nand g348 ( new_n499_, N116, N210 );
nand g349 ( new_n500_, N255, N260 );
nand g350 ( new_n501_, new_n499_, new_n500_ );
not g351 ( new_n502_, new_n501_ );
nand g352 ( new_n503_, new_n498_, new_n502_ );
nor g353 ( new_n504_, new_n497_, new_n503_ );
nand g354 ( new_n505_, new_n496_, new_n504_ );
nor g355 ( new_n506_, new_n495_, new_n505_ );
nand g356 ( N865, new_n493_, new_n506_ );
not g357 ( new_n508_, N177 );
not g358 ( new_n509_, keyIn_0_18 );
not g359 ( new_n510_, new_n261_ );
nor g360 ( new_n511_, new_n510_, N268 );
nand g361 ( new_n512_, new_n291_, new_n511_ );
not g362 ( new_n513_, new_n512_ );
nor g363 ( new_n514_, new_n513_, new_n509_ );
nand g364 ( new_n515_, new_n256_, N55 );
nor g365 ( new_n516_, new_n290_, new_n515_ );
not g366 ( new_n517_, new_n516_ );
nor g367 ( new_n518_, new_n517_, new_n253_ );
nand g368 ( new_n519_, N138, N152 );
not g369 ( new_n520_, new_n519_ );
nor g370 ( new_n521_, new_n518_, new_n520_ );
not g371 ( new_n522_, new_n521_ );
nor g372 ( new_n523_, new_n522_, new_n514_ );
nand g373 ( new_n524_, new_n282_, N106 );
not g374 ( new_n525_, new_n524_ );
nor g375 ( new_n526_, new_n512_, keyIn_0_18 );
nor g376 ( new_n527_, new_n525_, new_n526_ );
nand g377 ( new_n528_, new_n523_, new_n527_ );
not g378 ( new_n529_, new_n528_ );
nor g379 ( new_n530_, new_n529_, new_n508_ );
not g380 ( new_n531_, new_n530_ );
nand g381 ( new_n532_, new_n398_, new_n420_ );
not g382 ( new_n533_, keyIn_0_46 );
nand g383 ( new_n534_, new_n454_, new_n533_ );
xnor g384 ( new_n535_, new_n418_, keyIn_0_40 );
nand g385 ( new_n536_, new_n535_, keyIn_0_46 );
nand g386 ( new_n537_, new_n534_, new_n536_ );
nand g387 ( new_n538_, new_n532_, new_n537_ );
xnor g388 ( new_n539_, new_n538_, keyIn_0_54 );
nor g389 ( new_n540_, new_n528_, N177 );
not g390 ( new_n541_, new_n540_ );
nand g391 ( new_n542_, new_n539_, new_n541_ );
nand g392 ( new_n543_, new_n542_, new_n531_ );
not g393 ( new_n544_, keyIn_0_17 );
nor g394 ( new_n545_, new_n517_, new_n375_ );
nor g395 ( new_n546_, new_n545_, new_n544_ );
nand g396 ( new_n547_, N17, N138 );
nand g397 ( new_n548_, new_n512_, new_n547_ );
nor g398 ( new_n549_, new_n546_, new_n548_ );
not g399 ( new_n550_, new_n549_ );
nand g400 ( new_n551_, new_n545_, new_n544_ );
nand g401 ( new_n552_, new_n282_, N101 );
nand g402 ( new_n553_, new_n551_, new_n552_ );
nor g403 ( new_n554_, new_n550_, new_n553_ );
not g404 ( new_n555_, new_n554_ );
nor g405 ( new_n556_, new_n555_, N171 );
not g406 ( new_n557_, new_n556_ );
nand g407 ( new_n558_, new_n543_, new_n557_ );
nand g408 ( new_n559_, new_n555_, N171 );
xnor g409 ( new_n560_, new_n559_, keyIn_0_35 );
nand g410 ( new_n561_, new_n558_, new_n560_ );
not g411 ( new_n562_, N165 );
not g412 ( new_n563_, keyIn_0_21 );
nor g413 ( new_n564_, new_n517_, new_n360_ );
nor g414 ( new_n565_, new_n564_, new_n513_ );
not g415 ( new_n566_, new_n565_ );
nor g416 ( new_n567_, new_n566_, new_n563_ );
nor g417 ( new_n568_, new_n565_, keyIn_0_21 );
nand g418 ( new_n569_, new_n282_, N96 );
nand g419 ( new_n570_, N51, N138 );
nand g420 ( new_n571_, new_n569_, new_n570_ );
nor g421 ( new_n572_, new_n568_, new_n571_ );
not g422 ( new_n573_, new_n572_ );
nor g423 ( new_n574_, new_n573_, new_n567_ );
nand g424 ( new_n575_, new_n574_, new_n562_ );
nand g425 ( new_n576_, new_n561_, new_n575_ );
not g426 ( new_n577_, new_n574_ );
nand g427 ( new_n578_, new_n577_, N165 );
nand g428 ( new_n579_, new_n576_, new_n578_ );
not g429 ( new_n580_, keyIn_0_20 );
nand g430 ( new_n581_, new_n516_, N143 );
nand g431 ( new_n582_, new_n512_, new_n581_ );
not g432 ( new_n583_, new_n582_ );
nor g433 ( new_n584_, new_n583_, new_n580_ );
nor g434 ( new_n585_, new_n582_, keyIn_0_20 );
nand g435 ( new_n586_, new_n282_, N91 );
nand g436 ( new_n587_, N8, N138 );
nand g437 ( new_n588_, new_n586_, new_n587_ );
nor g438 ( new_n589_, new_n585_, new_n588_ );
not g439 ( new_n590_, new_n589_ );
nor g440 ( new_n591_, new_n590_, new_n584_ );
not g441 ( new_n592_, new_n591_ );
nor g442 ( new_n593_, new_n592_, N159 );
xnor g443 ( new_n594_, new_n593_, keyIn_0_33 );
not g444 ( new_n595_, new_n594_ );
nand g445 ( new_n596_, new_n579_, new_n595_ );
nand g446 ( new_n597_, new_n592_, N159 );
xnor g447 ( new_n598_, new_n597_, keyIn_0_43 );
nand g448 ( new_n599_, new_n596_, new_n598_ );
xnor g449 ( N866, new_n599_, keyIn_0_59 );
nor g450 ( new_n601_, new_n530_, new_n540_ );
nor g451 ( new_n602_, new_n539_, new_n601_ );
nand g452 ( new_n603_, new_n602_, keyIn_0_57 );
nor g453 ( new_n604_, new_n602_, keyIn_0_57 );
nand g454 ( new_n605_, new_n539_, new_n601_ );
nand g455 ( new_n606_, new_n605_, N219 );
nor g456 ( new_n607_, new_n604_, new_n606_ );
nand g457 ( new_n608_, new_n607_, new_n603_ );
nor g458 ( new_n609_, new_n343_, new_n508_ );
nand g459 ( new_n610_, new_n601_, N228 );
nor g460 ( new_n611_, new_n531_, new_n319_ );
nand g461 ( new_n612_, new_n528_, N246 );
nand g462 ( new_n613_, N101, N210 );
nand g463 ( new_n614_, new_n612_, new_n613_ );
nor g464 ( new_n615_, new_n611_, new_n614_ );
nand g465 ( new_n616_, new_n615_, new_n610_ );
nor g466 ( new_n617_, new_n616_, new_n609_ );
nand g467 ( new_n618_, new_n608_, new_n617_ );
xor g468 ( N874, new_n618_, keyIn_0_62 );
not g469 ( new_n620_, new_n597_ );
nor g470 ( new_n621_, new_n594_, new_n620_ );
nand g471 ( new_n622_, new_n579_, new_n621_ );
nor g472 ( new_n623_, new_n579_, new_n621_ );
nor g473 ( new_n624_, new_n623_, new_n431_ );
nand g474 ( new_n625_, new_n624_, new_n622_ );
nand g475 ( new_n626_, new_n441_, N159 );
nor g476 ( new_n627_, new_n591_, new_n324_ );
xnor g477 ( new_n628_, new_n627_, keyIn_0_34 );
nand g478 ( new_n629_, new_n626_, new_n628_ );
nor g479 ( new_n630_, new_n629_, keyIn_0_39 );
nand g480 ( new_n631_, new_n629_, keyIn_0_39 );
not g481 ( new_n632_, new_n621_ );
nor g482 ( new_n633_, new_n632_, new_n436_ );
nand g483 ( new_n634_, new_n620_, N237 );
not g484 ( new_n635_, new_n267_ );
nand g485 ( new_n636_, new_n635_, N210 );
nand g486 ( new_n637_, new_n634_, new_n636_ );
nor g487 ( new_n638_, new_n633_, new_n637_ );
nand g488 ( new_n639_, new_n638_, new_n631_ );
nor g489 ( new_n640_, new_n639_, new_n630_ );
nand g490 ( N878, new_n625_, new_n640_ );
not g491 ( new_n642_, keyIn_0_60 );
not g492 ( new_n643_, keyIn_0_54 );
xnor g493 ( new_n644_, new_n538_, new_n643_ );
nor g494 ( new_n645_, new_n644_, new_n540_ );
nand g495 ( new_n646_, new_n645_, new_n557_ );
not g496 ( new_n647_, new_n560_ );
nor g497 ( new_n648_, new_n647_, keyIn_0_44 );
nand g498 ( new_n649_, new_n647_, keyIn_0_44 );
nand g499 ( new_n650_, new_n557_, new_n530_ );
nand g500 ( new_n651_, new_n649_, new_n650_ );
nor g501 ( new_n652_, new_n651_, new_n648_ );
nand g502 ( new_n653_, new_n646_, new_n652_ );
nand g503 ( new_n654_, new_n578_, new_n575_ );
not g504 ( new_n655_, new_n654_ );
nor g505 ( new_n656_, new_n653_, new_n655_ );
nand g506 ( new_n657_, new_n656_, keyIn_0_58 );
nor g507 ( new_n658_, new_n656_, keyIn_0_58 );
nand g508 ( new_n659_, new_n653_, new_n655_ );
nand g509 ( new_n660_, new_n659_, N219 );
nor g510 ( new_n661_, new_n658_, new_n660_ );
nand g511 ( new_n662_, new_n661_, new_n657_ );
nand g512 ( new_n663_, N91, N210 );
xnor g513 ( new_n664_, new_n663_, keyIn_0_7 );
not g514 ( new_n665_, new_n664_ );
nand g515 ( new_n666_, new_n662_, new_n665_ );
not g516 ( new_n667_, new_n666_ );
nand g517 ( new_n668_, new_n667_, new_n642_ );
nand g518 ( new_n669_, new_n666_, keyIn_0_60 );
nor g519 ( new_n670_, new_n343_, new_n562_ );
nand g520 ( new_n671_, new_n655_, N228 );
nor g521 ( new_n672_, new_n578_, new_n319_ );
nor g522 ( new_n673_, new_n574_, new_n324_ );
nor g523 ( new_n674_, new_n672_, new_n673_ );
nand g524 ( new_n675_, new_n671_, new_n674_ );
nor g525 ( new_n676_, new_n675_, new_n670_ );
nand g526 ( new_n677_, new_n669_, new_n676_ );
not g527 ( new_n678_, new_n677_ );
nand g528 ( N879, new_n678_, new_n668_ );
not g529 ( new_n680_, keyIn_0_61 );
nor g530 ( new_n681_, new_n647_, new_n556_ );
nand g531 ( new_n682_, new_n543_, new_n681_ );
nor g532 ( new_n683_, new_n543_, new_n681_ );
nor g533 ( new_n684_, new_n683_, new_n431_ );
nand g534 ( new_n685_, new_n684_, new_n682_ );
nand g535 ( new_n686_, N96, N210 );
nand g536 ( new_n687_, new_n685_, new_n686_ );
xnor g537 ( new_n688_, new_n687_, new_n680_ );
nand g538 ( new_n689_, new_n681_, N228 );
nand g539 ( new_n690_, new_n555_, N246 );
nand g540 ( new_n691_, new_n689_, new_n690_ );
nor g541 ( new_n692_, new_n560_, new_n319_ );
nand g542 ( new_n693_, new_n692_, keyIn_0_45 );
nand g543 ( new_n694_, new_n441_, N171 );
not g544 ( new_n695_, keyIn_0_45 );
not g545 ( new_n696_, new_n692_ );
nand g546 ( new_n697_, new_n696_, new_n695_ );
nand g547 ( new_n698_, new_n697_, new_n694_ );
not g548 ( new_n699_, new_n698_ );
nand g549 ( new_n700_, new_n699_, new_n693_ );
nor g550 ( new_n701_, new_n700_, new_n691_ );
nand g551 ( new_n702_, new_n688_, new_n701_ );
xnor g552 ( N880, new_n702_, keyIn_0_63 );
endmodule