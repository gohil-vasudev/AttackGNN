module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n691_, new_n456_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n157_, new_n716_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n673_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n757_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

nand g000 ( new_n151_, N29, N42, N75 );
not g001 ( N388, new_n151_ );
nand g002 ( new_n153_, N29, N36, N80 );
not g003 ( N389, new_n153_ );
nand g004 ( new_n155_, N29, N36, N42 );
not g005 ( N390, new_n155_ );
nand g006 ( new_n157_, N85, N86 );
not g007 ( N391, new_n157_ );
nand g008 ( new_n159_, N1, N8 );
not g009 ( new_n160_, new_n159_ );
nand g010 ( new_n161_, new_n160_, N13, N17 );
not g011 ( N418, new_n161_ );
not g012 ( new_n163_, N13 );
not g013 ( new_n164_, N17 );
nand g014 ( new_n165_, N1, N26 );
nor g015 ( new_n166_, new_n165_, new_n163_, new_n164_ );
nand g016 ( N419, new_n166_, new_n155_ );
nand g017 ( N420, N59, N75, N80 );
nand g018 ( N421, N36, N59, N80 );
nand g019 ( N422, N36, N42, N59 );
not g020 ( new_n171_, N90 );
nor g021 ( new_n172_, N87, N88 );
nor g022 ( N423, new_n172_, new_n171_ );
nand g023 ( N446, new_n166_, N390 );
nand g024 ( new_n175_, N1, N26, N51 );
nand g025 ( new_n176_, new_n175_, keyIn_0_0 );
not g026 ( new_n177_, keyIn_0_0 );
nand g027 ( new_n178_, new_n177_, N1, N26, N51 );
nand g028 ( new_n179_, new_n176_, new_n178_ );
not g029 ( N447, new_n179_ );
nand g030 ( new_n181_, new_n160_, N13, N55 );
nand g031 ( new_n182_, N29, N68 );
nor g032 ( N448, new_n181_, new_n182_ );
not g033 ( new_n184_, N74 );
not g034 ( new_n185_, new_n181_ );
nand g035 ( new_n186_, new_n185_, N59, N68 );
nor g036 ( N449, new_n186_, new_n184_ );
not g037 ( new_n188_, N89 );
nor g038 ( N450, new_n172_, new_n188_ );
not g039 ( new_n190_, N130 );
not g040 ( new_n191_, N91 );
not g041 ( new_n192_, N96 );
nand g042 ( new_n193_, new_n191_, new_n192_ );
nand g043 ( new_n194_, N91, N96 );
nand g044 ( new_n195_, new_n193_, new_n194_ );
not g045 ( new_n196_, N101 );
not g046 ( new_n197_, N106 );
nand g047 ( new_n198_, new_n196_, new_n197_ );
nand g048 ( new_n199_, N101, N106 );
nand g049 ( new_n200_, new_n198_, new_n199_ );
nand g050 ( new_n201_, new_n195_, new_n200_ );
nand g051 ( new_n202_, new_n193_, new_n198_, new_n194_, new_n199_ );
nand g052 ( new_n203_, new_n201_, new_n202_ );
nand g053 ( new_n204_, new_n203_, new_n190_ );
nand g054 ( new_n205_, new_n201_, N130, new_n202_ );
nand g055 ( new_n206_, new_n204_, new_n205_ );
not g056 ( new_n207_, N111 );
not g057 ( new_n208_, N116 );
nand g058 ( new_n209_, new_n207_, new_n208_ );
nand g059 ( new_n210_, N111, N116 );
nand g060 ( new_n211_, new_n209_, new_n210_ );
not g061 ( new_n212_, N121 );
not g062 ( new_n213_, N126 );
nand g063 ( new_n214_, new_n212_, new_n213_ );
nand g064 ( new_n215_, N121, N126 );
nand g065 ( new_n216_, new_n214_, new_n215_ );
nand g066 ( new_n217_, new_n211_, new_n216_ );
nand g067 ( new_n218_, new_n209_, new_n214_, new_n210_, new_n215_ );
nand g068 ( new_n219_, new_n217_, new_n218_ );
nand g069 ( new_n220_, new_n219_, N135 );
not g070 ( new_n221_, N135 );
nand g071 ( new_n222_, new_n217_, new_n221_, new_n218_ );
nand g072 ( new_n223_, new_n220_, new_n222_ );
nand g073 ( new_n224_, new_n206_, new_n223_ );
nand g074 ( new_n225_, new_n204_, new_n220_, new_n205_, new_n222_ );
nand g075 ( N767, new_n224_, new_n225_ );
not g076 ( new_n227_, N159 );
not g077 ( new_n228_, N165 );
nand g078 ( new_n229_, new_n227_, new_n228_ );
nand g079 ( new_n230_, N159, N165 );
nand g080 ( new_n231_, new_n229_, new_n230_ );
not g081 ( new_n232_, N171 );
not g082 ( new_n233_, N177 );
nand g083 ( new_n234_, new_n232_, new_n233_ );
nand g084 ( new_n235_, N171, N177 );
nand g085 ( new_n236_, new_n234_, new_n235_ );
nand g086 ( new_n237_, new_n231_, new_n236_ );
nand g087 ( new_n238_, new_n229_, new_n234_, new_n230_, new_n235_ );
nand g088 ( new_n239_, new_n237_, new_n238_ );
nand g089 ( new_n240_, new_n239_, new_n190_ );
nand g090 ( new_n241_, new_n237_, N130, new_n238_ );
nand g091 ( new_n242_, new_n240_, new_n241_ );
not g092 ( new_n243_, N183 );
not g093 ( new_n244_, N189 );
nand g094 ( new_n245_, new_n243_, new_n244_ );
nand g095 ( new_n246_, N183, N189 );
nand g096 ( new_n247_, new_n245_, new_n246_ );
not g097 ( new_n248_, N195 );
not g098 ( new_n249_, N201 );
nand g099 ( new_n250_, new_n248_, new_n249_ );
nand g100 ( new_n251_, N195, N201 );
nand g101 ( new_n252_, new_n250_, new_n251_ );
nand g102 ( new_n253_, new_n247_, new_n252_ );
nand g103 ( new_n254_, new_n245_, new_n250_, new_n246_, new_n251_ );
nand g104 ( new_n255_, new_n253_, new_n254_ );
nand g105 ( new_n256_, new_n255_, N207 );
not g106 ( new_n257_, N207 );
nand g107 ( new_n258_, new_n253_, new_n257_, new_n254_ );
nand g108 ( new_n259_, new_n256_, new_n258_ );
nand g109 ( new_n260_, new_n242_, new_n259_ );
nand g110 ( new_n261_, new_n240_, new_n256_, new_n241_, new_n258_ );
nand g111 ( N768, new_n260_, new_n261_ );
not g112 ( new_n263_, keyIn_0_43 );
not g113 ( new_n264_, keyIn_0_21 );
not g114 ( new_n265_, keyIn_0_14 );
not g115 ( new_n266_, keyIn_0_8 );
nand g116 ( new_n267_, new_n179_, new_n266_ );
nand g117 ( new_n268_, new_n176_, keyIn_0_8, new_n178_ );
nand g118 ( new_n269_, new_n267_, new_n268_ );
nand g119 ( new_n270_, new_n269_, new_n265_ );
nand g120 ( new_n271_, new_n267_, keyIn_0_14, new_n268_ );
not g121 ( new_n272_, keyIn_0_13 );
not g122 ( new_n273_, keyIn_0_6 );
not g123 ( new_n274_, N42 );
nand g124 ( new_n275_, new_n164_, new_n274_ );
nand g125 ( new_n276_, new_n275_, new_n273_ );
nor g126 ( new_n277_, N17, N42 );
nand g127 ( new_n278_, new_n277_, keyIn_0_6 );
nand g128 ( new_n279_, new_n276_, new_n278_ );
nand g129 ( new_n280_, N17, N42 );
nand g130 ( new_n281_, new_n280_, keyIn_0_7 );
not g131 ( new_n282_, keyIn_0_7 );
nand g132 ( new_n283_, new_n282_, N17, N42 );
nand g133 ( new_n284_, new_n281_, new_n283_ );
nand g134 ( new_n285_, new_n279_, new_n284_ );
nand g135 ( new_n286_, new_n285_, new_n272_ );
not g136 ( new_n287_, new_n286_ );
nand g137 ( new_n288_, N59, N156 );
not g138 ( new_n289_, new_n288_ );
nand g139 ( new_n290_, new_n279_, keyIn_0_13, new_n284_ );
nand g140 ( new_n291_, new_n290_, new_n289_ );
nor g141 ( new_n292_, new_n287_, new_n291_ );
nand g142 ( new_n293_, new_n292_, keyIn_0_19, new_n270_, new_n271_ );
not g143 ( new_n294_, keyIn_0_1 );
nand g144 ( new_n295_, N1, N8, N17, N51 );
nand g145 ( new_n296_, new_n295_, new_n294_ );
nand g146 ( new_n297_, new_n160_, keyIn_0_1, N17, N51 );
nand g147 ( new_n298_, new_n297_, new_n296_ );
nand g148 ( new_n299_, new_n298_, keyIn_0_9 );
not g149 ( new_n300_, keyIn_0_9 );
nand g150 ( new_n301_, new_n297_, new_n300_, new_n296_ );
nand g151 ( new_n302_, new_n299_, new_n301_ );
not g152 ( new_n303_, keyIn_0_3 );
nand g153 ( new_n304_, N42, N59, N75 );
nand g154 ( new_n305_, new_n304_, new_n303_ );
nand g155 ( new_n306_, keyIn_0_3, N42, N59, N75 );
nand g156 ( new_n307_, new_n305_, new_n306_ );
nand g157 ( new_n308_, new_n307_, keyIn_0_11 );
not g158 ( new_n309_, keyIn_0_11 );
nand g159 ( new_n310_, new_n305_, new_n309_, new_n306_ );
nand g160 ( new_n311_, new_n308_, new_n310_ );
nand g161 ( new_n312_, new_n302_, new_n311_ );
nand g162 ( new_n313_, new_n312_, keyIn_0_15 );
not g163 ( new_n314_, keyIn_0_15 );
nand g164 ( new_n315_, new_n302_, new_n311_, new_n314_ );
nand g165 ( new_n316_, new_n313_, new_n315_ );
not g166 ( new_n317_, keyIn_0_19 );
not g167 ( new_n318_, new_n291_ );
nand g168 ( new_n319_, new_n318_, new_n270_, new_n271_, new_n286_ );
nand g169 ( new_n320_, new_n319_, new_n317_ );
nand g170 ( new_n321_, new_n320_, new_n316_, new_n293_ );
nand g171 ( new_n322_, new_n321_, new_n264_ );
nand g172 ( new_n323_, new_n320_, new_n316_, new_n293_, keyIn_0_21 );
nand g173 ( new_n324_, new_n322_, keyIn_0_31, N126, new_n323_ );
not g174 ( new_n325_, keyIn_0_20 );
not g175 ( new_n326_, keyIn_0_5 );
nand g176 ( new_n327_, new_n289_, new_n326_ );
nand g177 ( new_n328_, new_n288_, keyIn_0_5 );
nand g178 ( new_n329_, new_n327_, new_n328_ );
nand g179 ( new_n330_, new_n270_, N17, new_n271_, new_n329_ );
not g180 ( new_n331_, new_n330_ );
nand g181 ( new_n332_, new_n331_, new_n325_ );
nand g182 ( new_n333_, new_n330_, keyIn_0_20 );
nand g183 ( new_n334_, new_n332_, new_n333_ );
nand g184 ( new_n335_, new_n334_, keyIn_0_24, N1 );
not g185 ( new_n336_, keyIn_0_24 );
nand g186 ( new_n337_, new_n334_, N1 );
nand g187 ( new_n338_, new_n337_, new_n336_ );
nand g188 ( new_n339_, new_n338_, N153, new_n335_ );
not g189 ( new_n340_, keyIn_0_31 );
nand g190 ( new_n341_, new_n322_, N126, new_n323_ );
nand g191 ( new_n342_, new_n341_, new_n340_ );
nand g192 ( new_n343_, new_n342_, new_n339_, new_n324_ );
nand g193 ( new_n344_, new_n343_, keyIn_0_37 );
not g194 ( new_n345_, keyIn_0_37 );
nand g195 ( new_n346_, new_n342_, new_n339_, new_n345_, new_n324_ );
nand g196 ( new_n347_, new_n344_, new_n346_ );
not g197 ( new_n348_, keyIn_0_28 );
not g198 ( new_n349_, keyIn_0_18 );
nand g199 ( new_n350_, new_n270_, new_n271_ );
not g200 ( new_n351_, new_n350_ );
nand g201 ( new_n352_, N29, N75, N80 );
nand g202 ( new_n353_, new_n352_, keyIn_0_2 );
not g203 ( new_n354_, keyIn_0_2 );
nand g204 ( new_n355_, new_n354_, N29, N75, N80 );
nand g205 ( new_n356_, new_n353_, new_n355_ );
not g206 ( new_n357_, new_n356_ );
nand g207 ( new_n358_, new_n351_, N55, new_n357_ );
nor g208 ( new_n359_, new_n358_, new_n349_ );
nand g209 ( new_n360_, new_n358_, new_n349_ );
not g210 ( new_n361_, new_n360_ );
not g211 ( new_n362_, keyIn_0_12 );
not g212 ( new_n363_, N268 );
nor g213 ( new_n364_, new_n363_, keyIn_0_4 );
nand g214 ( new_n365_, new_n363_, keyIn_0_4 );
not g215 ( new_n366_, new_n365_ );
nor g216 ( new_n367_, new_n366_, new_n364_ );
not g217 ( new_n368_, new_n367_ );
nand g218 ( new_n369_, new_n368_, new_n362_ );
nand g219 ( new_n370_, new_n367_, keyIn_0_12 );
nand g220 ( new_n371_, new_n369_, new_n370_ );
nor g221 ( new_n372_, new_n361_, new_n359_, new_n371_ );
nand g222 ( new_n373_, new_n372_, new_n348_ );
not g223 ( new_n374_, new_n359_ );
nand g224 ( new_n375_, new_n374_, new_n360_, new_n369_, new_n370_ );
nand g225 ( new_n376_, new_n375_, keyIn_0_28 );
nand g226 ( new_n377_, new_n376_, new_n373_ );
nand g227 ( new_n378_, new_n347_, new_n377_ );
nand g228 ( new_n379_, new_n378_, new_n263_ );
nand g229 ( new_n380_, new_n347_, keyIn_0_43, new_n377_ );
nand g230 ( new_n381_, new_n379_, new_n380_ );
nand g231 ( new_n382_, new_n381_, N201 );
nand g232 ( new_n383_, new_n379_, new_n249_, new_n380_ );
nand g233 ( new_n384_, new_n382_, new_n383_ );
not g234 ( new_n385_, new_n384_ );
nand g235 ( new_n386_, new_n385_, N261 );
not g236 ( new_n387_, N261 );
nand g237 ( new_n388_, new_n384_, new_n387_ );
nand g238 ( new_n389_, new_n386_, N219, new_n388_ );
nand g239 ( new_n390_, new_n385_, N228 );
not g240 ( new_n391_, new_n390_ );
nand g241 ( new_n392_, new_n381_, N201, N237 );
nand g242 ( new_n393_, new_n381_, N246 );
not g243 ( new_n394_, N72 );
nor g244 ( new_n395_, new_n186_, new_n274_, new_n394_ );
nor g245 ( new_n396_, new_n395_, keyIn_0_10 );
nand g246 ( new_n397_, new_n395_, keyIn_0_10 );
nand g247 ( new_n398_, new_n397_, N73 );
nor g248 ( new_n399_, new_n398_, new_n396_ );
nand g249 ( new_n400_, new_n399_, N201 );
nand g250 ( new_n401_, N255, N267 );
nand g251 ( new_n402_, N121, N210 );
nand g252 ( new_n403_, new_n400_, new_n401_, new_n402_ );
not g253 ( new_n404_, new_n403_ );
nand g254 ( new_n405_, new_n392_, new_n393_, new_n404_ );
nor g255 ( new_n406_, new_n391_, new_n405_ );
nand g256 ( new_n407_, new_n406_, new_n389_ );
nand g257 ( new_n408_, new_n407_, keyIn_0_52 );
not g258 ( new_n409_, keyIn_0_52 );
nand g259 ( new_n410_, new_n406_, new_n409_, new_n389_ );
nand g260 ( N850, new_n408_, new_n410_ );
not g261 ( new_n412_, keyIn_0_57 );
not g262 ( new_n413_, keyIn_0_35 );
nand g263 ( new_n414_, new_n338_, N146, new_n335_ );
nand g264 ( new_n415_, new_n322_, N116, new_n323_ );
nand g265 ( new_n416_, new_n414_, new_n415_ );
nand g266 ( new_n417_, new_n416_, new_n413_ );
nand g267 ( new_n418_, new_n414_, keyIn_0_35, new_n415_ );
nand g268 ( new_n419_, new_n417_, new_n418_ );
nand g269 ( new_n420_, new_n372_, keyIn_0_26 );
not g270 ( new_n421_, keyIn_0_26 );
nand g271 ( new_n422_, new_n375_, new_n421_ );
nand g272 ( new_n423_, new_n422_, new_n420_ );
nand g273 ( new_n424_, new_n419_, new_n423_ );
nand g274 ( new_n425_, new_n424_, keyIn_0_41 );
not g275 ( new_n426_, keyIn_0_41 );
nand g276 ( new_n427_, new_n419_, new_n426_, new_n423_ );
nand g277 ( new_n428_, new_n425_, new_n244_, new_n427_ );
nand g278 ( new_n429_, new_n338_, N149, new_n335_ );
nand g279 ( new_n430_, new_n322_, N121, new_n323_ );
nand g280 ( new_n431_, new_n429_, keyIn_0_36, new_n430_ );
not g281 ( new_n432_, keyIn_0_36 );
nand g282 ( new_n433_, new_n429_, new_n430_ );
nand g283 ( new_n434_, new_n433_, new_n432_ );
nor g284 ( new_n435_, new_n372_, keyIn_0_27 );
not g285 ( new_n436_, keyIn_0_27 );
nor g286 ( new_n437_, new_n375_, new_n436_ );
nor g287 ( new_n438_, new_n437_, new_n435_ );
nand g288 ( new_n439_, new_n434_, new_n431_, new_n438_ );
nand g289 ( new_n440_, new_n439_, keyIn_0_42 );
not g290 ( new_n441_, keyIn_0_42 );
nand g291 ( new_n442_, new_n434_, new_n438_, new_n441_, new_n431_ );
nand g292 ( new_n443_, new_n440_, new_n248_, new_n442_ );
nand g293 ( new_n444_, new_n383_, N261, new_n428_, new_n443_ );
nand g294 ( new_n445_, new_n444_, keyIn_0_44 );
not g295 ( new_n446_, keyIn_0_44 );
nand g296 ( new_n447_, new_n428_, new_n443_ );
not g297 ( new_n448_, new_n447_ );
nand g298 ( new_n449_, new_n448_, new_n446_, N261, new_n383_ );
nand g299 ( new_n450_, new_n449_, new_n445_ );
nand g300 ( new_n451_, new_n440_, new_n442_ );
nand g301 ( new_n452_, new_n451_, N195 );
not g302 ( new_n453_, new_n452_ );
nand g303 ( new_n454_, new_n453_, new_n428_ );
nand g304 ( new_n455_, new_n454_, keyIn_0_45 );
not g305 ( new_n456_, keyIn_0_45 );
nand g306 ( new_n457_, new_n453_, new_n456_, new_n428_ );
nand g307 ( new_n458_, new_n455_, new_n457_ );
nand g308 ( new_n459_, new_n425_, new_n427_ );
nand g309 ( new_n460_, new_n459_, N189 );
not g310 ( new_n461_, keyIn_0_46 );
nor g311 ( new_n462_, new_n382_, new_n447_, new_n461_ );
nand g312 ( new_n463_, new_n381_, new_n428_, N201, new_n443_ );
nand g313 ( new_n464_, new_n463_, new_n461_ );
not g314 ( new_n465_, new_n464_ );
nor g315 ( new_n466_, new_n465_, new_n462_ );
nand g316 ( new_n467_, new_n466_, new_n450_, new_n458_, new_n460_ );
nand g317 ( new_n468_, new_n467_, keyIn_0_48 );
not g318 ( new_n469_, keyIn_0_48 );
nand g319 ( new_n470_, new_n458_, new_n460_ );
not g320 ( new_n471_, new_n470_ );
nand g321 ( new_n472_, new_n471_, new_n469_, new_n450_, new_n466_ );
nand g322 ( new_n473_, new_n468_, new_n472_ );
nand g323 ( new_n474_, new_n322_, new_n323_ );
not g324 ( new_n475_, new_n474_ );
nand g325 ( new_n476_, new_n475_, N111 );
nand g326 ( new_n477_, new_n338_, N143, new_n335_ );
nand g327 ( new_n478_, new_n476_, new_n477_ );
nand g328 ( new_n479_, new_n478_, keyIn_0_34 );
not g329 ( new_n480_, keyIn_0_34 );
nand g330 ( new_n481_, new_n476_, new_n480_, new_n477_ );
nand g331 ( new_n482_, new_n479_, new_n481_ );
nand g332 ( new_n483_, new_n372_, keyIn_0_25 );
not g333 ( new_n484_, keyIn_0_25 );
nand g334 ( new_n485_, new_n375_, new_n484_ );
nand g335 ( new_n486_, new_n485_, new_n483_ );
nand g336 ( new_n487_, new_n482_, new_n486_ );
nand g337 ( new_n488_, new_n487_, keyIn_0_40 );
not g338 ( new_n489_, keyIn_0_40 );
nand g339 ( new_n490_, new_n482_, new_n489_, new_n486_ );
nand g340 ( new_n491_, new_n488_, new_n490_ );
nand g341 ( new_n492_, new_n491_, N183 );
nand g342 ( new_n493_, new_n488_, new_n243_, new_n490_ );
nand g343 ( new_n494_, new_n492_, new_n493_ );
not g344 ( new_n495_, new_n494_ );
nand g345 ( new_n496_, new_n473_, new_n495_ );
nand g346 ( new_n497_, new_n468_, new_n472_, new_n494_ );
nand g347 ( new_n498_, new_n496_, N219, new_n497_ );
nand g348 ( new_n499_, new_n495_, N228 );
not g349 ( new_n500_, new_n499_ );
nand g350 ( new_n501_, new_n491_, N183, N237 );
nand g351 ( new_n502_, new_n491_, N246 );
nand g352 ( new_n503_, new_n399_, N183 );
nand g353 ( new_n504_, N106, N210 );
nand g354 ( new_n505_, new_n501_, new_n502_, new_n503_, new_n504_ );
nor g355 ( new_n506_, new_n500_, new_n505_ );
nand g356 ( new_n507_, new_n498_, new_n506_ );
nand g357 ( new_n508_, new_n507_, new_n412_ );
nand g358 ( new_n509_, new_n498_, keyIn_0_57, new_n506_ );
nand g359 ( N863, new_n508_, new_n509_ );
nand g360 ( new_n511_, new_n383_, N261 );
nand g361 ( new_n512_, new_n511_, new_n382_ );
nand g362 ( new_n513_, new_n512_, new_n443_ );
nand g363 ( new_n514_, new_n513_, new_n452_ );
nand g364 ( new_n515_, new_n514_, keyIn_0_49 );
not g365 ( new_n516_, keyIn_0_49 );
nand g366 ( new_n517_, new_n513_, new_n516_, new_n452_ );
nand g367 ( new_n518_, new_n515_, new_n517_ );
nand g368 ( new_n519_, new_n460_, new_n428_ );
not g369 ( new_n520_, new_n519_ );
nand g370 ( new_n521_, new_n518_, new_n520_ );
nand g371 ( new_n522_, new_n515_, new_n517_, new_n519_ );
nand g372 ( new_n523_, new_n521_, N219, new_n522_ );
nand g373 ( new_n524_, new_n520_, N228 );
not g374 ( new_n525_, new_n524_ );
nand g375 ( new_n526_, new_n459_, N189, N237 );
nand g376 ( new_n527_, new_n459_, N246 );
nand g377 ( new_n528_, new_n399_, N189 );
nand g378 ( new_n529_, N255, N259 );
nand g379 ( new_n530_, N111, N210 );
nand g380 ( new_n531_, new_n528_, new_n529_, new_n530_ );
not g381 ( new_n532_, new_n531_ );
nand g382 ( new_n533_, new_n526_, new_n527_, new_n532_ );
nor g383 ( new_n534_, new_n525_, new_n533_ );
nand g384 ( new_n535_, new_n523_, new_n534_ );
nand g385 ( new_n536_, new_n535_, keyIn_0_58 );
not g386 ( new_n537_, keyIn_0_58 );
nand g387 ( new_n538_, new_n523_, new_n537_, new_n534_ );
nand g388 ( N864, new_n536_, new_n538_ );
nand g389 ( new_n540_, new_n452_, new_n443_ );
not g390 ( new_n541_, new_n540_ );
nand g391 ( new_n542_, new_n512_, new_n541_ );
nand g392 ( new_n543_, new_n511_, new_n382_, new_n540_ );
nand g393 ( new_n544_, new_n542_, N219, new_n543_ );
nand g394 ( new_n545_, new_n541_, N228 );
not g395 ( new_n546_, new_n545_ );
nand g396 ( new_n547_, new_n453_, N237 );
nand g397 ( new_n548_, new_n451_, N246 );
nand g398 ( new_n549_, new_n399_, N195 );
nand g399 ( new_n550_, N255, N260 );
nand g400 ( new_n551_, N116, N210 );
nand g401 ( new_n552_, new_n549_, new_n550_, new_n551_ );
not g402 ( new_n553_, new_n552_ );
nand g403 ( new_n554_, new_n547_, new_n548_, new_n553_ );
nor g404 ( new_n555_, new_n546_, new_n554_ );
nand g405 ( new_n556_, new_n555_, new_n544_ );
nand g406 ( new_n557_, new_n556_, keyIn_0_59 );
not g407 ( new_n558_, keyIn_0_59 );
nand g408 ( new_n559_, new_n555_, new_n544_, new_n558_ );
nand g409 ( N865, new_n557_, new_n559_ );
not g410 ( new_n561_, keyIn_0_55 );
not g411 ( new_n562_, keyIn_0_54 );
not g412 ( new_n563_, keyIn_0_50 );
nand g413 ( new_n564_, new_n473_, new_n493_ );
nand g414 ( new_n565_, new_n564_, new_n563_ );
nand g415 ( new_n566_, new_n473_, keyIn_0_50, new_n493_ );
nand g416 ( new_n567_, new_n565_, new_n566_ );
nand g417 ( new_n568_, new_n567_, new_n492_ );
nand g418 ( new_n569_, new_n568_, keyIn_0_51 );
not g419 ( new_n570_, keyIn_0_51 );
nand g420 ( new_n571_, new_n567_, new_n570_, new_n492_ );
not g421 ( new_n572_, keyIn_0_38 );
not g422 ( new_n573_, keyIn_0_22 );
not g423 ( new_n574_, keyIn_0_17 );
nand g424 ( new_n575_, new_n351_, N17, new_n357_ );
nor g425 ( new_n576_, new_n575_, new_n574_ );
not g426 ( new_n577_, new_n576_ );
nand g427 ( new_n578_, new_n575_, new_n574_ );
nand g428 ( new_n579_, new_n577_, new_n367_, new_n578_ );
not g429 ( new_n580_, new_n579_ );
nand g430 ( new_n581_, new_n580_, new_n573_ );
nand g431 ( new_n582_, new_n579_, keyIn_0_22 );
nand g432 ( new_n583_, new_n581_, new_n582_ );
not g433 ( new_n584_, keyIn_0_16 );
nand g434 ( new_n585_, new_n351_, N55, new_n329_ );
nand g435 ( new_n586_, new_n585_, new_n584_ );
not g436 ( new_n587_, new_n586_ );
nor g437 ( new_n588_, new_n585_, new_n584_ );
nor g438 ( new_n589_, new_n587_, new_n588_ );
nand g439 ( new_n590_, new_n589_, N149 );
nand g440 ( new_n591_, new_n583_, new_n590_ );
nand g441 ( new_n592_, new_n591_, keyIn_0_29 );
not g442 ( new_n593_, keyIn_0_29 );
nand g443 ( new_n594_, new_n583_, new_n593_, new_n590_ );
nand g444 ( new_n595_, new_n592_, new_n594_ );
nand g445 ( new_n596_, new_n475_, N101 );
nand g446 ( new_n597_, N17, N138 );
nand g447 ( new_n598_, new_n596_, new_n597_ );
nand g448 ( new_n599_, new_n598_, keyIn_0_32 );
not g449 ( new_n600_, keyIn_0_32 );
nand g450 ( new_n601_, new_n596_, new_n600_, new_n597_ );
nand g451 ( new_n602_, new_n599_, new_n601_ );
nand g452 ( new_n603_, new_n595_, new_n602_ );
nand g453 ( new_n604_, new_n603_, new_n572_ );
nand g454 ( new_n605_, new_n595_, keyIn_0_38, new_n602_ );
nand g455 ( new_n606_, new_n604_, new_n232_, new_n605_ );
nand g456 ( new_n607_, new_n475_, N96 );
nand g457 ( new_n608_, new_n589_, N146 );
nand g458 ( new_n609_, N51, N138 );
nand g459 ( new_n610_, new_n608_, new_n579_, new_n609_ );
not g460 ( new_n611_, new_n610_ );
nand g461 ( new_n612_, new_n611_, new_n228_, new_n607_ );
nand g462 ( new_n613_, new_n606_, new_n612_ );
not g463 ( new_n614_, new_n613_ );
not g464 ( new_n615_, keyIn_0_39 );
not g465 ( new_n616_, keyIn_0_30 );
nand g466 ( new_n617_, new_n580_, keyIn_0_23 );
not g467 ( new_n618_, keyIn_0_23 );
nand g468 ( new_n619_, new_n579_, new_n618_ );
nand g469 ( new_n620_, new_n617_, new_n619_ );
nand g470 ( new_n621_, new_n589_, N153 );
nand g471 ( new_n622_, new_n620_, new_n621_ );
nand g472 ( new_n623_, new_n622_, new_n616_ );
nand g473 ( new_n624_, new_n620_, keyIn_0_30, new_n621_ );
nand g474 ( new_n625_, new_n623_, new_n624_ );
nand g475 ( new_n626_, new_n475_, N106 );
nand g476 ( new_n627_, N138, N152 );
nand g477 ( new_n628_, new_n626_, new_n627_ );
nand g478 ( new_n629_, new_n628_, keyIn_0_33 );
not g479 ( new_n630_, keyIn_0_33 );
nand g480 ( new_n631_, new_n626_, new_n630_, new_n627_ );
nand g481 ( new_n632_, new_n629_, new_n631_ );
nand g482 ( new_n633_, new_n625_, new_n632_ );
nand g483 ( new_n634_, new_n633_, new_n615_ );
nand g484 ( new_n635_, new_n625_, keyIn_0_39, new_n632_ );
nand g485 ( new_n636_, new_n634_, new_n233_, new_n635_ );
nand g486 ( new_n637_, new_n614_, new_n636_ );
not g487 ( new_n638_, new_n637_ );
nand g488 ( new_n639_, new_n569_, new_n562_, new_n571_, new_n638_ );
nand g489 ( new_n640_, new_n569_, new_n571_, new_n638_ );
nand g490 ( new_n641_, new_n640_, keyIn_0_54 );
not g491 ( new_n642_, keyIn_0_47 );
nand g492 ( new_n643_, new_n634_, new_n635_ );
nand g493 ( new_n644_, new_n643_, N177 );
not g494 ( new_n645_, new_n644_ );
nand g495 ( new_n646_, new_n614_, new_n645_ );
nor g496 ( new_n647_, new_n646_, new_n642_ );
nand g497 ( new_n648_, new_n646_, new_n642_ );
nand g498 ( new_n649_, new_n611_, new_n607_ );
nand g499 ( new_n650_, new_n649_, N165 );
nand g500 ( new_n651_, new_n604_, new_n605_ );
nand g501 ( new_n652_, new_n651_, N171 );
not g502 ( new_n653_, new_n652_ );
nand g503 ( new_n654_, new_n653_, new_n612_ );
nand g504 ( new_n655_, new_n648_, new_n650_, new_n654_ );
nor g505 ( new_n656_, new_n655_, new_n647_ );
nand g506 ( new_n657_, new_n641_, new_n639_, new_n656_ );
nand g507 ( new_n658_, new_n657_, new_n561_ );
nand g508 ( new_n659_, new_n641_, keyIn_0_55, new_n639_, new_n656_ );
nand g509 ( new_n660_, new_n658_, new_n659_ );
nand g510 ( new_n661_, new_n475_, N91 );
nand g511 ( new_n662_, new_n589_, N143 );
nand g512 ( new_n663_, N8, N138 );
nand g513 ( new_n664_, new_n662_, new_n579_, new_n663_ );
not g514 ( new_n665_, new_n664_ );
nand g515 ( new_n666_, new_n665_, new_n227_, new_n661_ );
nand g516 ( new_n667_, new_n660_, new_n666_ );
nand g517 ( new_n668_, new_n665_, new_n661_ );
nand g518 ( new_n669_, new_n668_, N159 );
nand g519 ( N866, new_n667_, new_n669_ );
nand g520 ( new_n671_, new_n569_, new_n571_ );
not g521 ( new_n672_, new_n671_ );
nand g522 ( new_n673_, new_n672_, new_n636_, new_n644_ );
nand g523 ( new_n674_, new_n644_, new_n636_ );
nand g524 ( new_n675_, new_n671_, new_n674_ );
nand g525 ( new_n676_, new_n673_, N219, new_n675_ );
nand g526 ( new_n677_, new_n644_, N228, new_n636_ );
not g527 ( new_n678_, new_n677_ );
nand g528 ( new_n679_, new_n645_, N237 );
nand g529 ( new_n680_, new_n643_, N246 );
nand g530 ( new_n681_, new_n399_, N177 );
nand g531 ( new_n682_, N101, N210 );
nand g532 ( new_n683_, new_n679_, new_n680_, new_n681_, new_n682_ );
nor g533 ( new_n684_, new_n683_, new_n678_ );
nand g534 ( new_n685_, new_n676_, new_n684_ );
nand g535 ( new_n686_, new_n685_, keyIn_0_60 );
not g536 ( new_n687_, keyIn_0_60 );
nand g537 ( new_n688_, new_n676_, new_n687_, new_n684_ );
nand g538 ( N874, new_n686_, new_n688_ );
nand g539 ( new_n690_, new_n669_, new_n666_ );
not g540 ( new_n691_, new_n690_ );
nand g541 ( new_n692_, new_n660_, new_n691_ );
nand g542 ( new_n693_, new_n658_, new_n659_, new_n690_ );
nand g543 ( new_n694_, new_n692_, N219, new_n693_ );
nand g544 ( new_n695_, new_n691_, N228 );
not g545 ( new_n696_, new_n695_ );
nand g546 ( new_n697_, new_n668_, N159, N237 );
nand g547 ( new_n698_, new_n668_, N246 );
nand g548 ( new_n699_, new_n371_, N210 );
nand g549 ( new_n700_, new_n399_, N159 );
nand g550 ( new_n701_, new_n697_, new_n698_, new_n699_, new_n700_ );
nor g551 ( new_n702_, new_n696_, new_n701_ );
nand g552 ( new_n703_, new_n694_, new_n702_ );
nand g553 ( new_n704_, new_n703_, keyIn_0_61 );
not g554 ( new_n705_, keyIn_0_61 );
nand g555 ( new_n706_, new_n694_, new_n705_, new_n702_ );
nand g556 ( N878, new_n704_, new_n706_ );
not g557 ( new_n708_, keyIn_0_62 );
not g558 ( new_n709_, keyIn_0_56 );
nand g559 ( new_n710_, new_n606_, new_n636_ );
not g560 ( new_n711_, new_n710_ );
nand g561 ( new_n712_, new_n569_, keyIn_0_53, new_n571_, new_n711_ );
not g562 ( new_n713_, keyIn_0_53 );
nand g563 ( new_n714_, new_n569_, new_n571_, new_n711_ );
nand g564 ( new_n715_, new_n714_, new_n713_ );
nand g565 ( new_n716_, new_n645_, new_n606_ );
nand g566 ( new_n717_, new_n716_, new_n652_ );
not g567 ( new_n718_, new_n717_ );
nand g568 ( new_n719_, new_n715_, new_n712_, new_n718_ );
nand g569 ( new_n720_, new_n719_, new_n709_ );
nand g570 ( new_n721_, new_n715_, keyIn_0_56, new_n712_, new_n718_ );
nand g571 ( new_n722_, new_n720_, new_n721_ );
nand g572 ( new_n723_, new_n650_, new_n612_ );
nand g573 ( new_n724_, new_n722_, new_n723_ );
not g574 ( new_n725_, new_n723_ );
nand g575 ( new_n726_, new_n720_, new_n721_, new_n725_ );
nand g576 ( new_n727_, new_n724_, N219, new_n726_ );
nand g577 ( new_n728_, new_n725_, N228 );
not g578 ( new_n729_, new_n728_ );
nand g579 ( new_n730_, new_n649_, N165, N237 );
nand g580 ( new_n731_, new_n649_, N246 );
nand g581 ( new_n732_, new_n399_, N165 );
nand g582 ( new_n733_, N91, N210 );
nand g583 ( new_n734_, new_n730_, new_n731_, new_n732_, new_n733_ );
nor g584 ( new_n735_, new_n729_, new_n734_ );
nand g585 ( new_n736_, new_n727_, new_n735_ );
nand g586 ( new_n737_, new_n736_, new_n708_ );
nand g587 ( new_n738_, new_n727_, keyIn_0_62, new_n735_ );
nand g588 ( N879, new_n737_, new_n738_ );
not g589 ( new_n740_, keyIn_0_63 );
nand g590 ( new_n741_, new_n672_, new_n636_ );
nand g591 ( new_n742_, new_n741_, new_n644_ );
nand g592 ( new_n743_, new_n652_, new_n606_ );
not g593 ( new_n744_, new_n743_ );
nand g594 ( new_n745_, new_n742_, new_n744_ );
nand g595 ( new_n746_, new_n741_, new_n644_, new_n743_ );
nand g596 ( new_n747_, new_n745_, N219, new_n746_ );
nand g597 ( new_n748_, new_n744_, N228 );
not g598 ( new_n749_, new_n748_ );
nand g599 ( new_n750_, new_n653_, N237 );
nand g600 ( new_n751_, new_n651_, N246 );
nand g601 ( new_n752_, new_n399_, N171 );
nand g602 ( new_n753_, N96, N210 );
nand g603 ( new_n754_, new_n750_, new_n751_, new_n752_, new_n753_ );
nor g604 ( new_n755_, new_n749_, new_n754_ );
nand g605 ( new_n756_, new_n747_, new_n755_ );
nand g606 ( new_n757_, new_n756_, new_n740_ );
nand g607 ( new_n758_, new_n747_, keyIn_0_63, new_n755_ );
nand g608 ( N880, new_n757_, new_n758_ );
endmodule