module add_mul_sub_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation_0_, 
        operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239;

  OR2_X1 U609 ( .A1(n593), .A2(n594), .ZN(Result_9_) );
  OR2_X1 U610 ( .A1(n595), .A2(n596), .ZN(n594) );
  AND2_X1 U611 ( .A1(n597), .A2(n598), .ZN(n596) );
  OR2_X1 U612 ( .A1(n599), .A2(n600), .ZN(n598) );
  OR2_X1 U613 ( .A1(n601), .A2(n602), .ZN(n600) );
  AND2_X1 U614 ( .A1(n603), .A2(n604), .ZN(n602) );
  INV_X1 U615 ( .A(n605), .ZN(n604) );
  AND2_X1 U616 ( .A1(n606), .A2(n607), .ZN(n601) );
  AND2_X1 U617 ( .A1(n608), .A2(n609), .ZN(n599) );
  INV_X1 U618 ( .A(n610), .ZN(n609) );
  AND2_X1 U619 ( .A1(n611), .A2(n612), .ZN(n595) );
  INV_X1 U620 ( .A(n597), .ZN(n612) );
  AND2_X1 U621 ( .A1(n613), .A2(n614), .ZN(n597) );
  OR2_X1 U622 ( .A1(a_1_), .A2(b_1_), .ZN(n613) );
  OR2_X1 U623 ( .A1(n615), .A2(n616), .ZN(n611) );
  OR2_X1 U624 ( .A1(n617), .A2(n618), .ZN(n616) );
  AND2_X1 U625 ( .A1(n603), .A2(n605), .ZN(n618) );
  AND2_X1 U626 ( .A1(n619), .A2(n606), .ZN(n617) );
  INV_X1 U627 ( .A(n607), .ZN(n619) );
  AND2_X1 U628 ( .A1(n608), .A2(n610), .ZN(n615) );
  AND2_X1 U629 ( .A1(n620), .A2(n621), .ZN(n593) );
  XNOR2_X1 U630 ( .A(n622), .B(n623), .ZN(n621) );
  XOR2_X1 U631 ( .A(n624), .B(n625), .Z(n623) );
  OR2_X1 U632 ( .A1(n626), .A2(n627), .ZN(Result_8_) );
  OR2_X1 U633 ( .A1(n628), .A2(n629), .ZN(n627) );
  AND2_X1 U634 ( .A1(n630), .A2(n631), .ZN(n629) );
  OR2_X1 U635 ( .A1(n632), .A2(n633), .ZN(n630) );
  OR2_X1 U636 ( .A1(n634), .A2(n635), .ZN(n633) );
  AND2_X1 U637 ( .A1(n636), .A2(n603), .ZN(n635) );
  INV_X1 U638 ( .A(n637), .ZN(n636) );
  AND2_X1 U639 ( .A1(n606), .A2(n638), .ZN(n634) );
  AND2_X1 U640 ( .A1(n639), .A2(n608), .ZN(n632) );
  INV_X1 U641 ( .A(n640), .ZN(n639) );
  AND2_X1 U642 ( .A1(n641), .A2(n642), .ZN(n628) );
  OR2_X1 U643 ( .A1(n643), .A2(n644), .ZN(n642) );
  OR2_X1 U644 ( .A1(n645), .A2(n646), .ZN(n644) );
  AND2_X1 U645 ( .A1(n603), .A2(n637), .ZN(n646) );
  AND2_X1 U646 ( .A1(n647), .A2(n606), .ZN(n645) );
  INV_X1 U647 ( .A(n638), .ZN(n647) );
  OR2_X1 U648 ( .A1(n648), .A2(n649), .ZN(n638) );
  AND2_X1 U649 ( .A1(n650), .A2(n651), .ZN(n649) );
  AND2_X1 U650 ( .A1(n607), .A2(n614), .ZN(n648) );
  OR2_X1 U651 ( .A1(n652), .A2(n653), .ZN(n607) );
  AND2_X1 U652 ( .A1(n654), .A2(n655), .ZN(n653) );
  AND2_X1 U653 ( .A1(n656), .A2(n657), .ZN(n652) );
  AND2_X1 U654 ( .A1(n608), .A2(n640), .ZN(n643) );
  INV_X1 U655 ( .A(n631), .ZN(n641) );
  OR2_X1 U656 ( .A1(n658), .A2(n659), .ZN(n631) );
  AND2_X1 U657 ( .A1(n620), .A2(n660), .ZN(n626) );
  XNOR2_X1 U658 ( .A(n661), .B(n662), .ZN(n660) );
  XOR2_X1 U659 ( .A(n663), .B(n664), .Z(n662) );
  OR2_X1 U660 ( .A1(n665), .A2(n666), .ZN(Result_7_) );
  AND2_X1 U661 ( .A1(n620), .A2(n667), .ZN(n665) );
  XOR2_X1 U662 ( .A(n668), .B(n669), .Z(n667) );
  OR2_X1 U663 ( .A1(n670), .A2(n666), .ZN(Result_6_) );
  AND2_X1 U664 ( .A1(n671), .A2(n620), .ZN(n670) );
  AND2_X1 U665 ( .A1(n672), .A2(n673), .ZN(n671) );
  OR2_X1 U666 ( .A1(n674), .A2(n675), .ZN(n672) );
  XOR2_X1 U667 ( .A(n676), .B(n677), .Z(n675) );
  INV_X1 U668 ( .A(n678), .ZN(n674) );
  OR2_X1 U669 ( .A1(n679), .A2(n666), .ZN(Result_5_) );
  AND2_X1 U670 ( .A1(n620), .A2(n680), .ZN(n679) );
  XOR2_X1 U671 ( .A(n681), .B(n682), .Z(n680) );
  AND2_X1 U672 ( .A1(n673), .A2(n683), .ZN(n682) );
  OR2_X1 U673 ( .A1(n684), .A2(n666), .ZN(Result_4_) );
  AND2_X1 U674 ( .A1(n685), .A2(n620), .ZN(n684) );
  XNOR2_X1 U675 ( .A(n686), .B(n687), .ZN(n685) );
  OR2_X1 U676 ( .A1(n688), .A2(n666), .ZN(Result_3_) );
  AND2_X1 U677 ( .A1(n620), .A2(n689), .ZN(n688) );
  XOR2_X1 U678 ( .A(n690), .B(n691), .Z(n689) );
  AND2_X1 U679 ( .A1(n692), .A2(n693), .ZN(n691) );
  OR2_X1 U680 ( .A1(n694), .A2(n695), .ZN(n693) );
  INV_X1 U681 ( .A(n696), .ZN(n692) );
  OR2_X1 U682 ( .A1(n697), .A2(n666), .ZN(Result_2_) );
  AND2_X1 U683 ( .A1(n698), .A2(n620), .ZN(n697) );
  XOR2_X1 U684 ( .A(n699), .B(n700), .Z(n698) );
  OR2_X1 U685 ( .A1(n701), .A2(n666), .ZN(Result_1_) );
  AND2_X1 U686 ( .A1(n620), .A2(n702), .ZN(n701) );
  XOR2_X1 U687 ( .A(n703), .B(n704), .Z(n702) );
  AND2_X1 U688 ( .A1(n705), .A2(n706), .ZN(n704) );
  OR2_X1 U689 ( .A1(n707), .A2(n708), .ZN(n706) );
  AND2_X1 U690 ( .A1(n709), .A2(n710), .ZN(n707) );
  INV_X1 U691 ( .A(n711), .ZN(n705) );
  OR2_X1 U692 ( .A1(n712), .A2(n713), .ZN(Result_15_) );
  AND2_X1 U693 ( .A1(n620), .A2(n714), .ZN(n713) );
  AND2_X1 U694 ( .A1(n715), .A2(n716), .ZN(n712) );
  OR2_X1 U695 ( .A1(n606), .A2(n717), .ZN(n716) );
  OR2_X1 U696 ( .A1(n608), .A2(n603), .ZN(n717) );
  OR2_X1 U697 ( .A1(n718), .A2(n719), .ZN(n715) );
  OR2_X1 U698 ( .A1(n720), .A2(n721), .ZN(Result_14_) );
  OR2_X1 U699 ( .A1(n722), .A2(n723), .ZN(n721) );
  AND2_X1 U700 ( .A1(n724), .A2(n725), .ZN(n723) );
  OR2_X1 U701 ( .A1(n726), .A2(n727), .ZN(n725) );
  OR2_X1 U702 ( .A1(n728), .A2(n729), .ZN(n727) );
  AND2_X1 U703 ( .A1(n603), .A2(n718), .ZN(n729) );
  AND2_X1 U704 ( .A1(n606), .A2(n714), .ZN(n728) );
  INV_X1 U705 ( .A(n730), .ZN(n714) );
  AND2_X1 U706 ( .A1(n608), .A2(n719), .ZN(n726) );
  INV_X1 U707 ( .A(n731), .ZN(n724) );
  AND2_X1 U708 ( .A1(n732), .A2(n731), .ZN(n722) );
  OR2_X1 U709 ( .A1(n733), .A2(n734), .ZN(n731) );
  OR2_X1 U710 ( .A1(n735), .A2(n736), .ZN(n732) );
  OR2_X1 U711 ( .A1(n737), .A2(n738), .ZN(n736) );
  AND2_X1 U712 ( .A1(n603), .A2(n739), .ZN(n738) );
  AND2_X1 U713 ( .A1(n606), .A2(n730), .ZN(n737) );
  AND2_X1 U714 ( .A1(n608), .A2(n740), .ZN(n735) );
  AND2_X1 U715 ( .A1(n620), .A2(n741), .ZN(n720) );
  OR2_X1 U716 ( .A1(n742), .A2(n743), .ZN(n741) );
  OR2_X1 U717 ( .A1(n744), .A2(n745), .ZN(n743) );
  AND2_X1 U718 ( .A1(n719), .A2(a_6_), .ZN(n745) );
  INV_X1 U719 ( .A(n740), .ZN(n719) );
  AND2_X1 U720 ( .A1(n734), .A2(a_7_), .ZN(n744) );
  INV_X1 U721 ( .A(n746), .ZN(n734) );
  OR2_X1 U722 ( .A1(n747), .A2(n748), .ZN(n742) );
  AND2_X1 U723 ( .A1(n718), .A2(b_6_), .ZN(n748) );
  AND2_X1 U724 ( .A1(n733), .A2(b_7_), .ZN(n747) );
  OR2_X1 U725 ( .A1(n749), .A2(n750), .ZN(Result_13_) );
  OR2_X1 U726 ( .A1(n751), .A2(n752), .ZN(n750) );
  AND2_X1 U727 ( .A1(n753), .A2(n754), .ZN(n752) );
  OR2_X1 U728 ( .A1(n755), .A2(n756), .ZN(n754) );
  OR2_X1 U729 ( .A1(n757), .A2(n758), .ZN(n756) );
  AND2_X1 U730 ( .A1(n603), .A2(n759), .ZN(n758) );
  AND2_X1 U731 ( .A1(n606), .A2(n760), .ZN(n757) );
  INV_X1 U732 ( .A(n761), .ZN(n760) );
  AND2_X1 U733 ( .A1(n608), .A2(n762), .ZN(n755) );
  INV_X1 U734 ( .A(n763), .ZN(n753) );
  AND2_X1 U735 ( .A1(n763), .A2(n764), .ZN(n751) );
  OR2_X1 U736 ( .A1(n765), .A2(n766), .ZN(n764) );
  OR2_X1 U737 ( .A1(n767), .A2(n768), .ZN(n766) );
  AND2_X1 U738 ( .A1(n603), .A2(n769), .ZN(n768) );
  INV_X1 U739 ( .A(n759), .ZN(n769) );
  AND2_X1 U740 ( .A1(n606), .A2(n761), .ZN(n767) );
  AND2_X1 U741 ( .A1(n608), .A2(n770), .ZN(n765) );
  XNOR2_X1 U742 ( .A(n771), .B(a_5_), .ZN(n763) );
  AND2_X1 U743 ( .A1(n620), .A2(n772), .ZN(n749) );
  XNOR2_X1 U744 ( .A(n773), .B(n774), .ZN(n772) );
  XOR2_X1 U745 ( .A(n775), .B(n776), .Z(n774) );
  OR2_X1 U746 ( .A1(n777), .A2(n778), .ZN(Result_12_) );
  OR2_X1 U747 ( .A1(n779), .A2(n780), .ZN(n778) );
  AND2_X1 U748 ( .A1(n781), .A2(n782), .ZN(n780) );
  OR2_X1 U749 ( .A1(n783), .A2(n784), .ZN(n782) );
  OR2_X1 U750 ( .A1(n785), .A2(n786), .ZN(n784) );
  AND2_X1 U751 ( .A1(n603), .A2(n787), .ZN(n786) );
  AND2_X1 U752 ( .A1(n788), .A2(n606), .ZN(n785) );
  INV_X1 U753 ( .A(n789), .ZN(n788) );
  AND2_X1 U754 ( .A1(n608), .A2(n790), .ZN(n783) );
  INV_X1 U755 ( .A(n791), .ZN(n781) );
  AND2_X1 U756 ( .A1(n791), .A2(n792), .ZN(n779) );
  OR2_X1 U757 ( .A1(n793), .A2(n794), .ZN(n792) );
  OR2_X1 U758 ( .A1(n795), .A2(n796), .ZN(n794) );
  AND2_X1 U759 ( .A1(n603), .A2(n797), .ZN(n796) );
  INV_X1 U760 ( .A(n787), .ZN(n797) );
  AND2_X1 U761 ( .A1(n606), .A2(n789), .ZN(n795) );
  AND2_X1 U762 ( .A1(n608), .A2(n798), .ZN(n793) );
  INV_X1 U763 ( .A(n790), .ZN(n798) );
  XNOR2_X1 U764 ( .A(n799), .B(a_4_), .ZN(n791) );
  AND2_X1 U765 ( .A1(n620), .A2(n800), .ZN(n777) );
  XNOR2_X1 U766 ( .A(n801), .B(n802), .ZN(n800) );
  XOR2_X1 U767 ( .A(n803), .B(n804), .Z(n802) );
  OR2_X1 U768 ( .A1(n805), .A2(n806), .ZN(Result_11_) );
  OR2_X1 U769 ( .A1(n807), .A2(n808), .ZN(n806) );
  AND2_X1 U770 ( .A1(n809), .A2(n810), .ZN(n808) );
  OR2_X1 U771 ( .A1(n811), .A2(n812), .ZN(n810) );
  OR2_X1 U772 ( .A1(n813), .A2(n814), .ZN(n812) );
  AND2_X1 U773 ( .A1(n603), .A2(n815), .ZN(n814) );
  AND2_X1 U774 ( .A1(n816), .A2(n606), .ZN(n813) );
  INV_X1 U775 ( .A(n817), .ZN(n816) );
  AND2_X1 U776 ( .A1(n608), .A2(n818), .ZN(n811) );
  INV_X1 U777 ( .A(n819), .ZN(n809) );
  AND2_X1 U778 ( .A1(n819), .A2(n820), .ZN(n807) );
  OR2_X1 U779 ( .A1(n821), .A2(n822), .ZN(n820) );
  OR2_X1 U780 ( .A1(n823), .A2(n824), .ZN(n822) );
  AND2_X1 U781 ( .A1(n603), .A2(n825), .ZN(n824) );
  INV_X1 U782 ( .A(n815), .ZN(n825) );
  AND2_X1 U783 ( .A1(n606), .A2(n817), .ZN(n823) );
  AND2_X1 U784 ( .A1(n608), .A2(n826), .ZN(n821) );
  INV_X1 U785 ( .A(n818), .ZN(n826) );
  XNOR2_X1 U786 ( .A(n827), .B(a_3_), .ZN(n819) );
  AND2_X1 U787 ( .A1(n620), .A2(n828), .ZN(n805) );
  XNOR2_X1 U788 ( .A(n829), .B(n830), .ZN(n828) );
  XOR2_X1 U789 ( .A(n831), .B(n832), .Z(n830) );
  OR2_X1 U790 ( .A1(n833), .A2(n834), .ZN(Result_10_) );
  OR2_X1 U791 ( .A1(n835), .A2(n836), .ZN(n834) );
  AND2_X1 U792 ( .A1(n837), .A2(n838), .ZN(n836) );
  OR2_X1 U793 ( .A1(n839), .A2(n840), .ZN(n838) );
  OR2_X1 U794 ( .A1(n841), .A2(n842), .ZN(n840) );
  AND2_X1 U795 ( .A1(n603), .A2(n843), .ZN(n842) );
  AND2_X1 U796 ( .A1(n844), .A2(n606), .ZN(n841) );
  INV_X1 U797 ( .A(n656), .ZN(n844) );
  AND2_X1 U798 ( .A1(n608), .A2(n845), .ZN(n839) );
  INV_X1 U799 ( .A(n846), .ZN(n837) );
  AND2_X1 U800 ( .A1(n846), .A2(n847), .ZN(n835) );
  OR2_X1 U801 ( .A1(n848), .A2(n849), .ZN(n847) );
  OR2_X1 U802 ( .A1(n850), .A2(n851), .ZN(n849) );
  AND2_X1 U803 ( .A1(n603), .A2(n852), .ZN(n851) );
  INV_X1 U804 ( .A(n843), .ZN(n852) );
  AND2_X1 U805 ( .A1(n606), .A2(n656), .ZN(n850) );
  OR2_X1 U806 ( .A1(n853), .A2(n854), .ZN(n656) );
  AND2_X1 U807 ( .A1(n855), .A2(n827), .ZN(n854) );
  AND2_X1 U808 ( .A1(n817), .A2(n856), .ZN(n853) );
  OR2_X1 U809 ( .A1(n857), .A2(n858), .ZN(n817) );
  AND2_X1 U810 ( .A1(n859), .A2(n799), .ZN(n858) );
  AND2_X1 U811 ( .A1(n789), .A2(n860), .ZN(n857) );
  OR2_X1 U812 ( .A1(n861), .A2(n862), .ZN(n789) );
  AND2_X1 U813 ( .A1(n863), .A2(n771), .ZN(n862) );
  AND2_X1 U814 ( .A1(n761), .A2(n864), .ZN(n861) );
  AND2_X1 U815 ( .A1(n865), .A2(n866), .ZN(n761) );
  OR2_X1 U816 ( .A1(n730), .A2(n867), .ZN(n865) );
  AND2_X1 U817 ( .A1(n868), .A2(n869), .ZN(n867) );
  AND2_X1 U818 ( .A1(n870), .A2(n871), .ZN(n606) );
  AND2_X1 U819 ( .A1(n608), .A2(n872), .ZN(n848) );
  INV_X1 U820 ( .A(n845), .ZN(n872) );
  XNOR2_X1 U821 ( .A(n655), .B(a_2_), .ZN(n846) );
  AND2_X1 U822 ( .A1(n620), .A2(n873), .ZN(n833) );
  XNOR2_X1 U823 ( .A(n874), .B(n875), .ZN(n873) );
  XOR2_X1 U824 ( .A(n876), .B(n877), .Z(n875) );
  OR2_X1 U825 ( .A1(n878), .A2(n666), .ZN(Result_0_) );
  OR2_X1 U826 ( .A1(n879), .A2(n880), .ZN(n666) );
  AND2_X1 U827 ( .A1(n608), .A2(n881), .ZN(n880) );
  OR2_X1 U828 ( .A1(n882), .A2(n659), .ZN(n881) );
  INV_X1 U829 ( .A(n883), .ZN(n659) );
  AND2_X1 U830 ( .A1(n640), .A2(n884), .ZN(n882) );
  OR2_X1 U831 ( .A1(n885), .A2(n886), .ZN(n640) );
  AND2_X1 U832 ( .A1(n610), .A2(n650), .ZN(n886) );
  AND2_X1 U833 ( .A1(b_1_), .A2(n887), .ZN(n885) );
  OR2_X1 U834 ( .A1(n650), .A2(n610), .ZN(n887) );
  OR2_X1 U835 ( .A1(n888), .A2(n889), .ZN(n610) );
  AND2_X1 U836 ( .A1(n845), .A2(n654), .ZN(n889) );
  AND2_X1 U837 ( .A1(b_2_), .A2(n890), .ZN(n888) );
  OR2_X1 U838 ( .A1(n654), .A2(n845), .ZN(n890) );
  OR2_X1 U839 ( .A1(n891), .A2(n892), .ZN(n845) );
  AND2_X1 U840 ( .A1(n818), .A2(n855), .ZN(n892) );
  AND2_X1 U841 ( .A1(b_3_), .A2(n893), .ZN(n891) );
  OR2_X1 U842 ( .A1(n855), .A2(n818), .ZN(n893) );
  OR2_X1 U843 ( .A1(n894), .A2(n895), .ZN(n818) );
  AND2_X1 U844 ( .A1(n790), .A2(n859), .ZN(n895) );
  AND2_X1 U845 ( .A1(b_4_), .A2(n896), .ZN(n894) );
  OR2_X1 U846 ( .A1(n859), .A2(n790), .ZN(n896) );
  OR2_X1 U847 ( .A1(n897), .A2(n898), .ZN(n790) );
  AND2_X1 U848 ( .A1(n762), .A2(n863), .ZN(n898) );
  AND2_X1 U849 ( .A1(b_5_), .A2(n899), .ZN(n897) );
  OR2_X1 U850 ( .A1(n863), .A2(n762), .ZN(n899) );
  INV_X1 U851 ( .A(n770), .ZN(n762) );
  AND2_X1 U852 ( .A1(n746), .A2(n900), .ZN(n770) );
  OR2_X1 U853 ( .A1(n740), .A2(n733), .ZN(n900) );
  OR2_X1 U854 ( .A1(a_7_), .A2(n901), .ZN(n740) );
  AND2_X1 U855 ( .A1(n871), .A2(operation_1_), .ZN(n608) );
  INV_X1 U856 ( .A(operation_0_), .ZN(n871) );
  AND2_X1 U857 ( .A1(n902), .A2(n603), .ZN(n879) );
  AND2_X1 U858 ( .A1(n870), .A2(operation_0_), .ZN(n603) );
  INV_X1 U859 ( .A(operation_1_), .ZN(n870) );
  AND2_X1 U860 ( .A1(n903), .A2(n883), .ZN(n902) );
  OR2_X1 U861 ( .A1(a_0_), .A2(n904), .ZN(n883) );
  OR2_X1 U862 ( .A1(n658), .A2(n637), .ZN(n903) );
  OR2_X1 U863 ( .A1(n905), .A2(n906), .ZN(n637) );
  AND2_X1 U864 ( .A1(a_1_), .A2(n605), .ZN(n906) );
  AND2_X1 U865 ( .A1(n907), .A2(n651), .ZN(n905) );
  OR2_X1 U866 ( .A1(a_1_), .A2(n605), .ZN(n907) );
  OR2_X1 U867 ( .A1(n908), .A2(n909), .ZN(n605) );
  AND2_X1 U868 ( .A1(a_2_), .A2(n843), .ZN(n909) );
  AND2_X1 U869 ( .A1(n910), .A2(n655), .ZN(n908) );
  OR2_X1 U870 ( .A1(a_2_), .A2(n843), .ZN(n910) );
  OR2_X1 U871 ( .A1(n911), .A2(n912), .ZN(n843) );
  AND2_X1 U872 ( .A1(a_3_), .A2(n815), .ZN(n912) );
  AND2_X1 U873 ( .A1(n913), .A2(n827), .ZN(n911) );
  OR2_X1 U874 ( .A1(a_3_), .A2(n815), .ZN(n913) );
  OR2_X1 U875 ( .A1(n914), .A2(n915), .ZN(n815) );
  AND2_X1 U876 ( .A1(a_4_), .A2(n787), .ZN(n915) );
  AND2_X1 U877 ( .A1(n916), .A2(n799), .ZN(n914) );
  OR2_X1 U878 ( .A1(a_4_), .A2(n787), .ZN(n916) );
  OR2_X1 U879 ( .A1(n917), .A2(n918), .ZN(n787) );
  AND2_X1 U880 ( .A1(a_5_), .A2(n759), .ZN(n918) );
  AND2_X1 U881 ( .A1(n919), .A2(n771), .ZN(n917) );
  OR2_X1 U882 ( .A1(a_5_), .A2(n759), .ZN(n919) );
  OR2_X1 U883 ( .A1(n920), .A2(n733), .ZN(n759) );
  AND2_X1 U884 ( .A1(n869), .A2(a_6_), .ZN(n733) );
  AND2_X1 U885 ( .A1(n718), .A2(n746), .ZN(n920) );
  OR2_X1 U886 ( .A1(a_6_), .A2(n869), .ZN(n746) );
  INV_X1 U887 ( .A(n739), .ZN(n718) );
  OR2_X1 U888 ( .A1(b_7_), .A2(n921), .ZN(n739) );
  INV_X1 U889 ( .A(n884), .ZN(n658) );
  OR2_X1 U890 ( .A1(b_0_), .A2(n922), .ZN(n884) );
  AND2_X1 U891 ( .A1(n620), .A2(n923), .ZN(n878) );
  OR2_X1 U892 ( .A1(n924), .A2(n925), .ZN(n923) );
  OR2_X1 U893 ( .A1(n711), .A2(n926), .ZN(n925) );
  AND2_X1 U894 ( .A1(n703), .A2(n708), .ZN(n926) );
  AND2_X1 U895 ( .A1(n699), .A2(n700), .ZN(n703) );
  XOR2_X1 U896 ( .A(n710), .B(n709), .Z(n700) );
  OR2_X1 U897 ( .A1(n927), .A2(n928), .ZN(n699) );
  INV_X1 U898 ( .A(n929), .ZN(n928) );
  OR2_X1 U899 ( .A1(n930), .A2(n696), .ZN(n927) );
  AND2_X1 U900 ( .A1(n694), .A2(n695), .ZN(n696) );
  AND2_X1 U901 ( .A1(n931), .A2(n932), .ZN(n695) );
  AND2_X1 U902 ( .A1(n690), .A2(n694), .ZN(n930) );
  AND2_X1 U903 ( .A1(n933), .A2(n929), .ZN(n694) );
  OR2_X1 U904 ( .A1(n934), .A2(n935), .ZN(n929) );
  INV_X1 U905 ( .A(n936), .ZN(n933) );
  AND2_X1 U906 ( .A1(n934), .A2(n935), .ZN(n936) );
  OR2_X1 U907 ( .A1(n937), .A2(n938), .ZN(n935) );
  AND2_X1 U908 ( .A1(n939), .A2(n940), .ZN(n938) );
  AND2_X1 U909 ( .A1(n941), .A2(n942), .ZN(n937) );
  OR2_X1 U910 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U911 ( .A(n943), .B(n944), .Z(n934) );
  XOR2_X1 U912 ( .A(n945), .B(n946), .Z(n944) );
  AND2_X1 U913 ( .A1(n947), .A2(n687), .ZN(n690) );
  XOR2_X1 U914 ( .A(n932), .B(n931), .Z(n687) );
  INV_X1 U915 ( .A(n948), .ZN(n931) );
  OR2_X1 U916 ( .A1(n949), .A2(n950), .ZN(n948) );
  AND2_X1 U917 ( .A1(n951), .A2(n952), .ZN(n950) );
  AND2_X1 U918 ( .A1(n953), .A2(n954), .ZN(n949) );
  OR2_X1 U919 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U920 ( .A(n955), .B(n941), .Z(n932) );
  XOR2_X1 U921 ( .A(n956), .B(n957), .Z(n941) );
  XOR2_X1 U922 ( .A(n958), .B(n959), .Z(n957) );
  XNOR2_X1 U923 ( .A(n940), .B(n939), .ZN(n955) );
  OR2_X1 U924 ( .A1(n960), .A2(n961), .ZN(n939) );
  AND2_X1 U925 ( .A1(n962), .A2(n963), .ZN(n961) );
  AND2_X1 U926 ( .A1(n964), .A2(n965), .ZN(n960) );
  OR2_X1 U927 ( .A1(n963), .A2(n962), .ZN(n965) );
  OR2_X1 U928 ( .A1(n827), .A2(n922), .ZN(n940) );
  INV_X1 U929 ( .A(n686), .ZN(n947) );
  AND2_X1 U930 ( .A1(n966), .A2(n967), .ZN(n686) );
  AND2_X1 U931 ( .A1(n968), .A2(n969), .ZN(n966) );
  OR2_X1 U932 ( .A1(n683), .A2(n681), .ZN(n969) );
  OR2_X1 U933 ( .A1(n673), .A2(n681), .ZN(n968) );
  OR2_X1 U934 ( .A1(n970), .A2(n971), .ZN(n681) );
  INV_X1 U935 ( .A(n967), .ZN(n971) );
  OR2_X1 U936 ( .A1(n972), .A2(n973), .ZN(n967) );
  AND2_X1 U937 ( .A1(n972), .A2(n973), .ZN(n970) );
  OR2_X1 U938 ( .A1(n974), .A2(n975), .ZN(n973) );
  AND2_X1 U939 ( .A1(n976), .A2(n977), .ZN(n975) );
  AND2_X1 U940 ( .A1(n978), .A2(n979), .ZN(n974) );
  OR2_X1 U941 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U942 ( .A(n953), .B(n980), .Z(n972) );
  XOR2_X1 U943 ( .A(n952), .B(n951), .Z(n980) );
  OR2_X1 U944 ( .A1(n799), .A2(n922), .ZN(n951) );
  OR2_X1 U945 ( .A1(n981), .A2(n982), .ZN(n952) );
  AND2_X1 U946 ( .A1(n983), .A2(n984), .ZN(n982) );
  AND2_X1 U947 ( .A1(n985), .A2(n986), .ZN(n981) );
  OR2_X1 U948 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U949 ( .A(n987), .B(n964), .ZN(n953) );
  XNOR2_X1 U950 ( .A(n988), .B(n989), .ZN(n964) );
  XNOR2_X1 U951 ( .A(n657), .B(n990), .ZN(n988) );
  XNOR2_X1 U952 ( .A(n963), .B(n962), .ZN(n987) );
  OR2_X1 U953 ( .A1(n991), .A2(n992), .ZN(n962) );
  AND2_X1 U954 ( .A1(n993), .A2(n994), .ZN(n992) );
  AND2_X1 U955 ( .A1(n995), .A2(n996), .ZN(n991) );
  OR2_X1 U956 ( .A1(n994), .A2(n993), .ZN(n996) );
  OR2_X1 U957 ( .A1(n827), .A2(n650), .ZN(n963) );
  OR2_X1 U958 ( .A1(n997), .A2(n678), .ZN(n673) );
  OR2_X1 U959 ( .A1(n669), .A2(n668), .ZN(n678) );
  OR2_X1 U960 ( .A1(n998), .A2(n999), .ZN(n668) );
  AND2_X1 U961 ( .A1(n664), .A2(n663), .ZN(n999) );
  AND2_X1 U962 ( .A1(n661), .A2(n1000), .ZN(n998) );
  OR2_X1 U963 ( .A1(n663), .A2(n664), .ZN(n1000) );
  OR2_X1 U964 ( .A1(n901), .A2(n922), .ZN(n664) );
  OR2_X1 U965 ( .A1(n1001), .A2(n1002), .ZN(n663) );
  AND2_X1 U966 ( .A1(n625), .A2(n624), .ZN(n1002) );
  AND2_X1 U967 ( .A1(n622), .A2(n1003), .ZN(n1001) );
  OR2_X1 U968 ( .A1(n624), .A2(n625), .ZN(n1003) );
  OR2_X1 U969 ( .A1(n901), .A2(n650), .ZN(n625) );
  OR2_X1 U970 ( .A1(n1004), .A2(n1005), .ZN(n624) );
  AND2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n1005) );
  AND2_X1 U972 ( .A1(n874), .A2(n1006), .ZN(n1004) );
  OR2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n1006) );
  OR2_X1 U974 ( .A1(n1007), .A2(n1008), .ZN(n876) );
  AND2_X1 U975 ( .A1(n832), .A2(n831), .ZN(n1008) );
  AND2_X1 U976 ( .A1(n829), .A2(n1009), .ZN(n1007) );
  OR2_X1 U977 ( .A1(n832), .A2(n831), .ZN(n1009) );
  OR2_X1 U978 ( .A1(n1010), .A2(n1011), .ZN(n831) );
  AND2_X1 U979 ( .A1(n804), .A2(n803), .ZN(n1011) );
  AND2_X1 U980 ( .A1(n801), .A2(n1012), .ZN(n1010) );
  OR2_X1 U981 ( .A1(n804), .A2(n803), .ZN(n1012) );
  OR2_X1 U982 ( .A1(n1013), .A2(n1014), .ZN(n803) );
  AND2_X1 U983 ( .A1(n776), .A2(n775), .ZN(n1014) );
  AND2_X1 U984 ( .A1(n773), .A2(n1015), .ZN(n1013) );
  OR2_X1 U985 ( .A1(n776), .A2(n775), .ZN(n1015) );
  OR2_X1 U986 ( .A1(n863), .A2(n901), .ZN(n775) );
  OR2_X1 U987 ( .A1(n866), .A2(n730), .ZN(n776) );
  OR2_X1 U988 ( .A1(n921), .A2(n901), .ZN(n730) );
  XNOR2_X1 U989 ( .A(n1016), .B(n866), .ZN(n773) );
  OR2_X1 U990 ( .A1(n868), .A2(n869), .ZN(n866) );
  OR2_X1 U991 ( .A1(n859), .A2(n901), .ZN(n804) );
  XNOR2_X1 U992 ( .A(n1017), .B(n1018), .ZN(n801) );
  XNOR2_X1 U993 ( .A(n1019), .B(n1020), .ZN(n1017) );
  OR2_X1 U994 ( .A1(n855), .A2(n901), .ZN(n832) );
  XOR2_X1 U995 ( .A(n1021), .B(n1022), .Z(n829) );
  XOR2_X1 U996 ( .A(n1023), .B(n1024), .Z(n1022) );
  OR2_X1 U997 ( .A1(n654), .A2(n901), .ZN(n877) );
  INV_X1 U998 ( .A(b_7_), .ZN(n901) );
  XOR2_X1 U999 ( .A(n1025), .B(n1026), .Z(n874) );
  XOR2_X1 U1000 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR2_X1 U1001 ( .A(n1029), .B(n1030), .Z(n622) );
  XOR2_X1 U1002 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR2_X1 U1003 ( .A(n1033), .B(n1034), .Z(n661) );
  XOR2_X1 U1004 ( .A(n1035), .B(n1036), .Z(n1034) );
  XOR2_X1 U1005 ( .A(n1037), .B(n1038), .Z(n669) );
  XOR2_X1 U1006 ( .A(n1039), .B(n1040), .Z(n1038) );
  OR2_X1 U1007 ( .A1(n1041), .A2(n1042), .ZN(n997) );
  AND2_X1 U1008 ( .A1(n676), .A2(n677), .ZN(n1042) );
  INV_X1 U1009 ( .A(n683), .ZN(n1041) );
  OR2_X1 U1010 ( .A1(n676), .A2(n677), .ZN(n683) );
  OR2_X1 U1011 ( .A1(n1043), .A2(n1044), .ZN(n677) );
  AND2_X1 U1012 ( .A1(n1040), .A2(n1039), .ZN(n1044) );
  AND2_X1 U1013 ( .A1(n1037), .A2(n1045), .ZN(n1043) );
  OR2_X1 U1014 ( .A1(n1039), .A2(n1040), .ZN(n1045) );
  OR2_X1 U1015 ( .A1(n869), .A2(n922), .ZN(n1040) );
  OR2_X1 U1016 ( .A1(n1046), .A2(n1047), .ZN(n1039) );
  AND2_X1 U1017 ( .A1(n1036), .A2(n1035), .ZN(n1047) );
  AND2_X1 U1018 ( .A1(n1033), .A2(n1048), .ZN(n1046) );
  OR2_X1 U1019 ( .A1(n1035), .A2(n1036), .ZN(n1048) );
  OR2_X1 U1020 ( .A1(n869), .A2(n650), .ZN(n1036) );
  OR2_X1 U1021 ( .A1(n1049), .A2(n1050), .ZN(n1035) );
  AND2_X1 U1022 ( .A1(n1032), .A2(n1031), .ZN(n1050) );
  AND2_X1 U1023 ( .A1(n1029), .A2(n1051), .ZN(n1049) );
  OR2_X1 U1024 ( .A1(n1031), .A2(n1032), .ZN(n1051) );
  OR2_X1 U1025 ( .A1(n869), .A2(n654), .ZN(n1032) );
  OR2_X1 U1026 ( .A1(n1052), .A2(n1053), .ZN(n1031) );
  AND2_X1 U1027 ( .A1(n1028), .A2(n1027), .ZN(n1053) );
  AND2_X1 U1028 ( .A1(n1025), .A2(n1054), .ZN(n1052) );
  OR2_X1 U1029 ( .A1(n1028), .A2(n1027), .ZN(n1054) );
  OR2_X1 U1030 ( .A1(n1055), .A2(n1056), .ZN(n1027) );
  AND2_X1 U1031 ( .A1(n1024), .A2(n1023), .ZN(n1056) );
  AND2_X1 U1032 ( .A1(n1021), .A2(n1057), .ZN(n1055) );
  OR2_X1 U1033 ( .A1(n1024), .A2(n1023), .ZN(n1057) );
  OR2_X1 U1034 ( .A1(n1058), .A2(n1059), .ZN(n1023) );
  AND2_X1 U1035 ( .A1(n1019), .A2(n1020), .ZN(n1059) );
  AND2_X1 U1036 ( .A1(n1018), .A2(n1060), .ZN(n1058) );
  OR2_X1 U1037 ( .A1(n1019), .A2(n1020), .ZN(n1060) );
  OR2_X1 U1038 ( .A1(n869), .A2(n1061), .ZN(n1020) );
  OR2_X1 U1039 ( .A1(n921), .A2(n1062), .ZN(n1061) );
  OR2_X1 U1040 ( .A1(n863), .A2(n869), .ZN(n1019) );
  XNOR2_X1 U1041 ( .A(n1063), .B(n1062), .ZN(n1018) );
  OR2_X1 U1042 ( .A1(n868), .A2(n771), .ZN(n1062) );
  OR2_X1 U1043 ( .A1(n921), .A2(n799), .ZN(n1063) );
  OR2_X1 U1044 ( .A1(n859), .A2(n869), .ZN(n1024) );
  XNOR2_X1 U1045 ( .A(n1064), .B(n1065), .ZN(n1021) );
  XNOR2_X1 U1046 ( .A(n1066), .B(n864), .ZN(n1064) );
  OR2_X1 U1047 ( .A1(n855), .A2(n869), .ZN(n1028) );
  INV_X1 U1048 ( .A(b_6_), .ZN(n869) );
  XOR2_X1 U1049 ( .A(n1067), .B(n1068), .Z(n1025) );
  XOR2_X1 U1050 ( .A(n1069), .B(n1070), .Z(n1068) );
  XOR2_X1 U1051 ( .A(n1071), .B(n1072), .Z(n1029) );
  XOR2_X1 U1052 ( .A(n1073), .B(n1074), .Z(n1072) );
  XOR2_X1 U1053 ( .A(n1075), .B(n1076), .Z(n1033) );
  XOR2_X1 U1054 ( .A(n1077), .B(n1078), .Z(n1076) );
  XOR2_X1 U1055 ( .A(n1079), .B(n1080), .Z(n1037) );
  XOR2_X1 U1056 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR2_X1 U1057 ( .A(n976), .B(n1083), .Z(n676) );
  XOR2_X1 U1058 ( .A(n979), .B(n977), .Z(n1083) );
  OR2_X1 U1059 ( .A1(n771), .A2(n922), .ZN(n977) );
  OR2_X1 U1060 ( .A1(n1084), .A2(n1085), .ZN(n979) );
  AND2_X1 U1061 ( .A1(n1082), .A2(n1081), .ZN(n1085) );
  AND2_X1 U1062 ( .A1(n1079), .A2(n1086), .ZN(n1084) );
  OR2_X1 U1063 ( .A1(n1081), .A2(n1082), .ZN(n1086) );
  OR2_X1 U1064 ( .A1(n771), .A2(n650), .ZN(n1082) );
  OR2_X1 U1065 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
  AND2_X1 U1066 ( .A1(n1078), .A2(n1077), .ZN(n1088) );
  AND2_X1 U1067 ( .A1(n1075), .A2(n1089), .ZN(n1087) );
  OR2_X1 U1068 ( .A1(n1077), .A2(n1078), .ZN(n1089) );
  OR2_X1 U1069 ( .A1(n771), .A2(n654), .ZN(n1078) );
  OR2_X1 U1070 ( .A1(n1090), .A2(n1091), .ZN(n1077) );
  AND2_X1 U1071 ( .A1(n1074), .A2(n1073), .ZN(n1091) );
  AND2_X1 U1072 ( .A1(n1071), .A2(n1092), .ZN(n1090) );
  OR2_X1 U1073 ( .A1(n1073), .A2(n1074), .ZN(n1092) );
  OR2_X1 U1074 ( .A1(n771), .A2(n855), .ZN(n1074) );
  OR2_X1 U1075 ( .A1(n1093), .A2(n1094), .ZN(n1073) );
  AND2_X1 U1076 ( .A1(n1070), .A2(n1069), .ZN(n1094) );
  AND2_X1 U1077 ( .A1(n1067), .A2(n1095), .ZN(n1093) );
  OR2_X1 U1078 ( .A1(n1070), .A2(n1069), .ZN(n1095) );
  OR2_X1 U1079 ( .A1(n1096), .A2(n1097), .ZN(n1069) );
  AND2_X1 U1080 ( .A1(n1065), .A2(n864), .ZN(n1097) );
  AND2_X1 U1081 ( .A1(n1098), .A2(n1066), .ZN(n1096) );
  OR2_X1 U1082 ( .A1(n1099), .A2(n1100), .ZN(n1066) );
  AND2_X1 U1083 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
  OR2_X1 U1084 ( .A1(n1065), .A2(n864), .ZN(n1098) );
  OR2_X1 U1085 ( .A1(n863), .A2(n771), .ZN(n864) );
  OR2_X1 U1086 ( .A1(n1102), .A2(n1016), .ZN(n1065) );
  OR2_X1 U1087 ( .A1(n921), .A2(n771), .ZN(n1016) );
  OR2_X1 U1088 ( .A1(n859), .A2(n771), .ZN(n1070) );
  INV_X1 U1089 ( .A(b_5_), .ZN(n771) );
  XNOR2_X1 U1090 ( .A(n1103), .B(n1104), .ZN(n1067) );
  XOR2_X1 U1091 ( .A(n1105), .B(n1100), .Z(n1103) );
  INV_X1 U1092 ( .A(n1106), .ZN(n1100) );
  XNOR2_X1 U1093 ( .A(n1107), .B(n1108), .ZN(n1071) );
  XNOR2_X1 U1094 ( .A(n860), .B(n1109), .ZN(n1107) );
  XOR2_X1 U1095 ( .A(n1110), .B(n1111), .Z(n1075) );
  XOR2_X1 U1096 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR2_X1 U1097 ( .A(n1114), .B(n1115), .Z(n1079) );
  XOR2_X1 U1098 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR2_X1 U1099 ( .A(n983), .B(n1118), .Z(n976) );
  XOR2_X1 U1100 ( .A(n986), .B(n984), .Z(n1118) );
  OR2_X1 U1101 ( .A1(n799), .A2(n650), .ZN(n984) );
  OR2_X1 U1102 ( .A1(n1119), .A2(n1120), .ZN(n986) );
  AND2_X1 U1103 ( .A1(n1117), .A2(n1116), .ZN(n1120) );
  AND2_X1 U1104 ( .A1(n1114), .A2(n1121), .ZN(n1119) );
  OR2_X1 U1105 ( .A1(n1116), .A2(n1117), .ZN(n1121) );
  OR2_X1 U1106 ( .A1(n799), .A2(n654), .ZN(n1117) );
  OR2_X1 U1107 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
  AND2_X1 U1108 ( .A1(n1113), .A2(n1112), .ZN(n1123) );
  AND2_X1 U1109 ( .A1(n1110), .A2(n1124), .ZN(n1122) );
  OR2_X1 U1110 ( .A1(n1112), .A2(n1113), .ZN(n1124) );
  OR2_X1 U1111 ( .A1(n799), .A2(n855), .ZN(n1113) );
  OR2_X1 U1112 ( .A1(n1125), .A2(n1126), .ZN(n1112) );
  AND2_X1 U1113 ( .A1(n1109), .A2(n860), .ZN(n1126) );
  AND2_X1 U1114 ( .A1(n1108), .A2(n1127), .ZN(n1125) );
  OR2_X1 U1115 ( .A1(n860), .A2(n1109), .ZN(n1127) );
  OR2_X1 U1116 ( .A1(n1128), .A2(n1129), .ZN(n1109) );
  AND2_X1 U1117 ( .A1(n1104), .A2(n1106), .ZN(n1129) );
  AND2_X1 U1118 ( .A1(n1130), .A2(n1105), .ZN(n1128) );
  OR2_X1 U1119 ( .A1(n1131), .A2(n1132), .ZN(n1105) );
  INV_X1 U1120 ( .A(n1133), .ZN(n1132) );
  AND2_X1 U1121 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
  OR2_X1 U1122 ( .A1(n1104), .A2(n1106), .ZN(n1130) );
  OR2_X1 U1123 ( .A1(n1101), .A2(n1102), .ZN(n1106) );
  OR2_X1 U1124 ( .A1(n868), .A2(n799), .ZN(n1102) );
  OR2_X1 U1125 ( .A1(n921), .A2(n827), .ZN(n1101) );
  OR2_X1 U1126 ( .A1(n863), .A2(n799), .ZN(n1104) );
  OR2_X1 U1127 ( .A1(n859), .A2(n799), .ZN(n860) );
  INV_X1 U1128 ( .A(b_4_), .ZN(n799) );
  XNOR2_X1 U1129 ( .A(n1136), .B(n1133), .ZN(n1108) );
  XNOR2_X1 U1130 ( .A(n1137), .B(n1138), .ZN(n1136) );
  XNOR2_X1 U1131 ( .A(n1139), .B(n1140), .ZN(n1110) );
  XNOR2_X1 U1132 ( .A(n1141), .B(n1142), .ZN(n1139) );
  XNOR2_X1 U1133 ( .A(n1143), .B(n1144), .ZN(n1114) );
  XNOR2_X1 U1134 ( .A(n856), .B(n1145), .ZN(n1143) );
  XNOR2_X1 U1135 ( .A(n1146), .B(n995), .ZN(n983) );
  XNOR2_X1 U1136 ( .A(n1147), .B(n1148), .ZN(n995) );
  XNOR2_X1 U1137 ( .A(n1149), .B(n1150), .ZN(n1147) );
  XNOR2_X1 U1138 ( .A(n994), .B(n993), .ZN(n1146) );
  OR2_X1 U1139 ( .A1(n1151), .A2(n1152), .ZN(n993) );
  AND2_X1 U1140 ( .A1(n1145), .A2(n856), .ZN(n1152) );
  AND2_X1 U1141 ( .A1(n1144), .A2(n1153), .ZN(n1151) );
  OR2_X1 U1142 ( .A1(n856), .A2(n1145), .ZN(n1153) );
  OR2_X1 U1143 ( .A1(n1154), .A2(n1155), .ZN(n1145) );
  AND2_X1 U1144 ( .A1(n1142), .A2(n1141), .ZN(n1155) );
  AND2_X1 U1145 ( .A1(n1140), .A2(n1156), .ZN(n1154) );
  OR2_X1 U1146 ( .A1(n1141), .A2(n1142), .ZN(n1156) );
  OR2_X1 U1147 ( .A1(n1157), .A2(n1158), .ZN(n1142) );
  AND2_X1 U1148 ( .A1(n1133), .A2(n1138), .ZN(n1158) );
  AND2_X1 U1149 ( .A1(n1159), .A2(n1137), .ZN(n1157) );
  OR2_X1 U1150 ( .A1(n1160), .A2(n1161), .ZN(n1137) );
  AND2_X1 U1151 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
  OR2_X1 U1152 ( .A1(n1138), .A2(n1133), .ZN(n1159) );
  OR2_X1 U1153 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
  OR2_X1 U1154 ( .A1(n921), .A2(n655), .ZN(n1135) );
  OR2_X1 U1155 ( .A1(n868), .A2(n827), .ZN(n1134) );
  OR2_X1 U1156 ( .A1(n827), .A2(n863), .ZN(n1138) );
  OR2_X1 U1157 ( .A1(n827), .A2(n859), .ZN(n1141) );
  XNOR2_X1 U1158 ( .A(n1164), .B(n1165), .ZN(n1140) );
  XOR2_X1 U1159 ( .A(n1166), .B(n1161), .Z(n1164) );
  INV_X1 U1160 ( .A(n1167), .ZN(n1161) );
  OR2_X1 U1161 ( .A1(n827), .A2(n855), .ZN(n856) );
  XOR2_X1 U1162 ( .A(n1168), .B(n1169), .Z(n1144) );
  XOR2_X1 U1163 ( .A(n1170), .B(n1171), .Z(n1169) );
  OR2_X1 U1164 ( .A1(n827), .A2(n654), .ZN(n994) );
  INV_X1 U1165 ( .A(b_3_), .ZN(n827) );
  AND2_X1 U1166 ( .A1(n709), .A2(n1172), .ZN(n711) );
  AND2_X1 U1167 ( .A1(n710), .A2(n708), .ZN(n1172) );
  XNOR2_X1 U1168 ( .A(n1173), .B(n1174), .ZN(n708) );
  OR2_X1 U1169 ( .A1(n904), .A2(n922), .ZN(n1173) );
  XNOR2_X1 U1170 ( .A(n1175), .B(n1176), .ZN(n710) );
  XOR2_X1 U1171 ( .A(n1177), .B(n1178), .Z(n1176) );
  INV_X1 U1172 ( .A(n1179), .ZN(n709) );
  OR2_X1 U1173 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
  AND2_X1 U1174 ( .A1(n946), .A2(n945), .ZN(n1181) );
  AND2_X1 U1175 ( .A1(n943), .A2(n1182), .ZN(n1180) );
  OR2_X1 U1176 ( .A1(n945), .A2(n946), .ZN(n1182) );
  OR2_X1 U1177 ( .A1(n655), .A2(n922), .ZN(n946) );
  OR2_X1 U1178 ( .A1(n1183), .A2(n1184), .ZN(n945) );
  AND2_X1 U1179 ( .A1(n959), .A2(n958), .ZN(n1184) );
  AND2_X1 U1180 ( .A1(n956), .A2(n1185), .ZN(n1183) );
  OR2_X1 U1181 ( .A1(n958), .A2(n959), .ZN(n1185) );
  OR2_X1 U1182 ( .A1(n655), .A2(n650), .ZN(n959) );
  OR2_X1 U1183 ( .A1(n1186), .A2(n1187), .ZN(n958) );
  AND2_X1 U1184 ( .A1(n990), .A2(n657), .ZN(n1187) );
  AND2_X1 U1185 ( .A1(n989), .A2(n1188), .ZN(n1186) );
  OR2_X1 U1186 ( .A1(n657), .A2(n990), .ZN(n1188) );
  OR2_X1 U1187 ( .A1(n1189), .A2(n1190), .ZN(n990) );
  AND2_X1 U1188 ( .A1(n1150), .A2(n1149), .ZN(n1190) );
  AND2_X1 U1189 ( .A1(n1148), .A2(n1191), .ZN(n1189) );
  OR2_X1 U1190 ( .A1(n1149), .A2(n1150), .ZN(n1191) );
  OR2_X1 U1191 ( .A1(n1192), .A2(n1193), .ZN(n1150) );
  AND2_X1 U1192 ( .A1(n1171), .A2(n1170), .ZN(n1193) );
  AND2_X1 U1193 ( .A1(n1168), .A2(n1194), .ZN(n1192) );
  OR2_X1 U1194 ( .A1(n1170), .A2(n1171), .ZN(n1194) );
  OR2_X1 U1195 ( .A1(n655), .A2(n859), .ZN(n1171) );
  OR2_X1 U1196 ( .A1(n1195), .A2(n1196), .ZN(n1170) );
  AND2_X1 U1197 ( .A1(n1165), .A2(n1167), .ZN(n1196) );
  AND2_X1 U1198 ( .A1(n1197), .A2(n1166), .ZN(n1195) );
  OR2_X1 U1199 ( .A1(n1198), .A2(n1199), .ZN(n1166) );
  AND2_X1 U1200 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
  OR2_X1 U1201 ( .A1(n1167), .A2(n1165), .ZN(n1197) );
  OR2_X1 U1202 ( .A1(n655), .A2(n863), .ZN(n1165) );
  OR2_X1 U1203 ( .A1(n1162), .A2(n1163), .ZN(n1167) );
  OR2_X1 U1204 ( .A1(n655), .A2(n868), .ZN(n1163) );
  OR2_X1 U1205 ( .A1(n921), .A2(n651), .ZN(n1162) );
  XOR2_X1 U1206 ( .A(n1202), .B(n1199), .Z(n1168) );
  INV_X1 U1207 ( .A(n1203), .ZN(n1199) );
  OR2_X1 U1208 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
  INV_X1 U1209 ( .A(n1206), .ZN(n1205) );
  AND2_X1 U1210 ( .A1(n1207), .A2(n1208), .ZN(n1204) );
  OR2_X1 U1211 ( .A1(n655), .A2(n855), .ZN(n1149) );
  XOR2_X1 U1212 ( .A(n1209), .B(n1210), .Z(n1148) );
  XOR2_X1 U1213 ( .A(n1211), .B(n1212), .Z(n1209) );
  OR2_X1 U1214 ( .A1(n655), .A2(n654), .ZN(n657) );
  INV_X1 U1215 ( .A(b_2_), .ZN(n655) );
  XOR2_X1 U1216 ( .A(n1213), .B(n1214), .Z(n989) );
  XOR2_X1 U1217 ( .A(n1215), .B(n1216), .Z(n1214) );
  XOR2_X1 U1218 ( .A(n1217), .B(n1218), .Z(n956) );
  XOR2_X1 U1219 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR2_X1 U1220 ( .A(n1221), .B(n1222), .ZN(n943) );
  XNOR2_X1 U1221 ( .A(n614), .B(n1223), .ZN(n1221) );
  AND2_X1 U1222 ( .A1(n1174), .A2(a_0_), .ZN(n924) );
  INV_X1 U1223 ( .A(n1224), .ZN(n1174) );
  OR2_X1 U1224 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
  AND2_X1 U1225 ( .A1(n1175), .A2(n1177), .ZN(n1226) );
  AND2_X1 U1226 ( .A1(n1227), .A2(n1178), .ZN(n1225) );
  OR2_X1 U1227 ( .A1(n651), .A2(n922), .ZN(n1178) );
  INV_X1 U1228 ( .A(a_0_), .ZN(n922) );
  OR2_X1 U1229 ( .A1(n1177), .A2(n1175), .ZN(n1227) );
  OR2_X1 U1230 ( .A1(n650), .A2(n904), .ZN(n1175) );
  OR2_X1 U1231 ( .A1(n1228), .A2(n1229), .ZN(n1177) );
  AND2_X1 U1232 ( .A1(n1222), .A2(n1223), .ZN(n1229) );
  AND2_X1 U1233 ( .A1(n1230), .A2(n614), .ZN(n1228) );
  OR2_X1 U1234 ( .A1(n651), .A2(n650), .ZN(n614) );
  INV_X1 U1235 ( .A(a_1_), .ZN(n650) );
  OR2_X1 U1236 ( .A1(n1223), .A2(n1222), .ZN(n1230) );
  OR2_X1 U1237 ( .A1(n654), .A2(n904), .ZN(n1222) );
  OR2_X1 U1238 ( .A1(n1231), .A2(n1232), .ZN(n1223) );
  AND2_X1 U1239 ( .A1(n1217), .A2(n1219), .ZN(n1232) );
  AND2_X1 U1240 ( .A1(n1233), .A2(n1220), .ZN(n1231) );
  OR2_X1 U1241 ( .A1(n855), .A2(n904), .ZN(n1220) );
  OR2_X1 U1242 ( .A1(n1219), .A2(n1217), .ZN(n1233) );
  OR2_X1 U1243 ( .A1(n651), .A2(n654), .ZN(n1217) );
  INV_X1 U1244 ( .A(a_2_), .ZN(n654) );
  OR2_X1 U1245 ( .A1(n1234), .A2(n1235), .ZN(n1219) );
  AND2_X1 U1246 ( .A1(n1213), .A2(n1215), .ZN(n1235) );
  AND2_X1 U1247 ( .A1(n1236), .A2(n1216), .ZN(n1234) );
  OR2_X1 U1248 ( .A1(n651), .A2(n855), .ZN(n1216) );
  INV_X1 U1249 ( .A(a_3_), .ZN(n855) );
  OR2_X1 U1250 ( .A1(n1215), .A2(n1213), .ZN(n1236) );
  OR2_X1 U1251 ( .A1(n859), .A2(n904), .ZN(n1213) );
  OR2_X1 U1252 ( .A1(n1237), .A2(n1238), .ZN(n1215) );
  AND2_X1 U1253 ( .A1(n1210), .A2(n1212), .ZN(n1238) );
  AND2_X1 U1254 ( .A1(n1211), .A2(n1239), .ZN(n1237) );
  OR2_X1 U1255 ( .A1(n1212), .A2(n1210), .ZN(n1239) );
  OR2_X1 U1256 ( .A1(n863), .A2(n904), .ZN(n1210) );
  OR2_X1 U1257 ( .A1(n651), .A2(n859), .ZN(n1212) );
  INV_X1 U1258 ( .A(a_4_), .ZN(n859) );
  AND2_X1 U1259 ( .A1(n1206), .A2(n1203), .ZN(n1211) );
  OR2_X1 U1260 ( .A1(n1201), .A2(n1200), .ZN(n1203) );
  OR2_X1 U1261 ( .A1(n921), .A2(n904), .ZN(n1200) );
  INV_X1 U1262 ( .A(a_7_), .ZN(n921) );
  OR2_X1 U1263 ( .A1(n868), .A2(n651), .ZN(n1201) );
  OR2_X1 U1264 ( .A1(n1208), .A2(n1207), .ZN(n1206) );
  OR2_X1 U1265 ( .A1(n868), .A2(n904), .ZN(n1207) );
  INV_X1 U1266 ( .A(b_0_), .ZN(n904) );
  INV_X1 U1267 ( .A(a_6_), .ZN(n868) );
  OR2_X1 U1268 ( .A1(n651), .A2(n863), .ZN(n1208) );
  INV_X1 U1269 ( .A(a_5_), .ZN(n863) );
  INV_X1 U1270 ( .A(b_1_), .ZN(n651) );
  AND2_X1 U1271 ( .A1(operation_0_), .A2(operation_1_), .ZN(n620) );
endmodule

