module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n172_, keyIn_0_45 );
not g001 ( new_n173_, N11 );
and g002 ( new_n174_, new_n173_, keyIn_0_2 );
not g003 ( new_n175_, N17 );
not g004 ( new_n176_, keyIn_0_2 );
and g005 ( new_n177_, new_n176_, N11 );
or g006 ( new_n178_, new_n177_, new_n175_ );
or g007 ( new_n179_, new_n178_, new_n174_ );
not g008 ( new_n180_, new_n179_ );
and g009 ( new_n181_, new_n180_, keyIn_0_21 );
not g010 ( new_n182_, keyIn_0_21 );
and g011 ( new_n183_, new_n179_, new_n182_ );
or g012 ( new_n184_, new_n181_, new_n183_ );
or g013 ( new_n185_, keyIn_0_14, N89 );
not g014 ( new_n186_, N95 );
and g015 ( new_n187_, keyIn_0_14, N89 );
or g016 ( new_n188_, new_n187_, new_n186_ );
not g017 ( new_n189_, new_n188_ );
and g018 ( new_n190_, new_n189_, new_n185_ );
not g019 ( new_n191_, new_n190_ );
or g020 ( new_n192_, new_n191_, keyIn_0_27 );
not g021 ( new_n193_, keyIn_0_27 );
or g022 ( new_n194_, new_n190_, new_n193_ );
and g023 ( new_n195_, new_n192_, new_n194_ );
not g024 ( new_n196_, N1 );
and g025 ( new_n197_, new_n196_, keyIn_0_0 );
not g026 ( new_n198_, new_n197_ );
or g027 ( new_n199_, new_n196_, keyIn_0_0 );
and g028 ( new_n200_, new_n199_, N4 );
and g029 ( new_n201_, new_n200_, new_n198_ );
not g030 ( new_n202_, new_n201_ );
and g031 ( new_n203_, new_n202_, keyIn_0_18 );
not g032 ( new_n204_, keyIn_0_18 );
and g033 ( new_n205_, new_n201_, new_n204_ );
or g034 ( new_n206_, new_n203_, new_n205_ );
and g035 ( new_n207_, new_n195_, new_n206_ );
and g036 ( new_n208_, new_n207_, new_n184_ );
not g037 ( new_n209_, keyIn_0_28 );
not g038 ( new_n210_, N102 );
and g039 ( new_n211_, new_n210_, keyIn_0_16 );
not g040 ( new_n212_, new_n211_ );
or g041 ( new_n213_, new_n210_, keyIn_0_16 );
and g042 ( new_n214_, new_n213_, N108 );
and g043 ( new_n215_, new_n214_, new_n212_ );
not g044 ( new_n216_, new_n215_ );
and g045 ( new_n217_, new_n216_, new_n209_ );
and g046 ( new_n218_, new_n215_, keyIn_0_28 );
or g047 ( new_n219_, new_n217_, new_n218_ );
not g048 ( new_n220_, keyIn_0_26 );
not g049 ( new_n221_, N76 );
and g050 ( new_n222_, new_n221_, keyIn_0_12 );
not g051 ( new_n223_, new_n222_ );
or g052 ( new_n224_, new_n221_, keyIn_0_12 );
and g053 ( new_n225_, new_n224_, N82 );
and g054 ( new_n226_, new_n225_, new_n223_ );
not g055 ( new_n227_, new_n226_ );
or g056 ( new_n228_, new_n227_, new_n220_ );
or g057 ( new_n229_, new_n226_, keyIn_0_26 );
and g058 ( new_n230_, new_n228_, new_n229_ );
and g059 ( new_n231_, new_n219_, new_n230_ );
not g060 ( new_n232_, N50 );
and g061 ( new_n233_, new_n232_, keyIn_0_8 );
not g062 ( new_n234_, N56 );
not g063 ( new_n235_, keyIn_0_8 );
and g064 ( new_n236_, new_n235_, N50 );
or g065 ( new_n237_, new_n236_, new_n234_ );
or g066 ( new_n238_, new_n237_, new_n233_ );
and g067 ( new_n239_, new_n238_, keyIn_0_24 );
not g068 ( new_n240_, keyIn_0_24 );
not g069 ( new_n241_, new_n233_ );
or g070 ( new_n242_, new_n232_, keyIn_0_8 );
and g071 ( new_n243_, new_n242_, N56 );
and g072 ( new_n244_, new_n243_, new_n241_ );
and g073 ( new_n245_, new_n244_, new_n240_ );
or g074 ( new_n246_, new_n239_, new_n245_ );
not g075 ( new_n247_, keyIn_0_25 );
not g076 ( new_n248_, N63 );
and g077 ( new_n249_, new_n248_, keyIn_0_10 );
not g078 ( new_n250_, N69 );
not g079 ( new_n251_, keyIn_0_10 );
and g080 ( new_n252_, new_n251_, N63 );
or g081 ( new_n253_, new_n252_, new_n250_ );
or g082 ( new_n254_, new_n253_, new_n249_ );
or g083 ( new_n255_, new_n254_, new_n247_ );
not g084 ( new_n256_, new_n249_ );
or g085 ( new_n257_, new_n248_, keyIn_0_10 );
and g086 ( new_n258_, new_n257_, N69 );
and g087 ( new_n259_, new_n258_, new_n256_ );
or g088 ( new_n260_, new_n259_, keyIn_0_25 );
and g089 ( new_n261_, new_n255_, new_n260_ );
and g090 ( new_n262_, new_n246_, new_n261_ );
not g091 ( new_n263_, keyIn_0_23 );
and g092 ( new_n264_, keyIn_0_6, N37 );
not g093 ( new_n265_, keyIn_0_6 );
not g094 ( new_n266_, N37 );
and g095 ( new_n267_, new_n265_, new_n266_ );
or g096 ( new_n268_, new_n267_, new_n264_ );
and g097 ( new_n269_, new_n268_, N43 );
and g098 ( new_n270_, new_n269_, new_n263_ );
not g099 ( new_n271_, N43 );
not g100 ( new_n272_, new_n264_ );
or g101 ( new_n273_, keyIn_0_6, N37 );
and g102 ( new_n274_, new_n272_, new_n273_ );
or g103 ( new_n275_, new_n274_, new_n271_ );
and g104 ( new_n276_, new_n275_, keyIn_0_23 );
or g105 ( new_n277_, new_n270_, new_n276_ );
not g106 ( new_n278_, keyIn_0_22 );
not g107 ( new_n279_, N24 );
and g108 ( new_n280_, new_n279_, keyIn_0_4 );
not g109 ( new_n281_, N30 );
not g110 ( new_n282_, keyIn_0_4 );
and g111 ( new_n283_, new_n282_, N24 );
or g112 ( new_n284_, new_n283_, new_n281_ );
or g113 ( new_n285_, new_n284_, new_n280_ );
and g114 ( new_n286_, new_n285_, new_n278_ );
not g115 ( new_n287_, new_n280_ );
or g116 ( new_n288_, new_n279_, keyIn_0_4 );
and g117 ( new_n289_, new_n288_, N30 );
and g118 ( new_n290_, new_n289_, new_n287_ );
and g119 ( new_n291_, new_n290_, keyIn_0_22 );
or g120 ( new_n292_, new_n286_, new_n291_ );
and g121 ( new_n293_, new_n277_, new_n292_ );
and g122 ( new_n294_, new_n293_, new_n262_ );
and g123 ( new_n295_, new_n294_, new_n231_ );
and g124 ( new_n296_, new_n295_, new_n208_ );
and g125 ( new_n297_, new_n296_, new_n172_ );
not g126 ( new_n298_, new_n297_ );
or g127 ( new_n299_, new_n296_, new_n172_ );
and g128 ( N223, new_n298_, new_n299_ );
not g129 ( new_n301_, keyIn_0_76 );
not g130 ( new_n302_, keyIn_0_60 );
not g131 ( new_n303_, keyIn_0_49 );
not g132 ( new_n304_, keyIn_0_46 );
or g133 ( new_n305_, N223, new_n304_ );
not g134 ( new_n306_, new_n296_ );
and g135 ( new_n307_, new_n306_, keyIn_0_45 );
or g136 ( new_n308_, new_n307_, new_n297_ );
or g137 ( new_n309_, new_n308_, keyIn_0_46 );
and g138 ( new_n310_, new_n309_, new_n305_ );
and g139 ( new_n311_, new_n310_, new_n184_ );
not g140 ( new_n312_, new_n311_ );
or g141 ( new_n313_, new_n310_, new_n184_ );
and g142 ( new_n314_, new_n312_, new_n313_ );
not g143 ( new_n315_, new_n314_ );
and g144 ( new_n316_, new_n315_, new_n303_ );
and g145 ( new_n317_, new_n314_, keyIn_0_49 );
or g146 ( new_n318_, new_n316_, new_n317_ );
not g147 ( new_n319_, N21 );
and g148 ( new_n320_, keyIn_0_3, N17 );
not g149 ( new_n321_, new_n320_ );
or g150 ( new_n322_, keyIn_0_3, N17 );
and g151 ( new_n323_, new_n321_, new_n322_ );
not g152 ( new_n324_, new_n323_ );
and g153 ( new_n325_, new_n324_, new_n319_ );
not g154 ( new_n326_, new_n325_ );
and g155 ( new_n327_, new_n326_, keyIn_0_29 );
not g156 ( new_n328_, new_n327_ );
or g157 ( new_n329_, new_n326_, keyIn_0_29 );
and g158 ( new_n330_, new_n328_, new_n329_ );
or g159 ( new_n331_, new_n318_, new_n330_ );
not g160 ( new_n332_, new_n331_ );
or g161 ( new_n333_, new_n332_, new_n302_ );
or g162 ( new_n334_, new_n331_, keyIn_0_60 );
and g163 ( new_n335_, new_n333_, new_n334_ );
not g164 ( new_n336_, keyIn_0_54 );
not g165 ( new_n337_, new_n230_ );
and g166 ( new_n338_, new_n308_, keyIn_0_46 );
and g167 ( new_n339_, N223, new_n304_ );
or g168 ( new_n340_, new_n338_, new_n339_ );
and g169 ( new_n341_, new_n340_, new_n337_ );
and g170 ( new_n342_, new_n310_, new_n230_ );
or g171 ( new_n343_, new_n341_, new_n342_ );
and g172 ( new_n344_, new_n343_, new_n336_ );
not g173 ( new_n345_, new_n344_ );
or g174 ( new_n346_, new_n343_, new_n336_ );
and g175 ( new_n347_, new_n345_, new_n346_ );
not g176 ( new_n348_, N86 );
and g177 ( new_n349_, keyIn_0_13, N82 );
not g178 ( new_n350_, new_n349_ );
or g179 ( new_n351_, keyIn_0_13, N82 );
and g180 ( new_n352_, new_n350_, new_n351_ );
and g181 ( new_n353_, new_n352_, new_n348_ );
not g182 ( new_n354_, new_n353_ );
and g183 ( new_n355_, new_n354_, keyIn_0_39 );
not g184 ( new_n356_, new_n355_ );
or g185 ( new_n357_, new_n354_, keyIn_0_39 );
and g186 ( new_n358_, new_n356_, new_n357_ );
not g187 ( new_n359_, new_n358_ );
and g188 ( new_n360_, new_n347_, new_n359_ );
not g189 ( new_n361_, new_n360_ );
or g190 ( new_n362_, new_n361_, keyIn_0_65 );
not g191 ( new_n363_, keyIn_0_65 );
or g192 ( new_n364_, new_n360_, new_n363_ );
and g193 ( new_n365_, new_n362_, new_n364_ );
not g194 ( new_n366_, new_n206_ );
and g195 ( new_n367_, new_n340_, new_n366_ );
and g196 ( new_n368_, new_n310_, new_n206_ );
or g197 ( new_n369_, new_n367_, new_n368_ );
and g198 ( new_n370_, new_n369_, keyIn_0_48 );
not g199 ( new_n371_, new_n370_ );
or g200 ( new_n372_, new_n369_, keyIn_0_48 );
and g201 ( new_n373_, new_n371_, new_n372_ );
not g202 ( new_n374_, N8 );
and g203 ( new_n375_, keyIn_0_1, N4 );
not g204 ( new_n376_, new_n375_ );
or g205 ( new_n377_, keyIn_0_1, N4 );
and g206 ( new_n378_, new_n376_, new_n377_ );
and g207 ( new_n379_, new_n378_, new_n374_ );
not g208 ( new_n380_, new_n379_ );
and g209 ( new_n381_, new_n380_, keyIn_0_19 );
not g210 ( new_n382_, new_n381_ );
or g211 ( new_n383_, new_n380_, keyIn_0_19 );
and g212 ( new_n384_, new_n382_, new_n383_ );
not g213 ( new_n385_, new_n384_ );
and g214 ( new_n386_, new_n373_, new_n385_ );
not g215 ( new_n387_, new_n386_ );
and g216 ( new_n388_, new_n387_, keyIn_0_58 );
not g217 ( new_n389_, keyIn_0_58 );
and g218 ( new_n390_, new_n386_, new_n389_ );
or g219 ( new_n391_, new_n388_, new_n390_ );
and g220 ( new_n392_, new_n365_, new_n391_ );
and g221 ( new_n393_, new_n392_, new_n335_ );
not g222 ( new_n394_, new_n246_ );
and g223 ( new_n395_, new_n340_, new_n394_ );
and g224 ( new_n396_, new_n310_, new_n246_ );
or g225 ( new_n397_, new_n395_, new_n396_ );
and g226 ( new_n398_, new_n397_, keyIn_0_52 );
not g227 ( new_n399_, new_n398_ );
or g228 ( new_n400_, new_n397_, keyIn_0_52 );
and g229 ( new_n401_, new_n399_, new_n400_ );
not g230 ( new_n402_, N60 );
and g231 ( new_n403_, new_n234_, keyIn_0_9 );
not g232 ( new_n404_, new_n403_ );
or g233 ( new_n405_, new_n234_, keyIn_0_9 );
and g234 ( new_n406_, new_n404_, new_n405_ );
not g235 ( new_n407_, new_n406_ );
and g236 ( new_n408_, new_n407_, new_n402_ );
not g237 ( new_n409_, new_n408_ );
and g238 ( new_n410_, new_n409_, keyIn_0_35 );
not g239 ( new_n411_, new_n410_ );
or g240 ( new_n412_, new_n409_, keyIn_0_35 );
and g241 ( new_n413_, new_n411_, new_n412_ );
not g242 ( new_n414_, new_n413_ );
and g243 ( new_n415_, new_n401_, new_n414_ );
not g244 ( new_n416_, new_n415_ );
or g245 ( new_n417_, new_n416_, keyIn_0_63 );
not g246 ( new_n418_, keyIn_0_63 );
or g247 ( new_n419_, new_n415_, new_n418_ );
and g248 ( new_n420_, new_n417_, new_n419_ );
not g249 ( new_n421_, new_n261_ );
and g250 ( new_n422_, new_n340_, new_n421_ );
and g251 ( new_n423_, new_n310_, new_n261_ );
or g252 ( new_n424_, new_n422_, new_n423_ );
and g253 ( new_n425_, new_n424_, keyIn_0_53 );
not g254 ( new_n426_, new_n425_ );
or g255 ( new_n427_, new_n424_, keyIn_0_53 );
and g256 ( new_n428_, new_n426_, new_n427_ );
not g257 ( new_n429_, N73 );
and g258 ( new_n430_, keyIn_0_11, N69 );
not g259 ( new_n431_, new_n430_ );
or g260 ( new_n432_, keyIn_0_11, N69 );
and g261 ( new_n433_, new_n431_, new_n432_ );
and g262 ( new_n434_, new_n433_, new_n429_ );
not g263 ( new_n435_, new_n434_ );
and g264 ( new_n436_, new_n435_, keyIn_0_37 );
not g265 ( new_n437_, new_n436_ );
or g266 ( new_n438_, new_n435_, keyIn_0_37 );
and g267 ( new_n439_, new_n437_, new_n438_ );
not g268 ( new_n440_, new_n439_ );
and g269 ( new_n441_, new_n428_, new_n440_ );
not g270 ( new_n442_, new_n441_ );
or g271 ( new_n443_, new_n442_, keyIn_0_64 );
not g272 ( new_n444_, keyIn_0_64 );
or g273 ( new_n445_, new_n441_, new_n444_ );
and g274 ( new_n446_, new_n443_, new_n445_ );
and g275 ( new_n447_, new_n420_, new_n446_ );
not g276 ( new_n448_, keyIn_0_66 );
not g277 ( new_n449_, new_n195_ );
and g278 ( new_n450_, new_n340_, new_n449_ );
and g279 ( new_n451_, new_n310_, new_n195_ );
or g280 ( new_n452_, new_n450_, new_n451_ );
and g281 ( new_n453_, new_n452_, keyIn_0_55 );
not g282 ( new_n454_, keyIn_0_55 );
or g283 ( new_n455_, new_n310_, new_n195_ );
or g284 ( new_n456_, new_n340_, new_n449_ );
and g285 ( new_n457_, new_n456_, new_n455_ );
and g286 ( new_n458_, new_n457_, new_n454_ );
or g287 ( new_n459_, new_n453_, new_n458_ );
not g288 ( new_n460_, keyIn_0_41 );
not g289 ( new_n461_, N99 );
and g290 ( new_n462_, keyIn_0_15, N95 );
not g291 ( new_n463_, new_n462_ );
or g292 ( new_n464_, keyIn_0_15, N95 );
and g293 ( new_n465_, new_n463_, new_n464_ );
not g294 ( new_n466_, new_n465_ );
and g295 ( new_n467_, new_n466_, new_n461_ );
not g296 ( new_n468_, new_n467_ );
and g297 ( new_n469_, new_n468_, new_n460_ );
and g298 ( new_n470_, new_n467_, keyIn_0_41 );
or g299 ( new_n471_, new_n469_, new_n470_ );
or g300 ( new_n472_, new_n459_, new_n471_ );
or g301 ( new_n473_, new_n472_, new_n448_ );
or g302 ( new_n474_, new_n457_, new_n454_ );
or g303 ( new_n475_, new_n452_, keyIn_0_55 );
and g304 ( new_n476_, new_n475_, new_n474_ );
not g305 ( new_n477_, new_n471_ );
and g306 ( new_n478_, new_n476_, new_n477_ );
or g307 ( new_n479_, new_n478_, keyIn_0_66 );
and g308 ( new_n480_, new_n473_, new_n479_ );
not g309 ( new_n481_, keyIn_0_56 );
not g310 ( new_n482_, new_n219_ );
and g311 ( new_n483_, new_n340_, new_n482_ );
and g312 ( new_n484_, new_n310_, new_n219_ );
or g313 ( new_n485_, new_n483_, new_n484_ );
or g314 ( new_n486_, new_n485_, new_n481_ );
or g315 ( new_n487_, new_n310_, new_n219_ );
or g316 ( new_n488_, new_n340_, new_n482_ );
and g317 ( new_n489_, new_n488_, new_n487_ );
or g318 ( new_n490_, new_n489_, keyIn_0_56 );
and g319 ( new_n491_, new_n486_, new_n490_ );
not g320 ( new_n492_, keyIn_0_43 );
not g321 ( new_n493_, N112 );
and g322 ( new_n494_, keyIn_0_17, N108 );
not g323 ( new_n495_, new_n494_ );
or g324 ( new_n496_, keyIn_0_17, N108 );
and g325 ( new_n497_, new_n495_, new_n496_ );
not g326 ( new_n498_, new_n497_ );
and g327 ( new_n499_, new_n498_, new_n493_ );
not g328 ( new_n500_, new_n499_ );
and g329 ( new_n501_, new_n500_, new_n492_ );
and g330 ( new_n502_, new_n499_, keyIn_0_43 );
or g331 ( new_n503_, new_n501_, new_n502_ );
or g332 ( new_n504_, new_n491_, new_n503_ );
or g333 ( new_n505_, new_n504_, keyIn_0_67 );
not g334 ( new_n506_, keyIn_0_67 );
and g335 ( new_n507_, new_n489_, keyIn_0_56 );
and g336 ( new_n508_, new_n485_, new_n481_ );
or g337 ( new_n509_, new_n508_, new_n507_ );
not g338 ( new_n510_, new_n503_ );
and g339 ( new_n511_, new_n509_, new_n510_ );
or g340 ( new_n512_, new_n511_, new_n506_ );
and g341 ( new_n513_, new_n505_, new_n512_ );
and g342 ( new_n514_, new_n480_, new_n513_ );
not g343 ( new_n515_, keyIn_0_61 );
not g344 ( new_n516_, keyIn_0_50 );
not g345 ( new_n517_, new_n292_ );
and g346 ( new_n518_, new_n340_, new_n517_ );
and g347 ( new_n519_, new_n310_, new_n292_ );
or g348 ( new_n520_, new_n518_, new_n519_ );
or g349 ( new_n521_, new_n520_, new_n516_ );
or g350 ( new_n522_, new_n310_, new_n292_ );
or g351 ( new_n523_, new_n340_, new_n517_ );
and g352 ( new_n524_, new_n523_, new_n522_ );
or g353 ( new_n525_, new_n524_, keyIn_0_50 );
and g354 ( new_n526_, new_n521_, new_n525_ );
not g355 ( new_n527_, keyIn_0_31 );
not g356 ( new_n528_, N34 );
and g357 ( new_n529_, keyIn_0_5, N30 );
not g358 ( new_n530_, new_n529_ );
or g359 ( new_n531_, keyIn_0_5, N30 );
and g360 ( new_n532_, new_n530_, new_n531_ );
and g361 ( new_n533_, new_n532_, new_n528_ );
not g362 ( new_n534_, new_n533_ );
and g363 ( new_n535_, new_n534_, new_n527_ );
and g364 ( new_n536_, new_n533_, keyIn_0_31 );
or g365 ( new_n537_, new_n535_, new_n536_ );
not g366 ( new_n538_, new_n537_ );
or g367 ( new_n539_, new_n526_, new_n538_ );
and g368 ( new_n540_, new_n539_, new_n515_ );
and g369 ( new_n541_, new_n524_, keyIn_0_50 );
and g370 ( new_n542_, new_n520_, new_n516_ );
or g371 ( new_n543_, new_n542_, new_n541_ );
and g372 ( new_n544_, new_n543_, new_n537_ );
and g373 ( new_n545_, new_n544_, keyIn_0_61 );
or g374 ( new_n546_, new_n540_, new_n545_ );
not g375 ( new_n547_, keyIn_0_62 );
not g376 ( new_n548_, keyIn_0_51 );
not g377 ( new_n549_, new_n277_ );
and g378 ( new_n550_, new_n340_, new_n549_ );
and g379 ( new_n551_, new_n310_, new_n277_ );
or g380 ( new_n552_, new_n550_, new_n551_ );
and g381 ( new_n553_, new_n552_, new_n548_ );
or g382 ( new_n554_, new_n310_, new_n277_ );
or g383 ( new_n555_, new_n340_, new_n549_ );
and g384 ( new_n556_, new_n555_, new_n554_ );
and g385 ( new_n557_, new_n556_, keyIn_0_51 );
or g386 ( new_n558_, new_n553_, new_n557_ );
not g387 ( new_n559_, keyIn_0_33 );
not g388 ( new_n560_, N47 );
and g389 ( new_n561_, keyIn_0_7, N43 );
not g390 ( new_n562_, new_n561_ );
or g391 ( new_n563_, keyIn_0_7, N43 );
and g392 ( new_n564_, new_n562_, new_n563_ );
not g393 ( new_n565_, new_n564_ );
and g394 ( new_n566_, new_n565_, new_n560_ );
not g395 ( new_n567_, new_n566_ );
and g396 ( new_n568_, new_n567_, new_n559_ );
and g397 ( new_n569_, new_n566_, keyIn_0_33 );
or g398 ( new_n570_, new_n568_, new_n569_ );
or g399 ( new_n571_, new_n558_, new_n570_ );
or g400 ( new_n572_, new_n571_, new_n547_ );
or g401 ( new_n573_, new_n556_, keyIn_0_51 );
or g402 ( new_n574_, new_n552_, new_n548_ );
and g403 ( new_n575_, new_n574_, new_n573_ );
not g404 ( new_n576_, new_n570_ );
and g405 ( new_n577_, new_n575_, new_n576_ );
or g406 ( new_n578_, new_n577_, keyIn_0_62 );
and g407 ( new_n579_, new_n572_, new_n578_ );
and g408 ( new_n580_, new_n546_, new_n579_ );
and g409 ( new_n581_, new_n580_, new_n514_ );
and g410 ( new_n582_, new_n581_, new_n447_ );
and g411 ( new_n583_, new_n582_, new_n393_ );
not g412 ( new_n584_, new_n583_ );
and g413 ( new_n585_, new_n584_, new_n301_ );
and g414 ( new_n586_, new_n583_, keyIn_0_76 );
or g415 ( N329, new_n585_, new_n586_ );
not g416 ( new_n588_, keyIn_0_107 );
not g417 ( new_n589_, keyIn_0_98 );
not g418 ( new_n590_, keyIn_0_86 );
and g419 ( new_n591_, N329, new_n590_ );
or g420 ( new_n592_, new_n583_, keyIn_0_76 );
not g421 ( new_n593_, new_n586_ );
and g422 ( new_n594_, new_n593_, new_n592_ );
and g423 ( new_n595_, new_n594_, keyIn_0_86 );
or g424 ( new_n596_, new_n591_, new_n595_ );
and g425 ( new_n597_, new_n596_, new_n391_ );
not g426 ( new_n598_, new_n391_ );
or g427 ( new_n599_, new_n594_, keyIn_0_86 );
or g428 ( new_n600_, N329, new_n590_ );
and g429 ( new_n601_, new_n600_, new_n599_ );
and g430 ( new_n602_, new_n601_, new_n598_ );
or g431 ( new_n603_, new_n597_, new_n602_ );
not g432 ( new_n604_, new_n603_ );
and g433 ( new_n605_, new_n604_, keyIn_0_88 );
not g434 ( new_n606_, keyIn_0_88 );
and g435 ( new_n607_, new_n603_, new_n606_ );
not g436 ( new_n608_, keyIn_0_59 );
not g437 ( new_n609_, N14 );
and g438 ( new_n610_, new_n378_, new_n609_ );
not g439 ( new_n611_, new_n610_ );
and g440 ( new_n612_, new_n611_, keyIn_0_20 );
not g441 ( new_n613_, new_n612_ );
or g442 ( new_n614_, new_n611_, keyIn_0_20 );
and g443 ( new_n615_, new_n613_, new_n614_ );
and g444 ( new_n616_, new_n373_, new_n615_ );
not g445 ( new_n617_, new_n616_ );
and g446 ( new_n618_, new_n617_, new_n608_ );
and g447 ( new_n619_, new_n616_, keyIn_0_59 );
or g448 ( new_n620_, new_n618_, new_n619_ );
and g449 ( new_n621_, new_n620_, keyIn_0_77 );
not g450 ( new_n622_, new_n621_ );
or g451 ( new_n623_, new_n620_, keyIn_0_77 );
and g452 ( new_n624_, new_n622_, new_n623_ );
not g453 ( new_n625_, new_n624_ );
or g454 ( new_n626_, new_n607_, new_n625_ );
or g455 ( new_n627_, new_n626_, new_n605_ );
not g456 ( new_n628_, new_n627_ );
and g457 ( new_n629_, new_n628_, new_n589_ );
and g458 ( new_n630_, new_n627_, keyIn_0_98 );
or g459 ( new_n631_, new_n629_, new_n630_ );
not g460 ( new_n632_, keyIn_0_90 );
and g461 ( new_n633_, new_n596_, new_n546_ );
not g462 ( new_n634_, new_n633_ );
or g463 ( new_n635_, new_n596_, new_n546_ );
and g464 ( new_n636_, new_n634_, new_n635_ );
and g465 ( new_n637_, new_n636_, new_n632_ );
not g466 ( new_n638_, new_n637_ );
or g467 ( new_n639_, new_n636_, new_n632_ );
not g468 ( new_n640_, keyIn_0_79 );
not g469 ( new_n641_, keyIn_0_32 );
not g470 ( new_n642_, N40 );
and g471 ( new_n643_, new_n532_, new_n642_ );
not g472 ( new_n644_, new_n643_ );
and g473 ( new_n645_, new_n644_, new_n641_ );
and g474 ( new_n646_, new_n643_, keyIn_0_32 );
or g475 ( new_n647_, new_n645_, new_n646_ );
and g476 ( new_n648_, new_n543_, new_n647_ );
not g477 ( new_n649_, new_n648_ );
and g478 ( new_n650_, new_n649_, keyIn_0_69 );
not g479 ( new_n651_, new_n650_ );
or g480 ( new_n652_, new_n649_, keyIn_0_69 );
and g481 ( new_n653_, new_n651_, new_n652_ );
not g482 ( new_n654_, new_n653_ );
and g483 ( new_n655_, new_n654_, new_n640_ );
and g484 ( new_n656_, new_n653_, keyIn_0_79 );
or g485 ( new_n657_, new_n655_, new_n656_ );
not g486 ( new_n658_, new_n657_ );
and g487 ( new_n659_, new_n639_, new_n658_ );
and g488 ( new_n660_, new_n659_, new_n638_ );
not g489 ( new_n661_, new_n660_ );
and g490 ( new_n662_, new_n661_, keyIn_0_100 );
not g491 ( new_n663_, keyIn_0_100 );
and g492 ( new_n664_, new_n660_, new_n663_ );
or g493 ( new_n665_, new_n662_, new_n664_ );
not g494 ( new_n666_, keyIn_0_102 );
and g495 ( new_n667_, new_n596_, new_n420_ );
not g496 ( new_n668_, new_n667_ );
or g497 ( new_n669_, new_n596_, new_n420_ );
and g498 ( new_n670_, new_n668_, new_n669_ );
and g499 ( new_n671_, new_n670_, keyIn_0_92 );
not g500 ( new_n672_, new_n671_ );
or g501 ( new_n673_, new_n670_, keyIn_0_92 );
not g502 ( new_n674_, keyIn_0_81 );
not g503 ( new_n675_, keyIn_0_71 );
not g504 ( new_n676_, new_n401_ );
not g505 ( new_n677_, N66 );
and g506 ( new_n678_, new_n407_, new_n677_ );
not g507 ( new_n679_, new_n678_ );
and g508 ( new_n680_, new_n679_, keyIn_0_36 );
not g509 ( new_n681_, new_n680_ );
or g510 ( new_n682_, new_n679_, keyIn_0_36 );
and g511 ( new_n683_, new_n681_, new_n682_ );
or g512 ( new_n684_, new_n676_, new_n683_ );
and g513 ( new_n685_, new_n684_, new_n675_ );
not g514 ( new_n686_, new_n685_ );
or g515 ( new_n687_, new_n684_, new_n675_ );
and g516 ( new_n688_, new_n686_, new_n687_ );
not g517 ( new_n689_, new_n688_ );
and g518 ( new_n690_, new_n689_, new_n674_ );
and g519 ( new_n691_, new_n688_, keyIn_0_81 );
or g520 ( new_n692_, new_n690_, new_n691_ );
and g521 ( new_n693_, new_n673_, new_n692_ );
and g522 ( new_n694_, new_n693_, new_n672_ );
not g523 ( new_n695_, new_n694_ );
and g524 ( new_n696_, new_n695_, new_n666_ );
and g525 ( new_n697_, new_n694_, keyIn_0_102 );
or g526 ( new_n698_, new_n696_, new_n697_ );
and g527 ( new_n699_, new_n665_, new_n698_ );
and g528 ( new_n700_, new_n699_, new_n631_ );
not g529 ( new_n701_, keyIn_0_99 );
and g530 ( new_n702_, new_n596_, new_n335_ );
not g531 ( new_n703_, new_n702_ );
or g532 ( new_n704_, new_n596_, new_n335_ );
and g533 ( new_n705_, new_n703_, new_n704_ );
and g534 ( new_n706_, new_n705_, keyIn_0_89 );
not g535 ( new_n707_, new_n706_ );
or g536 ( new_n708_, new_n705_, keyIn_0_89 );
and g537 ( new_n709_, new_n707_, new_n708_ );
not g538 ( new_n710_, new_n709_ );
not g539 ( new_n711_, keyIn_0_78 );
not g540 ( new_n712_, keyIn_0_68 );
not g541 ( new_n713_, new_n318_ );
not g542 ( new_n714_, N27 );
and g543 ( new_n715_, new_n324_, new_n714_ );
not g544 ( new_n716_, new_n715_ );
and g545 ( new_n717_, new_n716_, keyIn_0_30 );
not g546 ( new_n718_, new_n717_ );
or g547 ( new_n719_, new_n716_, keyIn_0_30 );
and g548 ( new_n720_, new_n718_, new_n719_ );
and g549 ( new_n721_, new_n713_, new_n720_ );
not g550 ( new_n722_, new_n721_ );
and g551 ( new_n723_, new_n722_, new_n712_ );
and g552 ( new_n724_, new_n721_, keyIn_0_68 );
or g553 ( new_n725_, new_n723_, new_n724_ );
and g554 ( new_n726_, new_n725_, new_n711_ );
not g555 ( new_n727_, new_n726_ );
or g556 ( new_n728_, new_n725_, new_n711_ );
and g557 ( new_n729_, new_n727_, new_n728_ );
not g558 ( new_n730_, new_n729_ );
and g559 ( new_n731_, new_n710_, new_n730_ );
or g560 ( new_n732_, new_n731_, new_n701_ );
not g561 ( new_n733_, keyIn_0_101 );
and g562 ( new_n734_, new_n596_, new_n579_ );
not g563 ( new_n735_, new_n734_ );
or g564 ( new_n736_, new_n596_, new_n579_ );
and g565 ( new_n737_, new_n735_, new_n736_ );
or g566 ( new_n738_, new_n737_, keyIn_0_91 );
not g567 ( new_n739_, new_n738_ );
and g568 ( new_n740_, new_n737_, keyIn_0_91 );
or g569 ( new_n741_, new_n739_, new_n740_ );
not g570 ( new_n742_, keyIn_0_80 );
not g571 ( new_n743_, N53 );
and g572 ( new_n744_, new_n565_, new_n743_ );
not g573 ( new_n745_, new_n744_ );
and g574 ( new_n746_, new_n745_, keyIn_0_34 );
not g575 ( new_n747_, new_n746_ );
or g576 ( new_n748_, new_n745_, keyIn_0_34 );
and g577 ( new_n749_, new_n747_, new_n748_ );
or g578 ( new_n750_, new_n558_, new_n749_ );
and g579 ( new_n751_, new_n750_, keyIn_0_70 );
not g580 ( new_n752_, new_n751_ );
or g581 ( new_n753_, new_n750_, keyIn_0_70 );
and g582 ( new_n754_, new_n752_, new_n753_ );
not g583 ( new_n755_, new_n754_ );
and g584 ( new_n756_, new_n755_, new_n742_ );
and g585 ( new_n757_, new_n754_, keyIn_0_80 );
or g586 ( new_n758_, new_n756_, new_n757_ );
and g587 ( new_n759_, new_n741_, new_n758_ );
or g588 ( new_n760_, new_n759_, new_n733_ );
and g589 ( new_n761_, new_n732_, new_n760_ );
or g590 ( new_n762_, new_n709_, new_n729_ );
or g591 ( new_n763_, new_n762_, keyIn_0_99 );
not g592 ( new_n764_, new_n740_ );
and g593 ( new_n765_, new_n764_, new_n738_ );
not g594 ( new_n766_, new_n758_ );
or g595 ( new_n767_, new_n765_, new_n766_ );
or g596 ( new_n768_, new_n767_, keyIn_0_101 );
and g597 ( new_n769_, new_n763_, new_n768_ );
and g598 ( new_n770_, new_n761_, new_n769_ );
and g599 ( new_n771_, new_n596_, new_n480_ );
not g600 ( new_n772_, new_n480_ );
and g601 ( new_n773_, new_n601_, new_n772_ );
or g602 ( new_n774_, new_n771_, new_n773_ );
or g603 ( new_n775_, new_n774_, keyIn_0_96 );
not g604 ( new_n776_, keyIn_0_96 );
or g605 ( new_n777_, new_n601_, new_n772_ );
or g606 ( new_n778_, new_n596_, new_n480_ );
and g607 ( new_n779_, new_n778_, new_n777_ );
or g608 ( new_n780_, new_n779_, new_n776_ );
and g609 ( new_n781_, new_n775_, new_n780_ );
not g610 ( new_n782_, keyIn_0_84 );
not g611 ( new_n783_, N105 );
and g612 ( new_n784_, new_n466_, new_n783_ );
not g613 ( new_n785_, new_n784_ );
and g614 ( new_n786_, new_n785_, keyIn_0_42 );
not g615 ( new_n787_, new_n786_ );
or g616 ( new_n788_, new_n785_, keyIn_0_42 );
and g617 ( new_n789_, new_n787_, new_n788_ );
and g618 ( new_n790_, new_n476_, new_n789_ );
not g619 ( new_n791_, new_n790_ );
and g620 ( new_n792_, new_n791_, keyIn_0_74 );
not g621 ( new_n793_, new_n792_ );
or g622 ( new_n794_, new_n791_, keyIn_0_74 );
and g623 ( new_n795_, new_n793_, new_n794_ );
not g624 ( new_n796_, new_n795_ );
and g625 ( new_n797_, new_n796_, new_n782_ );
and g626 ( new_n798_, new_n795_, keyIn_0_84 );
or g627 ( new_n799_, new_n797_, new_n798_ );
or g628 ( new_n800_, new_n781_, new_n799_ );
or g629 ( new_n801_, new_n800_, keyIn_0_105 );
not g630 ( new_n802_, keyIn_0_105 );
and g631 ( new_n803_, new_n779_, new_n776_ );
and g632 ( new_n804_, new_n774_, keyIn_0_96 );
or g633 ( new_n805_, new_n804_, new_n803_ );
not g634 ( new_n806_, new_n799_ );
and g635 ( new_n807_, new_n805_, new_n806_ );
or g636 ( new_n808_, new_n807_, new_n802_ );
and g637 ( new_n809_, new_n801_, new_n808_ );
not g638 ( new_n810_, new_n513_ );
or g639 ( new_n811_, new_n601_, new_n810_ );
or g640 ( new_n812_, new_n596_, new_n513_ );
and g641 ( new_n813_, new_n812_, new_n811_ );
and g642 ( new_n814_, new_n813_, keyIn_0_97 );
not g643 ( new_n815_, keyIn_0_97 );
and g644 ( new_n816_, new_n596_, new_n513_ );
and g645 ( new_n817_, new_n601_, new_n810_ );
or g646 ( new_n818_, new_n816_, new_n817_ );
and g647 ( new_n819_, new_n818_, new_n815_ );
not g648 ( new_n820_, N115 );
and g649 ( new_n821_, new_n498_, new_n820_ );
not g650 ( new_n822_, new_n821_ );
and g651 ( new_n823_, new_n822_, keyIn_0_44 );
not g652 ( new_n824_, new_n823_ );
or g653 ( new_n825_, new_n822_, keyIn_0_44 );
and g654 ( new_n826_, new_n824_, new_n825_ );
or g655 ( new_n827_, new_n491_, new_n826_ );
and g656 ( new_n828_, new_n827_, keyIn_0_75 );
not g657 ( new_n829_, new_n828_ );
or g658 ( new_n830_, new_n827_, keyIn_0_75 );
and g659 ( new_n831_, new_n829_, new_n830_ );
not g660 ( new_n832_, new_n831_ );
and g661 ( new_n833_, new_n832_, keyIn_0_85 );
not g662 ( new_n834_, new_n833_ );
or g663 ( new_n835_, new_n832_, keyIn_0_85 );
and g664 ( new_n836_, new_n834_, new_n835_ );
or g665 ( new_n837_, new_n819_, new_n836_ );
or g666 ( new_n838_, new_n837_, new_n814_ );
or g667 ( new_n839_, new_n838_, keyIn_0_106 );
not g668 ( new_n840_, keyIn_0_106 );
not g669 ( new_n841_, new_n814_ );
or g670 ( new_n842_, new_n813_, keyIn_0_97 );
not g671 ( new_n843_, new_n836_ );
and g672 ( new_n844_, new_n842_, new_n843_ );
and g673 ( new_n845_, new_n844_, new_n841_ );
or g674 ( new_n846_, new_n845_, new_n840_ );
and g675 ( new_n847_, new_n839_, new_n846_ );
and g676 ( new_n848_, new_n809_, new_n847_ );
not g677 ( new_n849_, keyIn_0_103 );
not g678 ( new_n850_, keyIn_0_93 );
and g679 ( new_n851_, new_n596_, new_n446_ );
not g680 ( new_n852_, new_n446_ );
and g681 ( new_n853_, new_n601_, new_n852_ );
or g682 ( new_n854_, new_n851_, new_n853_ );
or g683 ( new_n855_, new_n854_, new_n850_ );
or g684 ( new_n856_, new_n601_, new_n852_ );
or g685 ( new_n857_, new_n596_, new_n446_ );
and g686 ( new_n858_, new_n857_, new_n856_ );
or g687 ( new_n859_, new_n858_, keyIn_0_93 );
and g688 ( new_n860_, new_n855_, new_n859_ );
not g689 ( new_n861_, keyIn_0_82 );
not g690 ( new_n862_, new_n428_ );
not g691 ( new_n863_, N79 );
and g692 ( new_n864_, new_n433_, new_n863_ );
not g693 ( new_n865_, new_n864_ );
and g694 ( new_n866_, new_n865_, keyIn_0_38 );
not g695 ( new_n867_, new_n866_ );
or g696 ( new_n868_, new_n865_, keyIn_0_38 );
and g697 ( new_n869_, new_n867_, new_n868_ );
or g698 ( new_n870_, new_n862_, new_n869_ );
and g699 ( new_n871_, new_n870_, keyIn_0_72 );
not g700 ( new_n872_, new_n871_ );
or g701 ( new_n873_, new_n870_, keyIn_0_72 );
and g702 ( new_n874_, new_n872_, new_n873_ );
not g703 ( new_n875_, new_n874_ );
and g704 ( new_n876_, new_n875_, new_n861_ );
and g705 ( new_n877_, new_n874_, keyIn_0_82 );
or g706 ( new_n878_, new_n876_, new_n877_ );
or g707 ( new_n879_, new_n860_, new_n878_ );
or g708 ( new_n880_, new_n879_, new_n849_ );
not g709 ( new_n881_, keyIn_0_104 );
not g710 ( new_n882_, keyIn_0_94 );
and g711 ( new_n883_, new_n596_, new_n365_ );
not g712 ( new_n884_, new_n365_ );
and g713 ( new_n885_, new_n601_, new_n884_ );
or g714 ( new_n886_, new_n883_, new_n885_ );
or g715 ( new_n887_, new_n886_, new_n882_ );
or g716 ( new_n888_, new_n601_, new_n884_ );
or g717 ( new_n889_, new_n596_, new_n365_ );
and g718 ( new_n890_, new_n889_, new_n888_ );
or g719 ( new_n891_, new_n890_, keyIn_0_94 );
and g720 ( new_n892_, new_n887_, new_n891_ );
not g721 ( new_n893_, keyIn_0_83 );
not g722 ( new_n894_, new_n347_ );
not g723 ( new_n895_, N92 );
and g724 ( new_n896_, new_n352_, new_n895_ );
not g725 ( new_n897_, new_n896_ );
and g726 ( new_n898_, new_n897_, keyIn_0_40 );
not g727 ( new_n899_, new_n898_ );
or g728 ( new_n900_, new_n897_, keyIn_0_40 );
and g729 ( new_n901_, new_n899_, new_n900_ );
or g730 ( new_n902_, new_n894_, new_n901_ );
and g731 ( new_n903_, new_n902_, keyIn_0_73 );
not g732 ( new_n904_, new_n903_ );
or g733 ( new_n905_, new_n902_, keyIn_0_73 );
and g734 ( new_n906_, new_n904_, new_n905_ );
not g735 ( new_n907_, new_n906_ );
and g736 ( new_n908_, new_n907_, new_n893_ );
and g737 ( new_n909_, new_n906_, keyIn_0_83 );
or g738 ( new_n910_, new_n908_, new_n909_ );
or g739 ( new_n911_, new_n892_, new_n910_ );
or g740 ( new_n912_, new_n911_, new_n881_ );
and g741 ( new_n913_, new_n880_, new_n912_ );
and g742 ( new_n914_, new_n858_, keyIn_0_93 );
and g743 ( new_n915_, new_n854_, new_n850_ );
or g744 ( new_n916_, new_n915_, new_n914_ );
not g745 ( new_n917_, new_n878_ );
and g746 ( new_n918_, new_n916_, new_n917_ );
or g747 ( new_n919_, new_n918_, keyIn_0_103 );
and g748 ( new_n920_, new_n890_, keyIn_0_94 );
and g749 ( new_n921_, new_n886_, new_n882_ );
or g750 ( new_n922_, new_n921_, new_n920_ );
not g751 ( new_n923_, new_n910_ );
and g752 ( new_n924_, new_n922_, new_n923_ );
or g753 ( new_n925_, new_n924_, keyIn_0_104 );
and g754 ( new_n926_, new_n919_, new_n925_ );
and g755 ( new_n927_, new_n913_, new_n926_ );
and g756 ( new_n928_, new_n848_, new_n927_ );
and g757 ( new_n929_, new_n928_, new_n770_ );
and g758 ( new_n930_, new_n929_, new_n700_ );
not g759 ( new_n931_, new_n930_ );
and g760 ( new_n932_, new_n931_, new_n588_ );
and g761 ( new_n933_, new_n930_, keyIn_0_107 );
or g762 ( N370, new_n932_, new_n933_ );
not g763 ( new_n935_, keyIn_0_120 );
not g764 ( new_n936_, keyIn_0_113 );
or g765 ( new_n937_, new_n930_, keyIn_0_107 );
not g766 ( new_n938_, new_n933_ );
and g767 ( new_n939_, new_n938_, new_n937_ );
or g768 ( new_n940_, new_n939_, keyIn_0_108 );
not g769 ( new_n941_, keyIn_0_108 );
or g770 ( new_n942_, N370, new_n941_ );
and g771 ( new_n943_, new_n942_, new_n940_ );
or g772 ( new_n944_, new_n943_, new_n743_ );
or g773 ( new_n945_, new_n944_, keyIn_0_109 );
not g774 ( new_n946_, keyIn_0_109 );
and g775 ( new_n947_, N370, new_n941_ );
and g776 ( new_n948_, new_n939_, keyIn_0_108 );
or g777 ( new_n949_, new_n947_, new_n948_ );
and g778 ( new_n950_, new_n949_, N53 );
or g779 ( new_n951_, new_n950_, new_n946_ );
and g780 ( new_n952_, new_n945_, new_n951_ );
not g781 ( new_n953_, keyIn_0_95 );
and g782 ( new_n954_, N329, keyIn_0_87 );
not g783 ( new_n955_, new_n954_ );
or g784 ( new_n956_, N329, keyIn_0_87 );
and g785 ( new_n957_, new_n955_, new_n956_ );
not g786 ( new_n958_, new_n957_ );
and g787 ( new_n959_, new_n958_, N47 );
not g788 ( new_n960_, new_n959_ );
and g789 ( new_n961_, new_n960_, new_n953_ );
and g790 ( new_n962_, new_n959_, keyIn_0_95 );
or g791 ( new_n963_, new_n961_, new_n962_ );
and g792 ( new_n964_, N223, keyIn_0_47 );
not g793 ( new_n965_, new_n964_ );
or g794 ( new_n966_, N223, keyIn_0_47 );
and g795 ( new_n967_, new_n965_, new_n966_ );
and g796 ( new_n968_, new_n967_, N37 );
not g797 ( new_n969_, new_n968_ );
and g798 ( new_n970_, new_n969_, keyIn_0_57 );
not g799 ( new_n971_, new_n970_ );
or g800 ( new_n972_, new_n969_, keyIn_0_57 );
and g801 ( new_n973_, new_n971_, new_n972_ );
or g802 ( new_n974_, new_n973_, new_n271_ );
not g803 ( new_n975_, new_n974_ );
and g804 ( new_n976_, new_n963_, new_n975_ );
not g805 ( new_n977_, new_n976_ );
or g806 ( new_n978_, new_n952_, new_n977_ );
and g807 ( new_n979_, new_n978_, new_n936_ );
and g808 ( new_n980_, new_n950_, new_n946_ );
and g809 ( new_n981_, new_n944_, keyIn_0_109 );
or g810 ( new_n982_, new_n981_, new_n980_ );
and g811 ( new_n983_, new_n982_, new_n976_ );
and g812 ( new_n984_, new_n983_, keyIn_0_113 );
or g813 ( new_n985_, new_n979_, new_n984_ );
and g814 ( new_n986_, new_n949_, N66 );
and g815 ( new_n987_, new_n958_, N60 );
and g816 ( new_n988_, new_n967_, N50 );
or g817 ( new_n989_, new_n988_, new_n234_ );
or g818 ( new_n990_, new_n987_, new_n989_ );
or g819 ( new_n991_, new_n986_, new_n990_ );
not g820 ( new_n992_, new_n991_ );
and g821 ( new_n993_, new_n992_, keyIn_0_114 );
not g822 ( new_n994_, keyIn_0_114 );
and g823 ( new_n995_, new_n991_, new_n994_ );
or g824 ( new_n996_, new_n993_, new_n995_ );
not g825 ( new_n997_, new_n996_ );
and g826 ( new_n998_, new_n985_, new_n997_ );
not g827 ( new_n999_, keyIn_0_111 );
and g828 ( new_n1000_, new_n949_, N27 );
and g829 ( new_n1001_, new_n958_, N21 );
and g830 ( new_n1002_, new_n967_, N11 );
or g831 ( new_n1003_, new_n1002_, new_n175_ );
or g832 ( new_n1004_, new_n1001_, new_n1003_ );
or g833 ( new_n1005_, new_n1000_, new_n1004_ );
and g834 ( new_n1006_, new_n1005_, new_n999_ );
not g835 ( new_n1007_, new_n1006_ );
or g836 ( new_n1008_, new_n1005_, new_n999_ );
and g837 ( new_n1009_, new_n1007_, new_n1008_ );
and g838 ( new_n1010_, new_n949_, N40 );
and g839 ( new_n1011_, new_n958_, N34 );
and g840 ( new_n1012_, new_n967_, N24 );
or g841 ( new_n1013_, new_n1012_, new_n281_ );
or g842 ( new_n1014_, new_n1011_, new_n1013_ );
or g843 ( new_n1015_, new_n1010_, new_n1014_ );
and g844 ( new_n1016_, new_n1015_, keyIn_0_112 );
not g845 ( new_n1017_, new_n1016_ );
or g846 ( new_n1018_, new_n1015_, keyIn_0_112 );
and g847 ( new_n1019_, new_n1017_, new_n1018_ );
and g848 ( new_n1020_, new_n1009_, new_n1019_ );
not g849 ( new_n1021_, keyIn_0_117 );
and g850 ( new_n1022_, new_n949_, N105 );
and g851 ( new_n1023_, new_n958_, N99 );
and g852 ( new_n1024_, new_n967_, N89 );
or g853 ( new_n1025_, new_n1024_, new_n186_ );
or g854 ( new_n1026_, new_n1023_, new_n1025_ );
or g855 ( new_n1027_, new_n1022_, new_n1026_ );
and g856 ( new_n1028_, new_n1027_, new_n1021_ );
not g857 ( new_n1029_, new_n1028_ );
or g858 ( new_n1030_, new_n1027_, new_n1021_ );
and g859 ( new_n1031_, new_n1029_, new_n1030_ );
not g860 ( new_n1032_, new_n1031_ );
and g861 ( new_n1033_, new_n949_, N115 );
and g862 ( new_n1034_, new_n958_, N112 );
not g863 ( new_n1035_, N108 );
and g864 ( new_n1036_, new_n967_, N102 );
or g865 ( new_n1037_, new_n1036_, new_n1035_ );
or g866 ( new_n1038_, new_n1034_, new_n1037_ );
or g867 ( new_n1039_, new_n1033_, new_n1038_ );
not g868 ( new_n1040_, new_n1039_ );
and g869 ( new_n1041_, new_n1040_, keyIn_0_118 );
not g870 ( new_n1042_, keyIn_0_118 );
and g871 ( new_n1043_, new_n1039_, new_n1042_ );
or g872 ( new_n1044_, new_n1041_, new_n1043_ );
and g873 ( new_n1045_, new_n1032_, new_n1044_ );
not g874 ( new_n1046_, keyIn_0_115 );
and g875 ( new_n1047_, new_n949_, N79 );
and g876 ( new_n1048_, new_n958_, N73 );
and g877 ( new_n1049_, new_n967_, N63 );
or g878 ( new_n1050_, new_n1049_, new_n250_ );
or g879 ( new_n1051_, new_n1048_, new_n1050_ );
or g880 ( new_n1052_, new_n1047_, new_n1051_ );
not g881 ( new_n1053_, new_n1052_ );
or g882 ( new_n1054_, new_n1053_, new_n1046_ );
or g883 ( new_n1055_, new_n1052_, keyIn_0_115 );
and g884 ( new_n1056_, new_n1054_, new_n1055_ );
and g885 ( new_n1057_, new_n949_, N92 );
and g886 ( new_n1058_, new_n958_, N86 );
not g887 ( new_n1059_, N82 );
and g888 ( new_n1060_, new_n967_, N76 );
or g889 ( new_n1061_, new_n1060_, new_n1059_ );
or g890 ( new_n1062_, new_n1058_, new_n1061_ );
or g891 ( new_n1063_, new_n1057_, new_n1062_ );
and g892 ( new_n1064_, new_n1063_, keyIn_0_116 );
not g893 ( new_n1065_, new_n1064_ );
or g894 ( new_n1066_, new_n1063_, keyIn_0_116 );
and g895 ( new_n1067_, new_n1065_, new_n1066_ );
and g896 ( new_n1068_, new_n1056_, new_n1067_ );
and g897 ( new_n1069_, new_n1045_, new_n1068_ );
and g898 ( new_n1070_, new_n1069_, new_n1020_ );
and g899 ( new_n1071_, new_n1070_, new_n998_ );
and g900 ( new_n1072_, new_n1071_, keyIn_0_119 );
not g901 ( new_n1073_, new_n1072_ );
or g902 ( new_n1074_, new_n1071_, keyIn_0_119 );
not g903 ( new_n1075_, keyIn_0_110 );
and g904 ( new_n1076_, new_n949_, N14 );
and g905 ( new_n1077_, new_n958_, N8 );
not g906 ( new_n1078_, N4 );
and g907 ( new_n1079_, new_n967_, N1 );
or g908 ( new_n1080_, new_n1079_, new_n1078_ );
or g909 ( new_n1081_, new_n1077_, new_n1080_ );
or g910 ( new_n1082_, new_n1076_, new_n1081_ );
not g911 ( new_n1083_, new_n1082_ );
or g912 ( new_n1084_, new_n1083_, new_n1075_ );
or g913 ( new_n1085_, new_n1082_, keyIn_0_110 );
and g914 ( new_n1086_, new_n1084_, new_n1085_ );
and g915 ( new_n1087_, new_n1074_, new_n1086_ );
and g916 ( new_n1088_, new_n1087_, new_n1073_ );
and g917 ( new_n1089_, new_n1088_, new_n935_ );
not g918 ( new_n1090_, new_n1089_ );
or g919 ( new_n1091_, new_n1088_, new_n935_ );
and g920 ( N421, new_n1090_, new_n1091_ );
not g921 ( new_n1093_, keyIn_0_125 );
not g922 ( new_n1094_, keyIn_0_121 );
not g923 ( new_n1095_, new_n1019_ );
or g924 ( new_n1096_, new_n985_, new_n1095_ );
and g925 ( new_n1097_, new_n1096_, new_n1094_ );
or g926 ( new_n1098_, new_n983_, keyIn_0_113 );
or g927 ( new_n1099_, new_n978_, new_n936_ );
and g928 ( new_n1100_, new_n1099_, new_n1098_ );
and g929 ( new_n1101_, new_n1100_, new_n1019_ );
and g930 ( new_n1102_, new_n1101_, keyIn_0_121 );
or g931 ( new_n1103_, new_n1097_, new_n1102_ );
and g932 ( new_n1104_, new_n1020_, new_n997_ );
and g933 ( new_n1105_, new_n1103_, new_n1104_ );
not g934 ( new_n1106_, new_n1105_ );
and g935 ( new_n1107_, new_n1106_, new_n1093_ );
and g936 ( new_n1108_, new_n1105_, keyIn_0_125 );
or g937 ( N430, new_n1107_, new_n1108_ );
or g938 ( new_n1110_, new_n1100_, new_n996_ );
or g939 ( new_n1111_, new_n1095_, new_n1056_ );
or g940 ( new_n1112_, new_n1110_, new_n1111_ );
and g941 ( new_n1113_, new_n1112_, keyIn_0_122 );
not g942 ( new_n1114_, new_n1113_ );
or g943 ( new_n1115_, new_n1112_, keyIn_0_122 );
and g944 ( new_n1116_, new_n1114_, new_n1115_ );
not g945 ( new_n1117_, new_n1116_ );
not g946 ( new_n1118_, new_n1020_ );
or g947 ( new_n1119_, new_n1110_, new_n1067_ );
or g948 ( new_n1120_, new_n1119_, keyIn_0_123 );
not g949 ( new_n1121_, keyIn_0_123 );
not g950 ( new_n1122_, new_n1067_ );
and g951 ( new_n1123_, new_n998_, new_n1122_ );
or g952 ( new_n1124_, new_n1123_, new_n1121_ );
and g953 ( new_n1125_, new_n1120_, new_n1124_ );
or g954 ( new_n1126_, new_n1125_, new_n1118_ );
or g955 ( new_n1127_, new_n1126_, new_n1117_ );
or g956 ( new_n1128_, new_n1127_, keyIn_0_126 );
not g957 ( new_n1129_, keyIn_0_126 );
and g958 ( new_n1130_, new_n1123_, new_n1121_ );
and g959 ( new_n1131_, new_n1119_, keyIn_0_123 );
or g960 ( new_n1132_, new_n1131_, new_n1130_ );
and g961 ( new_n1133_, new_n1132_, new_n1020_ );
and g962 ( new_n1134_, new_n1133_, new_n1116_ );
or g963 ( new_n1135_, new_n1134_, new_n1129_ );
and g964 ( N431, new_n1128_, new_n1135_ );
not g965 ( new_n1137_, keyIn_0_127 );
and g966 ( new_n1138_, new_n1031_, new_n1067_ );
and g967 ( new_n1139_, new_n1138_, new_n1019_ );
and g968 ( new_n1140_, new_n1139_, new_n985_ );
not g969 ( new_n1141_, new_n1140_ );
and g970 ( new_n1142_, new_n1141_, keyIn_0_124 );
not g971 ( new_n1143_, new_n1142_ );
not g972 ( new_n1144_, keyIn_0_124 );
and g973 ( new_n1145_, new_n1140_, new_n1144_ );
not g974 ( new_n1146_, new_n1145_ );
and g975 ( new_n1147_, new_n1143_, new_n1146_ );
not g976 ( new_n1148_, new_n1009_ );
or g977 ( new_n1149_, new_n1101_, keyIn_0_121 );
or g978 ( new_n1150_, new_n1096_, new_n1094_ );
and g979 ( new_n1151_, new_n1150_, new_n1149_ );
or g980 ( new_n1152_, new_n1151_, new_n1148_ );
or g981 ( new_n1153_, new_n1152_, new_n1147_ );
or g982 ( new_n1154_, new_n1153_, new_n1117_ );
or g983 ( new_n1155_, new_n1154_, new_n1137_ );
or g984 ( new_n1156_, new_n1142_, new_n1145_ );
and g985 ( new_n1157_, new_n1103_, new_n1009_ );
and g986 ( new_n1158_, new_n1157_, new_n1156_ );
and g987 ( new_n1159_, new_n1158_, new_n1116_ );
or g988 ( new_n1160_, new_n1159_, keyIn_0_127 );
and g989 ( N432, new_n1155_, new_n1160_ );
endmodule