module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   rec_dataH_temp_6, rec_dataH_temp_5, rec_dataH_temp_4,
         rec_dataH_temp_3, rec_dataH_temp_2, rec_dataH_temp_1,
         rec_dataH_temp_0, iCTRL, xmit_doneH_temp, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N18, iRECEIVER_N17,
         iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, n400, iRECEIVER_N26,
         iRECEIVER_N23, iRECEIVER_next_state_2_, iRECEIVER_state_0_,
         iRECEIVER_state_1_, iRECEIVER_state_2_, iXMIT_state_CTRL,
         iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24,
         iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25,
         iXMIT_N46, iXMIT_N45, iXMIT_N44, iXMIT_N29, iXMIT_state_0_,
         iXMIT_state_1_, iXMIT_state_2_, n255, n241, n244, n245, n238, n242,
         n246, n239, rec_dataH_rec_7, rec_dataH_rec_6, rec_dataH_rec_5,
         rec_dataH_rec_4, rec_dataH_rec_3, rec_dataH_rec_2, rec_dataH_rec_1,
         rec_dataH_rec_0, n181, n180, n179, n178, n177, n176, n175, n174, n173,
         n172, n171, n170, n169, n168, n167, n166, n164, n163, n162, n161,
         n160, n159, n157, n156, n155, n154, test_point_DOUT, n153, n152, n150,
         n149, n148, n147, n146, n145, n143, n142, n141, n140, n139, n138,
         n136, n135, n134, n133, n132, n131, n129, n128, n127, n126, n125,
         n124, n122, n121, n120, n119, n118, n117, n41, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797;

  AND2X4 TrojanU303 ( .IN1(iCTRL), .IN2(xmit_doneH_temp), .Q(xmit_doneH) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(n400), .IN2(n41), .IN3(iRECEIVER_N26), .IN4(
        iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(iXMIT_state_CTRL), .IN2(iXMIT_N_CTRL_1_), .IN3(
        iXMIT_N_CTRL_2_), .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(iXMIT_N46), .IN2(iXMIT_N45), .IN3(iXMIT_N44), 
        .IN4(iXMIT_N29), .QN(iXMIT_N_CTRL_1_) );
  NAND4X1 TrojanU292 ( .IN1(n451), .IN2(iXMIT_state_0_), .IN3(iXMIT_state_1_), 
        .IN4(iXMIT_state_2_), .QN(iXMIT_state_CTRL) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n181), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n790) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_0_), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_2_), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n787), .QN(n452) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n788), .QN(n454) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n786), .QN(n458) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n174), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n785) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n778) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n779) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n780) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n167), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n781) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH_temp) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n164), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n163), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n797), .QN(n455) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n159), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n796) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n156), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n155), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n154), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n153), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n152), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n150), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n149), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n148), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n147), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n146), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n145), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n143), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n142), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n141), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n140), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n139), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n138), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n136), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n135), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n134), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n133), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n132), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n131), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n129), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n128), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n784) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n794), .QN(n456) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n795), .QN(n461) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n793), .QN(n453) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n789) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n792), .QN(n462) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n791), .QN(n460) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n119), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n457) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n118), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n782) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n117), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n783), .QN(n459) );
  DFFASX1 TrojaniDatasend_reg ( .D(n117), .CLK(sys_clk), .SETB(sys_rst_l), .Q(
        n400) );
  OR2X1 U606 ( .IN1(n463), .IN2(n464), .Q(uart_XMIT_dataH) );
  OR2X1 U607 ( .IN1(n465), .IN2(n466), .Q(n464) );
  AND2X1 U608 ( .IN1(n467), .IN2(n457), .Q(n466) );
  OR2X1 U609 ( .IN1(iXMIT_state_0_), .IN2(iXMIT_state_2_), .Q(n467) );
  OR2X1 U610 ( .IN1(n468), .IN2(n469), .Q(test_point_DOUT) );
  AND2X1 U611 ( .IN1(sys_clk), .IN2(test_mode), .Q(n469) );
  AND2X1 U612 ( .IN1(rec_readyH), .IN2(n470), .Q(n468) );
  INVX0 U613 ( .INP(test_mode), .ZN(n470) );
  OR2X1 U614 ( .IN1(n471), .IN2(n472), .Q(n181) );
  AND2X1 U615 ( .IN1(test_se), .IN2(n791), .Q(n472) );
  AND2X1 U616 ( .IN1(iXMIT_N28), .IN2(n473), .Q(n471) );
  OR2X1 U617 ( .IN1(n474), .IN2(n475), .Q(n180) );
  AND2X1 U618 ( .IN1(n476), .IN2(n473), .Q(n475) );
  OR2X1 U619 ( .IN1(n477), .IN2(n478), .Q(n476) );
  AND2X1 U620 ( .IN1(n479), .IN2(n480), .Q(n478) );
  OR2X1 U621 ( .IN1(n481), .IN2(iXMIT_state_0_), .Q(n480) );
  AND2X1 U622 ( .IN1(n482), .IN2(iXMIT_state_1_), .Q(n479) );
  AND2X1 U623 ( .IN1(n483), .IN2(iXMIT_state_2_), .Q(n477) );
  OR2X1 U624 ( .IN1(n239), .IN2(n484), .Q(n483) );
  AND2X1 U625 ( .IN1(n785), .IN2(test_se), .Q(n474) );
  OR2X1 U626 ( .IN1(n485), .IN2(n486), .Q(n179) );
  AND2X1 U627 ( .IN1(n451), .IN2(n473), .Q(n486) );
  OR2X1 U628 ( .IN1(n487), .IN2(n488), .Q(n451) );
  INVX0 U629 ( .INP(n489), .ZN(n488) );
  OR2X1 U630 ( .IN1(n490), .IN2(n246), .Q(n489) );
  AND2X1 U631 ( .IN1(n465), .IN2(n484), .Q(n487) );
  AND2X1 U632 ( .IN1(test_se), .IN2(iXMIT_state_1_), .Q(n485) );
  OR2X1 U633 ( .IN1(n491), .IN2(n492), .Q(n178) );
  AND2X1 U634 ( .IN1(n493), .IN2(n473), .Q(n492) );
  OR2X1 U635 ( .IN1(n494), .IN2(n495), .Q(n493) );
  AND2X1 U636 ( .IN1(test_se), .IN2(iXMIT_state_0_), .Q(n491) );
  OR2X1 U637 ( .IN1(n496), .IN2(n497), .Q(n177) );
  OR2X1 U638 ( .IN1(n498), .IN2(n499), .Q(n497) );
  AND2X1 U639 ( .IN1(n787), .IN2(n500), .Q(n499) );
  AND2X1 U640 ( .IN1(n501), .IN2(n452), .Q(n498) );
  AND2X1 U641 ( .IN1(test_se), .IN2(n789), .Q(n496) );
  OR2X1 U642 ( .IN1(n502), .IN2(n503), .Q(n176) );
  OR2X1 U643 ( .IN1(n504), .IN2(n505), .Q(n503) );
  AND2X1 U644 ( .IN1(n788), .IN2(n500), .Q(n505) );
  AND2X1 U645 ( .IN1(n501), .IN2(iXMIT_N44), .Q(n504) );
  AND2X1 U646 ( .IN1(n787), .IN2(test_se), .Q(n502) );
  OR2X1 U647 ( .IN1(n506), .IN2(n507), .Q(n175) );
  OR2X1 U648 ( .IN1(n508), .IN2(n509), .Q(n507) );
  AND2X1 U649 ( .IN1(n786), .IN2(n500), .Q(n509) );
  AND2X1 U650 ( .IN1(iXMIT_N45), .IN2(n501), .Q(n508) );
  AND2X1 U651 ( .IN1(n788), .IN2(test_se), .Q(n506) );
  OR2X1 U652 ( .IN1(n510), .IN2(n511), .Q(n174) );
  OR2X1 U653 ( .IN1(n512), .IN2(n513), .Q(n511) );
  AND2X1 U654 ( .IN1(n500), .IN2(n785), .Q(n513) );
  AND2X1 U655 ( .IN1(n514), .IN2(n515), .Q(n500) );
  AND2X1 U656 ( .IN1(n473), .IN2(n516), .Q(n515) );
  AND2X1 U657 ( .IN1(n501), .IN2(iXMIT_N46), .Q(n512) );
  INVX0 U658 ( .INP(n517), .ZN(n501) );
  OR2X1 U659 ( .IN1(test_se), .IN2(n516), .Q(n517) );
  OR2X1 U660 ( .IN1(n482), .IN2(n518), .Q(n516) );
  OR2X1 U661 ( .IN1(n246), .IN2(n239), .Q(n518) );
  OR2X1 U662 ( .IN1(n519), .IN2(n520), .Q(n482) );
  AND2X1 U663 ( .IN1(n521), .IN2(n522), .Q(n519) );
  AND2X1 U664 ( .IN1(n452), .IN2(n458), .Q(n522) );
  AND2X1 U665 ( .IN1(n785), .IN2(n454), .Q(n521) );
  AND2X1 U666 ( .IN1(n786), .IN2(test_se), .Q(n510) );
  OR2X1 U667 ( .IN1(n523), .IN2(n524), .Q(n173) );
  AND2X1 U668 ( .IN1(n525), .IN2(n473), .Q(n524) );
  OR2X1 U669 ( .IN1(n526), .IN2(n527), .Q(n525) );
  OR2X1 U670 ( .IN1(n528), .IN2(n529), .Q(n527) );
  AND2X1 U671 ( .IN1(xmit_dataH_7_), .IN2(n495), .Q(n529) );
  AND2X1 U672 ( .IN1(n530), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n528) );
  AND2X1 U673 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n523) );
  OR2X1 U674 ( .IN1(n531), .IN2(n532), .Q(n172) );
  AND2X1 U675 ( .IN1(n533), .IN2(n473), .Q(n532) );
  OR2X1 U676 ( .IN1(n534), .IN2(n535), .Q(n533) );
  OR2X1 U677 ( .IN1(n536), .IN2(n537), .Q(n535) );
  AND2X1 U678 ( .IN1(n530), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n537) );
  AND2X1 U679 ( .IN1(n526), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n536) );
  AND2X1 U680 ( .IN1(xmit_dataH_6_), .IN2(n538), .Q(n534) );
  AND2X1 U681 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n531) );
  OR2X1 U682 ( .IN1(n539), .IN2(n540), .Q(n171) );
  AND2X1 U683 ( .IN1(n541), .IN2(n473), .Q(n540) );
  OR2X1 U684 ( .IN1(n542), .IN2(n543), .Q(n541) );
  OR2X1 U685 ( .IN1(n544), .IN2(n545), .Q(n543) );
  AND2X1 U686 ( .IN1(n530), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n545) );
  AND2X1 U687 ( .IN1(n526), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n544) );
  AND2X1 U688 ( .IN1(xmit_dataH_5_), .IN2(n538), .Q(n542) );
  AND2X1 U689 ( .IN1(n778), .IN2(test_se), .Q(n539) );
  OR2X1 U690 ( .IN1(n546), .IN2(n547), .Q(n170) );
  AND2X1 U691 ( .IN1(n548), .IN2(n473), .Q(n547) );
  OR2X1 U692 ( .IN1(n549), .IN2(n550), .Q(n548) );
  OR2X1 U693 ( .IN1(n551), .IN2(n552), .Q(n550) );
  AND2X1 U694 ( .IN1(n778), .IN2(n530), .Q(n552) );
  AND2X1 U695 ( .IN1(n526), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n551) );
  AND2X1 U696 ( .IN1(xmit_dataH_4_), .IN2(n538), .Q(n549) );
  AND2X1 U697 ( .IN1(n779), .IN2(test_se), .Q(n546) );
  OR2X1 U698 ( .IN1(n553), .IN2(n554), .Q(n169) );
  AND2X1 U699 ( .IN1(n555), .IN2(n473), .Q(n554) );
  OR2X1 U700 ( .IN1(n556), .IN2(n557), .Q(n555) );
  OR2X1 U701 ( .IN1(n558), .IN2(n559), .Q(n557) );
  AND2X1 U702 ( .IN1(n779), .IN2(n530), .Q(n559) );
  AND2X1 U703 ( .IN1(n778), .IN2(n526), .Q(n558) );
  AND2X1 U704 ( .IN1(xmit_dataH_3_), .IN2(n538), .Q(n556) );
  AND2X1 U705 ( .IN1(n780), .IN2(test_se), .Q(n553) );
  OR2X1 U706 ( .IN1(n560), .IN2(n561), .Q(n168) );
  AND2X1 U707 ( .IN1(n562), .IN2(n473), .Q(n561) );
  OR2X1 U708 ( .IN1(n563), .IN2(n564), .Q(n562) );
  OR2X1 U709 ( .IN1(n565), .IN2(n566), .Q(n564) );
  AND2X1 U710 ( .IN1(n780), .IN2(n530), .Q(n566) );
  AND2X1 U711 ( .IN1(n779), .IN2(n526), .Q(n565) );
  AND2X1 U712 ( .IN1(xmit_dataH_2_), .IN2(n538), .Q(n563) );
  AND2X1 U713 ( .IN1(n781), .IN2(test_se), .Q(n560) );
  OR2X1 U714 ( .IN1(n567), .IN2(n568), .Q(n167) );
  AND2X1 U715 ( .IN1(n569), .IN2(n473), .Q(n568) );
  OR2X1 U716 ( .IN1(n570), .IN2(n571), .Q(n569) );
  OR2X1 U717 ( .IN1(n572), .IN2(n573), .Q(n571) );
  AND2X1 U718 ( .IN1(n781), .IN2(n530), .Q(n573) );
  AND2X1 U719 ( .IN1(n780), .IN2(n526), .Q(n572) );
  AND2X1 U720 ( .IN1(xmit_dataH_1_), .IN2(n538), .Q(n570) );
  AND2X1 U721 ( .IN1(test_se), .IN2(n457), .Q(n567) );
  OR2X1 U722 ( .IN1(n574), .IN2(n575), .Q(n166) );
  AND2X1 U723 ( .IN1(n576), .IN2(n473), .Q(n575) );
  OR2X1 U724 ( .IN1(n577), .IN2(n578), .Q(n576) );
  INVX0 U725 ( .INP(n514), .ZN(n578) );
  OR2X1 U726 ( .IN1(iXMIT_state_1_), .IN2(n579), .Q(n514) );
  OR2X1 U727 ( .IN1(xmitH), .IN2(iXMIT_state_2_), .Q(n579) );
  AND2X1 U728 ( .IN1(n481), .IN2(n465), .Q(n577) );
  AND2X1 U729 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n574) );
  OR2X1 U730 ( .IN1(n580), .IN2(n581), .Q(n164) );
  OR2X1 U731 ( .IN1(n582), .IN2(n583), .Q(n581) );
  AND2X1 U732 ( .IN1(n584), .IN2(n245), .Q(n583) );
  AND2X1 U733 ( .IN1(n585), .IN2(n473), .Q(n584) );
  OR2X1 U734 ( .IN1(n586), .IN2(n459), .Q(n585) );
  AND2X1 U735 ( .IN1(n587), .IN2(iRECEIVER_state_1_), .Q(n586) );
  AND2X1 U736 ( .IN1(n588), .IN2(iRECEIVER_state_0_), .Q(n582) );
  OR2X1 U737 ( .IN1(test_se), .IN2(n589), .Q(n588) );
  OR2X1 U738 ( .IN1(n590), .IN2(n591), .Q(n589) );
  AND2X1 U739 ( .IN1(n592), .IN2(n241), .Q(n591) );
  AND2X1 U740 ( .IN1(n238), .IN2(n459), .Q(n592) );
  AND2X1 U741 ( .IN1(n593), .IN2(iRECEIVER_state_1_), .Q(n590) );
  OR2X1 U742 ( .IN1(n594), .IN2(n595), .Q(n163) );
  AND2X1 U743 ( .IN1(n596), .IN2(n473), .Q(n595) );
  OR2X1 U744 ( .IN1(iRECEIVER_state_2_), .IN2(n597), .Q(n596) );
  OR2X1 U745 ( .IN1(n598), .IN2(n599), .Q(n597) );
  AND2X1 U746 ( .IN1(n600), .IN2(iRECEIVER_state_1_), .Q(n599) );
  OR2X1 U747 ( .IN1(n601), .IN2(n602), .Q(n600) );
  AND2X1 U748 ( .IN1(n603), .IN2(iRECEIVER_state_0_), .Q(n601) );
  OR2X1 U749 ( .IN1(n604), .IN2(n593), .Q(n603) );
  INVX0 U750 ( .INP(n605), .ZN(n593) );
  AND2X1 U751 ( .IN1(n606), .IN2(n607), .Q(n604) );
  AND2X1 U752 ( .IN1(n456), .IN2(n453), .Q(n607) );
  AND2X1 U753 ( .IN1(n784), .IN2(n461), .Q(n606) );
  AND2X1 U754 ( .IN1(n241), .IN2(n783), .Q(n598) );
  AND2X1 U755 ( .IN1(n784), .IN2(test_se), .Q(n594) );
  OR2X1 U756 ( .IN1(n608), .IN2(n609), .Q(n162) );
  AND2X1 U757 ( .IN1(test_si), .IN2(test_se), .Q(n609) );
  AND2X1 U758 ( .IN1(iRECEIVER_N20), .IN2(n473), .Q(n608) );
  OR2X1 U759 ( .IN1(n610), .IN2(n611), .Q(n161) );
  AND2X1 U760 ( .IN1(iRECEIVER_N21), .IN2(n473), .Q(n611) );
  AND2X1 U761 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n610) );
  OR2X1 U762 ( .IN1(n612), .IN2(n613), .Q(n160) );
  AND2X1 U763 ( .IN1(iRECEIVER_N22), .IN2(n473), .Q(n613) );
  AND2X1 U764 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n612) );
  OR2X1 U765 ( .IN1(n614), .IN2(n615), .Q(n159) );
  AND2X1 U766 ( .IN1(n797), .IN2(test_se), .Q(n615) );
  AND2X1 U767 ( .IN1(iRECEIVER_N23), .IN2(n473), .Q(n614) );
  OR2X1 U768 ( .IN1(n616), .IN2(iRECEIVER_next_state_2_), .Q(n157) );
  AND2X1 U769 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n616) );
  OR2X1 U770 ( .IN1(n617), .IN2(n618), .Q(n156) );
  AND2X1 U771 ( .IN1(n619), .IN2(n473), .Q(n618) );
  OR2X1 U772 ( .IN1(n620), .IN2(n621), .Q(n619) );
  AND2X1 U773 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n620)
         );
  AND2X1 U774 ( .IN1(n782), .IN2(test_se), .Q(n617) );
  OR2X1 U775 ( .IN1(n622), .IN2(n623), .Q(n155) );
  OR2X1 U776 ( .IN1(n624), .IN2(n625), .Q(n623) );
  AND2X1 U777 ( .IN1(n580), .IN2(n783), .Q(n625) );
  AND2X1 U778 ( .IN1(rec_dataH_rec_7), .IN2(n626), .Q(n624) );
  AND2X1 U779 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n622) );
  OR2X1 U780 ( .IN1(n627), .IN2(n628), .Q(n154) );
  AND2X1 U781 ( .IN1(rec_dataH_temp_6), .IN2(test_se), .Q(n628) );
  AND2X1 U782 ( .IN1(rec_dataH_rec_7), .IN2(n473), .Q(n627) );
  OR2X1 U783 ( .IN1(n629), .IN2(n630), .Q(n153) );
  AND2X1 U784 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n630) );
  AND2X1 U785 ( .IN1(test_so), .IN2(n473), .Q(n629) );
  OR2X1 U786 ( .IN1(n631), .IN2(n632), .Q(n152) );
  OR2X1 U787 ( .IN1(n633), .IN2(n634), .Q(n632) );
  AND2X1 U788 ( .IN1(n580), .IN2(rec_dataH_rec_7), .Q(n634) );
  AND2X1 U789 ( .IN1(rec_dataH_rec_6), .IN2(n626), .Q(n633) );
  AND2X1 U790 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n631) );
  OR2X1 U791 ( .IN1(n635), .IN2(n636), .Q(n150) );
  AND2X1 U792 ( .IN1(rec_dataH_temp_5), .IN2(test_se), .Q(n636) );
  AND2X1 U793 ( .IN1(rec_dataH_rec_6), .IN2(n473), .Q(n635) );
  OR2X1 U794 ( .IN1(n637), .IN2(n638), .Q(n149) );
  AND2X1 U795 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n638) );
  AND2X1 U796 ( .IN1(rec_dataH_temp_6), .IN2(n473), .Q(n637) );
  OR2X1 U797 ( .IN1(n639), .IN2(n640), .Q(n148) );
  OR2X1 U798 ( .IN1(n641), .IN2(n642), .Q(n640) );
  AND2X1 U799 ( .IN1(rec_dataH_rec_6), .IN2(n580), .Q(n642) );
  AND2X1 U800 ( .IN1(rec_dataH_rec_5), .IN2(n626), .Q(n641) );
  AND2X1 U801 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n639) );
  OR2X1 U802 ( .IN1(n643), .IN2(n644), .Q(n147) );
  AND2X1 U803 ( .IN1(rec_dataH_temp_4), .IN2(test_se), .Q(n644) );
  AND2X1 U804 ( .IN1(rec_dataH_rec_5), .IN2(n473), .Q(n643) );
  OR2X1 U805 ( .IN1(n645), .IN2(n646), .Q(n146) );
  AND2X1 U806 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n646) );
  AND2X1 U807 ( .IN1(rec_dataH_temp_5), .IN2(n473), .Q(n645) );
  OR2X1 U808 ( .IN1(n647), .IN2(n648), .Q(n145) );
  OR2X1 U809 ( .IN1(n649), .IN2(n650), .Q(n648) );
  AND2X1 U810 ( .IN1(rec_dataH_rec_5), .IN2(n580), .Q(n650) );
  AND2X1 U811 ( .IN1(rec_dataH_rec_4), .IN2(n626), .Q(n649) );
  AND2X1 U812 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n647) );
  OR2X1 U813 ( .IN1(n651), .IN2(n652), .Q(n143) );
  AND2X1 U814 ( .IN1(rec_dataH_temp_3), .IN2(test_se), .Q(n652) );
  AND2X1 U815 ( .IN1(rec_dataH_rec_4), .IN2(n473), .Q(n651) );
  OR2X1 U816 ( .IN1(n653), .IN2(n654), .Q(n142) );
  AND2X1 U817 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n654) );
  AND2X1 U818 ( .IN1(rec_dataH_temp_4), .IN2(n473), .Q(n653) );
  OR2X1 U819 ( .IN1(n655), .IN2(n656), .Q(n141) );
  OR2X1 U820 ( .IN1(n657), .IN2(n658), .Q(n656) );
  AND2X1 U821 ( .IN1(rec_dataH_rec_4), .IN2(n580), .Q(n658) );
  AND2X1 U822 ( .IN1(rec_dataH_rec_3), .IN2(n626), .Q(n657) );
  AND2X1 U823 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n655) );
  OR2X1 U824 ( .IN1(n659), .IN2(n660), .Q(n140) );
  AND2X1 U825 ( .IN1(rec_dataH_temp_2), .IN2(test_se), .Q(n660) );
  AND2X1 U826 ( .IN1(rec_dataH_rec_3), .IN2(n473), .Q(n659) );
  OR2X1 U827 ( .IN1(n661), .IN2(n662), .Q(n139) );
  AND2X1 U828 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n662) );
  AND2X1 U829 ( .IN1(rec_dataH_temp_3), .IN2(n473), .Q(n661) );
  OR2X1 U830 ( .IN1(n663), .IN2(n664), .Q(n138) );
  OR2X1 U831 ( .IN1(n665), .IN2(n666), .Q(n664) );
  AND2X1 U832 ( .IN1(rec_dataH_rec_3), .IN2(n580), .Q(n666) );
  AND2X1 U833 ( .IN1(rec_dataH_rec_2), .IN2(n626), .Q(n665) );
  AND2X1 U834 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n663) );
  OR2X1 U835 ( .IN1(n667), .IN2(n668), .Q(n136) );
  AND2X1 U836 ( .IN1(rec_dataH_temp_1), .IN2(test_se), .Q(n668) );
  AND2X1 U837 ( .IN1(rec_dataH_rec_2), .IN2(n473), .Q(n667) );
  OR2X1 U838 ( .IN1(n669), .IN2(n670), .Q(n135) );
  AND2X1 U839 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n670) );
  AND2X1 U840 ( .IN1(rec_dataH_temp_2), .IN2(n473), .Q(n669) );
  OR2X1 U841 ( .IN1(n671), .IN2(n672), .Q(n134) );
  OR2X1 U842 ( .IN1(n673), .IN2(n674), .Q(n672) );
  AND2X1 U843 ( .IN1(rec_dataH_rec_2), .IN2(n580), .Q(n674) );
  AND2X1 U844 ( .IN1(rec_dataH_rec_1), .IN2(n626), .Q(n673) );
  AND2X1 U845 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .Q(n671) );
  OR2X1 U846 ( .IN1(n675), .IN2(n676), .Q(n133) );
  AND2X1 U847 ( .IN1(rec_dataH_temp_0), .IN2(test_se), .Q(n676) );
  AND2X1 U848 ( .IN1(rec_dataH_rec_1), .IN2(n473), .Q(n675) );
  OR2X1 U849 ( .IN1(n677), .IN2(n678), .Q(n132) );
  AND2X1 U850 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n678) );
  AND2X1 U851 ( .IN1(rec_dataH_temp_1), .IN2(n473), .Q(n677) );
  OR2X1 U852 ( .IN1(n679), .IN2(n680), .Q(n131) );
  OR2X1 U853 ( .IN1(n681), .IN2(n682), .Q(n680) );
  AND2X1 U854 ( .IN1(rec_dataH_rec_1), .IN2(n580), .Q(n682) );
  AND2X1 U855 ( .IN1(rec_dataH_rec_0), .IN2(n626), .Q(n681) );
  AND2X1 U856 ( .IN1(n796), .IN2(test_se), .Q(n679) );
  OR2X1 U857 ( .IN1(n683), .IN2(n684), .Q(n129) );
  AND2X1 U858 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n684) );
  AND2X1 U859 ( .IN1(rec_dataH_rec_0), .IN2(n473), .Q(n683) );
  OR2X1 U860 ( .IN1(n685), .IN2(n686), .Q(n128) );
  AND2X1 U861 ( .IN1(xmit_doneH_temp), .IN2(test_se), .Q(n686) );
  AND2X1 U862 ( .IN1(rec_dataH_temp_0), .IN2(n473), .Q(n685) );
  OR2X1 U863 ( .IN1(n687), .IN2(n688), .Q(n127) );
  AND2X1 U864 ( .IN1(n784), .IN2(n689), .Q(n688) );
  OR2X1 U865 ( .IN1(n690), .IN2(n691), .Q(n689) );
  AND2X1 U866 ( .IN1(n580), .IN2(n692), .Q(n690) );
  OR2X1 U867 ( .IN1(n453), .IN2(n693), .Q(n692) );
  AND2X1 U868 ( .IN1(n793), .IN2(n694), .Q(n687) );
  OR2X1 U869 ( .IN1(n695), .IN2(test_se), .Q(n694) );
  AND2X1 U870 ( .IN1(n696), .IN2(n580), .Q(n695) );
  INVX0 U871 ( .INP(n697), .ZN(n696) );
  OR2X1 U872 ( .IN1(n693), .IN2(n784), .Q(n697) );
  OR2X1 U873 ( .IN1(n698), .IN2(n699), .Q(n126) );
  OR2X1 U874 ( .IN1(n700), .IN2(n701), .Q(n699) );
  AND2X1 U875 ( .IN1(n691), .IN2(n794), .Q(n701) );
  AND2X1 U876 ( .IN1(n580), .IN2(n456), .Q(n700) );
  AND2X1 U877 ( .IN1(test_se), .IN2(rec_readyH), .Q(n698) );
  OR2X1 U878 ( .IN1(n702), .IN2(n703), .Q(n125) );
  OR2X1 U879 ( .IN1(n704), .IN2(n705), .Q(n703) );
  AND2X1 U880 ( .IN1(n691), .IN2(n795), .Q(n705) );
  AND2X1 U881 ( .IN1(n580), .IN2(iRECEIVER_N26), .Q(n704) );
  AND2X1 U882 ( .IN1(test_se), .IN2(n794), .Q(n702) );
  OR2X1 U883 ( .IN1(n706), .IN2(n707), .Q(n124) );
  OR2X1 U884 ( .IN1(n708), .IN2(n709), .Q(n707) );
  AND2X1 U885 ( .IN1(n691), .IN2(n793), .Q(n709) );
  AND2X1 U886 ( .IN1(n710), .IN2(n626), .Q(n691) );
  AND2X1 U887 ( .IN1(n473), .IN2(n711), .Q(n626) );
  INVX0 U888 ( .INP(n712), .ZN(n711) );
  INVX0 U889 ( .INP(n621), .ZN(n710) );
  AND2X1 U890 ( .IN1(n241), .IN2(n713), .Q(n621) );
  AND2X1 U891 ( .IN1(n783), .IN2(n238), .Q(n713) );
  AND2X1 U892 ( .IN1(n580), .IN2(n41), .Q(n708) );
  OR2X1 U893 ( .IN1(n714), .IN2(n715), .Q(n41) );
  AND2X1 U894 ( .IN1(n716), .IN2(n453), .Q(n715) );
  AND2X1 U895 ( .IN1(n793), .IN2(n693), .Q(n714) );
  INVX0 U896 ( .INP(n716), .ZN(n693) );
  AND2X1 U897 ( .IN1(n795), .IN2(n794), .Q(n716) );
  AND2X1 U898 ( .IN1(n473), .IN2(n712), .Q(n580) );
  AND2X1 U899 ( .IN1(iRECEIVER_state_2_), .IN2(n245), .Q(n712) );
  AND2X1 U900 ( .IN1(test_se), .IN2(n795), .Q(n706) );
  OR2X1 U901 ( .IN1(n717), .IN2(n718), .Q(n122) );
  AND2X1 U902 ( .IN1(test_se), .IN2(n790), .Q(n718) );
  AND2X1 U903 ( .IN1(iXMIT_N29), .IN2(n473), .Q(n717) );
  OR2X1 U904 ( .IN1(n719), .IN2(n720), .Q(n121) );
  AND2X1 U905 ( .IN1(iXMIT_N26), .IN2(n473), .Q(n720) );
  AND2X1 U906 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n719) );
  OR2X1 U907 ( .IN1(n721), .IN2(n722), .Q(n120) );
  AND2X1 U908 ( .IN1(test_se), .IN2(n792), .Q(n722) );
  AND2X1 U909 ( .IN1(iXMIT_N27), .IN2(n473), .Q(n721) );
  OR2X1 U910 ( .IN1(n723), .IN2(n724), .Q(n119) );
  AND2X1 U911 ( .IN1(n725), .IN2(n473), .Q(n724) );
  OR2X1 U912 ( .IN1(n726), .IN2(n727), .Q(n725) );
  OR2X1 U913 ( .IN1(n728), .IN2(n729), .Q(n727) );
  AND2X1 U914 ( .IN1(n530), .IN2(n457), .Q(n729) );
  INVX0 U915 ( .INP(n495), .ZN(n530) );
  AND2X1 U916 ( .IN1(n781), .IN2(n526), .Q(n728) );
  AND2X1 U917 ( .IN1(n730), .IN2(n495), .Q(n526) );
  OR2X1 U918 ( .IN1(n731), .IN2(n538), .Q(n495) );
  AND2X1 U919 ( .IN1(n239), .IN2(iXMIT_state_2_), .Q(n731) );
  INVX0 U920 ( .INP(n538), .ZN(n730) );
  AND2X1 U921 ( .IN1(xmit_dataH_0_), .IN2(n538), .Q(n726) );
  AND2X1 U922 ( .IN1(xmitH), .IN2(n463), .Q(n538) );
  AND2X1 U923 ( .IN1(n242), .IN2(n246), .Q(n463) );
  AND2X1 U924 ( .IN1(test_se), .IN2(iXMIT_state_2_), .Q(n723) );
  OR2X1 U925 ( .IN1(n732), .IN2(n733), .Q(n118) );
  AND2X1 U926 ( .IN1(n783), .IN2(test_se), .Q(n733) );
  AND2X1 U927 ( .IN1(uart_REC_dataH), .IN2(n473), .Q(n732) );
  OR2X1 U928 ( .IN1(n734), .IN2(n735), .Q(n117) );
  AND2X1 U929 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n735) );
  AND2X1 U930 ( .IN1(n782), .IN2(n473), .Q(n734) );
  INVX0 U931 ( .INP(test_se), .ZN(n473) );
  OR2X1 U932 ( .IN1(n736), .IN2(n737), .Q(iXMIT_N46) );
  INVX0 U933 ( .INP(n738), .ZN(n737) );
  OR2X1 U934 ( .IN1(n739), .IN2(n785), .Q(n738) );
  AND2X1 U935 ( .IN1(n785), .IN2(n739), .Q(n736) );
  AND2X1 U936 ( .IN1(n739), .IN2(n740), .Q(iXMIT_N45) );
  OR2X1 U937 ( .IN1(n786), .IN2(n741), .Q(n740) );
  AND2X1 U938 ( .IN1(n787), .IN2(n788), .Q(n741) );
  OR2X1 U939 ( .IN1(n458), .IN2(n742), .Q(n739) );
  OR2X1 U940 ( .IN1(n452), .IN2(n454), .Q(n742) );
  OR2X1 U941 ( .IN1(n743), .IN2(n744), .Q(iXMIT_N44) );
  AND2X1 U942 ( .IN1(n788), .IN2(n452), .Q(n744) );
  AND2X1 U943 ( .IN1(n787), .IN2(n454), .Q(n743) );
  AND2X1 U944 ( .IN1(n745), .IN2(iXMIT_N25), .Q(iXMIT_N29) );
  AND2X1 U945 ( .IN1(n745), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U946 ( .IN1(n746), .IN2(n747), .Q(iXMIT_N27) );
  AND2X1 U947 ( .IN1(iXMIT_N26), .IN2(n791), .Q(n747) );
  AND2X1 U948 ( .IN1(n748), .IN2(n460), .Q(n746) );
  AND2X1 U949 ( .IN1(n792), .IN2(n745), .Q(n748) );
  AND2X1 U950 ( .IN1(n462), .IN2(n745), .Q(iXMIT_N26) );
  OR2X1 U951 ( .IN1(n465), .IN2(n494), .Q(n745) );
  AND2X1 U952 ( .IN1(n490), .IN2(iXMIT_state_1_), .Q(n494) );
  OR2X1 U953 ( .IN1(n239), .IN2(n520), .Q(n490) );
  OR2X1 U954 ( .IN1(n749), .IN2(n750), .Q(n520) );
  INVX0 U955 ( .INP(n751), .ZN(n750) );
  AND2X1 U956 ( .IN1(n790), .IN2(n789), .Q(n751) );
  OR2X1 U957 ( .IN1(n792), .IN2(n460), .Q(n749) );
  AND2X1 U958 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .Q(n465) );
  AND2X1 U959 ( .IN1(n484), .IN2(n752), .Q(iXMIT_N25) );
  OR2X1 U960 ( .IN1(n789), .IN2(n753), .Q(n752) );
  INVX0 U961 ( .INP(n481), .ZN(n484) );
  AND2X1 U962 ( .IN1(n753), .IN2(n789), .Q(n481) );
  AND2X1 U963 ( .IN1(n754), .IN2(n755), .Q(iXMIT_N24) );
  OR2X1 U964 ( .IN1(n790), .IN2(n756), .Q(n755) );
  INVX0 U965 ( .INP(n753), .ZN(n754) );
  AND2X1 U966 ( .IN1(n790), .IN2(n756), .Q(n753) );
  AND2X1 U967 ( .IN1(n792), .IN2(n791), .Q(n756) );
  AND2X1 U968 ( .IN1(n605), .IN2(n757), .Q(iRECEIVER_next_state_2_) );
  AND2X1 U969 ( .IN1(iRECEIVER_state_0_), .IN2(iRECEIVER_state_1_), .Q(n757)
         );
  OR2X1 U970 ( .IN1(n758), .IN2(n759), .Q(iRECEIVER_N26) );
  AND2X1 U971 ( .IN1(n795), .IN2(n456), .Q(n759) );
  AND2X1 U972 ( .IN1(n794), .IN2(n461), .Q(n758) );
  AND2X1 U973 ( .IN1(iRECEIVER_N19), .IN2(n760), .Q(iRECEIVER_N23) );
  AND2X1 U974 ( .IN1(n760), .IN2(iRECEIVER_N18), .Q(iRECEIVER_N22) );
  AND2X1 U975 ( .IN1(iRECEIVER_N17), .IN2(n760), .Q(iRECEIVER_N21) );
  AND2X1 U976 ( .IN1(n255), .IN2(n760), .Q(iRECEIVER_N20) );
  INVX0 U977 ( .INP(n761), .ZN(n760) );
  OR2X1 U978 ( .IN1(n762), .IN2(n763), .Q(n761) );
  OR2X1 U979 ( .IN1(n241), .IN2(iRECEIVER_state_2_), .Q(n763) );
  OR2X1 U980 ( .IN1(n764), .IN2(n765), .Q(n762) );
  AND2X1 U981 ( .IN1(n602), .IN2(n245), .Q(n765) );
  INVX0 U982 ( .INP(n587), .ZN(n602) );
  OR2X1 U983 ( .IN1(n766), .IN2(n767), .Q(n587) );
  OR2X1 U984 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(n455), .Q(n767) );
  OR2X1 U985 ( .IN1(n796), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n766) );
  AND2X1 U986 ( .IN1(n605), .IN2(iRECEIVER_state_0_), .Q(n764) );
  AND2X1 U987 ( .IN1(n768), .IN2(n769), .Q(n605) );
  AND2X1 U988 ( .IN1(n797), .IN2(n796), .Q(n769) );
  OR2X1 U989 ( .IN1(n770), .IN2(n771), .Q(iRECEIVER_N19) );
  INVX0 U990 ( .INP(n772), .ZN(n771) );
  OR2X1 U991 ( .IN1(n773), .IN2(n796), .Q(n772) );
  AND2X1 U992 ( .IN1(n796), .IN2(n773), .Q(n770) );
  AND2X1 U993 ( .IN1(n773), .IN2(n774), .Q(iRECEIVER_N18) );
  OR2X1 U994 ( .IN1(n797), .IN2(n775), .Q(n774) );
  AND2X1 U995 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .Q(n775) );
  OR2X1 U996 ( .IN1(n455), .IN2(n776), .Q(n773) );
  OR2X1 U997 ( .IN1(n255), .IN2(n244), .Q(n776) );
  OR2X1 U998 ( .IN1(n768), .IN2(n777), .Q(iRECEIVER_N17) );
  AND2X1 U999 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n777) );
  AND2X1 U1000 ( .IN1(n255), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n768) );
endmodule

