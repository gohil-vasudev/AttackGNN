module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n888_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n716_, new_n701_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n890_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n854_, new_n447_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n559_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n352_, new_n931_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n519_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n435_, new_n776_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n412_, new_n607_, new_n904_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n336_, new_n377_, new_n247_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n202_, keyIn_0_55 );
xnor g001 ( new_n203_, N65, N69 );
xor g002 ( new_n204_, new_n203_, keyIn_0_8 );
xnor g003 ( new_n205_, N73, N77 );
xnor g004 ( new_n206_, new_n205_, keyIn_0_9 );
xnor g005 ( new_n207_, new_n204_, new_n206_ );
xnor g006 ( new_n208_, new_n207_, keyIn_0_32 );
xnor g007 ( new_n209_, N81, N85 );
xnor g008 ( new_n210_, new_n209_, keyIn_0_10 );
xnor g009 ( new_n211_, N89, N93 );
xnor g010 ( new_n212_, new_n211_, keyIn_0_11 );
xnor g011 ( new_n213_, new_n210_, new_n212_ );
xnor g012 ( new_n214_, new_n213_, keyIn_0_33 );
xnor g013 ( new_n215_, new_n208_, new_n214_ );
xnor g014 ( new_n216_, new_n215_, keyIn_0_43 );
nand g015 ( new_n217_, N129, N137 );
xor g016 ( new_n218_, new_n216_, new_n217_ );
xnor g017 ( new_n219_, new_n218_, keyIn_0_47 );
xnor g018 ( new_n220_, N1, N17 );
xnor g019 ( new_n221_, N33, N49 );
xnor g020 ( new_n222_, new_n220_, new_n221_ );
not g021 ( new_n223_, new_n222_ );
nand g022 ( new_n224_, new_n219_, new_n223_ );
nand g023 ( new_n225_, new_n218_, keyIn_0_47 );
or g024 ( new_n226_, new_n218_, keyIn_0_47 );
nand g025 ( new_n227_, new_n226_, new_n225_, new_n222_ );
nand g026 ( new_n228_, new_n224_, new_n227_ );
nand g027 ( new_n229_, new_n228_, new_n202_ );
nand g028 ( new_n230_, new_n224_, new_n227_, keyIn_0_55 );
and g029 ( new_n231_, new_n229_, new_n230_ );
nand g030 ( new_n232_, new_n229_, new_n230_ );
xor g031 ( new_n233_, N97, N101 );
xnor g032 ( new_n234_, new_n233_, keyIn_0_12 );
not g033 ( new_n235_, keyIn_0_13 );
xnor g034 ( new_n236_, N105, N109 );
xnor g035 ( new_n237_, new_n236_, new_n235_ );
xnor g036 ( new_n238_, new_n234_, new_n237_ );
xnor g037 ( new_n239_, new_n238_, keyIn_0_34 );
xnor g038 ( new_n240_, new_n208_, new_n239_ );
xnor g039 ( new_n241_, new_n240_, keyIn_0_45 );
nand g040 ( new_n242_, N131, N137 );
xor g041 ( new_n243_, new_n242_, keyIn_0_16 );
not g042 ( new_n244_, new_n243_ );
xnor g043 ( new_n245_, new_n241_, new_n244_ );
nand g044 ( new_n246_, new_n245_, keyIn_0_49 );
or g045 ( new_n247_, new_n245_, keyIn_0_49 );
xor g046 ( new_n248_, N9, N25 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_21 );
xnor g048 ( new_n250_, N41, N57 );
xnor g049 ( new_n251_, new_n250_, keyIn_0_22 );
xnor g050 ( new_n252_, new_n249_, new_n251_ );
xor g051 ( new_n253_, new_n252_, keyIn_0_36 );
nand g052 ( new_n254_, new_n247_, new_n246_, new_n253_ );
nand g053 ( new_n255_, new_n247_, new_n246_ );
not g054 ( new_n256_, new_n253_ );
nand g055 ( new_n257_, new_n255_, new_n256_ );
nand g056 ( new_n258_, new_n257_, new_n254_ );
nand g057 ( new_n259_, new_n258_, keyIn_0_57 );
not g058 ( new_n260_, keyIn_0_57 );
nand g059 ( new_n261_, new_n257_, new_n260_, new_n254_ );
nand g060 ( new_n262_, new_n259_, new_n261_ );
not g061 ( new_n263_, keyIn_0_56 );
not g062 ( new_n264_, keyIn_0_35 );
not g063 ( new_n265_, keyIn_0_15 );
xnor g064 ( new_n266_, N121, N125 );
xnor g065 ( new_n267_, new_n266_, new_n265_ );
xnor g066 ( new_n268_, N113, N117 );
xnor g067 ( new_n269_, new_n268_, keyIn_0_14 );
xnor g068 ( new_n270_, new_n267_, new_n269_ );
xnor g069 ( new_n271_, new_n270_, new_n264_ );
xnor g070 ( new_n272_, new_n239_, new_n271_ );
xnor g071 ( new_n273_, new_n272_, keyIn_0_44 );
and g072 ( new_n274_, N130, N137 );
xnor g073 ( new_n275_, new_n273_, new_n274_ );
xnor g074 ( new_n276_, new_n275_, keyIn_0_48 );
xnor g075 ( new_n277_, N5, N21 );
xnor g076 ( new_n278_, N37, N53 );
xnor g077 ( new_n279_, new_n277_, new_n278_ );
not g078 ( new_n280_, new_n279_ );
nand g079 ( new_n281_, new_n276_, new_n280_ );
nand g080 ( new_n282_, new_n275_, keyIn_0_48 );
or g081 ( new_n283_, new_n275_, keyIn_0_48 );
nand g082 ( new_n284_, new_n283_, new_n282_, new_n279_ );
nand g083 ( new_n285_, new_n281_, new_n284_ );
nand g084 ( new_n286_, new_n285_, new_n263_ );
nand g085 ( new_n287_, new_n281_, new_n284_, keyIn_0_56 );
and g086 ( new_n288_, new_n286_, new_n287_ );
not g087 ( new_n289_, keyIn_0_50 );
xnor g088 ( new_n290_, new_n214_, new_n271_ );
xnor g089 ( new_n291_, new_n290_, keyIn_0_46 );
nand g090 ( new_n292_, N132, N137 );
xnor g091 ( new_n293_, new_n291_, new_n292_ );
nand g092 ( new_n294_, new_n293_, new_n289_ );
not g093 ( new_n295_, new_n292_ );
xnor g094 ( new_n296_, new_n291_, new_n295_ );
nand g095 ( new_n297_, new_n296_, keyIn_0_50 );
nand g096 ( new_n298_, new_n294_, new_n297_ );
xnor g097 ( new_n299_, N13, N29 );
xnor g098 ( new_n300_, new_n299_, keyIn_0_23 );
xnor g099 ( new_n301_, N45, N61 );
xnor g100 ( new_n302_, new_n300_, new_n301_ );
not g101 ( new_n303_, new_n302_ );
nand g102 ( new_n304_, new_n298_, new_n303_ );
nand g103 ( new_n305_, new_n294_, new_n297_, new_n302_ );
nand g104 ( new_n306_, new_n304_, keyIn_0_58, new_n305_ );
not g105 ( new_n307_, keyIn_0_58 );
nand g106 ( new_n308_, new_n304_, new_n305_ );
nand g107 ( new_n309_, new_n308_, new_n307_ );
nand g108 ( new_n310_, new_n309_, new_n306_ );
nand g109 ( new_n311_, new_n288_, new_n262_, new_n310_ );
and g110 ( new_n312_, new_n259_, new_n261_ );
nand g111 ( new_n313_, new_n310_, new_n286_, new_n287_ );
nand g112 ( new_n314_, new_n312_, new_n313_ );
nand g113 ( new_n315_, new_n286_, new_n287_ );
not g114 ( new_n316_, new_n310_ );
nand g115 ( new_n317_, new_n316_, new_n315_ );
nand g116 ( new_n318_, new_n314_, new_n311_, new_n232_, new_n317_ );
nor g117 ( new_n319_, new_n232_, new_n315_ );
nand g118 ( new_n320_, new_n259_, keyIn_0_63, new_n261_ );
not g119 ( new_n321_, keyIn_0_63 );
nand g120 ( new_n322_, new_n262_, new_n321_ );
nand g121 ( new_n323_, new_n319_, new_n322_, new_n310_, new_n320_ );
nand g122 ( new_n324_, new_n318_, new_n323_ );
not g123 ( new_n325_, keyIn_0_59 );
not g124 ( new_n326_, keyIn_0_39 );
not g125 ( new_n327_, keyIn_0_2 );
not g126 ( new_n328_, N17 );
not g127 ( new_n329_, N21 );
nand g128 ( new_n330_, new_n328_, new_n329_ );
nand g129 ( new_n331_, N17, N21 );
nand g130 ( new_n332_, new_n330_, new_n331_ );
nand g131 ( new_n333_, new_n332_, new_n327_ );
nand g132 ( new_n334_, new_n330_, keyIn_0_2, new_n331_ );
nand g133 ( new_n335_, new_n333_, new_n334_ );
or g134 ( new_n336_, N25, N29 );
nand g135 ( new_n337_, N25, N29 );
nand g136 ( new_n338_, new_n336_, new_n337_ );
nand g137 ( new_n339_, new_n338_, keyIn_0_3 );
not g138 ( new_n340_, keyIn_0_3 );
nand g139 ( new_n341_, new_n336_, new_n340_, new_n337_ );
nand g140 ( new_n342_, new_n339_, new_n341_ );
nand g141 ( new_n343_, new_n342_, new_n335_ );
nand g142 ( new_n344_, new_n339_, new_n333_, new_n334_, new_n341_ );
nand g143 ( new_n345_, new_n343_, new_n344_ );
nand g144 ( new_n346_, new_n345_, keyIn_0_29 );
not g145 ( new_n347_, keyIn_0_29 );
nand g146 ( new_n348_, new_n343_, new_n347_, new_n344_ );
nand g147 ( new_n349_, new_n346_, new_n348_ );
not g148 ( new_n350_, keyIn_0_0 );
or g149 ( new_n351_, N1, N5 );
nand g150 ( new_n352_, N1, N5 );
nand g151 ( new_n353_, new_n351_, new_n350_, new_n352_ );
nand g152 ( new_n354_, new_n351_, new_n352_ );
nand g153 ( new_n355_, new_n354_, keyIn_0_0 );
nand g154 ( new_n356_, new_n355_, new_n353_ );
not g155 ( new_n357_, keyIn_0_1 );
or g156 ( new_n358_, N9, N13 );
nand g157 ( new_n359_, N9, N13 );
nand g158 ( new_n360_, new_n358_, new_n357_, new_n359_ );
nand g159 ( new_n361_, new_n358_, new_n359_ );
nand g160 ( new_n362_, new_n361_, keyIn_0_1 );
nand g161 ( new_n363_, new_n362_, new_n360_ );
nand g162 ( new_n364_, new_n356_, new_n363_ );
nand g163 ( new_n365_, new_n355_, new_n362_, new_n353_, new_n360_ );
nand g164 ( new_n366_, new_n364_, new_n365_ );
nand g165 ( new_n367_, new_n366_, keyIn_0_28 );
not g166 ( new_n368_, keyIn_0_28 );
nand g167 ( new_n369_, new_n364_, new_n368_, new_n365_ );
nand g168 ( new_n370_, new_n367_, new_n369_ );
nand g169 ( new_n371_, new_n370_, new_n349_ );
nand g170 ( new_n372_, new_n367_, new_n346_, new_n348_, new_n369_ );
nand g171 ( new_n373_, new_n371_, new_n326_, new_n372_ );
nand g172 ( new_n374_, new_n371_, new_n372_ );
nand g173 ( new_n375_, new_n374_, keyIn_0_39 );
nand g174 ( new_n376_, new_n375_, new_n373_ );
nand g175 ( new_n377_, N133, N137 );
xor g176 ( new_n378_, new_n377_, keyIn_0_17 );
not g177 ( new_n379_, new_n378_ );
nand g178 ( new_n380_, new_n376_, new_n379_ );
nand g179 ( new_n381_, new_n375_, new_n373_, new_n378_ );
nand g180 ( new_n382_, new_n380_, new_n381_ );
nand g181 ( new_n383_, new_n382_, keyIn_0_51 );
not g182 ( new_n384_, keyIn_0_51 );
nand g183 ( new_n385_, new_n380_, new_n384_, new_n381_ );
nand g184 ( new_n386_, new_n383_, new_n385_ );
xnor g185 ( new_n387_, N65, N81 );
xnor g186 ( new_n388_, N97, N113 );
xor g187 ( new_n389_, new_n387_, new_n388_ );
not g188 ( new_n390_, new_n389_ );
nand g189 ( new_n391_, new_n386_, new_n390_ );
nand g190 ( new_n392_, new_n383_, new_n385_, new_n389_ );
nand g191 ( new_n393_, new_n391_, new_n392_ );
nand g192 ( new_n394_, new_n393_, new_n325_ );
nand g193 ( new_n395_, new_n391_, keyIn_0_59, new_n392_ );
nand g194 ( new_n396_, new_n394_, new_n395_ );
not g195 ( new_n397_, keyIn_0_60 );
not g196 ( new_n398_, keyIn_0_31 );
or g197 ( new_n399_, N49, N53 );
nand g198 ( new_n400_, N49, N53 );
nand g199 ( new_n401_, new_n399_, new_n400_ );
nand g200 ( new_n402_, new_n401_, keyIn_0_6 );
not g201 ( new_n403_, keyIn_0_6 );
nand g202 ( new_n404_, new_n399_, new_n403_, new_n400_ );
nand g203 ( new_n405_, new_n402_, new_n404_ );
xnor g204 ( new_n406_, N57, N61 );
nand g205 ( new_n407_, new_n406_, keyIn_0_7 );
not g206 ( new_n408_, keyIn_0_7 );
or g207 ( new_n409_, N57, N61 );
nand g208 ( new_n410_, N57, N61 );
nand g209 ( new_n411_, new_n409_, new_n408_, new_n410_ );
nand g210 ( new_n412_, new_n407_, new_n411_ );
nand g211 ( new_n413_, new_n405_, new_n412_ );
nand g212 ( new_n414_, new_n402_, new_n407_, new_n404_, new_n411_ );
nand g213 ( new_n415_, new_n413_, new_n414_ );
nand g214 ( new_n416_, new_n415_, new_n398_ );
nand g215 ( new_n417_, new_n413_, keyIn_0_31, new_n414_ );
not g216 ( new_n418_, keyIn_0_30 );
not g217 ( new_n419_, N33 );
not g218 ( new_n420_, N37 );
nand g219 ( new_n421_, new_n419_, new_n420_ );
nand g220 ( new_n422_, N33, N37 );
nand g221 ( new_n423_, new_n421_, keyIn_0_4, new_n422_ );
not g222 ( new_n424_, keyIn_0_4 );
nand g223 ( new_n425_, new_n421_, new_n422_ );
nand g224 ( new_n426_, new_n425_, new_n424_ );
nand g225 ( new_n427_, new_n426_, new_n423_ );
xnor g226 ( new_n428_, N41, N45 );
nand g227 ( new_n429_, new_n428_, keyIn_0_5 );
not g228 ( new_n430_, keyIn_0_5 );
nand g229 ( new_n431_, N41, N45 );
not g230 ( new_n432_, N41 );
not g231 ( new_n433_, N45 );
nand g232 ( new_n434_, new_n432_, new_n433_ );
nand g233 ( new_n435_, new_n434_, new_n430_, new_n431_ );
nand g234 ( new_n436_, new_n429_, new_n435_ );
nand g235 ( new_n437_, new_n427_, new_n436_ );
nand g236 ( new_n438_, new_n426_, new_n429_, new_n423_, new_n435_ );
nand g237 ( new_n439_, new_n437_, new_n438_ );
nand g238 ( new_n440_, new_n439_, new_n418_ );
nand g239 ( new_n441_, new_n437_, keyIn_0_30, new_n438_ );
nand g240 ( new_n442_, new_n416_, new_n440_, new_n417_, new_n441_ );
nand g241 ( new_n443_, new_n416_, new_n417_ );
nand g242 ( new_n444_, new_n440_, new_n441_ );
nand g243 ( new_n445_, new_n443_, new_n444_ );
nand g244 ( new_n446_, new_n445_, new_n442_ );
nand g245 ( new_n447_, new_n446_, keyIn_0_40 );
not g246 ( new_n448_, keyIn_0_40 );
nand g247 ( new_n449_, new_n445_, new_n448_, new_n442_ );
nand g248 ( new_n450_, new_n447_, new_n449_ );
nand g249 ( new_n451_, N134, N137 );
xor g250 ( new_n452_, new_n451_, keyIn_0_18 );
not g251 ( new_n453_, new_n452_ );
nand g252 ( new_n454_, new_n450_, new_n453_ );
nand g253 ( new_n455_, new_n447_, new_n449_, new_n452_ );
nand g254 ( new_n456_, new_n454_, new_n455_ );
nand g255 ( new_n457_, new_n456_, keyIn_0_52 );
not g256 ( new_n458_, keyIn_0_52 );
nand g257 ( new_n459_, new_n454_, new_n458_, new_n455_ );
nand g258 ( new_n460_, new_n457_, new_n459_ );
xor g259 ( new_n461_, N69, N85 );
xnor g260 ( new_n462_, new_n461_, keyIn_0_24 );
xnor g261 ( new_n463_, N101, N117 );
xnor g262 ( new_n464_, new_n463_, keyIn_0_25 );
xnor g263 ( new_n465_, new_n462_, new_n464_ );
xor g264 ( new_n466_, new_n465_, keyIn_0_37 );
not g265 ( new_n467_, new_n466_ );
nand g266 ( new_n468_, new_n460_, new_n467_ );
nand g267 ( new_n469_, new_n457_, new_n459_, new_n466_ );
nand g268 ( new_n470_, new_n468_, new_n469_ );
nand g269 ( new_n471_, new_n470_, new_n397_ );
nand g270 ( new_n472_, new_n468_, keyIn_0_60, new_n469_ );
nand g271 ( new_n473_, new_n471_, new_n472_ );
and g272 ( new_n474_, new_n396_, new_n473_ );
nand g273 ( new_n475_, new_n346_, new_n416_, new_n348_, new_n417_ );
nand g274 ( new_n476_, new_n349_, new_n443_ );
nand g275 ( new_n477_, new_n476_, new_n475_ );
nand g276 ( new_n478_, new_n477_, keyIn_0_42 );
not g277 ( new_n479_, keyIn_0_42 );
nand g278 ( new_n480_, new_n476_, new_n479_, new_n475_ );
nand g279 ( new_n481_, new_n478_, new_n480_ );
nand g280 ( new_n482_, N136, N137 );
xnor g281 ( new_n483_, new_n482_, keyIn_0_20 );
not g282 ( new_n484_, new_n483_ );
nand g283 ( new_n485_, new_n481_, new_n484_ );
nand g284 ( new_n486_, new_n478_, new_n480_, new_n483_ );
nand g285 ( new_n487_, new_n485_, new_n486_ );
nand g286 ( new_n488_, new_n487_, keyIn_0_54 );
not g287 ( new_n489_, keyIn_0_54 );
nand g288 ( new_n490_, new_n485_, new_n489_, new_n486_ );
nand g289 ( new_n491_, new_n488_, new_n490_ );
xnor g290 ( new_n492_, N77, N93 );
xnor g291 ( new_n493_, N109, N125 );
xnor g292 ( new_n494_, new_n492_, new_n493_ );
not g293 ( new_n495_, new_n494_ );
nand g294 ( new_n496_, new_n491_, new_n495_ );
nand g295 ( new_n497_, new_n488_, new_n490_, new_n494_ );
nand g296 ( new_n498_, new_n496_, new_n497_ );
nand g297 ( new_n499_, new_n498_, keyIn_0_62 );
not g298 ( new_n500_, keyIn_0_62 );
nand g299 ( new_n501_, new_n496_, new_n500_, new_n497_ );
and g300 ( new_n502_, new_n499_, new_n501_ );
not g301 ( new_n503_, keyIn_0_61 );
nand g302 ( new_n504_, new_n370_, new_n444_ );
nand g303 ( new_n505_, new_n367_, new_n440_, new_n369_, new_n441_ );
nand g304 ( new_n506_, new_n504_, new_n505_ );
nand g305 ( new_n507_, new_n506_, keyIn_0_41 );
not g306 ( new_n508_, keyIn_0_41 );
nand g307 ( new_n509_, new_n504_, new_n508_, new_n505_ );
nand g308 ( new_n510_, new_n507_, new_n509_ );
nand g309 ( new_n511_, N135, N137 );
xnor g310 ( new_n512_, new_n511_, keyIn_0_19 );
not g311 ( new_n513_, new_n512_ );
nand g312 ( new_n514_, new_n510_, new_n513_ );
nand g313 ( new_n515_, new_n507_, new_n509_, new_n512_ );
nand g314 ( new_n516_, new_n514_, new_n515_ );
nand g315 ( new_n517_, new_n516_, keyIn_0_53 );
not g316 ( new_n518_, keyIn_0_53 );
nand g317 ( new_n519_, new_n514_, new_n518_, new_n515_ );
nand g318 ( new_n520_, new_n517_, new_n519_ );
xor g319 ( new_n521_, N105, N121 );
xnor g320 ( new_n522_, new_n521_, keyIn_0_27 );
xnor g321 ( new_n523_, N73, N89 );
xnor g322 ( new_n524_, new_n523_, keyIn_0_26 );
xnor g323 ( new_n525_, new_n522_, new_n524_ );
xor g324 ( new_n526_, new_n525_, keyIn_0_38 );
not g325 ( new_n527_, new_n526_ );
nand g326 ( new_n528_, new_n520_, new_n527_ );
nand g327 ( new_n529_, new_n517_, new_n519_, new_n526_ );
nand g328 ( new_n530_, new_n528_, new_n529_ );
nand g329 ( new_n531_, new_n530_, new_n503_ );
nand g330 ( new_n532_, new_n528_, keyIn_0_61, new_n529_ );
nand g331 ( new_n533_, new_n531_, new_n532_ );
nor g332 ( new_n534_, new_n502_, new_n533_ );
and g333 ( new_n535_, new_n324_, new_n474_, new_n534_ );
nand g334 ( new_n536_, new_n535_, new_n231_ );
xnor g335 ( N724, new_n536_, N1 );
nand g336 ( new_n538_, new_n535_, new_n315_ );
xnor g337 ( N725, new_n538_, N5 );
nand g338 ( new_n540_, new_n535_, new_n312_ );
xnor g339 ( N726, new_n540_, N9 );
nand g340 ( new_n542_, new_n535_, new_n316_ );
xnor g341 ( N727, new_n542_, N13 );
not g342 ( new_n544_, keyIn_0_76 );
nand g343 ( new_n545_, new_n499_, new_n501_ );
not g344 ( new_n546_, new_n533_ );
nor g345 ( new_n547_, new_n546_, new_n545_ );
nand g346 ( new_n548_, new_n324_, new_n474_, new_n547_ );
nand g347 ( new_n549_, new_n548_, new_n544_ );
nand g348 ( new_n550_, new_n324_, keyIn_0_76, new_n474_, new_n547_ );
nand g349 ( new_n551_, new_n549_, new_n550_ );
nand g350 ( new_n552_, new_n551_, keyIn_0_82, new_n231_ );
not g351 ( new_n553_, keyIn_0_82 );
nand g352 ( new_n554_, new_n551_, new_n231_ );
nand g353 ( new_n555_, new_n554_, new_n553_ );
nand g354 ( new_n556_, new_n555_, new_n552_ );
nand g355 ( new_n557_, new_n556_, new_n328_ );
nand g356 ( new_n558_, new_n555_, N17, new_n552_ );
nand g357 ( new_n559_, new_n557_, new_n558_ );
nand g358 ( new_n560_, new_n559_, keyIn_0_105 );
not g359 ( new_n561_, keyIn_0_105 );
nand g360 ( new_n562_, new_n557_, new_n561_, new_n558_ );
nand g361 ( N728, new_n560_, new_n562_ );
not g362 ( new_n564_, keyIn_0_106 );
not g363 ( new_n565_, keyIn_0_83 );
nand g364 ( new_n566_, new_n551_, new_n565_, new_n315_ );
nand g365 ( new_n567_, new_n551_, new_n315_ );
nand g366 ( new_n568_, new_n567_, keyIn_0_83 );
nand g367 ( new_n569_, new_n568_, new_n566_ );
nand g368 ( new_n570_, new_n569_, N21 );
nand g369 ( new_n571_, new_n568_, new_n329_, new_n566_ );
nand g370 ( new_n572_, new_n570_, new_n571_ );
nand g371 ( new_n573_, new_n572_, new_n564_ );
nand g372 ( new_n574_, new_n570_, keyIn_0_106, new_n571_ );
nand g373 ( N729, new_n573_, new_n574_ );
nand g374 ( new_n576_, new_n551_, new_n312_ );
xnor g375 ( N730, new_n576_, N25 );
not g376 ( new_n578_, keyIn_0_107 );
nand g377 ( new_n579_, new_n551_, keyIn_0_84, new_n316_ );
not g378 ( new_n580_, keyIn_0_84 );
nand g379 ( new_n581_, new_n551_, new_n316_ );
nand g380 ( new_n582_, new_n581_, new_n580_ );
nand g381 ( new_n583_, new_n582_, new_n579_ );
nand g382 ( new_n584_, new_n583_, N29 );
not g383 ( new_n585_, N29 );
nand g384 ( new_n586_, new_n582_, new_n585_, new_n579_ );
nand g385 ( new_n587_, new_n584_, new_n586_ );
nand g386 ( new_n588_, new_n587_, new_n578_ );
nand g387 ( new_n589_, new_n584_, keyIn_0_107, new_n586_ );
nand g388 ( N731, new_n588_, new_n589_ );
not g389 ( new_n591_, keyIn_0_85 );
nand g390 ( new_n592_, new_n394_, new_n471_, new_n395_, new_n472_ );
nor g391 ( new_n593_, new_n592_, new_n502_, new_n533_ );
nand g392 ( new_n594_, new_n324_, keyIn_0_77, new_n593_ );
not g393 ( new_n595_, keyIn_0_77 );
nand g394 ( new_n596_, new_n324_, new_n593_ );
nand g395 ( new_n597_, new_n596_, new_n595_ );
nand g396 ( new_n598_, new_n597_, new_n594_ );
nand g397 ( new_n599_, new_n598_, new_n591_, new_n231_ );
nand g398 ( new_n600_, new_n598_, new_n231_ );
nand g399 ( new_n601_, new_n600_, keyIn_0_85 );
nand g400 ( new_n602_, new_n601_, new_n599_ );
nand g401 ( new_n603_, new_n602_, N33 );
nand g402 ( new_n604_, new_n601_, new_n419_, new_n599_ );
nand g403 ( new_n605_, new_n603_, new_n604_ );
nand g404 ( new_n606_, new_n605_, keyIn_0_108 );
not g405 ( new_n607_, keyIn_0_108 );
nand g406 ( new_n608_, new_n603_, new_n607_, new_n604_ );
nand g407 ( N732, new_n606_, new_n608_ );
not g408 ( new_n610_, keyIn_0_109 );
nand g409 ( new_n611_, new_n598_, keyIn_0_86, new_n315_ );
not g410 ( new_n612_, keyIn_0_86 );
nand g411 ( new_n613_, new_n598_, new_n315_ );
nand g412 ( new_n614_, new_n613_, new_n612_ );
nand g413 ( new_n615_, new_n614_, new_n611_ );
nand g414 ( new_n616_, new_n615_, N37 );
nand g415 ( new_n617_, new_n614_, new_n420_, new_n611_ );
nand g416 ( new_n618_, new_n616_, new_n617_ );
nand g417 ( new_n619_, new_n618_, new_n610_ );
nand g418 ( new_n620_, new_n616_, keyIn_0_109, new_n617_ );
nand g419 ( N733, new_n619_, new_n620_ );
nand g420 ( new_n622_, new_n598_, keyIn_0_87, new_n312_ );
not g421 ( new_n623_, keyIn_0_87 );
nand g422 ( new_n624_, new_n598_, new_n312_ );
nand g423 ( new_n625_, new_n624_, new_n623_ );
nand g424 ( new_n626_, new_n625_, new_n622_ );
nand g425 ( new_n627_, new_n626_, new_n432_ );
nand g426 ( new_n628_, new_n625_, N41, new_n622_ );
nand g427 ( new_n629_, new_n627_, new_n628_ );
nand g428 ( new_n630_, new_n629_, keyIn_0_110 );
not g429 ( new_n631_, keyIn_0_110 );
nand g430 ( new_n632_, new_n627_, new_n631_, new_n628_ );
nand g431 ( N734, new_n630_, new_n632_ );
nand g432 ( new_n634_, new_n598_, keyIn_0_88, new_n316_ );
not g433 ( new_n635_, keyIn_0_88 );
nand g434 ( new_n636_, new_n598_, new_n316_ );
nand g435 ( new_n637_, new_n636_, new_n635_ );
nand g436 ( new_n638_, new_n637_, new_n634_ );
nand g437 ( new_n639_, new_n638_, new_n433_ );
nand g438 ( new_n640_, new_n637_, N45, new_n634_ );
nand g439 ( new_n641_, new_n639_, new_n640_ );
nand g440 ( new_n642_, new_n641_, keyIn_0_111 );
not g441 ( new_n643_, keyIn_0_111 );
nand g442 ( new_n644_, new_n639_, new_n643_, new_n640_ );
nand g443 ( N735, new_n642_, new_n644_ );
not g444 ( new_n646_, new_n592_ );
and g445 ( new_n647_, new_n324_, new_n547_, new_n646_ );
nand g446 ( new_n648_, new_n647_, new_n231_ );
xnor g447 ( N736, new_n648_, N49 );
nand g448 ( new_n650_, new_n647_, new_n315_ );
xnor g449 ( N737, new_n650_, N53 );
nand g450 ( new_n652_, new_n647_, new_n312_ );
xnor g451 ( N738, new_n652_, N57 );
nand g452 ( new_n654_, new_n647_, new_n316_ );
xnor g453 ( N739, new_n654_, N61 );
not g454 ( new_n656_, N65 );
not g455 ( new_n657_, keyIn_0_89 );
not g456 ( new_n658_, keyIn_0_78 );
not g457 ( new_n659_, keyIn_0_75 );
not g458 ( new_n660_, keyIn_0_73 );
nand g459 ( new_n661_, new_n533_, keyIn_0_65 );
not g460 ( new_n662_, keyIn_0_65 );
nand g461 ( new_n663_, new_n531_, new_n662_, new_n532_ );
nand g462 ( new_n664_, new_n661_, new_n663_ );
nor g463 ( new_n665_, new_n592_, new_n502_ );
nand g464 ( new_n666_, new_n665_, new_n664_ );
nand g465 ( new_n667_, new_n666_, new_n660_ );
nand g466 ( new_n668_, new_n665_, new_n664_, keyIn_0_73 );
nand g467 ( new_n669_, new_n667_, new_n668_ );
not g468 ( new_n670_, keyIn_0_72 );
and g469 ( new_n671_, new_n471_, new_n472_ );
nor g470 ( new_n672_, new_n671_, new_n396_ );
nand g471 ( new_n673_, new_n534_, new_n672_, new_n670_ );
nand g472 ( new_n674_, new_n534_, new_n672_ );
nand g473 ( new_n675_, new_n674_, keyIn_0_72 );
nand g474 ( new_n676_, new_n675_, new_n673_ );
not g475 ( new_n677_, keyIn_0_64 );
nand g476 ( new_n678_, new_n533_, new_n677_ );
nand g477 ( new_n679_, new_n531_, keyIn_0_64, new_n532_ );
nand g478 ( new_n680_, new_n672_, new_n502_, new_n678_, new_n679_ );
nand g479 ( new_n681_, new_n680_, keyIn_0_71 );
not g480 ( new_n682_, keyIn_0_71 );
and g481 ( new_n683_, new_n678_, new_n502_ );
nand g482 ( new_n684_, new_n683_, new_n682_, new_n672_, new_n679_ );
nand g483 ( new_n685_, new_n681_, new_n684_ );
not g484 ( new_n686_, keyIn_0_66 );
nand g485 ( new_n687_, new_n531_, new_n686_, new_n532_ );
nand g486 ( new_n688_, new_n533_, keyIn_0_66 );
nand g487 ( new_n689_, new_n688_, new_n687_ );
and g488 ( new_n690_, new_n396_, new_n473_, new_n545_ );
nand g489 ( new_n691_, new_n689_, new_n690_ );
nand g490 ( new_n692_, new_n691_, keyIn_0_74 );
not g491 ( new_n693_, keyIn_0_74 );
nand g492 ( new_n694_, new_n689_, new_n690_, new_n693_ );
nand g493 ( new_n695_, new_n692_, new_n694_ );
nand g494 ( new_n696_, new_n685_, new_n669_, new_n695_, new_n676_ );
nand g495 ( new_n697_, new_n696_, new_n659_ );
and g496 ( new_n698_, new_n669_, new_n676_ );
and g497 ( new_n699_, new_n685_, new_n695_ );
nand g498 ( new_n700_, new_n699_, new_n698_, keyIn_0_75 );
nand g499 ( new_n701_, new_n700_, new_n697_ );
xnor g500 ( new_n702_, new_n315_, keyIn_0_67 );
nand g501 ( new_n703_, new_n231_, new_n312_, new_n310_ );
nor g502 ( new_n704_, new_n702_, new_n703_ );
nand g503 ( new_n705_, new_n701_, new_n704_ );
nand g504 ( new_n706_, new_n705_, new_n658_ );
nand g505 ( new_n707_, new_n701_, keyIn_0_78, new_n704_ );
nand g506 ( new_n708_, new_n706_, new_n707_ );
nand g507 ( new_n709_, new_n708_, new_n396_ );
nand g508 ( new_n710_, new_n709_, new_n657_ );
nand g509 ( new_n711_, new_n708_, keyIn_0_89, new_n396_ );
nand g510 ( new_n712_, new_n710_, new_n711_ );
nand g511 ( new_n713_, new_n712_, new_n656_ );
nand g512 ( new_n714_, new_n710_, N65, new_n711_ );
nand g513 ( new_n715_, new_n713_, new_n714_ );
nand g514 ( new_n716_, new_n715_, keyIn_0_112 );
not g515 ( new_n717_, keyIn_0_112 );
nand g516 ( new_n718_, new_n713_, new_n717_, new_n714_ );
nand g517 ( N740, new_n716_, new_n718_ );
not g518 ( new_n720_, keyIn_0_113 );
not g519 ( new_n721_, keyIn_0_90 );
nand g520 ( new_n722_, new_n708_, new_n671_ );
nand g521 ( new_n723_, new_n722_, new_n721_ );
nand g522 ( new_n724_, new_n708_, keyIn_0_90, new_n671_ );
nand g523 ( new_n725_, new_n723_, new_n724_ );
nand g524 ( new_n726_, new_n725_, N69 );
not g525 ( new_n727_, N69 );
nand g526 ( new_n728_, new_n723_, new_n727_, new_n724_ );
nand g527 ( new_n729_, new_n726_, new_n728_ );
nand g528 ( new_n730_, new_n729_, new_n720_ );
nand g529 ( new_n731_, new_n726_, keyIn_0_113, new_n728_ );
nand g530 ( N741, new_n730_, new_n731_ );
not g531 ( new_n733_, keyIn_0_114 );
not g532 ( new_n734_, keyIn_0_91 );
nand g533 ( new_n735_, new_n708_, new_n546_ );
nand g534 ( new_n736_, new_n735_, new_n734_ );
nand g535 ( new_n737_, new_n708_, keyIn_0_91, new_n546_ );
nand g536 ( new_n738_, new_n736_, new_n737_ );
nand g537 ( new_n739_, new_n738_, N73 );
not g538 ( new_n740_, N73 );
nand g539 ( new_n741_, new_n736_, new_n740_, new_n737_ );
nand g540 ( new_n742_, new_n739_, new_n741_ );
nand g541 ( new_n743_, new_n742_, new_n733_ );
nand g542 ( new_n744_, new_n739_, keyIn_0_114, new_n741_ );
nand g543 ( N742, new_n743_, new_n744_ );
not g544 ( new_n746_, keyIn_0_92 );
nand g545 ( new_n747_, new_n708_, new_n502_ );
nand g546 ( new_n748_, new_n747_, new_n746_ );
nand g547 ( new_n749_, new_n708_, keyIn_0_92, new_n502_ );
nand g548 ( new_n750_, new_n748_, new_n749_ );
nand g549 ( new_n751_, new_n750_, N77 );
not g550 ( new_n752_, N77 );
nand g551 ( new_n753_, new_n748_, new_n752_, new_n749_ );
nand g552 ( new_n754_, new_n751_, new_n753_ );
nand g553 ( new_n755_, new_n754_, keyIn_0_115 );
not g554 ( new_n756_, keyIn_0_115 );
nand g555 ( new_n757_, new_n751_, new_n756_, new_n753_ );
nand g556 ( N743, new_n755_, new_n757_ );
not g557 ( new_n759_, keyIn_0_116 );
not g558 ( new_n760_, keyIn_0_93 );
xnor g559 ( new_n761_, new_n262_, keyIn_0_68 );
nand g560 ( new_n762_, new_n319_, new_n316_ );
nor g561 ( new_n763_, new_n761_, new_n762_ );
nand g562 ( new_n764_, new_n701_, new_n763_ );
nand g563 ( new_n765_, new_n764_, keyIn_0_79 );
not g564 ( new_n766_, keyIn_0_79 );
nand g565 ( new_n767_, new_n701_, new_n763_, new_n766_ );
nand g566 ( new_n768_, new_n765_, new_n767_ );
nand g567 ( new_n769_, new_n768_, new_n396_ );
nand g568 ( new_n770_, new_n769_, new_n760_ );
nand g569 ( new_n771_, new_n768_, keyIn_0_93, new_n396_ );
nand g570 ( new_n772_, new_n770_, new_n771_ );
nand g571 ( new_n773_, new_n772_, N81 );
not g572 ( new_n774_, N81 );
nand g573 ( new_n775_, new_n770_, new_n774_, new_n771_ );
nand g574 ( new_n776_, new_n773_, new_n775_ );
nand g575 ( new_n777_, new_n776_, new_n759_ );
nand g576 ( new_n778_, new_n773_, keyIn_0_116, new_n775_ );
nand g577 ( N744, new_n777_, new_n778_ );
not g578 ( new_n780_, keyIn_0_94 );
nand g579 ( new_n781_, new_n768_, new_n671_ );
nand g580 ( new_n782_, new_n781_, new_n780_ );
nand g581 ( new_n783_, new_n768_, keyIn_0_94, new_n671_ );
nand g582 ( new_n784_, new_n782_, new_n783_ );
nand g583 ( new_n785_, new_n784_, N85 );
not g584 ( new_n786_, N85 );
nand g585 ( new_n787_, new_n782_, new_n786_, new_n783_ );
nand g586 ( new_n788_, new_n785_, new_n787_ );
nand g587 ( new_n789_, new_n788_, keyIn_0_117 );
not g588 ( new_n790_, keyIn_0_117 );
nand g589 ( new_n791_, new_n785_, new_n790_, new_n787_ );
nand g590 ( N745, new_n789_, new_n791_ );
not g591 ( new_n793_, keyIn_0_118 );
not g592 ( new_n794_, keyIn_0_95 );
nand g593 ( new_n795_, new_n768_, new_n546_ );
nand g594 ( new_n796_, new_n795_, new_n794_ );
nand g595 ( new_n797_, new_n768_, keyIn_0_95, new_n546_ );
nand g596 ( new_n798_, new_n796_, new_n797_ );
nand g597 ( new_n799_, new_n798_, N89 );
not g598 ( new_n800_, N89 );
nand g599 ( new_n801_, new_n796_, new_n800_, new_n797_ );
nand g600 ( new_n802_, new_n799_, new_n801_ );
nand g601 ( new_n803_, new_n802_, new_n793_ );
nand g602 ( new_n804_, new_n799_, keyIn_0_118, new_n801_ );
nand g603 ( N746, new_n803_, new_n804_ );
not g604 ( new_n806_, keyIn_0_119 );
not g605 ( new_n807_, keyIn_0_96 );
nand g606 ( new_n808_, new_n768_, new_n502_ );
nand g607 ( new_n809_, new_n808_, new_n807_ );
nand g608 ( new_n810_, new_n768_, keyIn_0_96, new_n502_ );
nand g609 ( new_n811_, new_n809_, new_n810_ );
nand g610 ( new_n812_, new_n811_, N93 );
not g611 ( new_n813_, N93 );
nand g612 ( new_n814_, new_n809_, new_n813_, new_n810_ );
nand g613 ( new_n815_, new_n812_, new_n814_ );
nand g614 ( new_n816_, new_n815_, new_n806_ );
nand g615 ( new_n817_, new_n812_, keyIn_0_119, new_n814_ );
nand g616 ( N747, new_n816_, new_n817_ );
not g617 ( new_n819_, keyIn_0_120 );
not g618 ( new_n820_, keyIn_0_80 );
nor g619 ( new_n821_, new_n231_, new_n288_, new_n262_, new_n316_ );
nand g620 ( new_n822_, new_n701_, new_n821_ );
nand g621 ( new_n823_, new_n822_, new_n820_ );
nand g622 ( new_n824_, new_n701_, keyIn_0_80, new_n821_ );
nand g623 ( new_n825_, new_n823_, new_n824_ );
nand g624 ( new_n826_, new_n825_, new_n396_ );
nand g625 ( new_n827_, new_n826_, keyIn_0_97 );
not g626 ( new_n828_, keyIn_0_97 );
nand g627 ( new_n829_, new_n825_, new_n828_, new_n396_ );
nand g628 ( new_n830_, new_n827_, new_n829_ );
nand g629 ( new_n831_, new_n830_, N97 );
not g630 ( new_n832_, N97 );
nand g631 ( new_n833_, new_n827_, new_n832_, new_n829_ );
nand g632 ( new_n834_, new_n831_, new_n833_ );
nand g633 ( new_n835_, new_n834_, new_n819_ );
nand g634 ( new_n836_, new_n831_, keyIn_0_120, new_n833_ );
nand g635 ( N748, new_n835_, new_n836_ );
not g636 ( new_n838_, keyIn_0_98 );
nand g637 ( new_n839_, new_n825_, new_n671_ );
nand g638 ( new_n840_, new_n839_, new_n838_ );
nand g639 ( new_n841_, new_n825_, keyIn_0_98, new_n671_ );
nand g640 ( new_n842_, new_n840_, new_n841_ );
nand g641 ( new_n843_, new_n842_, N101 );
not g642 ( new_n844_, N101 );
nand g643 ( new_n845_, new_n840_, new_n844_, new_n841_ );
nand g644 ( new_n846_, new_n843_, new_n845_ );
nand g645 ( new_n847_, new_n846_, keyIn_0_121 );
not g646 ( new_n848_, keyIn_0_121 );
nand g647 ( new_n849_, new_n843_, new_n848_, new_n845_ );
nand g648 ( N749, new_n847_, new_n849_ );
nand g649 ( new_n851_, new_n825_, new_n546_ );
nand g650 ( new_n852_, new_n851_, keyIn_0_99 );
not g651 ( new_n853_, keyIn_0_99 );
nand g652 ( new_n854_, new_n825_, new_n853_, new_n546_ );
nand g653 ( new_n855_, new_n852_, new_n854_ );
nand g654 ( new_n856_, new_n855_, N105 );
not g655 ( new_n857_, N105 );
nand g656 ( new_n858_, new_n852_, new_n857_, new_n854_ );
nand g657 ( new_n859_, new_n856_, new_n858_ );
nand g658 ( new_n860_, new_n859_, keyIn_0_122 );
not g659 ( new_n861_, keyIn_0_122 );
nand g660 ( new_n862_, new_n856_, new_n861_, new_n858_ );
nand g661 ( N750, new_n860_, new_n862_ );
not g662 ( new_n864_, keyIn_0_123 );
nand g663 ( new_n865_, new_n825_, new_n502_ );
nand g664 ( new_n866_, new_n865_, keyIn_0_100 );
not g665 ( new_n867_, keyIn_0_100 );
nand g666 ( new_n868_, new_n825_, new_n867_, new_n502_ );
nand g667 ( new_n869_, new_n866_, new_n868_ );
nand g668 ( new_n870_, new_n869_, N109 );
not g669 ( new_n871_, N109 );
nand g670 ( new_n872_, new_n866_, new_n871_, new_n868_ );
nand g671 ( new_n873_, new_n870_, new_n872_ );
nand g672 ( new_n874_, new_n873_, new_n864_ );
nand g673 ( new_n875_, new_n870_, keyIn_0_123, new_n872_ );
nand g674 ( N751, new_n874_, new_n875_ );
not g675 ( new_n877_, keyIn_0_101 );
not g676 ( new_n878_, keyIn_0_81 );
xnor g677 ( new_n879_, new_n262_, keyIn_0_70 );
nor g678 ( new_n880_, new_n231_, keyIn_0_69 );
nand g679 ( new_n881_, new_n229_, keyIn_0_69, new_n230_ );
nand g680 ( new_n882_, new_n881_, new_n315_, new_n316_ );
nor g681 ( new_n883_, new_n879_, new_n880_, new_n882_ );
nand g682 ( new_n884_, new_n701_, new_n883_ );
nand g683 ( new_n885_, new_n884_, new_n878_ );
nand g684 ( new_n886_, new_n701_, new_n883_, keyIn_0_81 );
nand g685 ( new_n887_, new_n885_, new_n886_ );
nand g686 ( new_n888_, new_n887_, new_n396_ );
nand g687 ( new_n889_, new_n888_, new_n877_ );
nand g688 ( new_n890_, new_n887_, keyIn_0_101, new_n396_ );
nand g689 ( new_n891_, new_n889_, new_n890_ );
nand g690 ( new_n892_, new_n891_, N113 );
not g691 ( new_n893_, N113 );
nand g692 ( new_n894_, new_n889_, new_n893_, new_n890_ );
nand g693 ( new_n895_, new_n892_, new_n894_ );
nand g694 ( new_n896_, new_n895_, keyIn_0_124 );
not g695 ( new_n897_, keyIn_0_124 );
nand g696 ( new_n898_, new_n892_, new_n897_, new_n894_ );
nand g697 ( N752, new_n896_, new_n898_ );
not g698 ( new_n900_, keyIn_0_125 );
not g699 ( new_n901_, keyIn_0_102 );
nand g700 ( new_n902_, new_n887_, new_n671_ );
nand g701 ( new_n903_, new_n902_, new_n901_ );
nand g702 ( new_n904_, new_n887_, keyIn_0_102, new_n671_ );
nand g703 ( new_n905_, new_n903_, new_n904_ );
nand g704 ( new_n906_, new_n905_, N117 );
not g705 ( new_n907_, N117 );
nand g706 ( new_n908_, new_n903_, new_n907_, new_n904_ );
nand g707 ( new_n909_, new_n906_, new_n908_ );
nand g708 ( new_n910_, new_n909_, new_n900_ );
nand g709 ( new_n911_, new_n906_, keyIn_0_125, new_n908_ );
nand g710 ( N753, new_n910_, new_n911_ );
not g711 ( new_n913_, N121 );
not g712 ( new_n914_, keyIn_0_103 );
nand g713 ( new_n915_, new_n887_, new_n546_ );
nand g714 ( new_n916_, new_n915_, new_n914_ );
nand g715 ( new_n917_, new_n887_, keyIn_0_103, new_n546_ );
nand g716 ( new_n918_, new_n916_, new_n917_ );
nand g717 ( new_n919_, new_n918_, new_n913_ );
nand g718 ( new_n920_, new_n916_, N121, new_n917_ );
nand g719 ( new_n921_, new_n919_, new_n920_ );
nand g720 ( new_n922_, new_n921_, keyIn_0_126 );
not g721 ( new_n923_, keyIn_0_126 );
nand g722 ( new_n924_, new_n919_, new_n923_, new_n920_ );
nand g723 ( N754, new_n922_, new_n924_ );
not g724 ( new_n926_, keyIn_0_127 );
not g725 ( new_n927_, keyIn_0_104 );
nand g726 ( new_n928_, new_n887_, new_n502_ );
nand g727 ( new_n929_, new_n928_, new_n927_ );
nand g728 ( new_n930_, new_n887_, keyIn_0_104, new_n502_ );
nand g729 ( new_n931_, new_n929_, new_n930_ );
nand g730 ( new_n932_, new_n931_, N125 );
not g731 ( new_n933_, N125 );
nand g732 ( new_n934_, new_n929_, new_n933_, new_n930_ );
nand g733 ( new_n935_, new_n932_, new_n934_ );
nand g734 ( new_n936_, new_n935_, new_n926_ );
nand g735 ( new_n937_, new_n932_, keyIn_0_127, new_n934_ );
nand g736 ( N755, new_n936_, new_n937_ );
endmodule