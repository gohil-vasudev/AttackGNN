module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g34435, g34788, g34839, g36, g44, g53, g54,
         g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751,
         g6753, g84, g90, g91, g92, g99, test_so10, test_so26, test_so35,
         test_so39, test_so42, test_so44, test_so46, test_so80, test_so86,
         test_so92, test_so100, g34783, n4896, n4895, n4837, n4921, n4920,
         n2787, n5045, g559, n4959, g33046, g5057, n5615, g34441, g2771, n5544,
         g33982, g1882, g34007, g2299, g24276, g4040, n5530, g30381, g2547,
         n5782, g30405, g3243, g25604, g452, g30416, g3542, g30466, g5232,
         g25736, g5813, g34617, g33974, g1744, g30505, g5909, g33554, g1802,
         n5536, g30432, g3554, g33064, g6219, n5385, g34881, g807, n5479,
         g6031, g24216, g847, n5709, g24232, n9367, g34733, g4172, g34882,
         g4372, g33026, g3512, g31867, n5471, g25668, g3490, n5454, g24344,
         n5432, g4235, g33966, g1600, g33550, g1714, n5460, g30393, g3155,
         n5366, g29248, g2236, g4571, g4555, g24274, g3698, g33973, g1736,
         g30360, g1968, n5664, g34460, g30494, g5607, g30384, g2657, n5316,
         g24340, n5439, g29223, g490, n5708, g26881, g311, n5317, g34252, g772,
         n5334, g30489, g5587, g29301, g6177, n5874, g6377, g33022, g3167,
         n5652, g30496, g5615, g33043, g4567, g29263, g30533, g6287, g24256,
         n5302, g34015, g2563, g34031, g4776, n5707, g34452, g4593, n5303,
         g34646, g6199, g34001, g2295, g25633, g1384, g24259, g1339, n5381,
         g33049, g5180, n5384, g34609, g2844, g31869, g1024, g30490, g30427,
         g3598, g21894, g4264, n5823, g33965, g767, n5333, g34645, g5853,
         g33571, g2089, g34267, g4933, g26971, g4521, n5752, g34644, g5507,
         g30534, g6291, g33535, g294, n5680, g30498, g25728, g25743, g25684,
         g3813, g25613, g562, g34438, g608, n5475, g24244, g1205, n5547,
         g30439, g3909, g30541, g6259, g30519, g5905, g25621, g921, g34807,
         g2955, g25599, g203, g24235, g34036, g4878, n5283, g30476, g5204,
         g30429, g3606, g32997, g1926, n5510, g33063, g6215, n5651, g30424,
         g3586, g32977, g291, n5679, g34026, g4674, n5440, g30420, g3570,
         g33560, g29226, g676, n5751, g25619, g843, g34455, g4332, n5540,
         g30457, g4153, g33625, g6336, n5592, g34790, g622, n5672, g30414,
         g3506, n5576, g26966, g4558, g25656, g3111, g30390, g25688, g34727,
         g939, g25594, g278, n5627, g26963, g4492, g34034, g4864, n5318,
         g33541, g1036, g28093, g24236, g1178, g30404, g3239, g28051, g718,
         g29303, g6195, n5741, g26917, g1135, n5328, g33624, g6395, n5396,
         g24337, g34911, g554, g33963, g496, g34627, g3853, g29282, g5134,
         n5807, g25676, g33013, g2485, n5509, g32981, g925, n5725, g34976,
         n9357, g30483, g5555, g32994, g1798, g28070, g34806, g2941, g30453,
         g3905, g33539, g763, n5332, g30526, g6255, g26951, g4375, g34035,
         g4871, n5443, g34636, g4722, g32978, g590, n5472, g30348, g1632,
         n5836, g24336, n5438, g3100, g24250, g29236, g1437, n5696, g29298,
         g6154, n5747, g1579, g30499, g5567, g33976, g1752, g32996, g1917,
         g30335, g744, n5470, g34637, g4737, n5867, g25694, g30528, g6267,
         g24251, g1442, g30521, g26960, g4477, n5849, g24239, g34259, g4643,
         n5382, g30474, g5264, n5703, g33016, g2610, g34643, g5160, g30510,
         g5933, g29239, g1454, n5866, g26897, g753, g34729, g1296, g34625,
         g3151, g34800, g24353, g6727, n5531, g33029, g3530, n5569, g4104,
         g24253, g1532, g24281, g33997, n9352, g34971, n9351, g34263, g4754,
         g24237, g1189, n5642, g33584, g2287, n5353, g24280, g4273, n5764,
         g26920, g1389, g33548, g29296, g5835, n5663, g30338, g1171, n5363,
         g21895, g4269, n5763, g33588, g2399, n5762, g34041, g4983, n5367,
         g30495, g5611, g29279, g4572, g25655, g3143, n5882, g34795, g2898,
         g24269, g3343, g30403, g3235, g33042, g30419, g3566, g34023, n9348,
         g28090, g4961, g34642, g4927, n5879, g30370, g2259, n5419, g34448,
         g2819, n5609, g26946, g5802, g34610, g2852, g24209, g417, n5358,
         g28047, g681, g24206, g437, g26891, g30504, g5901, g34798, g2886,
         g25669, g3494, n5889, g30480, g5511, n5575, g33027, g3518, n5645,
         g33972, g1604, g25697, g5092, g28099, g4831, g26947, g4382, g24350,
         g6386, g24210, g479, g30455, g3965, g28084, g33993, g2008, g736,
         g30444, g3933, g33537, g222, g25650, g3050, g25625, g1052, g30366,
         g2122, n5784, g33593, g2465, n5523, g30502, g5889, g33036, g4495,
         g25595, g34462, g33024, g3179, n5390, g33552, g1728, n5352, g34014,
         g2433, g29273, g3835, n5662, g25748, g6187, n5453, g34638, g4917,
         g30341, g1070, g26899, g822, n5422, g30336, g914, n5560, g5339,
         g26940, g4164, g25622, g34447, g2807, n5379, g33613, g4054, n5395,
         g25749, g6191, n5888, g25704, g5077, n5455, g33053, g5523, n5647,
         g3680, g30555, g6637, g25601, g174, n5402, g33971, g1682, g26892,
         g355, g1087, g26915, g1105, n5478, g33008, g30538, g6307, g3802,
         g25750, g6159, g30369, g2255, n5414, g34446, g2815, n5404, g29230,
         g911, n5559, g43, g33975, g1748, g30497, g5551, g30418, g3558, g25721,
         g5499, n5885, g34622, g30438, g3901, g34266, g4888, g30540, g6251,
         g32986, g1373, g25648, g33960, g157, n5678, g34442, g2783, n5403,
         g4281, g30421, g3574, g33573, g2112, g34730, g1283, g24205, g10122_Tj,
         g4297, n5698, g32979, g758, n5331, g34025, g4639, n5727, g25763,
         g6537, n5884, g30481, g5543, g30517, g5961, g30539, g6243, g34880,
         n9340, g24242, n5654, g30436, g29265, g3476, n5786, g32990, g1664,
         g24245, g1246, n5756, g30553, g6629, g26907, g246, n6008, g24278,
         g4049, g26955, g24282, g2932, g29276, g4575, g31894, g4098, n5350,
         g33037, g4498, g26894, g528, n5327, g34977, n5477, g25654, g3139,
         n5447, g33962, g34451, g4584, n5539, g34250, g142, n5724, g29295,
         g5831, g26905, g239, g25629, g1216, n5442, g34792, g2848, g25703,
         g5022, g32983, g1030, g30402, g3231, g25757, g1430, n9336, g33999,
         g2241, g1564, g25729, g6148, g30558, g6649, g34781, g110, g26901,
         g225, n5597, g26961, g33039, g4504, g33059, g5873, n5388, g31899,
         g5037, n5611, g33007, g2319, n5375, g25720, g5495, n5446, g21891,
         g30462, g5208, g30487, g5579, g33058, g5869, n5649, g24261, g1589,
         n5755, g25730, g5752, g30531, g6279, g30506, g34804, g2975, n5750,
         g25747, g6167, n5430, n5701, g33601, g2599, n5524, g26922, g1448,
         n5343, g29250, g2370, g30459, g5164, n5570, g1333, n5616, g33534,
         g153, n5677, g30543, g6549, n5571, g29275, g4087, n5480, g34030,
         g34980, g2984, g30451, g3961, g25627, g962, n5630, g34657, g101,
         g30552, g6625, g34979, n9332, g30337, g1018, g24254, g24277, g4045,
         g29237, g1467, n5693, g30378, g2461, n5840, g33019, n5300, g33623,
         g5990, n5589, g29235, g1256, n5558, g31902, g5029, n5601, g29306,
         g6519, n5806, g25689, g4169, n5729, g33978, g1816, g26970, g4369,
         g29278, g4578, g34253, g4459, n5765, g29272, g3831, n5872, g33595,
         g2514, g33610, g3288, n5400, g33589, g34605, g2145, n5307, g30350,
         g1700, n5417, g25611, g513, n5548, g2841, n5963, g33619, g5297, n5588,
         g34022, g2763, g34033, g4793, n5368, g34726, g952, g31870, g1263,
         n5674, g33985, g1950, g29283, g5138, n5871, g34003, g2307, g25677,
         g34463, g4664, g33006, g2223, g29292, g5808, n5749, g30557, g6645,
         g33989, g2016, g33033, g3873, n5387, n5699, g34005, g2315, g26932,
         g2811, g30516, g5957, g33575, g2047, g33032, g30486, g5575, g34974,
         n9327, g25678, g3752, g30440, g3917, DFF_480_n1, g1585, n5757, g26949,
         g4388, g30530, g6275, g30542, g6311, g25624, g1041, g30383, g33597,
         g2537, g34598, g26957, g4430, g26967, n9325, g28102, g4826, g30524,
         g6239, g26903, g232, g30475, g5268, g34647, g6545, g30377, n9324,
         g33553, g1772, n5504, g31903, g5052, n5607, g25715, g33984, g1890,
         g33602, g2629, n5521, g28045, g572, n5337, g34603, g2130, g33035,
         g4108, n5715, g4308, g24208, g475, g990, n5622, g31, n5469, g34970,
         n9322, g24213, g33614, g3990, n5594, g33060, g30362, g1992, g33023,
         g3171, n5603, g26898, g812, n5733, g25618, g832, g30518, g5897, g4570,
         n5702, g26959, g4455, g34801, g2902, g26884, g333, g25600, g168,
         n5606, g26933, g28066, g3684, g33612, g3639, n5591, g24268, g3338,
         n5527, g25716, g5406, g26906, g269, g24203, g401, g24346, g6040,
         g24207, g441, g25701, n5690, g29269, g3808, n5745, g9, n5468, g34255,
         g30450, g3957, g30456, g4093, n5340, g32991, g1760, n5602, g24348,
         n5437, g34249, g160, n5843, g30371, g2279, n5778, g29268, g3498,
         n5740, g29224, g586, n5336, g33017, g2619, n5508, g30339, g1183,
         n5599, g33967, g1608, g33559, g1779, g29255, g2652, g30368, g2193,
         n5839, g30375, g2393, n5421, g28052, g661, g28089, g4950, g33055,
         g5535, n5566, g30392, g2834, g30343, g1361, g30523, g6235, g24233,
         g1146, n5851, g33018, g32976, g150, n5676, g30349, g1696, n5628,
         g33067, g6555, g26900, g33034, g3881, n5564, g30551, g6621, g25667,
         g3470, n5424, g30452, g3897, g34719, g518, g538, g33607, g2606, n5311,
         g26923, g1472, n5290, g24211, g33050, g5188, n5567, g24341, g5689,
         n5529, g24201, g405, g30463, g5216, g6494, g34464, g4669, g24243,
         g996, g24335, g4531, g34611, g2860, g34262, g4743, g30546, g6593,
         g25591, g4411, g30347, g1413, g30556, g6641, g6, g33562, g1936, n5534,
         g55, g25610, g504, n5519, g33015, g2587, n5372, g31896, g4480, g34004,
         n9314, g30428, g30485, g5571, g30422, g3578, g25714, g29294, g5827,
         n5809, g30423, g3582, g30529, g6271, g34028, g4688, n5656, g33587,
         g2380, g30460, g5196, g30401, g3227, g33990, n9312, g29309, g6541,
         n5739, g30411, g3203, g33546, g1668, n5598, g28085, g4760, g26904,
         g262, g33556, g1840, n5451, g25722, g5467, g25605, g460, g33062,
         g6209, g26893, n5704, g28050, g655, g34626, g33583, g2204, n5620,
         g30472, g5256, g34454, g4608, n5274, g34850, g794, n5291, g4423,
         g24272, g3689, n5532, g5685, g24214, g703, n5821, g26909, g862, n5682,
         g30406, g3247, g33569, g2040, n5505, g34628, g4146, n5981, g34458,
         g4633, n5844, g24240, n5304, g34634, g4732, g25700, n5689, g29293,
         g5817, g33009, g2351, n5511, g33603, g2648, g24355, g6736, g34268,
         g4944, g25691, g4072, g26890, g3466, g28072, g4116, g31900, g5041,
         n5605, g26956, g4434, g29271, g3827, n5808, g29304, g6500, n5748,
         g29261, g3133, n5661, g28063, g3333, g979, n5320, g34027, g4681,
         g33961, g298, n5675, g33604, g32995, g1894, n5374, g34624, g2988,
         g30415, g3538, g33536, g301, g26888, n9306, DFF_709_n1, g28055, g827,
         n5728, g24238, g33600, g2555, n5351, g28105, g5011, g34721, g199,
         g29307, g6523, n5870, g30345, g34453, g4601, n5365, g32980, g854,
         g29238, g1484, n5865, g34639, g4922, g25695, g5080, n5893, g33057,
         g5863, g26969, g4581, n5670, g29253, g2518, g34021, g2567, g26895,
         g568, n5335, g30413, g3263, g30549, g6613, g24347, g25758, g6444,
         g34808, g2965, g30501, g5857, n5573, g33969, n9303, g34440, g890,
         n5305, g30433, g3562, g21900, g26921, g1404, g29270, g3817, n9302,
         g33038, g4501, g31865, g26926, g2724, n5301, g28083, g4704, g34797,
         g22, g2878, g30478, g5220, g34724, g617, n5339, g24212, g26883, g316,
         g32985, g1277, g25761, g6513, n5426, g26886, g336, n5824, g34796,
         g2882, g32982, g33561, g1906, n5503, g26880, g305, n5282, g34975, g8,
         g26931, g2799, g34641, g4912, g34629, g4157, n5983, g33598, g2541,
         n5461, g33576, g2153, n5356, g34720, g550, g26902, g255, g29244,
         g30468, g5240, g26924, g1478, n5289, g33031, g3863, g29245, g1959,
         g29266, g3480, n5868, g30559, g6653, g34794, g2864, g28087, g4894,
         g30435, g3857, n5572, g25609, g28057, g1002, g34439, g776, n5330, g28,
         n5324, g1236, g34260, g4646, n5712, g33012, g2476, g32989, g1657,
         n5525, g34006, g2375, g63, g358, g26910, g896, n5431, g28043, g33021,
         g3161, g29251, g2384, n5700, g34456, g4616, n5608, g26968, g4561,
         g33991, g2024, g3451, g26930, g2795, g34599, g613, n5474, g28082,
         g4527, g33557, g1844, g30511, g5937, g33045, g30379, g2523, n5281,
         g24267, n5436, g34020, g2643, g24249, g1489, n5850, g25592, g30382,
         n9295, g29285, g5156, n5734, n5526, n9294, g25662, g21896, g33563,
         g1955, g33622, g33582, g2273, n5458, g28086, g4771, g25744, g6098,
         g29262, g3147, n5738, g24270, g3347, g33581, g2269, g191, g24266,
         g2712, g34849, g626, n5288, g33618, g2729, g5357, n5393, g34038,
         g34032, g4709, n5518, g34803, g2927, g34459, g4340, n5653, g30509,
         g5929, g34640, g4907, g28069, g4035, g21899, g2946, g31868, g918,
         n5673, g26938, g4082, g25756, g30363, g30334, g577, n5294, g33970,
         g1620, g30391, g2831, g25615, g667, g33540, g930, n5731, g30445,
         g3937, g25617, g817, n5822, g24247, g1249, g24215, g837, n5562,
         g33964, g599, n5550, g25719, g5475, n5425, g29228, g30514, g5949,
         g33627, g6682, n5590, g24231, g904, g34615, g2873, n5488, g30356,
         g1854, n5785, g25696, g5084, n5681, g30493, g5603, n5726, g33594,
         g2495, n5522, g34009, g2437, g30365, g2102, n5666, g33004, g2208,
         g34018, g25685, g4064, n5416, g34040, g4899, n5517, g25639, g2719,
         n5465, g34029, g4785, n5361, g30488, g5583, g34600, g781, n5551,
         g29300, g6173, n5810, g34802, g2917, g25614, g686, g28058, g1252,
         n5554, g29225, g671, g33580, g30532, g6283, DFF_909_n1, g33054, g5527,
         n5389, g26962, g4489, g33564, g1974, n5450, g32984, g1270, n5716,
         g34039, g4966, n5706, g33065, g6227, n5568, g30443, g3929, g29291,
         g5503, n5737, g24279, g30508, g5925, g29232, g1124, n5692, g34269,
         g4955, g30464, g5224, g33988, g2012, g30522, g6203, n5574, g25708,
         g5120, g30374, g2389, n5631, g26953, g4438, g34008, g2429, g34444,
         g2787, n5610, g34731, g33606, g2675, n5457, g24334, g34265, g4836,
         n5713, g30340, g1199, g24257, n5401, g30482, g5547, g34604, g2138,
         n5275, g33591, g2338, n5310, g30525, g6247, g26929, g2791, g30448,
         g34602, g1291, n2549, g30513, g5945, g30469, g5244, g33608, g2759,
         g33626, g6741, n5398, g34725, g785, n5293, g30342, g1259, n5553,
         g29267, g3484, n5668, g25593, g209, n5595, g30548, g6609, g33052,
         g5517, g34012, g2449, g34017, n9281, DFF_961_n1, g24263, g2715, n5299,
         g26912, g936, n5557, g30364, g2098, n5280, g34254, g4462, n5671,
         g34251, g604, n5473, g30560, g6589, g33983, n9280, g24204, g429,
         g33980, g1870, g34631, g29243, g1825, g25623, g1008, n5321, g26950,
         g4392, n5710, g30431, g3546, g30467, g5236, g30353, g1768, n5834,
         g34467, g4854, g30442, g3925, g29305, g6509, g25616, g732, n5732,
         g29252, g2504, g4519, g4520, g33003, g2185, n5376, g34613, g37, g4031,
         g33570, g2070, n5535, g34734, g4176, g24275, n5435, g4405, g872,
         g29302, g6181, n5667, g24349, g34264, g4765, g30484, g5563, g25634,
         g1395, g33567, g1913, g33585, g2331, n5513, g30527, g6263, g34978,
         n9276, g30447, g3945, g347, n5860, g34256, g4473, g25630, g1266,
         g29290, g5489, n5660, g29227, g31872, g2748, n5516, g29287, g5471,
         g31897, g4540, g6723, g30562, g6605, g34011, n9274, g33996, g2173,
         g21898, g33014, g2491, g34465, g4849, g33995, g2169, g30372, n9273,
         g30545, g30389, g33590, g2407, n5459, g34616, g2868, g26927, g2767,
         g32992, g1783, n5596, g25631, g1312, n5466, g30477, g5212, g34632,
         g4245, g28046, g645, g4291, g26896, n5657, g25602, g26916, g1129,
         n5329, g33578, g2227, n5538, g33579, g2246, g30354, g1830, n5413,
         g30425, g3590, g24200, g392, g33544, g1592, n5362, g25764, g6505,
         g1221, g30507, g5921, g26889, g30333, g218, g32998, g1932, g32987,
         g1624, n5370, g25702, g5062, g29286, g5462, n5744, g34606, g2689,
         g33070, g6573, n5563, g29240, g1677, g32999, g2028, n5371, g33605,
         g2671, g24255, g26945, g33558, g1848, n5464, g25699, n5669, g29289,
         g5485, n5869, g30388, g2741, n5349, n5482, g29254, g2638, g28074,
         g4122, g34450, g4322, n5506, g30512, g5941, g33572, g2108, n5452, g25,
         g33551, g33538, g595, n5476, g33005, g2217, n5512, g24248, n9267,
         g33002, g2066, g24234, g1152, n5618, g30471, g5252, g34000, g2165,
         g34016, g2571, g33048, g5176, n5650, g25628, g26934, g2827, g34468,
         g4859, g24202, g424, g33542, g1274, n5730, n9265, n6006, g34445,
         g2803, n5545, g33555, g1821, g34013, g2509, g28091, g5073, g26919,
         n5556, g30554, g6633, g29281, g5124, g30537, g6303, g28092, g5069,
         g34732, g2994, n5634, g28049, g650, g33545, g1636, n5549, g30441,
         g3921, g29247, g24354, g6732, g25636, g1306, n5796, g26914, g1061,
         g25670, g3462, g33998, g2181, g25626, g956, n5341, g33977, g1756,
         g29297, g5849, n5736, g28071, g4112, g30387, n9262, g33577, g2197,
         n5514, g33592, g26913, g1046, g28044, g482, n5820, g26948, g4401,
         g30344, g1514, n5364, g26885, g329, n5766, g33069, g6565, n5386,
         g34621, g2950, g28059, g1345, g25762, g6533, n5445, g34633, g4727,
         g24352, g26925, g1536, g30446, g3941, g25597, g370, g24342, g5694,
         g30357, g1858, g26908, g446, g30399, g3219, g29242, g1811, g30547,
         g6601, g34010, g2441, g33986, g1874, g34257, g30544, g6581, g30561,
         g6597, g5008, g30430, g3610, g34799, g2890, g33565, g1978, g33968,
         g1612, g34843, g112, g34793, g2856, g33566, g1982, n5462, g30465,
         g28073, g4119, g24351, g6390, g30346, g1542, g21893, g4258, g4818,
         g31904, g5033, g34635, g4717, g25637, g1554, n5768, g29274, g3849,
         n5735, g30396, g3199, g25735, g34037, g4975, n5360, g34791, g790,
         n5292, g30520, g5913, g30358, g1902, n5837, g29299, g6163, g25690,
         g4125, g28096, g4821, n5880, g28088, g4939, g24241, n5392, g30397,
         g3207, g4483, g30409, g29284, g5142, n5658, g30470, g5248, g30367,
         g2126, g24273, g3694, g29288, g5481, n5805, g30359, g1964, n5315,
         g25698, g5097, n5753, g30398, g3215, n9255, n6005, g26952, g4427,
         g26928, g2779, n5694, g26954, g30351, g1720, n5780, g31871, g1367,
         g5112, g19, g26939, g4145, g33994, g2161, g25596, g376, n5633, g33586,
         g2361, n5537, g21901, DFF_1234_n1, g31866, g582, n5552, g33000, g2051,
         g26918, g1193, g30373, g2327, n5841, g28056, g907, n5555, g34601,
         g947, n5286, g30355, g1834, n5665, g30426, g3594, g34805, g2999,
         g34002, g2303, g28053, g29229, g723, n5826, g33620, g5703, n5397,
         g34722, g546, g33599, g2472, n5619, g30515, g5953, g25649, g33979,
         g1740, g30417, g3550, g3845, n5886, g33574, g2116, n5463, g30410,
         g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777, g33596,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g31895,
         g4417, g33068, g6561, n5646, g29233, g1141, n5691, g24258, n5655,
         g30376, g33549, g1710, g29308, g6527, n5659, g30408, g3255, g29241,
         g1691, g34620, g2936, g33621, g5644, n5593, g5152, n5883, g24339,
         g5352, g34443, g2775, n5378, g34619, g2922, g29234, g30503, g5893,
         g30550, g6617, g33001, g2060, n5507, g33040, g4512, g30492, g5599,
         g25664, g3401, g26944, g4366, g34614, g29260, g3129, n5861, g33047,
         g5170, g24298, g25733, g5821, n5429, g30536, g6299, g29246, g2079,
         g34261, g4698, g33611, g3703, n5399, g25638, g1559, n5441, g34728,
         n9247, g29222, g411, g25742, g30449, g3953, g34608, g2704, n5377,
         g24345, g6035, n5528, n9245, g25635, g1300, n5483, g25686, g4057,
         n5711, g30461, g5200, g34466, g4843, g31901, g5046, n5578, g29249,
         g2250, g26882, n5456, g33041, g33011, g2453, n5373, g25734, g5841,
         n5449, n5705, g34618, g2912, g33010, g2357, g31864, g164, n5561,
         g34630, g4253, n5484, g31898, g5016, n5369, g25653, g3119, n5423,
         g25632, g1351, n5322, g32988, g33616, g29280, g5115, n5743, g33609,
         g3352, n5604, g30563, g6657, g33044, g4552, g30437, g3893, g30412,
         g3211, g30491, g5595, g30434, g3614, g34612, g29259, g3125, n5781,
         g25681, g3821, n5428, g25687, g4141, n5612, g33617, g30479, g5272,
         g29256, g2735, n5600, g28054, g728, g30535, g6295, g30385, g2661,
         n5418, g30361, g1988, n5783, g25705, g24260, g1548, n5546, g29257,
         g3106, n5742, g34461, g4659, g34258, g4358, n5348, g32993, g1792,
         n5359, g33992, g2084, g30394, g3187, g34449, g4311, n5323, g34019,
         g2583, g18597, n9240, g29231, g1094, n5697, g25682, g21897, g4284,
         g30395, g3191, g21892, g4239, g4180, n5380, g28048, g691, n5520,
         g34723, g534, g25598, g385, n5632, g33987, g2004, g30380, g2527,
         n5420, g5456, g26965, n6007, g25706, g30458, g4507, n5846, g24338,
         g5348, g30400, g3223, g34623, g2970, g24343, g5698, g30473, g5260,
         g24252, g1521, g33028, g3522, n5383, g29258, g3115, g30407, g3251,
         g26958, g34457, g33568, g1996, n5355, g25663, g26964, g4515, g34735,
         g4300, g30352, n9236, g33543, g1379, g24271, n5433, g33981, g1878,
         g30500, g5619, g34649, g71, g29277, g25612, n5287, g28060, n2505,
         n2499, n2396, n2668, g72, n5960, n4689, n5961, n4708, n3593, n3595,
         n3574, n3576, n3517, n3519, n3628, n3630, n3555, n3557, n3646, n3648,
         n3536, n3538, n3611, n3613, n3765, n3505, n3525, n3635, n4888, n2595,
         n2527, n3524, n3005, n3623, n3549, n3799, n3033, n3622, n3587, n3586,
         n3605, n3604, n3568, n3567, n3548, n3512, n3511, n3531, n3530, n3641,
         n3640, n3131, n3111, n4537, n4201, n3745, n3684, n3274, n2982, n2706,
         n2649, n2556, n2509, n2487, n2427, n2423, n4826, n2421, n4172, n4173,
         n4190, n4191, n4388, n4210, n3951, n3774, n3842, n3808, n3908, n3984,
         n3875, n4015, n3446, n3914, n3406, n3780, n3481, n3957, n3426, n3848,
         n3491, n3990, n3416, n3814, n3436, n3881, n3502, n4022, n3501, n4027,
         n3407, n3785, n3482, n3962, n3427, n3853, n3437, n3886, n3417, n3819,
         n3492, n3995, n3447, n3919, n3682, n3272, n2980, n2704, n2647, n2554,
         n2507, n2485, n2425, n2419, n3743, n2405, n2760, n2552, n4198, n2404,
         n4962, n4948, n3195, n3116, n4945, n4525, n4518, n3281, n3277, n3276,
         n2989, n2991, n3687, n3279, n2710, n2707, n3174, n3362, n2644, n3115,
         n3833, n3023, n3933, n3729, n3664, n3662, n3673, n3671, n2607, n2790,
         n4490, n4178, n4514, n4196, n3736, n3741, n2598, n4804, n4811, n4814,
         n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145, n3164, n2422,
         n5121, n4037, n4034, n4039, n3972, n3969, n3929, n3926, n3863, n3860,
         n4003, n4002, n4032, n4035, n3797, n3792, n3790, n3795, n3891, n3893,
         n3827, n3826, n3896, n4007, n3931, n3793, n3924, n3831, n3829, n3927,
         n3974, n3898, n3970, n4000, n3865, n3861, n3824, n3894, n3967, n3858,
         n4005, n3395, n4956, n5026, n3941, n3733, n4798, n4805, n4175, n4193,
         n3738, n4721, n4523, n4524, n4526, n2573, n2577, n2563, n2567, n4938,
         n4913, n4714, n4516, n4517, n5111, n3730, n4305, n4283, n2608, n4447,
         n4448, n4402, n4403, n4425, n4426, n4436, n4437, n4391, n4392, n4379,
         n4380, n4414, n4415, n4458, n4459, n5016, n5014, n3064, n3065, n4535,
         n5112, n3675, counter_31, counter_30, counter_29, counter_28,
         counter_27, counter_26, counter_25, counter_24, counter_23,
         counter_22, counter_21, counter_20, counter_19, counter_18,
         counter_17, counter_16, counter_15, counter_14, counter_13,
         counter_12, counter_11, counter_10, counter_9, counter_8, counter_7,
         counter_6, counter_5, counter_4, counter_3, counter_2, counter_1,
         counter_0, carry_31, carry_30, carry_29, carry_28, carry_27, carry_26,
         carry_25, carry_24, carry_23, carry_22, carry_21, carry_20, carry_19,
         carry_18, carry_17, carry_16, carry_15, carry_14, carry_13, carry_12,
         carry_11, carry_10, carry_9, carry_8, carry_7, carry_6, carry_5,
         carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16, N17, N18, N19,
         N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87, n73, n86, n85,
         n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, n58, n59, n60,
         n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68, n69, n70, n71,
         n72, n55, n57, n92, n93, n115, n130, n141, n158, n178, g33959, n209,
         n217, n218, n223, n225, n227, n231, n232, g33533, n282, n297, n338,
         n342, n353, n388, n399, n463, n465, n470, n471, n517, n528, n549,
         n561, n562, n563, n564, n568, n580, n581, n705, n706, n719, n724,
         n729, n731, n735, n736, n764, n769, n788, n789, n790, n791, n794,
         n795, n797, n822, n837, n839, n843, n844, n865, n939, n943, n944,
         n945, n946, n985, n987, n997, n998, n1022, n1039, n1084, n1122, n1151,
         g25167, n1253, n1256, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1392, n1416, n1418, n1422, n1423, n1430, n1731, n1733, n1795,
         n8272, n8273, n8275, n8276, n8277, n8279, n8281, n8284, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8300, n8301, n8302, n8307, n8310,
         n8311, n8313, n8314, n8315, n8316, n8317, n8318, n8321, n8322, n8323,
         n8324, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8337,
         n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8354, n8356, n8358, n8359, n8360, n8361, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8373, n8374, n8375, n8378, n8379,
         n8381, n8382, n8411, n8412, n8413, n8414, n8415, n8416, n8419, n8506,
         n8507, n8511, n8512, n8513, n8514, n8515, n8516, n8521, n8522, n8523,
         n8524, n8525, n8526, n8537, n8540, n8541, n8542, n8543, n8544, n8545,
         n8547, n8548, n8551, n8552, n8553, n8555, n8572, n8573, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8688, n8689, n8690, n8691, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8733, n8734, n8735, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, g32975, n8806, n8807, n8808, n8809, n8810, n8811,
         g31860, n8813, g31862, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9241, n9242,
         n9243, n9244, n9246, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9256, n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9266, n9268,
         n9269, n9270, n9271, n9272, n9275, n9277, n9278, n9279, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9296, n9297, n9298, n9299, n9300, n9301, n9304, n9305, n9307, n9308,
         n9309, n9310, n9311, n9313, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9323, n9326, n9328, n9329, n9330, n9331, n9333, n9334, n9335,
         n9337, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9349, n9350, n9353, n9354, n9355, n9356, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, U5353_n1, U5355_n1, U5961_n1,
         U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1,
         U6100_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1,
         U6217_n1, U6218_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1,
         U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1,
         U6291_n1, U6292_n1, U6338_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1,
         U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1,
         U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1,
         U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1,
         U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1,
         U6373_n1, U6374_n1, U6375_n1, U6417_n1, U6446_n1, U6465_n1, U6497_n1,
         U6523_n1, U6542_n1, U6552_n1, U6553_n1, U6554_n1, U6555_n1, U6556_n1,
         U6559_n1, U6560_n1, U6561_n1, U6570_n1, U6911_n1, U6912_n1, U6917_n1,
         U6926_n1, U6927_n1, U6929_n1, U6931_n1, U6932_n1, U6933_n1, U6934_n1,
         U6935_n1, U6936_n1, U6937_n1, U6938_n1, U6939_n1, U6940_n1, U6941_n1,
         U6944_n1, U6950_n1, U6954_n1, U6955_n1, U6956_n1, U6957_n1, U7174_n1,
         U7248_n1, U7249_n1, U7402_n1, U7405_n1, U7413_n1, U7416_n1, U7427_n1,
         U7438_n1, U7449_n1, U7455_n1, U7464_n1, U7467_n1, U7482_n1, U7492_n1,
         U7513_n1, U7516_n1, U7549_n1, U7561_n1, U7574_n1, U7577_n1, U7585_n1,
         U7595_n1, U7614_n1, U7621_n1, U7629_n1, U7636_n1, U7639_n1, U7649_n1,
         U7652_n1, U7668_n1, U7673_n1, U7690_n1, U7707_n1, U7712_n1, U7792_n1,
         U7794_n1, U7895_n1, U7897_n1, U7977_n1, U8034_n1, U8036_n1, U8050_n1,
         U8055_n1, U8060_n1, U8070_n1, U8074_n1, U8088_n1, U8112_n1, U8113_n1,
         U8147_n1, U8165_n1, U8185_n1, U8192_n1, U8210_n1, U8223_n1, U8224_n1,
         U8281_n1, U8307_n1, U8974_n1, U8975_n1, U9065_n1, U9070_n1, U9075_n1,
         U9076_n1, U9080_n1, U9084_n1, U9085_n1, U9086_n1, U9090_n1, U9098_n1,
         U9099_n1, U9101_n1, U9107_n1, U9111_n1, U9116_n1, U9120_n1, U9124_n1,
         U9128_n1, U9132_n1, U9136_n1, U9315_n1, U9453_n1, U9825_n1, U9886_n1,
         U9927_n1, U9953_n1, U9957_n1, U9958_n1, U9968_n1, U9972_n1, U9992_n1,
         U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g27831 = g33533;
  assign g31863 = g25167;
  assign g26801 = g32975;
  assign g25114 = g31860;
  assign g25259 = g31862;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n8867), .CLK(n9171), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n8876), .CLK(n9180), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n8928), .CLK(n9232), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n8901), .CLK(n9205), .Q(
        g2299) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n8880), .CLK(n9184), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n8951), .CLK(n9260), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n8951), .CLK(n9260), .Q(g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n8960), .CLK(n9272), .Q(
        g3243) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n8892), .CLK(n9196), .Q(
        g452), .QN(n8419) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n8916), .CLK(n9220), .Q(
        g3542) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n8894), .CLK(n9198), .Q(
        g5232) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n8954), .CLK(n9264), .Q(
        g5813), .QN(n8694) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n8890), .CLK(n9194), .Q(
        test_so1), .QN(n8851) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n8907), .CLK(n9211), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n8897), .CLK(n9201), .Q(
        g5909) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n8963), .CLK(n9278), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n8916), .CLK(n9220), .Q(
        g3554) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n8954), .CLK(n9264), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n8948), .CLK(n9257), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n8948), .CLK(n9257), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n8892), .CLK(n9196), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n8920), .CLK(n9224), .Q(
        n9367) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n8894), .CLK(n9198), .Q(
        g4172) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n8923), .CLK(n9227), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n8923), .CLK(n9227), .Q(
        g3512), .QN(n8637) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n8943), .CLK(n9251), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n8924), .CLK(n9228), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n8883), .CLK(n9187), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n8966), .CLK(n9283), .Q(
        g4235), .QN(n8620) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n8875), .CLK(n9179), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n8919), .CLK(n9223), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n8950), .CLK(n9259), .Q(
        g14451), .QN(n8719) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n8956), .CLK(n9268), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n8904), .CLK(n9208), .Q(
        g2236), .QN(n8634) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n8898), .CLK(n9202), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n8873), .CLK(n9177), .Q(
        g3698), .QN(n8755) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n8907), .CLK(n9211), .Q(
        g1736) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n8928), .CLK(n9232), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n8944), .CLK(n9252), .Q(
        test_so3), .QN(n8842) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n8870), .CLK(n9174), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n8870), .CLK(n9174), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n8883), .CLK(n9187), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n8935), .CLK(n9241), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n8935), .CLK(n9241), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n8945), .CLK(n9253), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n8874), .CLK(n9178), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n8879), .CLK(n9183), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n8956), .CLK(n9268), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n8956), .CLK(n9268), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n8868), .CLK(n9172), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n8968), .CLK(n9285), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n8874), .CLK(n9178), .Q(
        test_so4), .QN(n8821) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n8899), .CLK(n9203), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n8885), .CLK(n9189), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n8929), .CLK(n9233), .Q(
        g2563) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n8949), .CLK(n9258), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n8958), .CLK(n9270), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n8958), .CLK(n9270), .Q(
        g6199) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n8901), .CLK(n9205), .Q(
        g2295) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n8920), .CLK(n9224), .Q(
        g1384), .QN(n8764) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n8932), .CLK(n9237), .Q(
        g1339), .QN(n5381) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n8930), .CLK(n9234), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n8886), .CLK(n9190), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n8922), .CLK(n9226), .Q(
        g1024), .QN(n8795) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n8870), .CLK(n9174), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n8915), .CLK(n9219), 
        .Q(g3598) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n8882), .CLK(n9186), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n8945), .CLK(n9253), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n8945), .CLK(n9253), .Q(
        g5853) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n8957), .CLK(n9269), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n8917), .CLK(n9221), .Q(
        g2089), .QN(n8328) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n8965), .CLK(n9282), .Q(
        g4933) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n8871), .CLK(n9175), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n8871), .CLK(n9175), .Q(
        g5507) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n8950), .CLK(n9259), .Q(
        g16656), .QN(n8718) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n8900), .CLK(n9204), .Q(
        g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n8884), .CLK(n9188), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n8973), .CLK(n9290), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n8954), .CLK(n9264), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n8878), .CLK(n9182), .Q(
        g9741), .QN(n8310) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n8878), .CLK(n9182), .Q(
        g3813), .QN(n8724) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n8878), .CLK(n9182), .Q(
        g562), .QN(n8281) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n8924), .CLK(n9228), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n8962), .CLK(n9277), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n8891), .CLK(n9195), .Q(
        g3909) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n8899), .CLK(n9203), .Q(
        g6259) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n8914), .CLK(n9218), .Q(
        g5905) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n8926), .CLK(n9230), .Q(
        g921), .QN(n8368) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n8867), .CLK(n9171), .Q(
        g2955), .QN(n8367) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n8909), .CLK(n9213), .Q(
        g203), .QN(n8672) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n8934), .CLK(n9239), .Q(
        test_so7), .QN(n8820) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n8939), .CLK(n9246), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n8958), .CLK(n9270), .Q(
        g5204) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n8958), .CLK(n9270), .Q(
        g17604), .QN(n8700) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n8916), .CLK(n9220), .Q(
        g3606) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n8946), .CLK(n9254), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n8954), .CLK(n9264), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n8916), .CLK(n9220), .Q(
        g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n8884), .CLK(n9188), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n8945), .CLK(n9253), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n8916), .CLK(n9220), .Q(
        g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n8925), .CLK(n9229), .Q(
        g9048), .QN(n8272) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n8925), .CLK(n9229), .Q(
        g17607), .QN(n8763) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n8963), .CLK(n9278), .Q(
        test_so8), .QN(n8827) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n8876), .CLK(n9180), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n8892), .CLK(n9196), .Q(
        g843), .QN(n8356) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n8955), .CLK(n9266), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n8894), .CLK(n9198), .Q(
        g4153) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n8894), .CLK(n9198), .Q(
        g17711), .QN(n8669) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n8879), .CLK(n9183), .Q(
        g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n8925), .CLK(n9229), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n8951), .CLK(n9260), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n8898), .CLK(n9202), .Q(
        g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n8943), .CLK(n9251), .Q(
        g17685), .QN(n8706) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n8956), .CLK(n9268), .Q(
        g3111), .QN(n8727) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n8904), .CLK(n9208), .Q(
        g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n8904), .CLK(n9208), .Q(
        test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n8970), .CLK(n9287), 
        .Q(g939) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n8889), .CLK(n9193), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n8889), .CLK(n9193), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n8939), .CLK(n9246), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n8900), .CLK(n9204), .Q(
        g1036), .QN(n8794) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n8900), .CLK(n9204), .Q(
        g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n8900), .CLK(n9204), .Q(
        g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n8959), .CLK(n9271), .Q(
        g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n8959), .CLK(n9271), .Q(
        g718), .QN(n8785) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n8959), .CLK(n9271), .Q(
        g6195), .QN(n5741) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n8907), .CLK(n9211), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n8956), .CLK(n9268), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n8911), .CLK(n9215), .Q(
        test_so10), .QN(n8828) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n8958), .CLK(n9270), 
        .Q(g554) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n8909), .CLK(n9213), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n8972), .CLK(n9289), .Q(
        g3853) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n8896), .CLK(n9200), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n8896), .CLK(n9200), .Q(
        g17404), .QN(n8733) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n8950), .CLK(n9259), .Q(
        g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n8950), .CLK(n9259), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n8970), .CLK(n9287), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n8867), .CLK(n9171), .Q(
        n9357) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n8868), .CLK(n9172), .Q(
        g5555) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n8906), .CLK(n9210), .Q(
        g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n8961), .CLK(n9275), .Q(
        g1798) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n8926), .CLK(n9230), .Q(
        test_so11), .QN(n8825) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n8891), .CLK(n9195), 
        .Q(g2941), .QN(n8526) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n8891), .CLK(n9195), .Q(
        g3905) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n8945), .CLK(n9253), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n8899), .CLK(n9203), .Q(
        g6255) );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(n8877), .CLK(n9181), .Q(
        g4375), .QN(n8277) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n8939), .CLK(n9246), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n8939), .CLK(n9246), .Q(
        g4722) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n8924), .CLK(n9228), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n8964), .CLK(n9279), .Q(
        g13099), .QN(n8716) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n8875), .CLK(n9179), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n8911), .CLK(n9215), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n8920), .CLK(n9224), .Q(
        g3100), .QN(n8324) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n8937), .CLK(n9243), .Q(
        test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n8947), .CLK(n9256), 
        .Q(g1437), .QN(n5696) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n8879), .CLK(n9183), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n8932), .CLK(n9237), .Q(
        g1579), .QN(n8360) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n8868), .CLK(n9172), .Q(
        g5567) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n8907), .CLK(n9211), .Q(
        g1752) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n8941), .CLK(n9249), .Q(
        g1917), .QN(n8779) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n8941), .CLK(n9249), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n8942), .CLK(n9250), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n8942), .CLK(n9250), .Q(
        g8132) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n8899), .CLK(n9203), .Q(
        g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n8899), .CLK(n9203), .Q(
        g16659), .QN(n8714) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n8937), .CLK(n9243), .Q(
        g1442), .QN(n8551) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n8898), .CLK(n9202), .Q(
        test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n8944), .CLK(n9252), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n8944), .CLK(n9252), .Q(
        g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n8944), .CLK(n9252), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n8895), .CLK(n9199), .Q(
        g5264) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n8943), .CLK(n9251), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n8943), .CLK(n9251), .Q(
        g2610), .QN(n8772) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n8943), .CLK(n9251), .Q(
        g5160) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n8914), .CLK(n9218), .Q(
        g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n8932), .CLK(n9237), .Q(
        g1454), .QN(n5866) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n8905), .CLK(n9209), .Q(
        g753), .QN(n8783) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n8905), .CLK(n9209), .Q(
        g1296), .QN(n8275) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n8905), .CLK(n9209), .Q(
        g3151) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n8890), .CLK(n9194), .Q(
        test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n8921), .CLK(n9225), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n8951), .CLK(n9260), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(n399), .SI(g3530), .SE(n8949), .CLK(n9258), .Q(
        g4104), .QN(n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n8885), .CLK(n9189), .Q(
        g1532), .QN(n8573) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n8885), .CLK(n9189), .Q(
        g9251), .QN(n8511) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n8904), .CLK(n9208), .Q(
        n9352) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n8878), .CLK(n9182), .Q(
        n9351) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n8878), .CLK(n9182), .Q(
        g4754) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n8900), .CLK(n9204), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n8901), .CLK(n9205), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n8882), .CLK(n9186), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n8920), .CLK(n9224), .Q(
        g1389), .QN(n8655) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n8962), .CLK(n9277), .Q(
        test_so15), .QN(n8862) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n8883), .CLK(n9187), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n8933), .CLK(n9238), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n8933), .CLK(n9238), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n8902), .CLK(n9206), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n8902), .CLK(n9206), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n8868), .CLK(n9172), .Q(
        g5611) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n8950), .CLK(n9259), .Q(
        g16627), .QN(n8720) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n8908), .CLK(n9212), .Q(
        g4572) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n8970), .CLK(n9287), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n8889), .CLK(n9193), .Q(
        g2898) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n8933), .CLK(n9238), .Q(
        g3343), .QN(n8411) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n8959), .CLK(n9271), .Q(
        g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n8968), .CLK(n9285), .Q(
        test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n8952), .CLK(n9261), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n8972), .CLK(n9289), .Q(
        n9348), .QN(n15422) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n8869), .CLK(n9173), .Q(
        g4961) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n8957), .CLK(n9269), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n8960), .CLK(n9272), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n8881), .CLK(n9185), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n8877), .CLK(n9181), .Q(
        g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n8878), .CLK(n9182), .Q(
        g5802), .QN(n8322) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n8886), .CLK(n9190), .Q(
        g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n8909), .CLK(n9213), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n8930), .CLK(n9234), .Q(
        g681), .QN(n8678) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n8912), .CLK(n9216), .Q(
        g437) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n8927), .CLK(n9231), .Q(
        test_so17), .QN(n8846) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n8915), .CLK(n9219), 
        .Q(g5901) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n8889), .CLK(n9193), .Q(
        g2886) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n8874), .CLK(n9178), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n8874), .CLK(n9178), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n8923), .CLK(n9227), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n8875), .CLK(n9179), .Q(
        g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n8867), .CLK(n9171), .Q(
        g5092), .QN(n8697) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n8898), .CLK(n9202), .Q(
        g4831) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n8936), .CLK(n9242), .Q(
        g4382) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n8956), .CLK(n9268), .Q(
        g6386), .QN(n8412) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n8909), .CLK(n9213), .Q(
        g479), .QN(n8358) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n8873), .CLK(n9177), .Q(
        g3965) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n8884), .CLK(n9188), .Q(
        test_so18) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n8918), .CLK(n9222), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n8940), .CLK(n9248), .Q(
        g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n8902), .CLK(n9206), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n8885), .CLK(n9189), .Q(
        g222) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n8920), .CLK(n9224), .Q(
        g3050) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n8920), .CLK(n9224), .Q(
        g1052) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n8920), .CLK(n9224), .Q(
        g17580), .QN(n8702) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n8941), .CLK(n9249), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n8913), .CLK(n9217), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n8913), .CLK(n9217), .Q(
        g5889) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n8908), .CLK(n9212), .Q(
        g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n8908), .CLK(n9212), .Q(
        g8719), .QN(n8690) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n8871), .CLK(n9175), .Q(
        test_so19), .QN(n8854) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n8955), .CLK(n9266), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n8963), .CLK(n9278), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n8880), .CLK(n9184), .Q(
        g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n8873), .CLK(n9177), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n8955), .CLK(n9266), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n8955), .CLK(n9266), .Q(
        g4917) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n8887), .CLK(n9191), .Q(
        g1070), .QN(n8792) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n8909), .CLK(n9213), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n8936), .CLK(n9242), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n8926), .CLK(n9230), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n8965), .CLK(n9282), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n8894), .CLK(n9198), .Q(
        g4164), .QN(n8516) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n8946), .CLK(n9254), .Q(
        test_so20) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n8881), .CLK(n9185), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n8961), .CLK(n9275), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n8879), .CLK(n9183), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n8879), .CLK(n9183), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n8879), .CLK(n9183), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n8923), .CLK(n9227), .Q(
        g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n8908), .CLK(n9212), .Q(
        g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n8963), .CLK(n9278), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n8875), .CLK(n9179), .Q(
        g1682), .QN(n8352) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n8962), .CLK(n9277), .Q(
        g355) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n8962), .CLK(n9277), .Q(
        g1087), .QN(n8543) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n8907), .CLK(n9211), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n8947), .CLK(n9256), .Q(
        test_so21), .QN(n8830) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n8900), .CLK(n9204), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n8950), .CLK(n9259), .Q(
        g3802), .QN(n8318) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n8959), .CLK(n9271), .Q(
        g6159), .QN(n8696) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n8959), .CLK(n9271), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n8881), .CLK(n9185), .Q(
        g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n8926), .CLK(n9230), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n8802), .SI(g911), .SE(n8879), .CLK(n9183), .Q(g43) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n8880), .CLK(n9184), .Q(
        g16775), .QN(n8666) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n8907), .CLK(n9211), .Q(
        g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n8874), .CLK(n9178), .Q(
        g5551) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n8916), .CLK(n9220), .Q(
        g3558) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n8961), .CLK(n9275), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n8890), .CLK(n9194), .Q(
        test_so22), .QN(n8850) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n8891), .CLK(n9195), 
        .Q(g3901) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n8972), .CLK(n9289), .Q(
        g4888) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n8899), .CLK(n9203), .Q(
        g6251) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n8943), .CLK(n9251), .Q(
        g17649), .QN(n8708) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n8920), .CLK(n9224), .Q(
        g1373), .QN(n8657) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n8920), .CLK(n9224), .Q(
        g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n8905), .CLK(n9209), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n8876), .CLK(n9180), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n8931), .CLK(n9235), .Q(
        g4281), .QN(n8541) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n8916), .CLK(n9220), .Q(
        g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n8971), .CLK(n9288), .Q(
        g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n8971), .CLK(n9288), .Q(
        g1283) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n8912), .CLK(n9216), .Q(
        test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n8882), .CLK(n9186), .Q(g4297), .QN(n8750) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n8883), .CLK(n9187), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n8887), .CLK(n9191), .Q(
        g13272), .QN(n8741) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n8943), .CLK(n9251), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(g34025), .SI(g758), .SE(n8943), .CLK(n9251), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n8885), .CLK(n9189), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n8885), .CLK(n9189), .Q(
        g5543) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n8885), .CLK(n9189), .Q(
        g8475), .QN(n8740) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n8898), .CLK(n9202), .Q(
        g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n8966), .CLK(n9283), .Q(
        g6243) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n8925), .CLK(n9229), .Q(
        n9340), .QN(n15421) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n8925), .CLK(n9229), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n8951), .CLK(n9260), .Q(
        test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n8970), .CLK(n9287), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n8919), .CLK(n9223), .Q(
        g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n8925), .CLK(n9229), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n8928), .CLK(n9232), .Q(
        g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n8912), .CLK(n9216), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n8880), .CLK(n9184), .Q(
        g4049), .QN(n8746) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n8969), .CLK(n9286), .Q(
        g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n8886), .CLK(n9190), .Q(
        g2932) );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(n8898), .CLK(n9202), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n8948), .CLK(n9257), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n8954), .CLK(n9264), .Q(
        g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n8962), .CLK(n9277), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n8867), .CLK(n9171), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n8970), .CLK(n9287), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n8909), .CLK(n9213), .Q(
        g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n8939), .CLK(n9246), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n8884), .CLK(n9188), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n8965), .CLK(n9282), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n8883), .CLK(n9187), .Q(
        g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n8913), .CLK(n9217), .Q(
        g239), .QN(n8659) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n8913), .CLK(n9217), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n8869), .CLK(n9173), .Q(
        g2848) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n8968), .CLK(n9285), .Q(
        g5022), .QN(n8767) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n8968), .CLK(n9285), .Q(
        g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n8922), .CLK(n9226), .Q(
        g1030), .QN(n8656) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n8923), .CLK(n9227), .Q(
        test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n8957), .CLK(n9269), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n8922), .CLK(n9226), .Q(
        g9817), .QN(n8313) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n8922), .CLK(n9226), .Q(
        g1430), .QN(n8544) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n8969), .CLK(n9286), .Q(
        n9336) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n8903), .CLK(n9207), .Q(
        g2241), .QN(n8351) );
  SDFFX1 DFF_375_Q_reg ( .D(n706), .SI(g2241), .SE(n8970), .CLK(n9287), .Q(
        g1564), .QN(n8729) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n8878), .CLK(n9182), .Q(
        g9680), .QN(n8321) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n8878), .CLK(n9182), 
        .Q(g6148), .QN(n8311) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n8967), .CLK(n9284), .Q(
        g6649) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n8919), .CLK(n9223), .Q(
        g110), .QN(n8800) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n8932), .CLK(n9237), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n8889), .CLK(n9193), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n8960), .CLK(n9272), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n8954), .CLK(n9264), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n8954), .CLK(n9264), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n8969), .CLK(n9286), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n8901), .CLK(n9205), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n8960), .CLK(n9272), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n8894), .CLK(n9198), .Q(
        g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n8894), .CLK(n9198), .Q(
        g5208) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n8868), .CLK(n9172), .Q(
        g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n8953), .CLK(n9263), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n8931), .CLK(n9235), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n8878), .CLK(n9182), .Q(
        g5752) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n8966), .CLK(n9283), .Q(
        g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n8914), .CLK(n9218), .Q(
        test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n8906), .CLK(n9210), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n8879), .CLK(n9183), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n8880), .CLK(n9184), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n8910), .CLK(n9214), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n8932), .CLK(n9237), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n8932), .CLK(n9237), .Q(
        g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n8947), .CLK(n9256), .Q(
        g2370), .QN(n8630) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n8947), .CLK(n9256), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n8947), .CLK(n9256), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n8905), .CLK(n9209), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n8949), .CLK(n9258), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n8949), .CLK(n9258), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n8949), .CLK(n9258), .Q(
        test_so29), .QN(n8836) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n8890), .CLK(n9194), 
        .Q(g2984) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n8872), .CLK(n9176), .Q(
        g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n8900), .CLK(n9204), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n8878), .CLK(n9182), .Q(
        g101), .QN(n8619) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n8878), .CLK(n9182), .Q(
        g8918) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n8952), .CLK(n9261), .Q(
        g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n8886), .CLK(n9190), .Q(
        n9332) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n8887), .CLK(n9191), .Q(
        g1018), .QN(n8653) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n8897), .CLK(n9201), .Q(
        g17320), .QN(n8735) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n8880), .CLK(n9184), .Q(
        g4045), .QN(n8416) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n8880), .CLK(n9184), .Q(
        g1467), .QN(n5693) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n8881), .CLK(n9185), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n8941), .CLK(n9249), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n8915), .CLK(n9219), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n8893), .CLK(n9197), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n8911), .CLK(n9215), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n8893), .CLK(n9197), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n8893), .CLK(n9197), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n8907), .CLK(n9211), .Q(
        g1816), .QN(n8300) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n8944), .CLK(n9252), .Q(
        g4369) );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(n8945), .CLK(n9253), .Q(
        g4578), .QN(n8775) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n8945), .CLK(n9253), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n8873), .CLK(n9177), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n8880), .CLK(n9184), .Q(
        g2514), .QN(n8330) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n8965), .CLK(n9282), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n8972), .CLK(n9289), .Q(
        test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n8875), .CLK(n9179), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n8919), .CLK(n9223), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n8935), .CLK(n9241), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n8904), .CLK(n9208), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n8896), .CLK(n9200), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n8941), .CLK(n9249), .Q(
        g2763), .QN(n8284) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n8949), .CLK(n9258), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n8949), .CLK(n9258), .Q(
        g952), .QN(n8276) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n8893), .CLK(n9197), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n8927), .CLK(n9231), .Q(
        g1950), .QN(n8350) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n8896), .CLK(n9200), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n8901), .CLK(n9205), .Q(
        g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n8938), .CLK(n9244), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n8871), .CLK(n9175), 
        .Q(g8398), .QN(n8317) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n8871), .CLK(n9175), .Q(
        g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n8904), .CLK(n9208), .Q(
        g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n8883), .CLK(n9187), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n8929), .CLK(n9233), .Q(
        g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n8918), .CLK(n9222), .Q(
        g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n8949), .CLK(n9258), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n8950), .CLK(n9259), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n8901), .CLK(n9205), .Q(
        g2315) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n8897), .CLK(n9201), .Q(
        g2811), .QN(n8295) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n8897), .CLK(n9201), .Q(
        g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n8921), .CLK(n9225), .Q(
        g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n8921), .CLK(n9225), .Q(
        test_so33), .QN(n8823) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n8943), .CLK(n9251), 
        .Q(g17760), .QN(n8665) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n8870), .CLK(n9174), .Q(
        g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n8871), .CLK(n9175), .Q(
        n9327) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n8871), .CLK(n9175), .Q(
        g3752) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n8902), .CLK(n9206), .Q(
        g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n8931), .CLK(n9235), 
        .Q(g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n8931), .CLK(n9235), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n8936), .CLK(n9242), .Q(
        g4388), .QN(n8731) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n8900), .CLK(n9204), .Q(
        g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n8900), .CLK(n9204), .Q(
        g6311) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n8900), .CLK(n9204), .Q(
        g8916) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n8900), .CLK(n9204), .Q(
        g1041), .QN(n8765) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n8910), .CLK(n9214), .Q(
        test_so34), .QN(n8856) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n8910), .CLK(n9214), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n8877), .CLK(n9181), .Q(
        g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n8877), .CLK(n9181), .Q(
        g4430), .QN(n8728) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n8898), .CLK(n9202), .Q(
        n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n8898), .CLK(n9202), .Q(
        g4826), .QN(n8337) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n8899), .CLK(n9203), .Q(
        g6239) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n8906), .CLK(n9210), .Q(
        g232), .QN(n8658) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n8895), .CLK(n9199), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n8895), .CLK(n9199), .Q(
        g6545) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n8888), .CLK(n9192), .Q(
        n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n8888), .CLK(n9192), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n8912), .CLK(n9216), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n8912), .CLK(n9216), .Q(
        test_so35), .QN(n8315) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n8928), .CLK(n9232), 
        .Q(g1890) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n8962), .CLK(n9277), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n8927), .CLK(n9231), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n8927), .CLK(n9231), .Q(
        g2130) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n8948), .CLK(n9257), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n8949), .CLK(n9258), .Q(
        g4308), .QN(n8542) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n8912), .CLK(n9216), .Q(
        g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n8933), .CLK(n9238), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n8933), .CLK(n9238), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n8869), .CLK(n9173), .Q(
        n9322) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(n8869), .CLK(n9173), .Q(
        g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n8869), .CLK(n9173), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n8954), .CLK(n9264), .Q(
        test_so36), .QN(n8832) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n8928), .CLK(n9232), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n8928), .CLK(n9232), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n8892), .CLK(n9196), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n8909), .CLK(n9213), .Q(
        g832), .QN(n8545) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n8914), .CLK(n9218), .Q(
        g5897) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n8914), .CLK(n9218), .Q(
        g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n8898), .CLK(n9202), .Q(
        g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n8938), .CLK(n9244), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n8938), .CLK(n9244), .Q(
        g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n8890), .CLK(n9194), .Q(
        g2902), .QN(n8365) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n8962), .CLK(n9277), .Q(
        g333) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n8963), .CLK(n9278), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n8881), .CLK(n9185), .Q(
        test_so37) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n8971), .CLK(n9288), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n8870), .CLK(n9174), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n8932), .CLK(n9237), .Q(
        g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n8932), .CLK(n9237), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n8912), .CLK(n9216), .Q(
        g5406) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n8912), .CLK(n9216), .Q(
        g269), .QN(n8660) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n8912), .CLK(n9216), .Q(
        g401) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n8912), .CLK(n9216), .Q(
        g6040), .QN(n8413) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n8912), .CLK(n9216), .Q(
        g441) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n8911), .CLK(n9215), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n8873), .CLK(n9177), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n8873), .CLK(n9177), .Q(
        g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n8944), .CLK(n9252), .Q(
        test_so38), .QN(n8838) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n8891), .CLK(n9195), 
        .Q(g3957) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n8948), .CLK(n9257), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n8888), .CLK(n9192), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n8943), .CLK(n9251), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n8905), .CLK(n9209), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n8965), .CLK(n9282), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n8924), .CLK(n9228), .Q(
        g3498), .QN(n5740) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n8924), .CLK(n9228), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n8906), .CLK(n9210), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n8906), .CLK(n9210), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n8933), .CLK(n9238), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n8875), .CLK(n9179), .Q(
        g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n8942), .CLK(n9250), .Q(
        test_so39), .QN(n8649) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n8943), .CLK(n9251), 
        .Q(g17577), .QN(n8703) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n8963), .CLK(n9278), .Q(
        g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n8972), .CLK(n9289), .Q(
        g2652), .QN(n8622) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n8897), .CLK(n9201), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n8902), .CLK(n9206), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n8960), .CLK(n9272), .Q(
        g661), .QN(n8381) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n8870), .CLK(n9174), .Q(
        g4950) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n8870), .CLK(n9174), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n8881), .CLK(n9185), .Q(
        g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n8882), .CLK(n9186), .Q(
        g1361), .QN(n8654) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n8955), .CLK(n9266), .Q(
        g6235) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n8955), .CLK(n9266), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n8906), .CLK(n9210), .Q(
        test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n8905), .CLK(n9209), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n8919), .CLK(n9223), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n8952), .CLK(n9261), .Q(
        g6555), .QN(n8643) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n8906), .CLK(n9210), .Q(
        g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n8950), .CLK(n9259), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n8908), .CLK(n9212), .Q(
        g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n8874), .CLK(n9178), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n8903), .CLK(n9207), .Q(
        g3897) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n8967), .CLK(n9284), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n8910), .CLK(n9214), .Q(
        g2606), .QN(n5311) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n8880), .CLK(n9184), .Q(
        g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n8877), .CLK(n9181), .Q(
        test_so41) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n8930), .CLK(n9234), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n8883), .CLK(n9187), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n8933), .CLK(n9238), .Q(
        g13259), .QN(n8748) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n8933), .CLK(n9238), .Q(
        g405), .QN(n8674) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n8895), .CLK(n9199), .Q(
        g5216) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n8952), .CLK(n9261), .Q(
        g6494), .QN(n8314) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n8871), .CLK(n9175), .Q(
        g4669) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n8946), .CLK(n9254), .Q(
        g996), .QN(n8373) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n8871), .CLK(n9175), .Q(
        g4531), .QN(n8742) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n8886), .CLK(n9190), .Q(
        g2860) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n8884), .CLK(n9188), .Q(
        g4743) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n8929), .CLK(n9233), .Q(
        g6593) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n8929), .CLK(n9233), .Q(
        test_so42), .QN(n8547) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n8877), .CLK(n9181), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n8882), .CLK(n9186), .Q(
        g1413), .QN(n8791) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n8944), .CLK(n9252), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n8944), .CLK(n9252), .Q(
        g13039), .QN(n8704) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n8952), .CLK(n9261), .Q(
        g6641) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n8952), .CLK(n9261), .Q(
        g6) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n8935), .CLK(n9241), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n8801), .SI(g1936), .SE(n8935), .CLK(n9241), .Q(
        g55), .QN(n8273) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n8935), .CLK(n9241), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n8910), .CLK(n9214), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n8953), .CLK(n9263), .Q(
        g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n8901), .CLK(n9205), .Q(
        n9314) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n8916), .CLK(n9220), .Q(
        test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n8874), .CLK(n9178), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n8917), .CLK(n9221), .Q(
        g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n8917), .CLK(n9221), .Q(
        g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n8915), .CLK(n9219), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n8915), .CLK(n9219), .Q(
        g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n8899), .CLK(n9203), .Q(
        g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n8946), .CLK(n9254), .Q(
        g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n8901), .CLK(n9205), .Q(
        g2380), .QN(n8329) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n8953), .CLK(n9263), .Q(
        g5196) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n8960), .CLK(n9272), .Q(
        g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n8918), .CLK(n9222), .Q(
        n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n8918), .CLK(n9222), .Q(
        g14518), .QN(n8713) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n8918), .CLK(n9222), .Q(
        test_so44), .QN(n8841) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n8934), .CLK(n9239), 
        .Q(g6541), .QN(n5739) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n8959), .CLK(n9271), .Q(
        g3203) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n8962), .CLK(n9277), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n8913), .CLK(n9217), .Q(
        g4760) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n8913), .CLK(n9217), .Q(
        g262), .QN(n8662) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n8963), .CLK(n9278), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n8891), .CLK(n9195), .Q(
        g5467), .QN(n8725) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n8891), .CLK(n9195), .Q(
        g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n8954), .CLK(n9264), .Q(
        g6209), .QN(n8641) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n8927), .CLK(n9231), .Q(
        g29211), .QN(n8688) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n8927), .CLK(n9231), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n8930), .CLK(n9234), .Q(
        g655), .QN(n8784) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n8931), .CLK(n9235), .Q(
        test_so45) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n8897), .CLK(n9201), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n8947), .CLK(n9256), .Q(
        g5256) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n8948), .CLK(n9257), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n8948), .CLK(n9257), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n8968), .CLK(n9285), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n8968), .CLK(n9285), .Q(
        g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n8923), .CLK(n9227), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n8972), .CLK(n9289), .Q(
        g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n8892), .CLK(n9196), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n8892), .CLK(n9196), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n8957), .CLK(n9269), .Q(
        g3247) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n8921), .CLK(n9225), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n8921), .CLK(n9225), .Q(
        test_so46) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n8894), .CLK(n9198), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n8944), .CLK(n9252), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n8933), .CLK(n9238), .Q(
        g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n8938), .CLK(n9244), .Q(
        g4732) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n8938), .CLK(n9244), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n8883), .CLK(n9187), .Q(
        g5817), .QN(n8782) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n8947), .CLK(n9256), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n8929), .CLK(n9233), .Q(
        g2648), .QN(n8333) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n8971), .CLK(n9288), .Q(
        g6736), .QN(n8753) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n8869), .CLK(n9173), .Q(
        g4944) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n8926), .CLK(n9230), .Q(
        g4072) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n8926), .CLK(n9230), .Q(
        g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n8967), .CLK(n9284), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(n178), .SI(test_si48), .SE(n8874), .CLK(n9178), 
        .Q(g3466), .QN(n8760) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n8893), .CLK(n9197), .Q(
        g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n8969), .CLK(n9286), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n8969), .CLK(n9286), .Q(
        g4434), .QN(n8343) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n8970), .CLK(n9287), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n8904), .CLK(n9208), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n8958), .CLK(n9270), .Q(
        g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n8922), .CLK(n9226), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n8922), .CLK(n9226), .Q(
        g3333), .QN(n8340) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n8922), .CLK(n9226), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n8946), .CLK(n9254), .Q(
        g4681), .QN(n8553) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n8884), .CLK(n9188), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n8962), .CLK(n9277), .Q(
        test_so48), .QN(n8860) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n8934), .CLK(n9239), 
        .Q(g8789), .QN(n8652) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n8928), .CLK(n9232), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n8886), .CLK(n9190), .Q(
        g2988) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n8952), .CLK(n9261), .Q(
        g3538) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n8905), .CLK(n9209), .Q(
        g301) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n8905), .CLK(n9209), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n8909), .CLK(n9213), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n8913), .CLK(n9217), .Q(
        g17291), .QN(n8699) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n8962), .CLK(n9277), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n8908), .CLK(n9212), .Q(
        g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n8885), .CLK(n9189), .Q(
        g199) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n8885), .CLK(n9189), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n8937), .CLK(n9243), .Q(
        test_so49), .QN(n8819) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n8958), .CLK(n9270), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n8892), .CLK(n9196), .Q(
        g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n8957), .CLK(n9269), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n8957), .CLK(n9269), .Q(
        g4922) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n8867), .CLK(n9171), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n8953), .CLK(n9263), .Q(
        g5863), .QN(n8638) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n8953), .CLK(n9263), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n8953), .CLK(n9263), .Q(
        g2518), .QN(n8624) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n8929), .CLK(n9233), .Q(
        g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n8927), .CLK(n9231), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n8928), .CLK(n9232), .Q(
        g3263) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n8928), .CLK(n9232), .Q(
        g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n8957), .CLK(n9269), .Q(
        test_so50), .QN(n8844) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n8971), .CLK(n9288), 
        .Q(g6444) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n8906), .CLK(n9210), .Q(
        g2965), .QN(n8366) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n8953), .CLK(n9263), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n8875), .CLK(n9179), .Q(
        n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n8889), .CLK(n9193), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n8925), .CLK(n9229), .Q(
        g17646), .QN(n8761) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n8916), .CLK(n9220), .Q(
        g3562) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n8882), .CLK(n9186), .Q(
        g10122_Tj), .QN(n8749) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n8910), .CLK(n9214), 
        .Q(g1404), .QN(n8757) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n8873), .CLK(n9177), .Q(
        g3817), .QN(n8759) );
  SDFFX1 DFF_743_Q_reg ( .D(n8806), .SI(g3817), .SE(n8884), .CLK(n9188), .Q(
        n9302) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n8884), .CLK(n9188), .Q(
        g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n8884), .CLK(n9188), .Q(
        test_so51), .QN(n8855) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n8940), .CLK(n9248), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n8896), .CLK(n9200), .Q(
        g4704) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n8889), .CLK(n9193), .Q(
        g2878) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n8895), .CLK(n9199), .Q(
        g5220) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n8924), .CLK(n9228), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n8925), .CLK(n9229), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n8937), .CLK(n9243), .Q(
        g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n8893), .CLK(n9197), .Q(
        g1277) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n8893), .CLK(n9197), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n8935), .CLK(n9241), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n8889), .CLK(n9193), .Q(
        g2882) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n8970), .CLK(n9287), .Q(
        test_so52) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n8934), .CLK(n9239), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n8935), .CLK(n9241), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n8886), .CLK(n9190), .Q(g8) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n8897), .CLK(n9201), .Q(
        g2799), .QN(n8292) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n8932), .CLK(n9237), .Q(
        g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n8932), .CLK(n9237), .Q(
        g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n8957), .CLK(n9269), .Q(
        g4912) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n8894), .CLK(n9198), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n8911), .CLK(n9215), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n8964), .CLK(n9279), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n8877), .CLK(n9181), .Q(
        g550), .QN(n8537) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n8906), .CLK(n9210), .Q(
        g255), .QN(n8661) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n8967), .CLK(n9284), .Q(
        test_so53), .QN(n8849) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n8947), .CLK(n9256), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n8947), .CLK(n9256), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n8949), .CLK(n9258), .Q(
        g3863), .QN(n8639) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n8967), .CLK(n9284), .Q(
        g1959), .QN(n8625) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n8874), .CLK(n9178), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n8908), .CLK(n9212), .Q(
        g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n8965), .CLK(n9282), .Q(
        g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n8889), .CLK(n9193), .Q(
        g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n8902), .CLK(n9206), .Q(
        g4894) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n8902), .CLK(n9206), .Q(
        g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n8902), .CLK(n9206), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n8902), .CLK(n9206), .Q(
        g16693), .QN(n8712) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n8962), .CLK(n9277), .Q(
        test_so54) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n8887), .CLK(n9191), 
        .Q(g1002), .QN(n8796) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n8945), .CLK(n9253), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n8945), .CLK(n9253), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n8945), .CLK(n9253), .Q(
        g1236), .QN(n8359) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n8945), .CLK(n9253), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n8951), .CLK(n9260), .Q(
        g2476), .QN(n8773) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n8919), .CLK(n9223), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n8901), .CLK(n9205), .Q(
        g2375), .QN(n8349) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n8871), .CLK(n9175), .Q(
        g63), .QN(n8675) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n8883), .CLK(n9187), .Q(
        g17739), .QN(n8667) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n8908), .CLK(n9212), .Q(
        g358), .QN(n8788) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n8889), .CLK(n9193), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n8973), .CLK(n9290), .Q(
        test_so55), .QN(n8847) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n8956), .CLK(n9268), 
        .Q(g3161), .QN(n8644) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n8961), .CLK(n9275), .Q(
        g2384), .QN(n8629) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n8921), .CLK(n9225), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n8958), .CLK(n9270), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n8898), .CLK(n9202), .Q(
        g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n8918), .CLK(n9222), .Q(
        g2024) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n8951), .CLK(n9260), .Q(
        g3451), .QN(n8302) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n8876), .CLK(n9180), .Q(
        g2795), .QN(n8293) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n8924), .CLK(n9228), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n8872), .CLK(n9176), .Q(
        g4527), .QN(n8514) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n8888), .CLK(n9192), .Q(
        g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n8914), .CLK(n9218), .Q(
        g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n8969), .CLK(n9286), .Q(
        test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n8953), .CLK(n9263), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n8938), .CLK(n9244), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n8929), .CLK(n9233), .Q(
        g2643), .QN(n8348) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n8937), .CLK(n9243), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n8964), .CLK(n9279), .Q(
        g8358), .QN(n8374) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n8911), .CLK(n9215), .Q(
        n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n8911), .CLK(n9215), .Q(
        g5156), .QN(n5734) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n8925), .CLK(n9229), .Q(
        g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n8925), .CLK(n9229), .Q(
        n9294) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n8951), .CLK(n9260), .Q(
        g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n8931), .CLK(n9235), .Q(
        g8839), .QN(n8513) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n8927), .CLK(n9231), .Q(
        g1955), .QN(n8326) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n8958), .CLK(n9270), .Q(
        test_so57), .QN(n8835) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n8965), .CLK(n9282), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n8965), .CLK(n9282), .Q(
        g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n8971), .CLK(n9288), .Q(
        g4771) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n8878), .CLK(n9182), .Q(
        g6098) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n8956), .CLK(n9268), .Q(
        g3147), .QN(n5738) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n8932), .CLK(n9237), .Q(
        g3347), .QN(n8743) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n8964), .CLK(n9279), .Q(
        g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n8964), .CLK(n9279), .Q(
        g191), .QN(n8375) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n8964), .CLK(n9279), .Q(
        g2712), .QN(n8751) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n8925), .CLK(n9229), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n8896), .CLK(n9200), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n8940), .CLK(n9248), .Q(
        test_so58), .QN(n8837) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n8915), .CLK(n9219), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n8915), .CLK(n9219), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n8890), .CLK(n9194), .Q(
        g2927), .QN(n8363) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n8938), .CLK(n9244), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n8897), .CLK(n9201), .Q(
        g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n8957), .CLK(n9269), .Q(
        g4907) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n8957), .CLK(n9269), .Q(
        g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n8961), .CLK(n9275), .Q(
        g4035), .QN(n8341) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n8931), .CLK(n9235), .Q(
        g2946) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n8926), .CLK(n9230), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n8926), .CLK(n9230), .Q(
        g4082), .QN(n8677) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n8952), .CLK(n9261), .Q(
        g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n8918), .CLK(n9222), .Q(
        test_so59), .QN(n8857) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n8924), .CLK(n9228), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n8875), .CLK(n9179), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n8876), .CLK(n9180), .Q(
        g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n8876), .CLK(n9180), .Q(
        g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n8970), .CLK(n9287), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n8903), .CLK(n9207), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n8909), .CLK(n9213), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n8910), .CLK(n9214), .Q(
        g1249), .QN(n8770) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n8892), .CLK(n9196), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n8950), .CLK(n9259), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n8924), .CLK(n9228), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n8869), .CLK(n9173), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n8941), .CLK(n9249), .Q(
        test_so60), .QN(n8853) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n8914), .CLK(n9218), 
        .Q(g5949) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n8902), .CLK(n9206), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n8925), .CLK(n9229), .Q(
        g904), .QN(n8771) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n8886), .CLK(n9190), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n8961), .CLK(n9275), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n8867), .CLK(n9171), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n8874), .CLK(n9178), .Q(
        g5603) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n8872), .CLK(n9176), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n8971), .CLK(n9288), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n8881), .CLK(n9185), .Q(
        g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n8919), .CLK(n9223), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n8919), .CLK(n9223), .Q(
        g2208), .QN(n8721) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n8910), .CLK(n9214), .Q(
        test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n8893), .CLK(n9197), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n8940), .CLK(n9248), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n8940), .CLK(n9248), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n8949), .CLK(n9258), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n8868), .CLK(n9172), .Q(
        g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n8946), .CLK(n9254), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n8956), .CLK(n9268), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n8956), .CLK(n9268), .Q(
        g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n8890), .CLK(n9194), .Q(
        g2917), .QN(n8364) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n8892), .CLK(n9196), .Q(
        g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n8893), .CLK(n9197), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n8876), .CLK(n9180), .Q(
        g671), .QN(n8307) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n8964), .CLK(n9279), .Q(
        test_so62), .QN(n8861) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n8899), .CLK(n9203), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n8942), .CLK(n9250), .Q(
        g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n8942), .CLK(n9250), .Q(
        g17519), .QN(n8705) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n8942), .CLK(n9250), .Q(
        g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n8879), .CLK(n9183), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n8960), .CLK(n9272), .Q(
        g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n8963), .CLK(n9278), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n8893), .CLK(n9197), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n8940), .CLK(n9248), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n8954), .CLK(n9264), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n8891), .CLK(n9195), .Q(
        g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n8891), .CLK(n9195), .Q(
        g5503), .QN(n5737) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n8872), .CLK(n9176), .Q(
        test_so63) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n8915), .CLK(n9219), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n8934), .CLK(n9239), .Q(
        g1124), .QN(n5692) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n8869), .CLK(n9173), .Q(
        g4955) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n8947), .CLK(n9256), .Q(
        g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n8918), .CLK(n9222), .Q(
        g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n8954), .CLK(n9264), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n8911), .CLK(n9215), .Q(
        g5120), .QN(n8726) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n8911), .CLK(n9215), .Q(
        g17674), .QN(n8670) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n8901), .CLK(n9205), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n8968), .CLK(n9285), .Q(
        g4438) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n8880), .CLK(n9184), .Q(
        g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n8876), .CLK(n9180), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n8971), .CLK(n9288), .Q(
        test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n8870), .CLK(n9174), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n8939), .CLK(n9246), .Q(
        g18881) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n8939), .CLK(n9246), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n8887), .CLK(n9191), .Q(
        g1199), .QN(n8379) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n8887), .CLK(n9191), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n8875), .CLK(n9179), .Q(
        g5547) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n8875), .CLK(n9179), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n8950), .CLK(n9259), .Q(
        g16744), .QN(n8663) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n8966), .CLK(n9283), .Q(
        g2338), .QN(n5310) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n8966), .CLK(n9283), .Q(
        g8919) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n8899), .CLK(n9203), .Q(
        g6247) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n8876), .CLK(n9180), .Q(
        g2791), .QN(n8294) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n8902), .CLK(n9206), .Q(
        test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n8867), .CLK(n9171), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n8897), .CLK(n9201), .Q(
        g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n8930), .CLK(n9234), .Q(
        g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n8941), .CLK(n9249), .Q(
        g2759), .QN(n8793) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n8902), .CLK(n9206), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n8946), .CLK(n9254), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n8893), .CLK(n9197), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n8874), .CLK(n9178), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n8929), .CLK(n9233), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n8952), .CLK(n9261), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n8957), .CLK(n9269), .Q(
        g5517), .QN(n8640) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n8881), .CLK(n9185), .Q(
        g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n8910), .CLK(n9214), .Q(
        test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n8939), .CLK(n9246), 
        .Q(n9281), .QN(DFF_961_n1) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n8904), .CLK(n9208), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n8926), .CLK(n9230), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n8918), .CLK(n9222), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n8944), .CLK(n9252), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n8924), .CLK(n9228), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n8952), .CLK(n9261), .Q(
        g6589) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n8928), .CLK(n9232), .Q(
        n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n8942), .CLK(n9250), .Q(
        g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n8964), .CLK(n9279), .Q(
        g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n8912), .CLK(n9216), .Q(
        g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n8927), .CLK(n9231), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n8927), .CLK(n9231), .Q(
        test_so67) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n8972), .CLK(n9289), 
        .Q(g1825), .QN(n8631) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n8887), .CLK(n9191), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n8936), .CLK(n9242), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n8936), .CLK(n9242), 
        .Q(g8283), .QN(n8683) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n8916), .CLK(n9220), .Q(
        g3546) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n8895), .CLK(n9199), .Q(
        g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n8888), .CLK(n9192), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n8939), .CLK(n9246), .Q(
        g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n8891), .CLK(n9195), .Q(
        g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n8905), .CLK(n9209), .Q(
        g6509), .QN(n8737) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n8905), .CLK(n9209), .Q(
        g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n8951), .CLK(n9260), .Q(
        g2504), .QN(n8623) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n8951), .CLK(n9260), .Q(
        test_so68), .QN(n8824) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n8872), .CLK(n9176), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n8872), .CLK(n9176), .Q(
        g8917) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n8941), .CLK(n9249), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n8917), .CLK(n9221), .Q(
        g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n8917), .CLK(n9221), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n8917), .CLK(n9221), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n8942), .CLK(n9250), .Q(
        g8235), .QN(n8681) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n8894), .CLK(n9198), .Q(
        g4176) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n8880), .CLK(n9184), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n8936), .CLK(n9242), .Q(
        g4405) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n8936), .CLK(n9242), .Q(
        g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n8879), .CLK(n9183), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n8956), .CLK(n9268), .Q(
        test_so69), .QN(n8829) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n8879), .CLK(n9183), 
        .Q(g4765) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n8868), .CLK(n9172), .Q(
        g5563) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n8951), .CLK(n9260), .Q(
        g1395) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n8934), .CLK(n9239), .Q(
        g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n8966), .CLK(n9283), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n8966), .CLK(n9283), .Q(
        g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n8872), .CLK(n9176), .Q(
        n9276) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n8872), .CLK(n9176), .Q(
        g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n8926), .CLK(n9230), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n8944), .CLK(n9252), .Q(
        g4473), .QN(n8752) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n8944), .CLK(n9252), .Q(
        g1266), .QN(n8369) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n8960), .CLK(n9272), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n8877), .CLK(n9181), .Q(
        test_so70), .QN(n8852) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n8941), .CLK(n9249), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n8869), .CLK(n9173), .Q(
        g5471), .QN(n8780) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n8968), .CLK(n9285), .Q(
        g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n8969), .CLK(n9286), .Q(
        g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n8969), .CLK(n9286), .Q(
        g6605) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n8881), .CLK(n9185), .Q(
        n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n8904), .CLK(n9208), .Q(
        g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n8931), .CLK(n9235), .Q(
        g9019), .QN(n8512) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n8951), .CLK(n9260), .Q(
        g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n8939), .CLK(n9246), .Q(
        g4849), .QN(n8766) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n8903), .CLK(n9207), .Q(
        g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n8904), .CLK(n9208), .Q(
        n9273) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n8904), .CLK(n9208), .Q(
        test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n8888), .CLK(n9192), 
        .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n8888), .CLK(n9192), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n8886), .CLK(n9190), .Q(
        g2868), .QN(n8680) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n8876), .CLK(n9180), .Q(
        g2767), .QN(n8297) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n8961), .CLK(n9275), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n8961), .CLK(n9275), .Q(
        g16718), .QN(n8664) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n8932), .CLK(n9237), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n8930), .CLK(n9234), .Q(
        g5212) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n8930), .CLK(n9234), .Q(
        g4245) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n8930), .CLK(n9234), .Q(
        g645) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n8931), .CLK(n9235), .Q(
        g4291), .QN(n8540) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n8963), .CLK(n9278), .Q(
        g29212), .QN(n5657) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n8963), .CLK(n9278), 
        .Q(test_so72), .QN(n8834) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n8934), .CLK(n9239), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n8934), .CLK(n9239), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n8934), .CLK(n9239), .Q(
        g8788), .QN(n8651) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n8903), .CLK(n9207), .Q(
        g2246), .QN(n8332) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n8888), .CLK(n9192), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n8916), .CLK(n9220), .Q(
        g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n8892), .CLK(n9196), .Q(
        g392), .QN(n8673) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n8962), .CLK(n9277), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n8934), .CLK(n9239), .Q(
        g6505), .QN(n8695) );
  SDFFX1 DFF_1057_Q_reg ( .D(n297), .SI(g6505), .SE(n8934), .CLK(n9239), .Q(
        g1221), .QN(n8730) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n8914), .CLK(n9218), .Q(
        g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n8906), .CLK(n9210), .Q(
        g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n8972), .CLK(n9289), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n8929), .CLK(
        n9233), .Q(g218), .QN(n8548) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n8946), .CLK(n9254), .Q(
        g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n8946), .CLK(n9254), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n8911), .CLK(n9215), .Q(
        g5062), .QN(n8768) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n8868), .CLK(n9172), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n8868), .CLK(n9172), .Q(
        g2689) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n8952), .CLK(n9261), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n8919), .CLK(n9223), .Q(
        g1677), .QN(n8628) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n8918), .CLK(n9222), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n8870), .CLK(n9174), .Q(
        g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n8931), .CLK(n9235), .Q(
        g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n8936), .CLK(n9242), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n8801), .SI(g7243), .SE(n8963), .CLK(n9278), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n8888), .CLK(n9192), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n8867), .CLK(n9171), .Q(
        g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n8867), .CLK(n9171), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n8940), .CLK(n9248), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n8940), .CLK(n9248), .Q(
        g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n8972), .CLK(n9289), 
        .Q(g2638), .QN(n8621) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n8894), .CLK(n9198), .Q(
        g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n8955), .CLK(n9266), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n8915), .CLK(n9219), .Q(
        g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n8915), .CLK(n9219), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n8915), .CLK(n9219), .Q(
        g13068), .QN(n8762) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n8915), .CLK(n9219), .Q(
        g25), .QN(n8679) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n8913), .CLK(n9217), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n8924), .CLK(n9228), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n8904), .CLK(n9208), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n8887), .CLK(n9191), .Q(
        n9267) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n8887), .CLK(n9191), .Q(
        g2066) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n8955), .CLK(n9266), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n8895), .CLK(n9199), .Q(
        g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n8903), .CLK(n9207), .Q(
        g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n8929), .CLK(n9233), .Q(
        g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n8929), .CLK(n9233), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n8936), .CLK(n9242), .Q(
        g8403), .QN(n8684) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n8936), .CLK(n9242), .Q(
        g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n8913), .CLK(n9217), 
        .Q(test_so76), .QN(n8839) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n8881), .CLK(n9185), 
        .Q(g2827), .QN(n8296) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n8906), .CLK(n9210), .Q(
        g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n8939), .CLK(n9246), 
        .Q(g4859) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n8940), .CLK(n9248), .Q(
        g424) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n8893), .CLK(n9197), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n8897), .CLK(n9201), .Q(
        g17423), .QN(n8734) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n8946), .CLK(n9254), 
        .Q(n9265), .QN(n6006) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n8881), .CLK(n9185), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n8907), .CLK(n9211), .Q(
        g1821), .QN(n8327) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n8880), .CLK(n9184), .Q(
        g2509), .QN(n8347) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n8969), .CLK(n9286), .Q(
        g5073), .QN(n8722) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n8972), .CLK(n9289), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n8942), .CLK(n9250), 
        .Q(g8353), .QN(n8682) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n8942), .CLK(n9250), .Q(
        g13085), .QN(n8707) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n8967), .CLK(n9284), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n8895), .CLK(n9199), .Q(
        g5124), .QN(n8787) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n8918), .CLK(n9222), 
        .Q(g17400), .QN(n8698) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n8899), .CLK(n9203), 
        .Q(g6303) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n8867), .CLK(n9171), .Q(
        g5069), .QN(n8344) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n8886), .CLK(n9190), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n8930), .CLK(n9234), .Q(
        g650) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n8913), .CLK(n9217), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n8903), .CLK(n9207), .Q(
        g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n8941), .CLK(n9249), .Q(
        test_so78), .QN(n8833) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n8971), .CLK(n9288), 
        .Q(g6732), .QN(n8506) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n8885), .CLK(n9189), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n8920), .CLK(n9224), .Q(
        g1061), .QN(n8756) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n8970), .CLK(n9287), .Q(
        g3462), .QN(n8723) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n8903), .CLK(n9207), .Q(
        g2181) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n8921), .CLK(n9225), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n8907), .CLK(n9211), .Q(
        g1756) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n8954), .CLK(n9264), .Q(
        g5849), .QN(n5736) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n8970), .CLK(n9287), .Q(
        g4112) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n8870), .CLK(n9174), .Q(
        n9262) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n8897), .CLK(n9201), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n8972), .CLK(n9289), .Q(
        test_so79), .QN(n8826) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n8900), .CLK(n9204), 
        .Q(g1046), .QN(n8572) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n8935), .CLK(n9241), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n8937), .CLK(n9243), .Q(
        g4401), .QN(n8342) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n8937), .CLK(n9243), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n8937), .CLK(n9243), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n8937), .CLK(n9243), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n8890), .CLK(n9194), .Q(
        g2950), .QN(n8524) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n8882), .CLK(n9186), .Q(
        g1345), .QN(n8799) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n8937), .CLK(n9243), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n8937), .CLK(n9243), .Q(
        g14421), .QN(n8710) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n8938), .CLK(n9244), 
        .Q(g4727) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n8921), .CLK(n9225), .Q(
        test_so80), .QN(n8840) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n8882), .CLK(n9186), 
        .Q(g1536), .QN(n8279) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n8891), .CLK(n9195), .Q(
        g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n8908), .CLK(n9212), .Q(
        g370), .QN(n8636) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n8884), .CLK(n9188), .Q(
        g5694), .QN(n8415) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n8888), .CLK(n9192), .Q(
        g1858) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n8888), .CLK(n9192), .Q(
        g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n8959), .CLK(n9271), .Q(
        g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n8908), .CLK(n9212), .Q(
        g1811), .QN(n8632) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n8908), .CLK(n9212), .Q(
        g6601) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n8881), .CLK(n9185), .Q(
        g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n8927), .CLK(n9231), .Q(
        g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n8938), .CLK(n9244), .Q(
        test_so81), .QN(n8822) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n8952), .CLK(n9261), 
        .Q(g6581) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n8929), .CLK(n9233), .Q(
        g6597) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n8936), .CLK(n9242), .Q(
        g5008) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n8917), .CLK(n9221), .Q(
        g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n8886), .CLK(n9190), .Q(
        g2890) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n8964), .CLK(n9279), .Q(
        g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n8875), .CLK(n9179), .Q(
        g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n8913), .CLK(n9217), .Q(
        g112), .QN(n8671) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n8870), .CLK(n9174), .Q(
        g2856) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n8964), .CLK(n9279), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n8964), .CLK(n9279), .Q(
        g17722), .QN(n8715) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n8930), .CLK(n9234), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n8894), .CLK(n9198), 
        .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n8956), .CLK(n9268), .Q(
        g6390), .QN(n8744) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n8882), .CLK(n9186), .Q(
        g1542), .QN(n8378) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n8882), .CLK(n9186), .Q(
        g4258), .QN(n8758) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n8942), .CLK(n9250), .Q(
        g4818) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n8911), .CLK(n9215), .Q(
        g5033), .QN(n8739) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n8938), .CLK(n9244), .Q(
        g4717) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n8971), .CLK(n9288), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n8921), .CLK(n9225), .Q(
        g3849), .QN(n5735) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n8921), .CLK(n9225), .Q(
        g17778), .QN(n8668) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n8959), .CLK(n9271), 
        .Q(g3199) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n8973), .CLK(n9290), .Q(
        test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n8940), .CLK(n9248), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n8946), .CLK(n9254), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n8897), .CLK(n9201), .Q(
        g5913) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n8928), .CLK(n9232), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n8879), .CLK(n9183), .Q(
        g6163), .QN(n8781) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n8914), .CLK(n9218), .Q(
        g4125), .QN(n8555) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n8914), .CLK(n9218), .Q(
        g4821), .QN(n5880) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n8933), .CLK(n9238), .Q(
        g4939) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n8933), .CLK(n9238), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n8960), .CLK(n9272), 
        .Q(g3207) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n8960), .CLK(n9272), .Q(
        g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n8928), .CLK(n9232), .Q(
        test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n8896), .CLK(n9200), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n8895), .CLK(n9199), .Q(
        g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n8873), .CLK(n9177), .Q(
        g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n8873), .CLK(n9177), .Q(
        g3694), .QN(n8414) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n8869), .CLK(n9173), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n8869), .CLK(n9173), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n8867), .CLK(n9171), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n8957), .CLK(n9269), .Q(
        g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n8968), .CLK(n9285), .Q(
        g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n8968), .CLK(n9285), 
        .Q(n9255), .QN(n6005) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n8877), .CLK(n9181), .Q(
        g4427), .QN(n8647) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n8877), .CLK(n9181), .Q(
        test_so85) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n8876), .CLK(n9180), 
        .Q(g2779), .QN(n8291) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n8942), .CLK(n9250), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n8967), .CLK(n9284), .Q(
        g7245) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n8967), .CLK(n9284), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n8967), .CLK(n9284), .Q(
        g1367), .QN(n8798) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n8967), .CLK(n9284), .Q(
        g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n8968), .CLK(n9285), .Q(
        g19), .QN(n8777) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n8968), .CLK(n9285), .Q(
        g4145), .QN(n8515) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n8903), .CLK(n9207), .Q(
        g2161) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n8909), .CLK(n9213), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n8966), .CLK(n9283), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n8931), .CLK(n9235), .Q(
        test_so86), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n8924), .CLK(n9228), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n8941), .CLK(n9249), .Q(
        g2051), .QN(n8778) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n8887), .CLK(n9191), .Q(
        g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n8901), .CLK(n9205), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n8926), .CLK(n9230), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n8926), .CLK(n9230), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n8888), .CLK(n9192), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n8917), .CLK(n9221), .Q(
        g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n8886), .CLK(n9190), .Q(
        g2999) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n8901), .CLK(n9205), .Q(
        g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n8921), .CLK(n9225), .Q(
        g17688), .QN(n8717) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n8930), .CLK(n9234), 
        .Q(test_so87), .QN(n8845) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n8909), .CLK(n9213), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n8955), .CLK(n9266), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n8967), .CLK(n9284), .Q(
        g546) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n8913), .CLK(n9217), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n8914), .CLK(n9218), .Q(
        g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n8971), .CLK(n9288), .Q(
        g8277), .QN(n8323) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n8907), .CLK(n9211), .Q(
        g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n8916), .CLK(n9220), .Q(
        g3550) );
  SDFFX1 DFF_1260_Q_reg ( .D(n568), .SI(g3550), .SE(n8873), .CLK(n9177), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n8873), .CLK(n9177), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n8958), .CLK(n9270), .Q(
        g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n8958), .CLK(n9270), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n8891), .CLK(n9195), 
        .Q(g3913) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n8889), .CLK(n9193), .Q(
        g10306), .QN(n8691) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n8875), .CLK(n9179), 
        .Q(g1687), .QN(n8331) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n8910), .CLK(n9214), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n8910), .CLK(n9214), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n8935), .CLK(n9241), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n8935), .CLK(n9241), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n8936), .CLK(n9242), .Q(
        g4417), .QN(n8790) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n8949), .CLK(n9258), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n8920), .CLK(n9224), .Q(
        g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n8910), .CLK(n9214), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n8947), .CLK(n9256), 
        .Q(test_so89), .QN(n8863) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n8919), .CLK(n9223), 
        .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n8885), .CLK(n9189), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n8960), .CLK(n9272), .Q(
        g3255) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n8919), .CLK(n9223), .Q(
        g1691), .QN(n8627) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n8890), .CLK(n9194), .Q(
        g2936), .QN(n8525) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n8884), .CLK(n9188), .Q(
        g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(n227), .SI(g5644), .SE(n8896), .CLK(n9200), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n8896), .CLK(n9200), .Q(
        g5352), .QN(n8774) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n8896), .CLK(n9200), .Q(
        g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n8876), .CLK(n9180), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n8890), .CLK(n9194), .Q(
        g2922), .QN(n8523) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n8907), .CLK(n9211), .Q(
        test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n8914), .CLK(n9218), 
        .Q(g5893) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n8961), .CLK(n9275), .Q(
        g16603), .QN(n8711) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n8967), .CLK(n9284), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n8887), .CLK(n9191), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n8972), .CLK(n9289), .Q(
        g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n8868), .CLK(n9172), .Q(
        g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n8923), .CLK(n9227), .Q(
        g3401) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n8923), .CLK(n9227), .Q(
        g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n8923), .CLK(n9227), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n8923), .CLK(n9227), 
        .Q(g29214) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n8922), .CLK(n9226), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n8965), .CLK(n9282), .Q(
        test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n8953), .CLK(n9263), 
        .Q(g5170), .QN(n8642) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n8953), .CLK(n9263), .Q(
        g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n8883), .CLK(n9187), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n8899), .CLK(n9203), .Q(
        g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n8933), .CLK(n9238), .Q(
        g8416), .QN(n8747) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n8887), .CLK(n9191), .Q(
        g2079), .QN(n8626) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n8896), .CLK(n9200), .Q(
        g4698) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n8874), .CLK(n9178), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n8970), .CLK(n9287), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n8971), .CLK(n9288), .Q(
        n9247) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n8892), .CLK(n9196), .Q(
        g411) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n8955), .CLK(n9266), .Q(
        test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n8903), .CLK(n9207), 
        .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n8903), .CLK(n9207), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n8948), .CLK(n9257), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n8948), .CLK(n9257), .Q(
        n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n8948), .CLK(n9257), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n8948), .CLK(n9257), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n8961), .CLK(n9275), .Q(
        g5200) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n8939), .CLK(n9246), .Q(
        g4843), .QN(n8689) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n8911), .CLK(n9215), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n8941), .CLK(n9249), .Q(
        g2250), .QN(n8633) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n8937), .CLK(n9243), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n8969), .CLK(n9286), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n8950), .CLK(n9259), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n8883), .CLK(n9187), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n8883), .CLK(n9187), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n8890), .CLK(n9194), 
        .Q(g2912), .QN(n8522) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n8947), .CLK(n9256), .Q(
        g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n8966), .CLK(n9283), .Q(
        g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n8905), .CLK(n9209), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n8872), .CLK(n9176), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n8969), .CLK(n9286), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n8922), .CLK(n9226), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n8882), .CLK(n9186), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n8946), .CLK(n9254), .Q(
        test_so94), .QN(n8831) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n8872), .CLK(n9176), 
        .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n8895), .CLK(n9199), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n8965), .CLK(n9282), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n8908), .CLK(n9212), .Q(
        g6657) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n8969), .CLK(n9286), .Q(
        g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n8903), .CLK(n9207), .Q(
        g3893) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n8960), .CLK(n9272), .Q(
        g3211) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n8958), .CLK(n9270), .Q(
        g13049), .QN(n8701) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n8961), .CLK(n9275), 
        .Q(g16624), .QN(n8709) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n8868), .CLK(n9172), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n8917), .CLK(n9221), .Q(
        g3614) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n8917), .CLK(n9221), .Q(
        test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n8965), .CLK(n9282), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n8965), .CLK(n9282), .Q(
        g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n8873), .CLK(n9177), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n8948), .CLK(n9257), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n8898), .CLK(n9202), .Q(
        g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n8895), .CLK(n9199), .Q(
        g5272) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n8940), .CLK(n9248), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n8892), .CLK(n9196), .Q(
        g728), .QN(n8382) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n8966), .CLK(n9283), .Q(
        g6295) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n8870), .CLK(n9174), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n8964), .CLK(n9279), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n8895), .CLK(n9199), .Q(
        test_so96), .QN(n8848) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n8922), .CLK(n9226), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n8922), .CLK(n9226), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n8871), .CLK(n9175), .Q(
        g4659), .QN(n8769) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n8871), .CLK(n9175), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n8961), .CLK(n9275), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n8917), .CLK(n9221), .Q(
        g2084), .QN(n8346) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n8955), .CLK(n9266), .Q(
        g3187) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n8955), .CLK(n9266), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n8966), .CLK(n9283), .Q(
        g2583) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n8906), .CLK(n9210), .Q(
        n9240) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n8907), .CLK(n9211), .Q(
        g1094), .QN(n5697) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n8921), .CLK(n9225), .Q(
        test_so97), .QN(n8858) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n8931), .CLK(n9235), 
        .Q(g4284), .QN(n8361) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n8959), .CLK(n9271), .Q(
        g3191) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n8882), .CLK(n9186), .Q(
        g4239), .QN(n8354) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n8934), .CLK(n9239), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n8877), .CLK(n9181), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n8877), .CLK(n9181), .Q(
        g534) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n8909), .CLK(n9213), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n8918), .CLK(n9222), .Q(
        g2004) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n8953), .CLK(n9263), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n8953), .CLK(n9263), .Q(
        g5456), .QN(n8316) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n8889), .CLK(n9193), .Q(
        n6007), .QN(n8648) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n8966), .CLK(n9283), .Q(
        test_so98), .QN(n8859) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n8945), .CLK(n9253), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n8896), .CLK(n9200), .Q(
        g5348), .QN(n8507) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n8959), .CLK(n9271), .Q(
        g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n8890), .CLK(n9194), .Q(
        g2970), .QN(n8521) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n8884), .CLK(n9188), .Q(
        g5698), .QN(n8754) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n8930), .CLK(n9234), .Q(
        g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n8885), .CLK(n9189), .Q(
        g1521) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n8923), .CLK(n9227), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n8922), .CLK(n9226), .Q(
        g3115), .QN(n8738) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n8959), .CLK(n9271), .Q(
        g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n8938), .CLK(n9244), .Q(
        g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n8938), .CLK(n9244), 
        .Q(test_so99), .QN(n8843) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n8917), .CLK(n9221), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n8923), .CLK(n9227), .Q(
        g8342), .QN(n8301) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n8872), .CLK(n9176), .Q(
        g4515), .QN(n8552) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n8943), .CLK(n9251), .Q(
        g8787), .QN(n8650) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n8872), .CLK(n9176), .Q(
        g4300) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n8919), .CLK(n9223), .Q(
        n9236) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n8920), .CLK(n9224), .Q(
        g1379), .QN(n8797) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n8950), .CLK(n9259), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n8927), .CLK(n9231), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n8868), .CLK(n9172), .Q(
        g5619) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n8869), .CLK(n9173), .Q(
        g71), .QN(n8618) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n8898), .CLK(n9202), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1430), .SI(g4704), .SE(n8963), .CLK(n9278), .Q(
        g22), .QN(n8789) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n8935), .CLK(n9241), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n8940), .CLK(n9248), .Q(
        g2729), .QN(n8676) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n8866), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n8865), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n8866), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n8865), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n8866), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n8865), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n8866), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n8865), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n8866), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n8865), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n8866), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n8865), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n8866), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n8865), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n8866), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n8865), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n8866), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n8865), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n8866), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n8865), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n8866), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n8865), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n282), .IN2(n549), .IN3(n353), .IN4(n58), .QN(n87)
         );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n282), .IN2(n549), .IN3(n353), .IN4(n59), .QN(n37)
         );
  NAND3X0 Trojan_U17 ( .IN1(n141), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n3279), .IN3(n8803), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U8791 ( .INP(n87), .ZN(n8864) );
  INVX0 U8792 ( .INP(n8864), .ZN(n8865) );
  INVX0 U8793 ( .INP(n8864), .ZN(n8866) );
  NBUFFX2 U8794 ( .INP(n8995), .Z(n8868) );
  NBUFFX2 U8795 ( .INP(n8995), .Z(n8867) );
  NBUFFX2 U8796 ( .INP(n8991), .Z(n8888) );
  NBUFFX2 U8797 ( .INP(n8981), .Z(n8938) );
  NBUFFX2 U8798 ( .INP(n8990), .Z(n8893) );
  NBUFFX2 U8799 ( .INP(n8994), .Z(n8872) );
  NBUFFX2 U8800 ( .INP(n8986), .Z(n8910) );
  NBUFFX2 U8801 ( .INP(n8978), .Z(n8953) );
  NBUFFX2 U8802 ( .INP(n8975), .Z(n8967) );
  NBUFFX2 U8803 ( .INP(n8988), .Z(n8903) );
  NBUFFX2 U8804 ( .INP(n8982), .Z(n8931) );
  NBUFFX2 U8805 ( .INP(n8991), .Z(n8887) );
  NBUFFX2 U8806 ( .INP(n8986), .Z(n8913) );
  NBUFFX2 U8807 ( .INP(n8980), .Z(n8940) );
  NBUFFX2 U8808 ( .INP(n8985), .Z(n8918) );
  NBUFFX2 U8809 ( .INP(n8981), .Z(n8936) );
  NBUFFX2 U8810 ( .INP(n8983), .Z(n8927) );
  NBUFFX2 U8811 ( .INP(n8986), .Z(n8912) );
  NBUFFX2 U8812 ( .INP(n8992), .Z(n8881) );
  NBUFFX2 U8813 ( .INP(n8994), .Z(n8869) );
  NBUFFX2 U8814 ( .INP(n8978), .Z(n8952) );
  NBUFFX2 U8815 ( .INP(n8987), .Z(n8908) );
  NBUFFX2 U8816 ( .INP(n8988), .Z(n8902) );
  NBUFFX2 U8817 ( .INP(n8982), .Z(n8933) );
  NBUFFX2 U8818 ( .INP(n8984), .Z(n8921) );
  NBUFFX2 U8819 ( .INP(n8987), .Z(n8905) );
  NBUFFX2 U8820 ( .INP(n8989), .Z(n8895) );
  NBUFFX2 U8821 ( .INP(n8980), .Z(n8942) );
  NBUFFX2 U8822 ( .INP(n8980), .Z(n8941) );
  NBUFFX2 U8823 ( .INP(n8979), .Z(n8947) );
  NBUFFX2 U8824 ( .INP(n8981), .Z(n8937) );
  NBUFFX2 U8825 ( .INP(n8975), .Z(n8964) );
  NBUFFX2 U8826 ( .INP(n8993), .Z(n8877) );
  NBUFFX2 U8827 ( .INP(n8976), .Z(n8961) );
  NBUFFX2 U8828 ( .INP(n8987), .Z(n8906) );
  NBUFFX2 U8829 ( .INP(n8989), .Z(n8896) );
  NBUFFX2 U8830 ( .INP(n8986), .Z(n8911) );
  NBUFFX2 U8831 ( .INP(n8976), .Z(n8959) );
  NBUFFX2 U8832 ( .INP(n8990), .Z(n8889) );
  NBUFFX2 U8833 ( .INP(n8977), .Z(n8955) );
  NBUFFX2 U8834 ( .INP(n8983), .Z(n8925) );
  NBUFFX2 U8835 ( .INP(n8979), .Z(n8946) );
  NBUFFX2 U8836 ( .INP(n8980), .Z(n8939) );
  NBUFFX2 U8837 ( .INP(n8981), .Z(n8934) );
  NBUFFX2 U8838 ( .INP(n8986), .Z(n8909) );
  NBUFFX2 U8839 ( .INP(n8983), .Z(n8926) );
  NBUFFX2 U8840 ( .INP(n8985), .Z(n8914) );
  NBUFFX2 U8841 ( .INP(n8990), .Z(n8891) );
  NBUFFX2 U8842 ( .INP(n8976), .Z(n8962) );
  NBUFFX2 U8843 ( .INP(n8993), .Z(n8878) );
  NBUFFX2 U8844 ( .INP(n8991), .Z(n8884) );
  NBUFFX2 U8845 ( .INP(n8988), .Z(n8900) );
  NBUFFX2 U8846 ( .INP(n8994), .Z(n8871) );
  NBUFFX2 U8847 ( .INP(n8975), .Z(n8965) );
  NBUFFX2 U8848 ( .INP(n8985), .Z(n8917) );
  NBUFFX2 U8849 ( .INP(n8977), .Z(n8957) );
  NBUFFX2 U8850 ( .INP(n8992), .Z(n8882) );
  NBUFFX2 U8851 ( .INP(n8985), .Z(n8915) );
  NBUFFX2 U8852 ( .INP(n8984), .Z(n8922) );
  NBUFFX2 U8853 ( .INP(n8991), .Z(n8886) );
  NBUFFX2 U8854 ( .INP(n8982), .Z(n8930) );
  NBUFFX2 U8855 ( .INP(n8982), .Z(n8932) );
  NBUFFX2 U8856 ( .INP(n8977), .Z(n8958) );
  NBUFFX2 U8857 ( .INP(n8978), .Z(n8949) );
  NBUFFX2 U8858 ( .INP(n8982), .Z(n8929) );
  NBUFFX2 U8859 ( .INP(n8991), .Z(n8885) );
  NBUFFX2 U8860 ( .INP(n8988), .Z(n8899) );
  NBUFFX2 U8861 ( .INP(n8975), .Z(n8968) );
  NBUFFX2 U8862 ( .INP(n8992), .Z(n8879) );
  NBUFFX2 U8863 ( .INP(n8993), .Z(n8874) );
  NBUFFX2 U8864 ( .INP(n8979), .Z(n8945) );
  NBUFFX2 U8865 ( .INP(n8981), .Z(n8935) );
  NBUFFX2 U8866 ( .INP(n8994), .Z(n8870) );
  NBUFFX2 U8867 ( .INP(n8979), .Z(n8944) );
  NBUFFX2 U8868 ( .INP(n8994), .Z(n8873) );
  NBUFFX2 U8869 ( .INP(n8989), .Z(n8898) );
  NBUFFX2 U8870 ( .INP(n8987), .Z(n8904) );
  NBUFFX2 U8871 ( .INP(n8977), .Z(n8956) );
  NBUFFX2 U8872 ( .INP(n8978), .Z(n8950) );
  NBUFFX2 U8873 ( .INP(n8984), .Z(n8919) );
  NBUFFX2 U8874 ( .INP(n8993), .Z(n8875) );
  NBUFFX2 U8875 ( .INP(n8975), .Z(n8966) );
  NBUFFX2 U8876 ( .INP(n8992), .Z(n8883) );
  NBUFFX2 U8877 ( .INP(n8983), .Z(n8924) );
  NBUFFX2 U8878 ( .INP(n8980), .Z(n8943) );
  NBUFFX2 U8879 ( .INP(n8984), .Z(n8923) );
  NBUFFX2 U8880 ( .INP(n8984), .Z(n8920) );
  NBUFFX2 U8881 ( .INP(n8979), .Z(n8948) );
  NBUFFX2 U8882 ( .INP(n8976), .Z(n8963) );
  NBUFFX2 U8883 ( .INP(n8989), .Z(n8897) );
  NBUFFX2 U8884 ( .INP(n8987), .Z(n8907) );
  NBUFFX2 U8885 ( .INP(n8990), .Z(n8890) );
  NBUFFX2 U8886 ( .INP(n8977), .Z(n8954) );
  NBUFFX2 U8887 ( .INP(n8989), .Z(n8894) );
  NBUFFX2 U8888 ( .INP(n8985), .Z(n8916) );
  NBUFFX2 U8889 ( .INP(n8990), .Z(n8892) );
  NBUFFX2 U8890 ( .INP(n8976), .Z(n8960) );
  NBUFFX2 U8891 ( .INP(n8978), .Z(n8951) );
  NBUFFX2 U8892 ( .INP(n8992), .Z(n8880) );
  NBUFFX2 U8893 ( .INP(n8988), .Z(n8901) );
  NBUFFX2 U8894 ( .INP(n8983), .Z(n8928) );
  NBUFFX2 U8895 ( .INP(n8993), .Z(n8876) );
  NBUFFX2 U8896 ( .INP(n9319), .Z(n9172) );
  NBUFFX2 U8897 ( .INP(n9319), .Z(n9171) );
  NBUFFX2 U8898 ( .INP(n9315), .Z(n9192) );
  NBUFFX2 U8899 ( .INP(n9300), .Z(n9244) );
  NBUFFX2 U8900 ( .INP(n9313), .Z(n9197) );
  NBUFFX2 U8901 ( .INP(n9318), .Z(n9176) );
  NBUFFX2 U8902 ( .INP(n9308), .Z(n9214) );
  NBUFFX2 U8903 ( .INP(n9297), .Z(n9263) );
  NBUFFX2 U8904 ( .INP(n9292), .Z(n9284) );
  NBUFFX2 U8905 ( .INP(n9310), .Z(n9207) );
  NBUFFX2 U8906 ( .INP(n9301), .Z(n9235) );
  NBUFFX2 U8907 ( .INP(n9315), .Z(n9191) );
  NBUFFX2 U8908 ( .INP(n9308), .Z(n9217) );
  NBUFFX2 U8909 ( .INP(n9299), .Z(n9248) );
  NBUFFX2 U8910 ( .INP(n9307), .Z(n9222) );
  NBUFFX2 U8911 ( .INP(n9300), .Z(n9242) );
  NBUFFX2 U8912 ( .INP(n9304), .Z(n9231) );
  NBUFFX2 U8913 ( .INP(n9308), .Z(n9216) );
  NBUFFX2 U8914 ( .INP(n9316), .Z(n9185) );
  NBUFFX2 U8915 ( .INP(n9318), .Z(n9173) );
  NBUFFX2 U8916 ( .INP(n9297), .Z(n9261) );
  NBUFFX2 U8917 ( .INP(n9309), .Z(n9212) );
  NBUFFX2 U8918 ( .INP(n9310), .Z(n9206) );
  NBUFFX2 U8919 ( .INP(n9301), .Z(n9238) );
  NBUFFX2 U8920 ( .INP(n9305), .Z(n9225) );
  NBUFFX2 U8921 ( .INP(n9309), .Z(n9209) );
  NBUFFX2 U8922 ( .INP(n9311), .Z(n9199) );
  NBUFFX2 U8923 ( .INP(n9299), .Z(n9250) );
  NBUFFX2 U8924 ( .INP(n9299), .Z(n9249) );
  NBUFFX2 U8925 ( .INP(n9298), .Z(n9256) );
  NBUFFX2 U8926 ( .INP(n9300), .Z(n9243) );
  NBUFFX2 U8927 ( .INP(n9292), .Z(n9279) );
  NBUFFX2 U8928 ( .INP(n9317), .Z(n9181) );
  NBUFFX2 U8929 ( .INP(n9293), .Z(n9275) );
  NBUFFX2 U8930 ( .INP(n9309), .Z(n9210) );
  NBUFFX2 U8931 ( .INP(n9311), .Z(n9200) );
  NBUFFX2 U8932 ( .INP(n9308), .Z(n9215) );
  NBUFFX2 U8933 ( .INP(n9293), .Z(n9271) );
  NBUFFX2 U8934 ( .INP(n9313), .Z(n9193) );
  NBUFFX2 U8935 ( .INP(n9296), .Z(n9266) );
  NBUFFX2 U8936 ( .INP(n9304), .Z(n9229) );
  NBUFFX2 U8937 ( .INP(n9298), .Z(n9254) );
  NBUFFX2 U8938 ( .INP(n9299), .Z(n9246) );
  NBUFFX2 U8939 ( .INP(n9300), .Z(n9239) );
  NBUFFX2 U8940 ( .INP(n9308), .Z(n9213) );
  NBUFFX2 U8941 ( .INP(n9304), .Z(n9230) );
  NBUFFX2 U8942 ( .INP(n9307), .Z(n9218) );
  NBUFFX2 U8943 ( .INP(n9313), .Z(n9195) );
  NBUFFX2 U8944 ( .INP(n9293), .Z(n9277) );
  NBUFFX2 U8945 ( .INP(n9317), .Z(n9182) );
  NBUFFX2 U8946 ( .INP(n9315), .Z(n9188) );
  NBUFFX2 U8947 ( .INP(n9310), .Z(n9204) );
  NBUFFX2 U8948 ( .INP(n9318), .Z(n9175) );
  NBUFFX2 U8949 ( .INP(n9292), .Z(n9282) );
  NBUFFX2 U8950 ( .INP(n9307), .Z(n9221) );
  NBUFFX2 U8951 ( .INP(n9296), .Z(n9269) );
  NBUFFX2 U8952 ( .INP(n9316), .Z(n9186) );
  NBUFFX2 U8953 ( .INP(n9307), .Z(n9219) );
  NBUFFX2 U8954 ( .INP(n9305), .Z(n9226) );
  NBUFFX2 U8955 ( .INP(n9315), .Z(n9190) );
  NBUFFX2 U8956 ( .INP(n9301), .Z(n9234) );
  NBUFFX2 U8957 ( .INP(n9301), .Z(n9237) );
  NBUFFX2 U8958 ( .INP(n9296), .Z(n9270) );
  NBUFFX2 U8959 ( .INP(n9297), .Z(n9258) );
  NBUFFX2 U8960 ( .INP(n9301), .Z(n9233) );
  NBUFFX2 U8961 ( .INP(n9315), .Z(n9189) );
  NBUFFX2 U8962 ( .INP(n9310), .Z(n9203) );
  NBUFFX2 U8963 ( .INP(n9292), .Z(n9285) );
  NBUFFX2 U8964 ( .INP(n9316), .Z(n9183) );
  NBUFFX2 U8965 ( .INP(n9317), .Z(n9178) );
  NBUFFX2 U8966 ( .INP(n9298), .Z(n9253) );
  NBUFFX2 U8967 ( .INP(n9300), .Z(n9241) );
  NBUFFX2 U8968 ( .INP(n9318), .Z(n9174) );
  NBUFFX2 U8969 ( .INP(n9298), .Z(n9252) );
  NBUFFX2 U8970 ( .INP(n9318), .Z(n9177) );
  NBUFFX2 U8971 ( .INP(n9311), .Z(n9202) );
  NBUFFX2 U8972 ( .INP(n9309), .Z(n9208) );
  NBUFFX2 U8973 ( .INP(n9296), .Z(n9268) );
  NBUFFX2 U8976 ( .INP(n9297), .Z(n9259) );
  NBUFFX2 U8977 ( .INP(n9305), .Z(n9223) );
  NBUFFX2 U8978 ( .INP(n9317), .Z(n9179) );
  NBUFFX2 U8979 ( .INP(n9292), .Z(n9283) );
  NBUFFX2 U8980 ( .INP(n9316), .Z(n9187) );
  NBUFFX2 U8981 ( .INP(n9304), .Z(n9228) );
  NBUFFX2 U8982 ( .INP(n9299), .Z(n9251) );
  NBUFFX2 U8983 ( .INP(n9305), .Z(n9227) );
  NBUFFX2 U8984 ( .INP(n9305), .Z(n9224) );
  NBUFFX2 U8985 ( .INP(n9298), .Z(n9257) );
  NBUFFX2 U8986 ( .INP(n9293), .Z(n9278) );
  NBUFFX2 U8987 ( .INP(n9311), .Z(n9201) );
  NBUFFX2 U8988 ( .INP(n9309), .Z(n9211) );
  NBUFFX2 U8989 ( .INP(n9313), .Z(n9194) );
  NBUFFX2 U8990 ( .INP(n9296), .Z(n9264) );
  NBUFFX2 U8991 ( .INP(n9311), .Z(n9198) );
  NBUFFX2 U8992 ( .INP(n9307), .Z(n9220) );
  NBUFFX2 U8993 ( .INP(n9313), .Z(n9196) );
  NBUFFX2 U8994 ( .INP(n9293), .Z(n9272) );
  NBUFFX2 U8995 ( .INP(n9297), .Z(n9260) );
  NBUFFX2 U8996 ( .INP(n9316), .Z(n9184) );
  NBUFFX2 U8997 ( .INP(n9310), .Z(n9205) );
  NBUFFX2 U8998 ( .INP(n9304), .Z(n9232) );
  NBUFFX2 U8999 ( .INP(n9317), .Z(n9180) );
  NBUFFX2 U9000 ( .INP(n8974), .Z(n8969) );
  NBUFFX2 U9001 ( .INP(n8974), .Z(n8971) );
  NBUFFX2 U9002 ( .INP(n8974), .Z(n8972) );
  NBUFFX2 U9003 ( .INP(n8974), .Z(n8970) );
  NBUFFX2 U9004 ( .INP(n9291), .Z(n9286) );
  NBUFFX2 U9005 ( .INP(n9291), .Z(n9288) );
  NBUFFX2 U9006 ( .INP(n9291), .Z(n9289) );
  NBUFFX2 U9007 ( .INP(n9291), .Z(n9287) );
  NBUFFX2 U9008 ( .INP(n8974), .Z(n8973) );
  NBUFFX2 U9009 ( .INP(n9291), .Z(n9290) );
  NBUFFX2 U9010 ( .INP(n9003), .Z(n8974) );
  NBUFFX2 U9011 ( .INP(n9002), .Z(n8975) );
  NBUFFX2 U9012 ( .INP(n9002), .Z(n8976) );
  NBUFFX2 U9013 ( .INP(n9002), .Z(n8977) );
  NBUFFX2 U9014 ( .INP(n9001), .Z(n8978) );
  NBUFFX2 U9015 ( .INP(n9001), .Z(n8979) );
  NBUFFX2 U9016 ( .INP(n9001), .Z(n8980) );
  NBUFFX2 U9017 ( .INP(n9000), .Z(n8981) );
  NBUFFX2 U9018 ( .INP(n9000), .Z(n8982) );
  NBUFFX2 U9019 ( .INP(n9000), .Z(n8983) );
  NBUFFX2 U9020 ( .INP(n8999), .Z(n8984) );
  NBUFFX2 U9021 ( .INP(n8999), .Z(n8985) );
  NBUFFX2 U9022 ( .INP(n8999), .Z(n8986) );
  NBUFFX2 U9023 ( .INP(n8998), .Z(n8987) );
  NBUFFX2 U9024 ( .INP(n8998), .Z(n8988) );
  NBUFFX2 U9025 ( .INP(n8998), .Z(n8989) );
  NBUFFX2 U9026 ( .INP(n8997), .Z(n8990) );
  NBUFFX2 U9027 ( .INP(n8997), .Z(n8991) );
  NBUFFX2 U9028 ( .INP(n8997), .Z(n8992) );
  NBUFFX2 U9029 ( .INP(n8996), .Z(n8993) );
  NBUFFX2 U9030 ( .INP(n8996), .Z(n8994) );
  NBUFFX2 U9031 ( .INP(n8996), .Z(n8995) );
  NBUFFX2 U9032 ( .INP(n9006), .Z(n8996) );
  NBUFFX2 U9033 ( .INP(n9006), .Z(n8997) );
  NBUFFX2 U9034 ( .INP(n9005), .Z(n8998) );
  NBUFFX2 U9035 ( .INP(n9005), .Z(n8999) );
  NBUFFX2 U9036 ( .INP(n9005), .Z(n9000) );
  NBUFFX2 U9037 ( .INP(n9004), .Z(n9001) );
  NBUFFX2 U9038 ( .INP(n9004), .Z(n9002) );
  NBUFFX2 U9039 ( .INP(n9004), .Z(n9003) );
  NBUFFX2 U9040 ( .INP(test_se), .Z(n9004) );
  NBUFFX2 U9041 ( .INP(test_se), .Z(n9005) );
  NBUFFX2 U9042 ( .INP(test_se), .Z(n9006) );
  NBUFFX2 U9043 ( .INP(n9108), .Z(n9007) );
  NBUFFX2 U9044 ( .INP(n9107), .Z(n9008) );
  NBUFFX2 U9045 ( .INP(n9107), .Z(n9009) );
  NBUFFX2 U9046 ( .INP(n9107), .Z(n9010) );
  NBUFFX2 U9047 ( .INP(n9106), .Z(n9011) );
  NBUFFX2 U9048 ( .INP(n9106), .Z(n9012) );
  NBUFFX2 U9049 ( .INP(n9106), .Z(n9013) );
  NBUFFX2 U9050 ( .INP(n9105), .Z(n9014) );
  NBUFFX2 U9051 ( .INP(n9105), .Z(n9015) );
  NBUFFX2 U9052 ( .INP(n9105), .Z(n9016) );
  NBUFFX2 U9053 ( .INP(n9104), .Z(n9017) );
  NBUFFX2 U9054 ( .INP(n9104), .Z(n9018) );
  NBUFFX2 U9055 ( .INP(n9104), .Z(n9019) );
  NBUFFX2 U9056 ( .INP(n9103), .Z(n9020) );
  NBUFFX2 U9057 ( .INP(n9103), .Z(n9021) );
  NBUFFX2 U9058 ( .INP(n9103), .Z(n9022) );
  NBUFFX2 U9059 ( .INP(n9102), .Z(n9023) );
  NBUFFX2 U9060 ( .INP(n9102), .Z(n9024) );
  NBUFFX2 U9061 ( .INP(n9102), .Z(n9025) );
  NBUFFX2 U9062 ( .INP(n9101), .Z(n9026) );
  NBUFFX2 U9063 ( .INP(n9101), .Z(n9027) );
  NBUFFX2 U9064 ( .INP(n9101), .Z(n9028) );
  NBUFFX2 U9066 ( .INP(n9100), .Z(n9029) );
  NBUFFX2 U9067 ( .INP(n9100), .Z(n9030) );
  NBUFFX2 U9068 ( .INP(n9100), .Z(n9031) );
  NBUFFX2 U9069 ( .INP(n9099), .Z(n9032) );
  NBUFFX2 U9071 ( .INP(n9099), .Z(n9033) );
  NBUFFX2 U9072 ( .INP(n9099), .Z(n9034) );
  NBUFFX2 U9073 ( .INP(n9098), .Z(n9035) );
  NBUFFX2 U9074 ( .INP(n9098), .Z(n9036) );
  NBUFFX2 U9077 ( .INP(n9098), .Z(n9037) );
  NBUFFX2 U9078 ( .INP(n9097), .Z(n9038) );
  NBUFFX2 U9079 ( .INP(n9097), .Z(n9039) );
  NBUFFX2 U9081 ( .INP(n9097), .Z(n9040) );
  NBUFFX2 U9082 ( .INP(n9096), .Z(n9041) );
  NBUFFX2 U9083 ( .INP(n9096), .Z(n9042) );
  NBUFFX2 U9087 ( .INP(n9096), .Z(n9043) );
  NBUFFX2 U9088 ( .INP(n9095), .Z(n9044) );
  NBUFFX2 U9089 ( .INP(n9095), .Z(n9045) );
  NBUFFX2 U9091 ( .INP(n9095), .Z(n9046) );
  NBUFFX2 U9092 ( .INP(n9094), .Z(n9047) );
  NBUFFX2 U9093 ( .INP(n9094), .Z(n9048) );
  NBUFFX2 U9094 ( .INP(n9094), .Z(n9049) );
  NBUFFX2 U9095 ( .INP(n9093), .Z(n9050) );
  NBUFFX2 U9096 ( .INP(n9093), .Z(n9051) );
  NBUFFX2 U9097 ( .INP(n9093), .Z(n9052) );
  NBUFFX2 U9100 ( .INP(n9092), .Z(n9053) );
  NBUFFX2 U9102 ( .INP(n9092), .Z(n9054) );
  NBUFFX2 U9103 ( .INP(n9092), .Z(n9055) );
  NBUFFX2 U9104 ( .INP(n9091), .Z(n9056) );
  NBUFFX2 U9105 ( .INP(n9091), .Z(n9057) );
  NBUFFX2 U9106 ( .INP(n9091), .Z(n9058) );
  NBUFFX2 U9108 ( .INP(n9090), .Z(n9059) );
  NBUFFX2 U9109 ( .INP(n9090), .Z(n9060) );
  NBUFFX2 U9110 ( .INP(n9090), .Z(n9061) );
  NBUFFX2 U9112 ( .INP(n9089), .Z(n9062) );
  NBUFFX2 U9113 ( .INP(n9089), .Z(n9063) );
  NBUFFX2 U9114 ( .INP(n9089), .Z(n9064) );
  NBUFFX2 U9115 ( .INP(n9088), .Z(n9065) );
  NBUFFX2 U9117 ( .INP(n9088), .Z(n9066) );
  NBUFFX2 U9118 ( .INP(n9088), .Z(n9067) );
  NBUFFX2 U9119 ( .INP(n9087), .Z(n9068) );
  NBUFFX2 U9121 ( .INP(n9087), .Z(n9069) );
  NBUFFX2 U9122 ( .INP(n9087), .Z(n9070) );
  NBUFFX2 U9123 ( .INP(n9086), .Z(n9071) );
  NBUFFX2 U9125 ( .INP(n9086), .Z(n9072) );
  NBUFFX2 U9126 ( .INP(n9086), .Z(n9073) );
  NBUFFX2 U9127 ( .INP(n9085), .Z(n9074) );
  NBUFFX2 U9129 ( .INP(n9085), .Z(n9075) );
  NBUFFX2 U9130 ( .INP(n9085), .Z(n9076) );
  NBUFFX2 U9131 ( .INP(n9084), .Z(n9077) );
  NBUFFX2 U9133 ( .INP(n9084), .Z(n9078) );
  NBUFFX2 U9134 ( .INP(n9084), .Z(n9079) );
  NBUFFX2 U9135 ( .INP(n9083), .Z(n9080) );
  NBUFFX2 U9137 ( .INP(n9083), .Z(n9081) );
  NBUFFX2 U9138 ( .INP(n9083), .Z(n9082) );
  NBUFFX2 U9139 ( .INP(n9117), .Z(n9083) );
  NBUFFX2 U9140 ( .INP(n9117), .Z(n9084) );
  NBUFFX2 U9141 ( .INP(n9116), .Z(n9085) );
  NBUFFX2 U9142 ( .INP(n9116), .Z(n9086) );
  NBUFFX2 U9143 ( .INP(n9116), .Z(n9087) );
  NBUFFX2 U9144 ( .INP(n9115), .Z(n9088) );
  NBUFFX2 U9145 ( .INP(n9115), .Z(n9089) );
  NBUFFX2 U9146 ( .INP(n9115), .Z(n9090) );
  NBUFFX2 U9147 ( .INP(n9114), .Z(n9091) );
  NBUFFX2 U9148 ( .INP(n9114), .Z(n9092) );
  NBUFFX2 U9149 ( .INP(n9114), .Z(n9093) );
  NBUFFX2 U9150 ( .INP(n9113), .Z(n9094) );
  NBUFFX2 U9151 ( .INP(n9113), .Z(n9095) );
  NBUFFX2 U9152 ( .INP(n9113), .Z(n9096) );
  NBUFFX2 U9153 ( .INP(n9112), .Z(n9097) );
  NBUFFX2 U9154 ( .INP(n9112), .Z(n9098) );
  NBUFFX2 U9155 ( .INP(n9112), .Z(n9099) );
  NBUFFX2 U9156 ( .INP(n9111), .Z(n9100) );
  NBUFFX2 U9157 ( .INP(n9111), .Z(n9101) );
  NBUFFX2 U9158 ( .INP(n9111), .Z(n9102) );
  NBUFFX2 U9159 ( .INP(n9110), .Z(n9103) );
  NBUFFX2 U9160 ( .INP(n9110), .Z(n9104) );
  NBUFFX2 U9161 ( .INP(n9110), .Z(n9105) );
  NBUFFX2 U9162 ( .INP(n9109), .Z(n9106) );
  NBUFFX2 U9163 ( .INP(n9109), .Z(n9107) );
  NBUFFX2 U9164 ( .INP(n9109), .Z(n9108) );
  NBUFFX2 U9165 ( .INP(n9120), .Z(n9109) );
  NBUFFX2 U9166 ( .INP(n9120), .Z(n9110) );
  NBUFFX2 U9167 ( .INP(n9120), .Z(n9111) );
  NBUFFX2 U9168 ( .INP(n9119), .Z(n9112) );
  NBUFFX2 U9169 ( .INP(n9119), .Z(n9113) );
  NBUFFX2 U9170 ( .INP(n9119), .Z(n9114) );
  NBUFFX2 U9171 ( .INP(n9118), .Z(n9115) );
  NBUFFX2 U9172 ( .INP(n9118), .Z(n9116) );
  NBUFFX2 U9173 ( .INP(n9118), .Z(n9117) );
  NBUFFX2 U9174 ( .INP(g35), .Z(n9118) );
  NBUFFX2 U9175 ( .INP(g35), .Z(n9119) );
  NBUFFX2 U9176 ( .INP(g35), .Z(n9120) );
  INVX0 U9177 ( .INP(n9008), .ZN(n9121) );
  INVX0 U9178 ( .INP(n9008), .ZN(n9122) );
  INVX0 U9179 ( .INP(n9008), .ZN(n9123) );
  INVX0 U9180 ( .INP(n9009), .ZN(n9124) );
  INVX0 U9181 ( .INP(n9009), .ZN(n9125) );
  INVX0 U9182 ( .INP(n9009), .ZN(n9126) );
  INVX0 U9183 ( .INP(n9009), .ZN(n9127) );
  INVX0 U9184 ( .INP(n9010), .ZN(n9128) );
  INVX0 U9185 ( .INP(n9009), .ZN(n9129) );
  INVX0 U9186 ( .INP(n9009), .ZN(n9130) );
  INVX0 U9187 ( .INP(n9009), .ZN(n9131) );
  INVX0 U9188 ( .INP(n9009), .ZN(n9132) );
  INVX0 U9189 ( .INP(n9010), .ZN(n9133) );
  INVX0 U9190 ( .INP(n9010), .ZN(n9134) );
  INVX0 U9191 ( .INP(n9010), .ZN(n9135) );
  INVX0 U9192 ( .INP(n9010), .ZN(n9136) );
  INVX0 U9193 ( .INP(n9010), .ZN(n9137) );
  INVX0 U9194 ( .INP(n9010), .ZN(n9138) );
  INVX0 U9195 ( .INP(n9010), .ZN(n9139) );
  INVX0 U9196 ( .INP(n9010), .ZN(n9140) );
  INVX0 U9197 ( .INP(n9011), .ZN(n9141) );
  INVX0 U9198 ( .INP(n9011), .ZN(n9142) );
  INVX0 U9199 ( .INP(n9011), .ZN(n9143) );
  INVX0 U9200 ( .INP(n9011), .ZN(n9144) );
  INVX0 U9201 ( .INP(n9011), .ZN(n9145) );
  INVX0 U9202 ( .INP(n9011), .ZN(n9146) );
  INVX0 U9203 ( .INP(n9011), .ZN(n9147) );
  INVX0 U9204 ( .INP(n9011), .ZN(n9148) );
  INVX0 U9205 ( .INP(n9011), .ZN(n9149) );
  INVX0 U9206 ( .INP(n9012), .ZN(n9150) );
  INVX0 U9207 ( .INP(n9012), .ZN(n9151) );
  INVX0 U9208 ( .INP(n9012), .ZN(n9152) );
  INVX0 U9209 ( .INP(n9012), .ZN(n9153) );
  INVX0 U9210 ( .INP(n9012), .ZN(n9154) );
  INVX0 U9211 ( .INP(n9012), .ZN(n9155) );
  INVX0 U9212 ( .INP(n9012), .ZN(n9156) );
  INVX0 U9213 ( .INP(n9012), .ZN(n9157) );
  INVX0 U9214 ( .INP(n9013), .ZN(n9158) );
  INVX0 U9215 ( .INP(n9013), .ZN(n9159) );
  INVX0 U9216 ( .INP(n9013), .ZN(n9160) );
  INVX0 U9217 ( .INP(n9013), .ZN(n9161) );
  INVX0 U9218 ( .INP(n9013), .ZN(n9162) );
  INVX0 U9219 ( .INP(n9013), .ZN(n9163) );
  INVX0 U9220 ( .INP(n9013), .ZN(n9164) );
  INVX0 U9221 ( .INP(n9014), .ZN(n9165) );
  INVX0 U9222 ( .INP(n9013), .ZN(n9166) );
  INVX0 U9223 ( .INP(n9014), .ZN(n9167) );
  INVX0 U9224 ( .INP(n9012), .ZN(n9168) );
  INVX0 U9225 ( .INP(n9013), .ZN(n9169) );
  INVX0 U9226 ( .INP(n9014), .ZN(n9170) );
  NBUFFX2 U9227 ( .INP(n9331), .Z(n9291) );
  NBUFFX2 U9228 ( .INP(n9330), .Z(n9292) );
  NBUFFX2 U9229 ( .INP(n9330), .Z(n9293) );
  NBUFFX2 U9230 ( .INP(n9330), .Z(n9296) );
  NBUFFX2 U9231 ( .INP(n9329), .Z(n9297) );
  NBUFFX2 U9232 ( .INP(n9329), .Z(n9298) );
  NBUFFX2 U9233 ( .INP(n9329), .Z(n9299) );
  NBUFFX2 U9234 ( .INP(n9328), .Z(n9300) );
  NBUFFX2 U9235 ( .INP(n9328), .Z(n9301) );
  NBUFFX2 U9236 ( .INP(n9328), .Z(n9304) );
  NBUFFX2 U9237 ( .INP(n9326), .Z(n9305) );
  NBUFFX2 U9238 ( .INP(n9326), .Z(n9307) );
  NBUFFX2 U9239 ( .INP(n9326), .Z(n9308) );
  NBUFFX2 U9240 ( .INP(n9323), .Z(n9309) );
  NBUFFX2 U9241 ( .INP(n9323), .Z(n9310) );
  NBUFFX2 U9242 ( .INP(n9323), .Z(n9311) );
  NBUFFX2 U9243 ( .INP(n9321), .Z(n9313) );
  NBUFFX2 U9244 ( .INP(n9321), .Z(n9315) );
  NBUFFX2 U9245 ( .INP(n9321), .Z(n9316) );
  NBUFFX2 U9246 ( .INP(n9320), .Z(n9317) );
  NBUFFX2 U9247 ( .INP(n9320), .Z(n9318) );
  NBUFFX2 U9248 ( .INP(n9320), .Z(n9319) );
  NBUFFX2 U9249 ( .INP(n9335), .Z(n9320) );
  NBUFFX2 U9250 ( .INP(n9335), .Z(n9321) );
  NBUFFX2 U9251 ( .INP(n9334), .Z(n9323) );
  NBUFFX2 U9252 ( .INP(n9334), .Z(n9326) );
  NBUFFX2 U9253 ( .INP(n9334), .Z(n9328) );
  NBUFFX2 U9254 ( .INP(n9333), .Z(n9329) );
  NBUFFX2 U9255 ( .INP(n9333), .Z(n9330) );
  NBUFFX2 U9256 ( .INP(n9333), .Z(n9331) );
  NBUFFX2 U9257 ( .INP(CK), .Z(n9333) );
  NBUFFX2 U9258 ( .INP(CK), .Z(n9334) );
  NBUFFX2 U9259 ( .INP(CK), .Z(n9335) );
  AND3X1 U9260 ( .IN1(n9337), .IN2(n9338), .IN3(n9339), .Q(n8802) );
  INVX0 U9261 ( .INP(n9341), .ZN(n865) );
  INVX0 U9262 ( .INP(n9342), .ZN(n795) );
  INVX0 U9263 ( .INP(n9343), .ZN(n791) );
  INVX0 U9264 ( .INP(n9344), .ZN(n789) );
  OR3X1 U9265 ( .IN1(n9345), .IN2(n9346), .IN3(n9347), .Q(n706) );
  AND2X1 U9266 ( .IN1(n9349), .IN2(n8729), .Q(n9347) );
  INVX0 U9267 ( .INP(n9350), .ZN(n9349) );
  AND2X1 U9268 ( .IN1(n9143), .IN2(g1548), .Q(n9346) );
  AND3X1 U9269 ( .IN1(n9350), .IN2(g1564), .IN3(n9064), .Q(n9345) );
  OR4X1 U9270 ( .IN1(n9353), .IN2(n9354), .IN3(n9355), .IN4(n9356), .Q(n5961)
         );
  AND2X1 U9271 ( .IN1(n8507), .IN2(n9358), .Q(n9356) );
  AND2X1 U9272 ( .IN1(n9359), .IN2(g5348), .Q(n9355) );
  AND2X1 U9273 ( .IN1(n8774), .IN2(n9360), .Q(n9354) );
  AND2X1 U9274 ( .IN1(g31860), .IN2(g5352), .Q(n9353) );
  OR4X1 U9275 ( .IN1(n9361), .IN2(n9362), .IN3(n9363), .IN4(n9364), .Q(n5960)
         );
  AND2X1 U9276 ( .IN1(n8753), .IN2(n9365), .Q(n9364) );
  AND2X1 U9277 ( .IN1(n9366), .IN2(g6736), .Q(n9363) );
  AND2X1 U9278 ( .IN1(n8506), .IN2(n9368), .Q(n9362) );
  AND2X1 U9279 ( .IN1(n9369), .IN2(g6732), .Q(n9361) );
  INVX0 U9280 ( .INP(n9370), .ZN(n581) );
  INVX0 U9281 ( .INP(n9371), .ZN(n580) );
  OR3X1 U9282 ( .IN1(n9372), .IN2(n9373), .IN3(n9374), .Q(n568) );
  AND2X1 U9283 ( .IN1(n9375), .IN2(g3845), .Q(n9374) );
  AND4X1 U9284 ( .IN1(n9376), .IN2(n9081), .IN3(n5662), .IN4(n8858), .Q(n9373)
         );
  AND2X1 U9285 ( .IN1(test_so97), .IN2(n9377), .Q(n9372) );
  OR2X1 U9286 ( .IN1(n9130), .IN2(n9378), .Q(n9377) );
  AND2X1 U9287 ( .IN1(n9376), .IN2(g3835), .Q(n9378) );
  INVX0 U9288 ( .INP(n9379), .ZN(n4921) );
  INVX0 U9289 ( .INP(n9380), .ZN(n4896) );
  OR2X1 U9290 ( .IN1(n8628), .IN2(n9381), .Q(n4459) );
  OR2X1 U9291 ( .IN1(n8632), .IN2(n9382), .Q(n4448) );
  OR2X1 U9292 ( .IN1(n9383), .IN2(n8849), .Q(n4437) );
  OR2X1 U9293 ( .IN1(n8626), .IN2(n9384), .Q(n4426) );
  OR2X1 U9294 ( .IN1(n8634), .IN2(n9385), .Q(n4415) );
  OR2X1 U9295 ( .IN1(n8630), .IN2(n9386), .Q(n4403) );
  OR2X1 U9296 ( .IN1(n8623), .IN2(n9387), .Q(n4392) );
  OR2X1 U9297 ( .IN1(n8621), .IN2(n9388), .Q(n4380) );
  OR4X1 U9298 ( .IN1(n9389), .IN2(n9390), .IN3(n9391), .IN4(n9392), .Q(n4305)
         );
  OR2X1 U9299 ( .IN1(n9393), .IN2(n9394), .Q(n9392) );
  AND2X1 U9300 ( .IN1(g4646), .IN2(g29220), .Q(n9394) );
  AND2X1 U9301 ( .IN1(n5880), .IN2(g4674), .Q(n9393) );
  AND2X1 U9302 ( .IN1(g4831), .IN2(g4681), .Q(n9391) );
  AND3X1 U9303 ( .IN1(n9395), .IN2(n9396), .IN3(n5656), .Q(n9390) );
  OR3X1 U9304 ( .IN1(n9397), .IN2(n9398), .IN3(n9399), .Q(n9396) );
  AND3X1 U9305 ( .IN1(n9400), .IN2(n9401), .IN3(n5707), .Q(n9399) );
  OR2X1 U9306 ( .IN1(n5368), .IN2(g34657), .Q(n9401) );
  OR2X1 U9307 ( .IN1(n9402), .IN2(g4793), .Q(n9400) );
  AND2X1 U9308 ( .IN1(n9403), .IN2(n8836), .Q(n9402) );
  OR3X1 U9309 ( .IN1(n9404), .IN2(n9405), .IN3(n9406), .Q(n9403) );
  AND2X1 U9310 ( .IN1(n9407), .IN2(n5867), .Q(n9406) );
  AND2X1 U9311 ( .IN1(n9408), .IN2(n9409), .Q(n9398) );
  OR2X1 U9312 ( .IN1(n9410), .IN2(n9411), .Q(n9409) );
  AND2X1 U9313 ( .IN1(n9412), .IN2(g34657), .Q(n9411) );
  INVX0 U9314 ( .INP(n9413), .ZN(n9410) );
  OR2X1 U9316 ( .IN1(n9412), .IN2(g34657), .Q(n9413) );
  INVX0 U9317 ( .INP(n9414), .ZN(n9412) );
  OR4X1 U9318 ( .IN1(n9415), .IN2(n9416), .IN3(n9417), .IN4(n9418), .Q(n9414)
         );
  AND2X1 U9319 ( .IN1(n9407), .IN2(g4727), .Q(n9418) );
  AND3X1 U9320 ( .IN1(n5361), .IN2(g4722), .IN3(n5518), .Q(n9417) );
  AND2X1 U9321 ( .IN1(n9404), .IN2(g4717), .Q(n9416) );
  AND2X1 U9322 ( .IN1(n9405), .IN2(g4732), .Q(n9415) );
  AND2X1 U9323 ( .IN1(n8337), .IN2(g4688), .Q(n9389) );
  OR4X1 U9324 ( .IN1(n9419), .IN2(n9420), .IN3(n9421), .IN4(n9422), .Q(n4283)
         );
  OR2X1 U9325 ( .IN1(n9423), .IN2(n9424), .Q(n9422) );
  AND2X1 U9326 ( .IN1(g4871), .IN2(g3684), .Q(n9424) );
  AND2X1 U9327 ( .IN1(n8340), .IN2(g4864), .Q(n9423) );
  AND2X1 U9328 ( .IN1(g4836), .IN2(g5011), .Q(n9421) );
  AND3X1 U9329 ( .IN1(n9425), .IN2(n9426), .IN3(n5283), .Q(n9420) );
  OR3X1 U9330 ( .IN1(n9427), .IN2(n9428), .IN3(n9429), .Q(n9426) );
  AND3X1 U9331 ( .IN1(n9430), .IN2(n9431), .IN3(n5706), .Q(n9429) );
  OR2X1 U9332 ( .IN1(n5367), .IN2(g34649), .Q(n9431) );
  OR2X1 U9333 ( .IN1(n9432), .IN2(g4983), .Q(n9430) );
  AND2X1 U9334 ( .IN1(n9433), .IN2(n8837), .Q(n9432) );
  OR3X1 U9335 ( .IN1(n9434), .IN2(n9435), .IN3(n9436), .Q(n9433) );
  AND2X1 U9336 ( .IN1(n9437), .IN2(n5879), .Q(n9436) );
  AND2X1 U9337 ( .IN1(n9438), .IN2(n9439), .Q(n9428) );
  OR2X1 U9338 ( .IN1(n9440), .IN2(n9441), .Q(n9439) );
  AND2X1 U9339 ( .IN1(n9442), .IN2(g34649), .Q(n9441) );
  INVX0 U9340 ( .INP(n9443), .ZN(n9440) );
  OR2X1 U9341 ( .IN1(n9442), .IN2(g34649), .Q(n9443) );
  INVX0 U9342 ( .INP(n9444), .ZN(n9442) );
  OR4X1 U9343 ( .IN1(n9445), .IN2(n9446), .IN3(n9447), .IN4(n9448), .Q(n9444)
         );
  AND2X1 U9344 ( .IN1(n9437), .IN2(g4917), .Q(n9448) );
  AND3X1 U9345 ( .IN1(n5360), .IN2(g4912), .IN3(n5517), .Q(n9447) );
  AND2X1 U9346 ( .IN1(n9434), .IN2(g4907), .Q(n9446) );
  AND2X1 U9347 ( .IN1(n9435), .IN2(g4922), .Q(n9445) );
  AND2X1 U9348 ( .IN1(n8341), .IN2(g4878), .Q(n9419) );
  INVX0 U9349 ( .INP(n9449), .ZN(n4210) );
  AND3X1 U9350 ( .IN1(n5652), .IN2(n5366), .IN3(n8644), .Q(n4034) );
  AND3X1 U9351 ( .IN1(n5645), .IN2(n5576), .IN3(n8637), .Q(n4002) );
  INVX0 U9352 ( .INP(n9450), .ZN(n399) );
  AND2X1 U9353 ( .IN1(n3064), .IN2(n9451), .Q(n9450) );
  OR2X1 U9354 ( .IN1(n5715), .IN2(n9452), .Q(n9451) );
  AND2X1 U9355 ( .IN1(n9453), .IN2(n9026), .Q(n9452) );
  OR2X1 U9356 ( .IN1(g4104), .IN2(n9454), .Q(n9453) );
  AND3X1 U9357 ( .IN1(n5572), .IN2(n8823), .IN3(n8639), .Q(n3969) );
  AND4X1 U9358 ( .IN1(n9337), .IN2(n9338), .IN3(n2760), .IN4(g43), .Q(n3933)
         );
  AND3X1 U9359 ( .IN1(n5650), .IN2(n5570), .IN3(n8642), .Q(n3926) );
  AND3X1 U9360 ( .IN1(n5647), .IN2(n5575), .IN3(n8640), .Q(n3893) );
  AND3X1 U9361 ( .IN1(n5649), .IN2(n5573), .IN3(n8638), .Q(n3860) );
  AND3X1 U9362 ( .IN1(n5651), .IN2(n5574), .IN3(n8641), .Q(n3826) );
  AND3X1 U9363 ( .IN1(n5646), .IN2(n5571), .IN3(n8643), .Q(n3792) );
  OR4X1 U9364 ( .IN1(g691), .IN2(g417), .IN3(n9455), .IN4(n9456), .Q(n3675) );
  AND2X1 U9365 ( .IN1(n9457), .IN2(g392), .Q(n9456) );
  OR3X1 U9366 ( .IN1(n9458), .IN2(n9459), .IN3(g441), .Q(n9457) );
  AND2X1 U9367 ( .IN1(n8419), .IN2(n8834), .Q(n9459) );
  AND2X1 U9368 ( .IN1(test_so72), .IN2(g452), .Q(n9458) );
  AND2X1 U9369 ( .IN1(n8673), .IN2(n9460), .Q(n9455) );
  OR3X1 U9370 ( .IN1(n9461), .IN2(n9462), .IN3(g411), .Q(n9460) );
  AND2X1 U9371 ( .IN1(n5402), .IN2(n8834), .Q(n9462) );
  AND2X1 U9372 ( .IN1(test_so72), .IN2(g174), .Q(n9461) );
  OR2X1 U9373 ( .IN1(n5349), .IN2(n9463), .Q(n3635) );
  OR2X1 U9374 ( .IN1(n9464), .IN2(n9465), .Q(n353) );
  INVX0 U9375 ( .INP(n9466), .ZN(n9465) );
  INVX0 U9376 ( .INP(n9467), .ZN(n342) );
  INVX0 U9377 ( .INP(n9468), .ZN(n338) );
  AND2X1 U9378 ( .IN1(n9469), .IN2(n9470), .Q(n3174) );
  OR2X1 U9379 ( .IN1(n9471), .IN2(n9472), .Q(n9470) );
  AND2X1 U9380 ( .IN1(g73), .IN2(g490), .Q(n9472) );
  AND2X1 U9381 ( .IN1(n5708), .IN2(n9473), .Q(n9471) );
  OR2X1 U9382 ( .IN1(n9474), .IN2(n9475), .Q(n9469) );
  AND2X1 U9383 ( .IN1(n5820), .IN2(n9476), .Q(n9475) );
  AND2X1 U9384 ( .IN1(g72), .IN2(g482), .Q(n9474) );
  AND2X1 U9385 ( .IN1(n2760), .IN2(n9302), .Q(n3084) );
  OR3X1 U9386 ( .IN1(n8693), .IN2(n9121), .IN3(n9477), .Q(n3065) );
  AND2X1 U9387 ( .IN1(n9478), .IN2(g4108), .Q(n9477) );
  OR3X1 U9388 ( .IN1(n9479), .IN2(n9480), .IN3(n9481), .Q(n297) );
  AND2X1 U9389 ( .IN1(n8730), .IN2(n9482), .Q(n9481) );
  INVX0 U9390 ( .INP(n9483), .ZN(n9482) );
  AND2X1 U9391 ( .IN1(n9161), .IN2(g1205), .Q(n9480) );
  AND3X1 U9392 ( .IN1(n9483), .IN2(g1221), .IN3(n9066), .Q(n9479) );
  OR2X1 U9393 ( .IN1(n9484), .IN2(n9485), .Q(n2608) );
  AND2X1 U9394 ( .IN1(n2607), .IN2(g4311), .Q(n9485) );
  AND2X1 U9395 ( .IN1(n5323), .IN2(n9486), .Q(n9484) );
  INVX0 U9396 ( .INP(n2607), .ZN(n9486) );
  AND2X1 U9397 ( .IN1(n9466), .IN2(g34971), .Q(n2396) );
  OR3X1 U9398 ( .IN1(n9487), .IN2(n9488), .IN3(n9489), .Q(n227) );
  AND2X1 U9399 ( .IN1(n9490), .IN2(g5152), .Q(n9489) );
  AND4X1 U9400 ( .IN1(g32975), .IN2(n9081), .IN3(n5658), .IN4(n8859), .Q(n9488) );
  AND2X1 U9401 ( .IN1(test_so98), .IN2(n9491), .Q(n9487) );
  OR2X1 U9402 ( .IN1(n9130), .IN2(n9492), .Q(n9491) );
  AND2X1 U9403 ( .IN1(g32975), .IN2(g5142), .Q(n9492) );
  INVX0 U9404 ( .INP(n9493), .ZN(n218) );
  INVX0 U9405 ( .INP(n9494), .ZN(n217) );
  INVX0 U9406 ( .INP(n9495), .ZN(n209) );
  OR3X1 U9407 ( .IN1(n9496), .IN2(n9497), .IN3(n9498), .Q(n178) );
  INVX0 U9408 ( .INP(n9499), .ZN(n9498) );
  OR2X1 U9409 ( .IN1(n9500), .IN2(n9501), .Q(n9499) );
  AND3X1 U9410 ( .IN1(n9502), .IN2(g3462), .IN3(n8821), .Q(n9497) );
  AND2X1 U9411 ( .IN1(test_so4), .IN2(n9503), .Q(n9496) );
  OR2X1 U9412 ( .IN1(n9131), .IN2(n9504), .Q(n9503) );
  AND2X1 U9413 ( .IN1(n8723), .IN2(n9501), .Q(n9504) );
  INVX0 U9414 ( .INP(n9505), .ZN(n1731) );
  INVX0 U9415 ( .INP(n9506), .ZN(n1373) );
  INVX0 U9416 ( .INP(n9507), .ZN(n1371) );
  INVX0 U9417 ( .INP(n9508), .ZN(n1369) );
  INVX0 U9418 ( .INP(n9509), .ZN(n1367) );
  INVX0 U9419 ( .INP(n9510), .ZN(n1122) );
  INVX0 U9420 ( .INP(n9511), .ZN(n1039) );
  OR2X1 U9421 ( .IN1(n9512), .IN2(n9513), .Q(g34980) );
  AND2X1 U9422 ( .IN1(n9514), .IN2(n9026), .Q(n9513) );
  OR2X1 U9423 ( .IN1(n9515), .IN2(g2984), .Q(n9514) );
  AND4X1 U9424 ( .IN1(n8801), .IN2(n9516), .IN3(n9517), .IN4(n9518), .Q(n9515)
         );
  AND2X1 U9425 ( .IN1(test_so14), .IN2(n9138), .Q(n9512) );
  OR2X1 U9426 ( .IN1(n8789), .IN2(n8801), .Q(g34972) );
  OR2X1 U9427 ( .IN1(n9519), .IN2(n9520), .Q(n8801) );
  INVX0 U9428 ( .INP(n9521), .ZN(n9520) );
  OR2X1 U9429 ( .IN1(n9522), .IN2(n9523), .Q(n9521) );
  AND2X1 U9430 ( .IN1(n9523), .IN2(n9522), .Q(n9519) );
  AND2X1 U9431 ( .IN1(n9524), .IN2(n9525), .Q(n9522) );
  INVX0 U9432 ( .INP(n9526), .ZN(n9525) );
  AND2X1 U9433 ( .IN1(n9527), .IN2(n9528), .Q(n9526) );
  OR2X1 U9434 ( .IN1(n9528), .IN2(n9527), .Q(n9524) );
  OR2X1 U9435 ( .IN1(n9529), .IN2(n9530), .Q(n9527) );
  AND2X1 U9436 ( .IN1(g34975), .IN2(n9531), .Q(n9530) );
  INVX0 U9437 ( .INP(g34974), .ZN(n9531) );
  AND2X1 U9438 ( .IN1(g34974), .IN2(n9532), .Q(n9529) );
  INVX0 U9439 ( .INP(g34975), .ZN(n9532) );
  OR2X1 U9440 ( .IN1(n9533), .IN2(n8273), .Q(n9528) );
  AND2X1 U9441 ( .IN1(g54), .IN2(n9518), .Q(n9533) );
  INVX0 U9442 ( .INP(g56), .ZN(n9518) );
  OR2X1 U9443 ( .IN1(n9534), .IN2(n9535), .Q(n9523) );
  AND2X1 U9444 ( .IN1(n9536), .IN2(g34970), .Q(n9535) );
  INVX0 U9445 ( .INP(n9537), .ZN(n9534) );
  OR2X1 U9446 ( .IN1(n9536), .IN2(g34970), .Q(n9537) );
  OR2X1 U9447 ( .IN1(n9538), .IN2(n9539), .Q(n9536) );
  AND2X1 U9448 ( .IN1(n9540), .IN2(n9541), .Q(n9539) );
  INVX0 U9449 ( .INP(g34971), .ZN(n9541) );
  AND2X1 U9450 ( .IN1(n9542), .IN2(g34971), .Q(n9538) );
  INVX0 U9451 ( .INP(n9540), .ZN(n9542) );
  OR2X1 U9452 ( .IN1(n9543), .IN2(n9544), .Q(n9540) );
  AND3X1 U9454 ( .IN1(n9545), .IN2(n9546), .IN3(n9547), .Q(n9544) );
  OR2X1 U9455 ( .IN1(n9548), .IN2(n9549), .Q(n9547) );
  AND2X1 U9456 ( .IN1(g34977), .IN2(n9550), .Q(n9549) );
  AND2X1 U9457 ( .IN1(g34976), .IN2(n9551), .Q(n9548) );
  OR2X1 U9458 ( .IN1(g34979), .IN2(n9552), .Q(n9546) );
  OR2X1 U9459 ( .IN1(g34978), .IN2(n9464), .Q(n9545) );
  AND3X1 U9460 ( .IN1(n9553), .IN2(n9554), .IN3(n9555), .Q(n9543) );
  OR2X1 U9461 ( .IN1(n9556), .IN2(n9557), .Q(n9555) );
  AND2X1 U9462 ( .IN1(g34979), .IN2(n9552), .Q(n9557) );
  INVX0 U9463 ( .INP(g34978), .ZN(n9552) );
  AND2X1 U9464 ( .IN1(g34978), .IN2(n9464), .Q(n9556) );
  INVX0 U9465 ( .INP(g34979), .ZN(n9464) );
  OR2X1 U9466 ( .IN1(g34977), .IN2(n9550), .Q(n9554) );
  INVX0 U9467 ( .INP(g34976), .ZN(n9550) );
  OR2X1 U9468 ( .IN1(g34976), .IN2(n9551), .Q(n9553) );
  INVX0 U9469 ( .INP(g34977), .ZN(n9551) );
  OR2X1 U9470 ( .IN1(n8789), .IN2(g34979), .Q(g34927) );
  OR4X1 U9471 ( .IN1(n9558), .IN2(n9559), .IN3(n9560), .IN4(n9561), .Q(g34979)
         );
  OR4X1 U9472 ( .IN1(n9562), .IN2(n9563), .IN3(n9564), .IN4(n9565), .Q(n9561)
         );
  AND2X1 U9473 ( .IN1(n9566), .IN2(n9332), .Q(n9565) );
  AND2X1 U9474 ( .IN1(n9567), .IN2(g1283), .Q(n9564) );
  AND2X1 U9475 ( .IN1(n9568), .IN2(g2138), .Q(n9563) );
  AND2X1 U9476 ( .IN1(n9569), .IN2(g2697), .Q(n9562) );
  OR2X1 U9477 ( .IN1(n9570), .IN2(n9571), .Q(n9560) );
  AND2X1 U9478 ( .IN1(test_so67), .IN2(n9572), .Q(n9571) );
  AND2X1 U9479 ( .IN1(n9573), .IN2(g4146), .Q(n9570) );
  AND2X1 U9480 ( .IN1(n9574), .IN2(g939), .Q(n9559) );
  AND2X1 U9481 ( .IN1(n1430), .IN2(n9575), .Q(n9558) );
  OR4X1 U9482 ( .IN1(n9576), .IN2(n9577), .IN3(n9578), .IN4(n9579), .Q(n9575)
         );
  OR4X1 U9483 ( .IN1(n9580), .IN2(n9581), .IN3(n9582), .IN4(n9583), .Q(n9579)
         );
  OR3X1 U9484 ( .IN1(n9584), .IN2(n9585), .IN3(n9586), .Q(n9583) );
  AND2X1 U9485 ( .IN1(test_so14), .IN2(n9466), .Q(n9586) );
  AND2X1 U9486 ( .IN1(g92), .IN2(n9587), .Q(n9585) );
  AND2X1 U9487 ( .IN1(g127), .IN2(n9588), .Q(n9584) );
  AND2X1 U9488 ( .IN1(n9589), .IN2(g744), .Q(n9582) );
  AND2X1 U9489 ( .IN1(n9590), .IN2(g2886), .Q(n9581) );
  AND2X1 U9490 ( .IN1(n9591), .IN2(g785), .Q(n9580) );
  OR3X1 U9491 ( .IN1(n9592), .IN2(n9593), .IN3(n9594), .Q(n9578) );
  AND2X1 U9492 ( .IN1(n9595), .IN2(g2975), .Q(n9594) );
  AND2X1 U9493 ( .IN1(n9596), .IN2(g2970), .Q(n9593) );
  AND2X1 U9494 ( .IN1(n9597), .IN2(g604), .Q(n9592) );
  OR2X1 U9495 ( .IN1(n9598), .IN2(n9599), .Q(n9577) );
  AND2X1 U9496 ( .IN1(n9600), .IN2(g568), .Q(n9599) );
  AND2X1 U9497 ( .IN1(g29221), .IN2(n9601), .Q(n9598) );
  OR2X1 U9498 ( .IN1(n8789), .IN2(g34978), .Q(g34925) );
  OR4X1 U9499 ( .IN1(n9602), .IN2(n9603), .IN3(n9604), .IN4(n9605), .Q(g34978)
         );
  OR4X1 U9500 ( .IN1(n9606), .IN2(n9607), .IN3(n9608), .IN4(n9609), .Q(n9605)
         );
  AND2X1 U9501 ( .IN1(n9566), .IN2(n9276), .Q(n9609) );
  AND2X1 U9502 ( .IN1(n8275), .IN2(n9567), .Q(n9608) );
  AND2X1 U9503 ( .IN1(n9568), .IN2(g2130), .Q(n9607) );
  AND2X1 U9504 ( .IN1(n9569), .IN2(g2689), .Q(n9606) );
  OR2X1 U9505 ( .IN1(n9610), .IN2(n9611), .Q(n9604) );
  AND2X1 U9506 ( .IN1(n9572), .IN2(g4253), .Q(n9611) );
  AND2X1 U9507 ( .IN1(n9573), .IN2(g4176), .Q(n9610) );
  AND2X1 U9508 ( .IN1(n8276), .IN2(n9574), .Q(n9603) );
  AND2X1 U9509 ( .IN1(n1430), .IN2(n9612), .Q(n9602) );
  OR4X1 U9510 ( .IN1(n9613), .IN2(n9576), .IN3(n9614), .IN4(n9615), .Q(n9612)
         );
  OR4X1 U9511 ( .IN1(n9616), .IN2(n9617), .IN3(n9618), .IN4(n9619), .Q(n9615)
         );
  OR3X1 U9512 ( .IN1(n9620), .IN2(n9621), .IN3(n9622), .Q(n9619) );
  AND2X1 U9513 ( .IN1(n9591), .IN2(g790), .Q(n9622) );
  AND2X1 U9514 ( .IN1(n9587), .IN2(g29214), .Q(n9621) );
  AND2X1 U9515 ( .IN1(n9588), .IN2(g2873), .Q(n9620) );
  AND2X1 U9516 ( .IN1(n9597), .IN2(g608), .Q(n9618) );
  AND2X1 U9517 ( .IN1(test_so2), .IN2(n9589), .Q(n9617) );
  AND2X1 U9518 ( .IN1(n9590), .IN2(g2878), .Q(n9616) );
  OR3X1 U9519 ( .IN1(n9623), .IN2(n9624), .IN3(n9625), .Q(n9614) );
  AND2X1 U9520 ( .IN1(n8537), .IN2(n9601), .Q(n9625) );
  AND2X1 U9521 ( .IN1(n9595), .IN2(g2965), .Q(n9624) );
  AND2X1 U9522 ( .IN1(test_so22), .IN2(n9596), .Q(n9623) );
  AND2X1 U9523 ( .IN1(n9600), .IN2(g572), .Q(n9613) );
  OR2X1 U9524 ( .IN1(n8789), .IN2(g34977), .Q(g34923) );
  OR4X1 U9525 ( .IN1(n9626), .IN2(n9627), .IN3(n9628), .IN4(n9629), .Q(g34977)
         );
  OR4X1 U9526 ( .IN1(n9630), .IN2(n9576), .IN3(n9631), .IN4(n9632), .Q(n9629)
         );
  AND2X1 U9527 ( .IN1(n5867), .IN2(n9633), .Q(n9632) );
  AND2X1 U9528 ( .IN1(n9566), .IN2(n9245), .Q(n9631) );
  AND2X1 U9529 ( .IN1(n5879), .IN2(n9634), .Q(n9630) );
  OR3X1 U9530 ( .IN1(n9635), .IN2(n9636), .IN3(n9637), .Q(n9628) );
  AND2X1 U9531 ( .IN1(n1430), .IN2(n9638), .Q(n9637) );
  OR4X1 U9532 ( .IN1(n9639), .IN2(n9640), .IN3(n9641), .IN4(n9642), .Q(n9638)
         );
  OR4X1 U9533 ( .IN1(n9643), .IN2(n9644), .IN3(n9645), .IN4(n9646), .Q(n9642)
         );
  OR3X1 U9534 ( .IN1(n9647), .IN2(n9648), .IN3(n9649), .Q(n9646) );
  AND2X1 U9535 ( .IN1(g37), .IN2(n9587), .Q(n9649) );
  AND2X1 U9536 ( .IN1(n9588), .IN2(g2868), .Q(n9648) );
  AND2X1 U9537 ( .IN1(n9589), .IN2(g758), .Q(n9645) );
  AND2X1 U9538 ( .IN1(n9590), .IN2(g2882), .Q(n9644) );
  AND2X1 U9539 ( .IN1(n9591), .IN2(g794), .Q(n9643) );
  OR3X1 U9540 ( .IN1(n9650), .IN2(n9651), .IN3(n9652), .Q(n9641) );
  AND2X1 U9541 ( .IN1(n9595), .IN2(g2955), .Q(n9652) );
  AND2X1 U9542 ( .IN1(n9596), .IN2(g2950), .Q(n9651) );
  AND2X1 U9543 ( .IN1(n9597), .IN2(g613), .Q(n9650) );
  AND2X1 U9544 ( .IN1(n9600), .IN2(g586), .Q(n9640) );
  AND2X1 U9545 ( .IN1(n9601), .IN2(g534), .Q(n9639) );
  AND2X1 U9546 ( .IN1(n9572), .IN2(g4300), .Q(n9636) );
  AND2X1 U9547 ( .IN1(n9573), .IN2(g4172), .Q(n9635) );
  AND2X1 U9548 ( .IN1(n9567), .IN2(g1291), .Q(n9627) );
  AND2X1 U9549 ( .IN1(n9574), .IN2(g947), .Q(n9626) );
  OR2X1 U9550 ( .IN1(n8789), .IN2(g34976), .Q(g34921) );
  OR4X1 U9551 ( .IN1(n9653), .IN2(n9654), .IN3(n9655), .IN4(n9656), .Q(g34976)
         );
  OR4X1 U9552 ( .IN1(n9657), .IN2(n9576), .IN3(n9658), .IN4(n9659), .Q(n9656)
         );
  AND2X1 U9553 ( .IN1(n9633), .IN2(g4722), .Q(n9659) );
  AND2X1 U9554 ( .IN1(n9568), .IN2(g5160), .Q(n9658) );
  AND2X1 U9555 ( .IN1(n9634), .IN2(g4912), .Q(n9657) );
  OR3X1 U9556 ( .IN1(n9660), .IN2(n9661), .IN3(n9662), .Q(n9655) );
  AND2X1 U9557 ( .IN1(n1430), .IN2(n9663), .Q(n9662) );
  OR4X1 U9558 ( .IN1(n9664), .IN2(n9665), .IN3(n9666), .IN4(n9667), .Q(n9663)
         );
  OR4X1 U9559 ( .IN1(n9668), .IN2(n9669), .IN3(n9670), .IN4(n9671), .Q(n9667)
         );
  OR3X1 U9560 ( .IN1(n9647), .IN2(n9672), .IN3(n9673), .Q(n9671) );
  AND2X1 U9561 ( .IN1(n9591), .IN2(g807), .Q(n9673) );
  AND2X1 U9562 ( .IN1(n9588), .IN2(g2988), .Q(n9672) );
  AND2X1 U9563 ( .IN1(n9597), .IN2(g617), .Q(n9670) );
  AND2X1 U9564 ( .IN1(n9589), .IN2(g763), .Q(n9669) );
  AND2X1 U9565 ( .IN1(n9590), .IN2(g2898), .Q(n9668) );
  OR3X1 U9566 ( .IN1(n9674), .IN2(n9675), .IN3(n9676), .Q(n9666) );
  AND2X1 U9567 ( .IN1(n9595), .IN2(g2941), .Q(n9676) );
  AND2X1 U9568 ( .IN1(test_so95), .IN2(n9677), .Q(n9675) );
  AND2X1 U9569 ( .IN1(n9596), .IN2(g2936), .Q(n9674) );
  AND2X1 U9570 ( .IN1(n9600), .IN2(g577), .Q(n9665) );
  AND2X1 U9571 ( .IN1(test_so41), .IN2(n9601), .Q(n9664) );
  AND2X1 U9572 ( .IN1(n9678), .IN2(g1135), .Q(n9661) );
  AND2X1 U9573 ( .IN1(n9679), .IN2(g1478), .Q(n9660) );
  AND2X1 U9574 ( .IN1(n9569), .IN2(g6545), .Q(n9654) );
  AND2X1 U9575 ( .IN1(n9566), .IN2(n9357), .Q(n9653) );
  OR2X1 U9576 ( .IN1(n8789), .IN2(g34975), .Q(g34919) );
  OR4X1 U9577 ( .IN1(n9680), .IN2(n9681), .IN3(n9682), .IN4(n9683), .Q(g34975)
         );
  OR4X1 U9578 ( .IN1(n9684), .IN2(n9576), .IN3(n9685), .IN4(n9686), .Q(n9683)
         );
  AND2X1 U9579 ( .IN1(n9633), .IN2(g4717), .Q(n9686) );
  AND2X1 U9580 ( .IN1(n9568), .IN2(g5507), .Q(n9685) );
  AND2X1 U9581 ( .IN1(n9634), .IN2(g4907), .Q(n9684) );
  OR3X1 U9582 ( .IN1(n9687), .IN2(n9688), .IN3(n9689), .Q(n9682) );
  AND2X1 U9583 ( .IN1(n1430), .IN2(n9690), .Q(n9689) );
  OR4X1 U9584 ( .IN1(n9691), .IN2(n9692), .IN3(n9693), .IN4(n9694), .Q(n9690)
         );
  OR4X1 U9585 ( .IN1(n9695), .IN2(n9696), .IN3(n9697), .IN4(n9698), .Q(n9694)
         );
  OR2X1 U9586 ( .IN1(n9699), .IN2(n9700), .Q(n9698) );
  AND2X1 U9587 ( .IN1(n9591), .IN2(g554), .Q(n9700) );
  AND2X1 U9588 ( .IN1(n5634), .IN2(n9588), .Q(n9699) );
  AND2X1 U9589 ( .IN1(n9590), .IN2(g2864), .Q(n9697) );
  AND2X1 U9590 ( .IN1(n9597), .IN2(g622), .Q(n9696) );
  AND2X1 U9591 ( .IN1(n9589), .IN2(g767), .Q(n9695) );
  OR3X1 U9592 ( .IN1(n9701), .IN2(n9702), .IN3(n9703), .Q(n9693) );
  AND2X1 U9593 ( .IN1(n9595), .IN2(g2927), .Q(n9703) );
  AND2X1 U9594 ( .IN1(n9677), .IN2(g2860), .Q(n9702) );
  AND2X1 U9595 ( .IN1(n9596), .IN2(g2922), .Q(n9701) );
  AND2X1 U9596 ( .IN1(n9600), .IN2(g582), .Q(n9692) );
  AND2X1 U9597 ( .IN1(n9601), .IN2(g546), .Q(n9691) );
  AND2X1 U9598 ( .IN1(n9678), .IN2(g1105), .Q(n9688) );
  AND2X1 U9599 ( .IN1(n9679), .IN2(g1448), .Q(n9687) );
  AND2X1 U9600 ( .IN1(n9569), .IN2(g3151), .Q(n9681) );
  AND2X1 U9601 ( .IN1(n9566), .IN2(n9294), .Q(n9680) );
  OR2X1 U9602 ( .IN1(n8789), .IN2(g34974), .Q(g34917) );
  OR4X1 U9603 ( .IN1(n9704), .IN2(n9705), .IN3(n9706), .IN4(n9707), .Q(g34974)
         );
  OR4X1 U9604 ( .IN1(n9708), .IN2(n9709), .IN3(n9710), .IN4(n9711), .Q(n9707)
         );
  AND2X1 U9605 ( .IN1(n9568), .IN2(g5853), .Q(n9711) );
  AND2X1 U9606 ( .IN1(test_so45), .IN2(n9569), .Q(n9710) );
  AND2X1 U9607 ( .IN1(n9634), .IN2(g4922), .Q(n9709) );
  AND2X1 U9608 ( .IN1(n9633), .IN2(g4732), .Q(n9708) );
  OR3X1 U9609 ( .IN1(n9712), .IN2(n9713), .IN3(n9714), .Q(n9706) );
  AND2X1 U9610 ( .IN1(n9678), .IN2(g1129), .Q(n9714) );
  AND2X1 U9611 ( .IN1(n9679), .IN2(g1472), .Q(n9713) );
  AND2X1 U9612 ( .IN1(n9566), .IN2(n9327), .Q(n9705) );
  AND2X1 U9613 ( .IN1(n1430), .IN2(n9715), .Q(n9704) );
  OR2X1 U9614 ( .IN1(n9716), .IN2(n9717), .Q(n9715) );
  OR4X1 U9615 ( .IN1(n9718), .IN2(n9719), .IN3(n9720), .IN4(n9721), .Q(n9717)
         );
  AND2X1 U9616 ( .IN1(n9677), .IN2(g2852), .Q(n9721) );
  AND2X1 U9617 ( .IN1(n9596), .IN2(g2912), .Q(n9720) );
  AND2X1 U9618 ( .IN1(n9600), .IN2(g590), .Q(n9719) );
  AND2X1 U9619 ( .IN1(n9595), .IN2(g2917), .Q(n9718) );
  OR4X1 U9620 ( .IN1(n9722), .IN2(n9723), .IN3(n9724), .IN4(n9725), .Q(n9716)
         );
  AND2X1 U9621 ( .IN1(n9590), .IN2(g2856), .Q(n9725) );
  AND2X1 U9622 ( .IN1(n9588), .IN2(g2999), .Q(n9724) );
  AND2X1 U9623 ( .IN1(n9597), .IN2(g626), .Q(n9723) );
  AND2X1 U9624 ( .IN1(n9589), .IN2(g772), .Q(n9722) );
  OR2X1 U9625 ( .IN1(n8789), .IN2(g34971), .Q(g34915) );
  OR4X1 U9626 ( .IN1(n9726), .IN2(n9727), .IN3(n9728), .IN4(n9729), .Q(g34971)
         );
  OR4X1 U9627 ( .IN1(n9730), .IN2(n9731), .IN3(n9732), .IN4(n9733), .Q(n9729)
         );
  AND2X1 U9628 ( .IN1(n9566), .IN2(n9351), .Q(n9733) );
  AND2X1 U9629 ( .IN1(test_so64), .IN2(n9567), .Q(n9732) );
  AND2X1 U9630 ( .IN1(n9568), .IN2(g2145), .Q(n9731) );
  AND2X1 U9631 ( .IN1(n9569), .IN2(g2704), .Q(n9730) );
  OR2X1 U9632 ( .IN1(n9734), .IN2(n9735), .Q(n9728) );
  AND2X1 U9633 ( .IN1(n9572), .IN2(g4245), .Q(n9735) );
  AND2X1 U9634 ( .IN1(n9736), .IN2(n9737), .Q(n9572) );
  AND2X1 U9635 ( .IN1(n9573), .IN2(g4157), .Q(n9734) );
  AND2X1 U9636 ( .IN1(n1430), .IN2(n9677), .Q(n9573) );
  AND2X1 U9637 ( .IN1(n9574), .IN2(n9247), .Q(n9727) );
  AND2X1 U9638 ( .IN1(n1430), .IN2(n9738), .Q(n9726) );
  OR4X1 U9639 ( .IN1(n9739), .IN2(n9576), .IN3(n9740), .IN4(n9741), .Q(n9738)
         );
  OR4X1 U9640 ( .IN1(n9742), .IN2(n9743), .IN3(n9744), .IN4(n9745), .Q(n9741)
         );
  OR2X1 U9641 ( .IN1(n9647), .IN2(n9746), .Q(n9745) );
  AND2X1 U9642 ( .IN1(n9588), .IN2(g2890), .Q(n9746) );
  AND2X1 U9643 ( .IN1(n9747), .IN2(n9736), .Q(n9588) );
  AND4X1 U9644 ( .IN1(g28), .IN2(n9748), .IN3(n5477), .IN4(g19), .Q(n9647) );
  AND2X1 U9645 ( .IN1(g100), .IN2(n9587), .Q(n9744) );
  AND3X1 U9646 ( .IN1(g28), .IN2(n9749), .IN3(n9747), .Q(n9587) );
  AND2X1 U9647 ( .IN1(n9591), .IN2(g781), .Q(n9743) );
  AND2X1 U9648 ( .IN1(n9466), .IN2(g2984), .Q(n9742) );
  AND4X1 U9649 ( .IN1(test_so25), .IN2(n9748), .IN3(n5324), .IN4(n8777), .Q(
        n9466) );
  OR3X1 U9650 ( .IN1(n9750), .IN2(n9751), .IN3(n9752), .Q(n9740) );
  AND2X1 U9651 ( .IN1(n9601), .IN2(g199), .Q(n9752) );
  AND2X1 U9652 ( .IN1(n9597), .IN2(g599), .Q(n9751) );
  AND2X1 U9653 ( .IN1(test_so60), .IN2(n9589), .Q(n9750) );
  OR2X1 U9654 ( .IN1(n9753), .IN2(n9712), .Q(n9576) );
  AND2X1 U9655 ( .IN1(n9591), .IN2(n9754), .Q(n9753) );
  AND2X1 U9656 ( .IN1(n9755), .IN2(n9736), .Q(n9591) );
  AND2X1 U9657 ( .IN1(n9600), .IN2(g562), .Q(n9739) );
  OR2X1 U9658 ( .IN1(n8789), .IN2(g34970), .Q(g34913) );
  OR4X1 U9659 ( .IN1(n9756), .IN2(n9757), .IN3(n9758), .IN4(n9759), .Q(g34970)
         );
  OR4X1 U9660 ( .IN1(n9760), .IN2(n9761), .IN3(n9762), .IN4(n9763), .Q(n9759)
         );
  AND2X1 U9661 ( .IN1(n1430), .IN2(n9764), .Q(n9763) );
  OR2X1 U9662 ( .IN1(n9765), .IN2(n9766), .Q(n9764) );
  OR4X1 U9663 ( .IN1(n9767), .IN2(n9768), .IN3(n9769), .IN4(n9770), .Q(n9766)
         );
  AND2X1 U9664 ( .IN1(n9595), .IN2(g2902), .Q(n9770) );
  AND3X1 U9665 ( .IN1(n5324), .IN2(n9771), .IN3(n9748), .Q(n9595) );
  AND2X1 U9666 ( .IN1(n9677), .IN2(g2844), .Q(n9769) );
  AND3X1 U9667 ( .IN1(g9), .IN2(n9772), .IN3(n9771), .Q(n9677) );
  AND2X1 U9668 ( .IN1(n9600), .IN2(g595), .Q(n9768) );
  AND2X1 U9669 ( .IN1(n9601), .IN2(g538), .Q(n9767) );
  AND2X1 U9670 ( .IN1(n9772), .IN2(n9755), .Q(n9601) );
  OR4X1 U9671 ( .IN1(n9773), .IN2(n9774), .IN3(n9775), .IN4(n9776), .Q(n9765)
         );
  AND2X1 U9672 ( .IN1(n9589), .IN2(g776), .Q(n9776) );
  AND2X1 U9673 ( .IN1(n9590), .IN2(g2848), .Q(n9775) );
  AND3X1 U9674 ( .IN1(g9), .IN2(n9771), .IN3(n9736), .Q(n9590) );
  AND2X1 U9675 ( .IN1(test_so1), .IN2(n9596), .Q(n9774) );
  AND3X1 U9676 ( .IN1(g28), .IN2(n9771), .IN3(n9748), .Q(n9596) );
  AND4X1 U9677 ( .IN1(n3395), .IN2(test_so85), .IN3(g8), .IN4(g9), .Q(n9748)
         );
  AND2X1 U9678 ( .IN1(n9597), .IN2(n9340), .Q(n9773) );
  AND2X1 U9679 ( .IN1(n9568), .IN2(g6199), .Q(n9762) );
  AND2X1 U9680 ( .IN1(n9772), .IN2(n9737), .Q(n9568) );
  AND2X1 U9681 ( .IN1(n9634), .IN2(g4917), .Q(n9761) );
  AND3X1 U9682 ( .IN1(n1430), .IN2(n9736), .IN3(n2527), .Q(n9634) );
  AND2X1 U9683 ( .IN1(n9633), .IN2(g4727), .Q(n9760) );
  AND3X1 U9684 ( .IN1(n1430), .IN2(n9772), .IN3(n2527), .Q(n9633) );
  OR3X1 U9685 ( .IN1(n9712), .IN2(n9777), .IN3(n9778), .Q(n9758) );
  AND2X1 U9686 ( .IN1(n9678), .IN2(g956), .Q(n9778) );
  AND2X1 U9687 ( .IN1(n9574), .IN2(n5286), .Q(n9678) );
  AND3X1 U9688 ( .IN1(n1430), .IN2(n2552), .IN3(n9736), .Q(n9574) );
  AND3X1 U9689 ( .IN1(g28), .IN2(n9779), .IN3(n5469), .Q(n9736) );
  AND2X1 U9690 ( .IN1(n9679), .IN2(g1300), .Q(n9777) );
  AND2X1 U9691 ( .IN1(n9567), .IN2(n2549), .Q(n9679) );
  AND3X1 U9692 ( .IN1(n1430), .IN2(n9772), .IN3(n9747), .Q(n9567) );
  AND3X1 U9693 ( .IN1(n8777), .IN2(n5468), .IN3(test_so25), .Q(n9747) );
  AND2X1 U9694 ( .IN1(n9780), .IN2(n9754), .Q(n9712) );
  AND2X1 U9695 ( .IN1(n9159), .IN2(n1430), .Q(n9754) );
  OR3X1 U9696 ( .IN1(n9597), .IN2(n9600), .IN3(n9589), .Q(n9780) );
  AND3X1 U9697 ( .IN1(g28), .IN2(n9749), .IN3(n9755), .Q(n9589) );
  AND2X1 U9698 ( .IN1(n9771), .IN2(n5468), .Q(n9755) );
  AND2X1 U9699 ( .IN1(n5477), .IN2(n8777), .Q(n9771) );
  AND3X1 U9700 ( .IN1(n9749), .IN2(n2552), .IN3(n5324), .Q(n9600) );
  AND2X1 U9701 ( .IN1(n2552), .IN2(n9772), .Q(n9597) );
  AND3X1 U9702 ( .IN1(n9779), .IN2(n5324), .IN3(n5469), .Q(n9772) );
  INVX0 U9703 ( .INP(n9781), .ZN(n9779) );
  AND2X1 U9704 ( .IN1(n9569), .IN2(g3853), .Q(n9757) );
  AND3X1 U9705 ( .IN1(n9749), .IN2(n5324), .IN3(n9737), .Q(n9569) );
  AND4X1 U9706 ( .IN1(g9), .IN2(n1430), .IN3(n5477), .IN4(g19), .Q(n9737) );
  INVX0 U9707 ( .INP(n9782), .ZN(n1430) );
  INVX0 U9708 ( .INP(n9783), .ZN(n9749) );
  OR2X1 U9709 ( .IN1(n5469), .IN2(n9781), .Q(n9783) );
  OR3X1 U9710 ( .IN1(test_so85), .IN2(g8), .IN3(g6), .Q(n9781) );
  AND2X1 U9711 ( .IN1(n9566), .IN2(n9322), .Q(n9756) );
  AND2X1 U9712 ( .IN1(n9516), .IN2(n9782), .Q(n9566) );
  OR4X1 U9713 ( .IN1(g53), .IN2(n9517), .IN3(g56), .IN4(n9784), .Q(n9782) );
  OR2X1 U9714 ( .IN1(test_so74), .IN2(g57), .Q(n9784) );
  INVX0 U9715 ( .INP(g54), .ZN(n9517) );
  INVX0 U9716 ( .INP(g53), .ZN(n9516) );
  OR2X1 U9717 ( .IN1(n9785), .IN2(n9786), .Q(g34911) );
  AND2X1 U9718 ( .IN1(n2404), .IN2(g554), .Q(n9786) );
  AND2X1 U9719 ( .IN1(n9787), .IN2(g807), .Q(n9785) );
  OR2X1 U9720 ( .IN1(n2405), .IN2(n9122), .Q(n9787) );
  OR2X1 U9721 ( .IN1(n9788), .IN2(n9789), .Q(g34882) );
  AND2X1 U9722 ( .IN1(n9790), .IN2(n9026), .Q(n9789) );
  OR3X1 U9723 ( .IN1(n9791), .IN2(n9792), .IN3(n9793), .Q(n9790) );
  AND3X1 U9724 ( .IN1(n5653), .IN2(n9794), .IN3(n9795), .Q(n9793) );
  OR2X1 U9725 ( .IN1(g4358), .IN2(n9796), .Q(n9794) );
  AND3X1 U9726 ( .IN1(n9796), .IN2(n8822), .IN3(n5348), .Q(n9792) );
  OR4X1 U9727 ( .IN1(test_so81), .IN2(g4340), .IN3(n9797), .IN4(n9798), .Q(
        n9796) );
  AND3X1 U9728 ( .IN1(n5506), .IN2(g4311), .IN3(g4332), .Q(n9798) );
  AND2X1 U9729 ( .IN1(n5540), .IN2(n9799), .Q(n9797) );
  OR3X1 U9730 ( .IN1(n9800), .IN2(n9801), .IN3(n9802), .Q(n9799) );
  AND3X1 U9731 ( .IN1(g90), .IN2(n5634), .IN3(n5506), .Q(n9801) );
  AND2X1 U9732 ( .IN1(n8552), .IN2(g4322), .Q(n9800) );
  AND3X1 U9733 ( .IN1(test_so81), .IN2(g4340), .IN3(g4358), .Q(n9791) );
  AND2X1 U9734 ( .IN1(n9156), .IN2(g4366), .Q(n9788) );
  OR3X1 U9735 ( .IN1(n9803), .IN2(n9804), .IN3(n9805), .Q(g34881) );
  AND2X1 U9736 ( .IN1(n9156), .IN2(g794), .Q(n9805) );
  AND2X1 U9737 ( .IN1(n2405), .IN2(n5479), .Q(n9804) );
  AND3X1 U9738 ( .IN1(n2404), .IN2(n9806), .IN3(g807), .Q(n9803) );
  INVX0 U9739 ( .INP(n2405), .ZN(n9806) );
  OR3X1 U9740 ( .IN1(n9807), .IN2(n9808), .IN3(n9809), .Q(g34880) );
  AND2X1 U9741 ( .IN1(n9156), .IN2(g626), .Q(n9809) );
  AND2X1 U9742 ( .IN1(n2422), .IN2(n15421), .Q(n9808) );
  AND3X1 U9743 ( .IN1(n2421), .IN2(n9810), .IN3(n9340), .Q(n9807) );
  INVX0 U9744 ( .INP(n2422), .ZN(n9810) );
  OR3X1 U9745 ( .IN1(n9811), .IN2(n9812), .IN3(n9813), .Q(g34850) );
  AND2X1 U9746 ( .IN1(n9156), .IN2(g790), .Q(n9813) );
  AND2X1 U9747 ( .IN1(n2419), .IN2(n5291), .Q(n9812) );
  AND3X1 U9748 ( .IN1(n2404), .IN2(n9814), .IN3(g794), .Q(n9811) );
  INVX0 U9749 ( .INP(n2419), .ZN(n9814) );
  OR3X1 U9750 ( .IN1(n9815), .IN2(n9816), .IN3(n9817), .Q(g34849) );
  AND2X1 U9751 ( .IN1(n9156), .IN2(g622), .Q(n9817) );
  AND2X1 U9752 ( .IN1(n2423), .IN2(n5288), .Q(n9816) );
  AND3X1 U9753 ( .IN1(n2421), .IN2(n9818), .IN3(g626), .Q(n9815) );
  INVX0 U9754 ( .INP(n2423), .ZN(n9818) );
  AND2X1 U9755 ( .IN1(n9819), .IN2(g4369), .Q(g34839) );
  OR3X1 U9756 ( .IN1(n9820), .IN2(n9821), .IN3(g4366), .Q(n9819) );
  AND2X1 U9757 ( .IN1(n9822), .IN2(g4332), .Q(n9821) );
  OR3X1 U9758 ( .IN1(n9823), .IN2(g4311), .IN3(n9824), .Q(n9822) );
  AND2X1 U9759 ( .IN1(n5540), .IN2(n9825), .Q(n9820) );
  OR3X1 U9760 ( .IN1(g73), .IN2(n9823), .IN3(g4311), .Q(n9825) );
  INVX0 U9761 ( .INP(n9826), .ZN(n9823) );
  OR2X1 U9762 ( .IN1(n9827), .IN2(n9828), .Q(g34808) );
  AND2X1 U9763 ( .IN1(n9829), .IN2(n9026), .Q(n9828) );
  OR3X1 U9764 ( .IN1(n9830), .IN2(n9831), .IN3(g2965), .Q(n9829) );
  AND2X1 U9765 ( .IN1(n9157), .IN2(g2955), .Q(n9827) );
  OR2X1 U9766 ( .IN1(n9832), .IN2(n9833), .Q(g34807) );
  AND2X1 U9767 ( .IN1(n9834), .IN2(n9027), .Q(n9833) );
  OR4X1 U9768 ( .IN1(n9835), .IN2(n9836), .IN3(n9837), .IN4(n9838), .Q(n9834)
         );
  OR3X1 U9769 ( .IN1(n9839), .IN2(g2955), .IN3(g2946), .Q(n9838) );
  AND2X1 U9770 ( .IN1(n9157), .IN2(g2941), .Q(n9832) );
  OR2X1 U9771 ( .IN1(n9840), .IN2(n9841), .Q(g34806) );
  AND2X1 U9772 ( .IN1(n9842), .IN2(n9027), .Q(n9841) );
  OR3X1 U9773 ( .IN1(g2941), .IN2(g4072), .IN3(g4153), .Q(n9842) );
  AND2X1 U9774 ( .IN1(n9157), .IN2(g2927), .Q(n9840) );
  AND2X1 U9775 ( .IN1(n9843), .IN2(n9027), .Q(g34805) );
  OR2X1 U9776 ( .IN1(g2932), .IN2(g2999), .Q(n9843) );
  OR2X1 U9777 ( .IN1(n9844), .IN2(n9845), .Q(g34804) );
  AND2X1 U9778 ( .IN1(n9846), .IN2(n9028), .Q(n9845) );
  OR3X1 U9779 ( .IN1(n5796), .IN2(n5630), .IN3(g2975), .Q(n9846) );
  AND2X1 U9780 ( .IN1(n9157), .IN2(g2965), .Q(n9844) );
  OR2X1 U9781 ( .IN1(n9847), .IN2(n9848), .Q(g34803) );
  AND2X1 U9782 ( .IN1(n9849), .IN2(n9028), .Q(n9848) );
  OR3X1 U9783 ( .IN1(g2932), .IN2(n9850), .IN3(g2927), .Q(n9849) );
  AND2X1 U9784 ( .IN1(n9157), .IN2(g2917), .Q(n9847) );
  OR2X1 U9785 ( .IN1(n9851), .IN2(n9852), .Q(g34802) );
  AND2X1 U9786 ( .IN1(n9853), .IN2(n9028), .Q(n9852) );
  OR3X1 U9787 ( .IN1(n9854), .IN2(n9855), .IN3(g2917), .Q(n9853) );
  AND2X1 U9788 ( .IN1(n9157), .IN2(g2902), .Q(n9851) );
  OR2X1 U9789 ( .IN1(n9856), .IN2(n9857), .Q(g34801) );
  AND2X1 U9790 ( .IN1(n9858), .IN2(n9028), .Q(n9857) );
  OR4X1 U9791 ( .IN1(g2902), .IN2(g301), .IN3(n5520), .IN4(g209), .Q(n9858) );
  AND2X1 U9792 ( .IN1(n9157), .IN2(g2970), .Q(n9856) );
  OR2X1 U9793 ( .IN1(n9859), .IN2(n9860), .Q(g34800) );
  AND2X1 U9794 ( .IN1(n9861), .IN2(n9028), .Q(n9860) );
  OR2X1 U9795 ( .IN1(test_so14), .IN2(test_so74), .Q(n9861) );
  AND2X1 U9796 ( .IN1(n9157), .IN2(g2886), .Q(n9859) );
  OR2X1 U9797 ( .IN1(n9862), .IN2(n9863), .Q(g34799) );
  AND2X1 U9798 ( .IN1(n9864), .IN2(n9028), .Q(n9863) );
  OR2X1 U9799 ( .IN1(n9850), .IN2(g2890), .Q(n9864) );
  INVX0 U9800 ( .INP(g44), .ZN(n9850) );
  AND2X1 U9801 ( .IN1(n9157), .IN2(g2873), .Q(n9862) );
  OR2X1 U9802 ( .IN1(n9865), .IN2(n9866), .Q(g34798) );
  AND2X1 U9803 ( .IN1(n9867), .IN2(n9028), .Q(n9866) );
  OR2X1 U9804 ( .IN1(g2946), .IN2(g2886), .Q(n9867) );
  AND2X1 U9805 ( .IN1(n9157), .IN2(g2878), .Q(n9865) );
  OR2X1 U9806 ( .IN1(n9868), .IN2(n9869), .Q(g34797) );
  AND2X1 U9807 ( .IN1(n9870), .IN2(n9028), .Q(n9869) );
  OR2X1 U9808 ( .IN1(n9831), .IN2(g2878), .Q(n9870) );
  INVX0 U9809 ( .INP(g91), .ZN(n9831) );
  AND2X1 U9810 ( .IN1(n9157), .IN2(g2882), .Q(n9868) );
  OR2X1 U9811 ( .IN1(n9871), .IN2(n9872), .Q(g34796) );
  AND2X1 U9812 ( .IN1(n9873), .IN2(n9029), .Q(n9872) );
  OR2X1 U9813 ( .IN1(n9830), .IN2(g2882), .Q(n9873) );
  OR2X1 U9814 ( .IN1(n9874), .IN2(n9875), .Q(n9830) );
  AND2X1 U9815 ( .IN1(n9157), .IN2(g2898), .Q(n9871) );
  OR2X1 U9816 ( .IN1(n9876), .IN2(n9877), .Q(g34795) );
  AND2X1 U9817 ( .IN1(n9878), .IN2(n9029), .Q(n9877) );
  OR2X1 U9818 ( .IN1(n9836), .IN2(g2898), .Q(n9878) );
  INVX0 U9819 ( .INP(n9879), .ZN(n9836) );
  AND4X1 U9820 ( .IN1(n9880), .IN2(n9881), .IN3(n9882), .IN4(n9883), .Q(n9879)
         );
  AND2X1 U9821 ( .IN1(n5861), .IN2(n5882), .Q(n9883) );
  AND2X1 U9822 ( .IN1(n9157), .IN2(g2864), .Q(n9876) );
  OR2X1 U9823 ( .IN1(n9884), .IN2(n9885), .Q(g34794) );
  AND2X1 U9824 ( .IN1(n9886), .IN2(n9029), .Q(n9885) );
  OR2X1 U9826 ( .IN1(n9837), .IN2(g2864), .Q(n9886) );
  INVX0 U9827 ( .INP(n9887), .ZN(n9837) );
  AND3X1 U9828 ( .IN1(n9888), .IN2(n9889), .IN3(n9890), .Q(n9887) );
  AND2X1 U9829 ( .IN1(n9157), .IN2(g2856), .Q(n9884) );
  OR2X1 U9830 ( .IN1(n9891), .IN2(n9892), .Q(g34793) );
  AND2X1 U9831 ( .IN1(n9893), .IN2(n9029), .Q(n9892) );
  OR2X1 U9832 ( .IN1(n9835), .IN2(g2856), .Q(n9893) );
  OR2X1 U9833 ( .IN1(n9894), .IN2(n9895), .Q(n9835) );
  AND2X1 U9834 ( .IN1(n9157), .IN2(g2848), .Q(n9891) );
  OR2X1 U9835 ( .IN1(n9896), .IN2(n9897), .Q(g34792) );
  AND2X1 U9836 ( .IN1(n9898), .IN2(n9029), .Q(n9897) );
  OR2X1 U9837 ( .IN1(n9839), .IN2(g2848), .Q(n9898) );
  INVX0 U9838 ( .INP(n9899), .ZN(n9839) );
  AND2X1 U9839 ( .IN1(n9900), .IN2(n9901), .Q(n9899) );
  AND2X1 U9840 ( .IN1(n9157), .IN2(g29214), .Q(n9896) );
  OR3X1 U9841 ( .IN1(n9902), .IN2(n9903), .IN3(n9904), .Q(g34791) );
  AND2X1 U9842 ( .IN1(n9157), .IN2(g785), .Q(n9904) );
  AND2X1 U9843 ( .IN1(n2425), .IN2(n5292), .Q(n9903) );
  AND3X1 U9844 ( .IN1(n2404), .IN2(n9905), .IN3(g790), .Q(n9902) );
  INVX0 U9845 ( .INP(n2425), .ZN(n9905) );
  OR3X1 U9846 ( .IN1(n9906), .IN2(n9907), .IN3(n9908), .Q(g34790) );
  AND2X1 U9847 ( .IN1(n9157), .IN2(g617), .Q(n9908) );
  AND2X1 U9848 ( .IN1(n2427), .IN2(n5672), .Q(n9907) );
  AND3X1 U9849 ( .IN1(n2421), .IN2(n9909), .IN3(g622), .Q(n9906) );
  INVX0 U9850 ( .INP(n2427), .ZN(n9909) );
  AND2X1 U9851 ( .IN1(n9910), .IN2(g890), .Q(g34788) );
  OR2X1 U9852 ( .IN1(n8358), .IN2(n9911), .Q(n9910) );
  INVX0 U9853 ( .INP(n3195), .ZN(n9911) );
  OR2X1 U9854 ( .IN1(n9912), .IN2(n9913), .Q(g34783) );
  AND3X1 U9855 ( .IN1(n9914), .IN2(n9915), .IN3(n9916), .Q(n9913) );
  AND3X1 U9856 ( .IN1(n9917), .IN2(n9918), .IN3(n9919), .Q(n9912) );
  OR2X1 U9857 ( .IN1(n9920), .IN2(n9921), .Q(g34735) );
  AND2X1 U9858 ( .IN1(n9922), .IN2(n9029), .Q(n9921) );
  OR2X1 U9859 ( .IN1(test_so63), .IN2(g4300), .Q(n9922) );
  AND2X1 U9860 ( .IN1(n9157), .IN2(g4297), .Q(n9920) );
  OR2X1 U9861 ( .IN1(n9923), .IN2(n9924), .Q(g34734) );
  AND2X1 U9862 ( .IN1(n9925), .IN2(n9029), .Q(n9924) );
  OR2X1 U9863 ( .IN1(g4072), .IN2(g4176), .Q(n9925) );
  AND2X1 U9864 ( .IN1(n9157), .IN2(g4172), .Q(n9923) );
  AND2X1 U9865 ( .IN1(n9926), .IN2(n9030), .Q(g34733) );
  OR2X1 U9866 ( .IN1(g4153), .IN2(g4172), .Q(n9926) );
  OR2X1 U9867 ( .IN1(n9927), .IN2(n9928), .Q(g34732) );
  AND2X1 U9868 ( .IN1(n9157), .IN2(g2999), .Q(n9928) );
  AND2X1 U9869 ( .IN1(n9039), .IN2(g2994), .Q(n9927) );
  OR2X1 U9870 ( .IN1(n9929), .IN2(n9930), .Q(g34731) );
  AND2X1 U9871 ( .IN1(n9931), .IN2(n9030), .Q(n9930) );
  OR2X1 U9872 ( .IN1(test_so64), .IN2(n9854), .Q(n9931) );
  AND2X1 U9873 ( .IN1(n9157), .IN2(g1283), .Q(n9929) );
  OR2X1 U9874 ( .IN1(n9932), .IN2(n9933), .Q(g34730) );
  AND2X1 U9875 ( .IN1(n9934), .IN2(n9030), .Q(n9933) );
  OR2X1 U9876 ( .IN1(g1283), .IN2(g1277), .Q(n9934) );
  AND2X1 U9877 ( .IN1(n9158), .IN2(g1296), .Q(n9932) );
  OR3X1 U9878 ( .IN1(n9935), .IN2(n9936), .IN3(n2499), .Q(g34729) );
  AND2X1 U9879 ( .IN1(n9158), .IN2(g1291), .Q(n9936) );
  AND2X1 U9880 ( .IN1(n5796), .IN2(n9031), .Q(n9935) );
  OR2X1 U9881 ( .IN1(n9937), .IN2(n9938), .Q(g34728) );
  AND2X1 U9882 ( .IN1(n9939), .IN2(n9031), .Q(n9938) );
  OR2X1 U9883 ( .IN1(n9855), .IN2(n9247), .Q(n9939) );
  AND2X1 U9884 ( .IN1(n9158), .IN2(g939), .Q(n9937) );
  OR2X1 U9885 ( .IN1(n9940), .IN2(n9941), .Q(g34727) );
  AND2X1 U9887 ( .IN1(n9942), .IN2(n9030), .Q(n9941) );
  OR2X1 U9888 ( .IN1(test_so52), .IN2(g939), .Q(n9942) );
  AND2X1 U9889 ( .IN1(n9158), .IN2(g952), .Q(n9940) );
  OR3X1 U9890 ( .IN1(n9943), .IN2(n9944), .IN3(n2505), .Q(g34726) );
  AND2X1 U9891 ( .IN1(n9158), .IN2(g947), .Q(n9944) );
  AND2X1 U9892 ( .IN1(n5630), .IN2(n9030), .Q(n9943) );
  OR3X1 U9893 ( .IN1(n9945), .IN2(n9946), .IN3(n9947), .Q(g34725) );
  AND2X1 U9894 ( .IN1(n9158), .IN2(g781), .Q(n9947) );
  AND2X1 U9895 ( .IN1(n2485), .IN2(n5293), .Q(n9946) );
  AND3X1 U9896 ( .IN1(n2404), .IN2(n9948), .IN3(g785), .Q(n9945) );
  INVX0 U9897 ( .INP(n2485), .ZN(n9948) );
  OR3X1 U9898 ( .IN1(n9949), .IN2(n9950), .IN3(n9951), .Q(g34724) );
  AND2X1 U9899 ( .IN1(n9158), .IN2(g613), .Q(n9951) );
  AND2X1 U9900 ( .IN1(n2487), .IN2(n5339), .Q(n9950) );
  AND3X1 U9901 ( .IN1(n2421), .IN2(n9952), .IN3(g617), .Q(n9949) );
  INVX0 U9902 ( .INP(n2487), .ZN(n9952) );
  OR2X1 U9903 ( .IN1(n9953), .IN2(n9954), .Q(g34723) );
  AND2X1 U9904 ( .IN1(n9955), .IN2(n9031), .Q(n9954) );
  OR2X1 U9905 ( .IN1(g301), .IN2(g534), .Q(n9955) );
  AND2X1 U9906 ( .IN1(test_so41), .IN2(n9138), .Q(n9953) );
  OR2X1 U9907 ( .IN1(n9956), .IN2(n9957), .Q(g34722) );
  AND2X1 U9908 ( .IN1(n9958), .IN2(n9032), .Q(n9957) );
  OR2X1 U9909 ( .IN1(n5520), .IN2(g546), .Q(n9958) );
  AND2X1 U9910 ( .IN1(n9158), .IN2(g538), .Q(n9956) );
  OR2X1 U9911 ( .IN1(n9959), .IN2(n9960), .Q(g34721) );
  AND2X1 U9912 ( .IN1(n9961), .IN2(n9031), .Q(n9960) );
  OR2X1 U9913 ( .IN1(g199), .IN2(g222), .Q(n9961) );
  AND2X1 U9914 ( .IN1(g29221), .IN2(n9138), .Q(n9959) );
  OR2X1 U9915 ( .IN1(n9962), .IN2(n9963), .Q(g34720) );
  AND2X1 U9916 ( .IN1(n9964), .IN2(n9031), .Q(n9963) );
  OR2X1 U9917 ( .IN1(n5657), .IN2(g550), .Q(n9964) );
  AND2X1 U9918 ( .IN1(n9158), .IN2(g534), .Q(n9962) );
  AND2X1 U9919 ( .IN1(n9965), .IN2(n9031), .Q(g34719) );
  OR2X1 U9920 ( .IN1(g209), .IN2(g538), .Q(n9965) );
  AND2X1 U9921 ( .IN1(n9036), .IN2(g6545), .Q(g34647) );
  AND2X1 U9922 ( .IN1(n9036), .IN2(g6199), .Q(g34646) );
  AND2X1 U9923 ( .IN1(n9036), .IN2(g5853), .Q(g34645) );
  AND2X1 U9924 ( .IN1(n9035), .IN2(g5507), .Q(g34644) );
  AND2X1 U9925 ( .IN1(n9035), .IN2(g5160), .Q(g34643) );
  OR2X1 U9926 ( .IN1(n9966), .IN2(n9967), .Q(g34642) );
  AND2X1 U9928 ( .IN1(n9158), .IN2(g4912), .Q(n9967) );
  AND2X1 U9929 ( .IN1(n9035), .IN2(g4927), .Q(n9966) );
  OR2X1 U9930 ( .IN1(n9968), .IN2(n9969), .Q(g34641) );
  AND2X1 U9931 ( .IN1(n9158), .IN2(g4907), .Q(n9969) );
  AND2X1 U9932 ( .IN1(n9035), .IN2(g4912), .Q(n9968) );
  OR2X1 U9933 ( .IN1(n9970), .IN2(n9971), .Q(g34640) );
  AND2X1 U9934 ( .IN1(n9158), .IN2(g4922), .Q(n9971) );
  AND2X1 U9935 ( .IN1(n9034), .IN2(g4907), .Q(n9970) );
  OR2X1 U9936 ( .IN1(n9972), .IN2(n9973), .Q(g34639) );
  AND2X1 U9937 ( .IN1(n9158), .IN2(g4917), .Q(n9973) );
  AND2X1 U9938 ( .IN1(n9033), .IN2(g4922), .Q(n9972) );
  AND2X1 U9939 ( .IN1(n9032), .IN2(g4917), .Q(g34638) );
  OR2X1 U9940 ( .IN1(n9974), .IN2(n9975), .Q(g34637) );
  AND2X1 U9941 ( .IN1(n9158), .IN2(g4722), .Q(n9975) );
  AND2X1 U9942 ( .IN1(n9033), .IN2(g4737), .Q(n9974) );
  OR2X1 U9943 ( .IN1(n9976), .IN2(n9977), .Q(g34636) );
  AND2X1 U9944 ( .IN1(n9158), .IN2(g4717), .Q(n9977) );
  AND2X1 U9945 ( .IN1(n9032), .IN2(g4722), .Q(n9976) );
  OR2X1 U9946 ( .IN1(n9978), .IN2(n9979), .Q(g34635) );
  AND2X1 U9947 ( .IN1(n9158), .IN2(g4732), .Q(n9979) );
  AND2X1 U9948 ( .IN1(n9035), .IN2(g4717), .Q(n9978) );
  OR2X1 U9949 ( .IN1(n9980), .IN2(n9981), .Q(g34634) );
  AND2X1 U9950 ( .IN1(n9158), .IN2(g4727), .Q(n9981) );
  AND2X1 U9951 ( .IN1(n9032), .IN2(g4732), .Q(n9980) );
  AND2X1 U9952 ( .IN1(n9040), .IN2(g4727), .Q(g34633) );
  OR2X1 U9954 ( .IN1(n9982), .IN2(n9983), .Q(g34632) );
  AND2X1 U9955 ( .IN1(test_so67), .IN2(n9139), .Q(n9983) );
  AND2X1 U9956 ( .IN1(n9032), .IN2(g4245), .Q(n9982) );
  OR2X1 U9959 ( .IN1(n9984), .IN2(n9985), .Q(g34631) );
  AND2X1 U9960 ( .IN1(n9158), .IN2(g4253), .Q(n9985) );
  AND2X1 U9961 ( .IN1(test_so67), .IN2(n9015), .Q(n9984) );
  OR2X1 U9962 ( .IN1(n9986), .IN2(n9987), .Q(g34630) );
  AND2X1 U9963 ( .IN1(n9158), .IN2(g4300), .Q(n9987) );
  AND2X1 U9964 ( .IN1(n9032), .IN2(g4253), .Q(n9986) );
  OR2X1 U9965 ( .IN1(n9988), .IN2(n9989), .Q(g34629) );
  AND2X1 U9966 ( .IN1(n9158), .IN2(g4146), .Q(n9989) );
  AND2X1 U9967 ( .IN1(n9033), .IN2(g4157), .Q(n9988) );
  OR2X1 U9969 ( .IN1(n9990), .IN2(n9991), .Q(g34628) );
  AND2X1 U9970 ( .IN1(n9158), .IN2(g4176), .Q(n9991) );
  AND2X1 U9971 ( .IN1(n9034), .IN2(g4146), .Q(n9990) );
  AND2X1 U9973 ( .IN1(n9033), .IN2(g3853), .Q(g34627) );
  AND2X1 U9974 ( .IN1(test_so45), .IN2(n9014), .Q(g34626) );
  AND2X1 U9975 ( .IN1(n9035), .IN2(g3151), .Q(g34625) );
  OR2X1 U9976 ( .IN1(n9992), .IN2(n9993), .Q(g34624) );
  AND2X1 U9977 ( .IN1(n9158), .IN2(g2994), .Q(n9993) );
  AND2X1 U9978 ( .IN1(n9034), .IN2(g2988), .Q(n9992) );
  OR2X1 U9979 ( .IN1(n9994), .IN2(n9995), .Q(g34623) );
  AND2X1 U9980 ( .IN1(test_so22), .IN2(n9140), .Q(n9995) );
  AND2X1 U9981 ( .IN1(n9033), .IN2(g2970), .Q(n9994) );
  OR2X1 U9982 ( .IN1(n9996), .IN2(n9997), .Q(g34622) );
  AND2X1 U9983 ( .IN1(n9159), .IN2(g2950), .Q(n9997) );
  AND2X1 U9984 ( .IN1(test_so22), .IN2(n9015), .Q(n9996) );
  OR2X1 U9985 ( .IN1(n9998), .IN2(n9999), .Q(g34621) );
  AND2X1 U9986 ( .IN1(n9159), .IN2(g2936), .Q(n9999) );
  AND2X1 U9987 ( .IN1(n9034), .IN2(g2950), .Q(n9998) );
  OR2X1 U9988 ( .IN1(n10000), .IN2(n10001), .Q(g34620) );
  AND2X1 U9989 ( .IN1(n9159), .IN2(g2922), .Q(n10001) );
  AND2X1 U9990 ( .IN1(n9034), .IN2(g2936), .Q(n10000) );
  OR2X1 U9991 ( .IN1(n10002), .IN2(n10003), .Q(g34619) );
  AND2X1 U9993 ( .IN1(n9159), .IN2(g2912), .Q(n10003) );
  AND2X1 U9994 ( .IN1(n9034), .IN2(g2922), .Q(n10002) );
  OR2X1 U9995 ( .IN1(n10004), .IN2(n10005), .Q(g34618) );
  AND2X1 U9996 ( .IN1(test_so1), .IN2(n9140), .Q(n10005) );
  AND2X1 U9997 ( .IN1(n9034), .IN2(g2912), .Q(n10004) );
  OR2X1 U9998 ( .IN1(n10006), .IN2(n10007), .Q(g34617) );
  AND2X1 U9999 ( .IN1(n9159), .IN2(g2984), .Q(n10007) );
  AND2X1 U10000 ( .IN1(test_so1), .IN2(n9015), .Q(n10006) );
  OR2X1 U10001 ( .IN1(n10008), .IN2(n10009), .Q(g34616) );
  AND2X1 U10002 ( .IN1(n9159), .IN2(g2988), .Q(n10009) );
  AND2X1 U10003 ( .IN1(n9036), .IN2(g2868), .Q(n10008) );
  OR2X1 U10004 ( .IN1(n10010), .IN2(n10011), .Q(g34615) );
  AND2X1 U10005 ( .IN1(n9159), .IN2(g2868), .Q(n10011) );
  AND2X1 U10006 ( .IN1(n9036), .IN2(g2873), .Q(n10010) );
  OR2X1 U10007 ( .IN1(n10012), .IN2(n10013), .Q(g34614) );
  AND2X1 U10008 ( .IN1(g37), .IN2(n9140), .Q(n10013) );
  AND2X1 U10009 ( .IN1(n9037), .IN2(g29214), .Q(n10012) );
  OR2X1 U10010 ( .IN1(n10014), .IN2(n10015), .Q(g34613) );
  AND2X1 U10011 ( .IN1(g37), .IN2(n9016), .Q(n10015) );
  AND2X1 U10012 ( .IN1(test_so95), .IN2(n9139), .Q(n10014) );
  OR2X1 U10013 ( .IN1(n10016), .IN2(n10017), .Q(g34612) );
  AND2X1 U10014 ( .IN1(n9159), .IN2(g2860), .Q(n10017) );
  AND2X1 U10015 ( .IN1(test_so95), .IN2(n9016), .Q(n10016) );
  OR2X1 U10016 ( .IN1(n10018), .IN2(n10019), .Q(g34611) );
  AND2X1 U10017 ( .IN1(n9159), .IN2(g2852), .Q(n10019) );
  AND2X1 U10018 ( .IN1(n9037), .IN2(g2860), .Q(n10018) );
  OR2X1 U10019 ( .IN1(n10020), .IN2(n10021), .Q(g34610) );
  AND2X1 U10020 ( .IN1(n9159), .IN2(g2844), .Q(n10021) );
  AND2X1 U10021 ( .IN1(n9037), .IN2(g2852), .Q(n10020) );
  OR2X1 U10022 ( .IN1(n10022), .IN2(n10023), .Q(g34609) );
  AND2X1 U10023 ( .IN1(n9159), .IN2(g2890), .Q(n10023) );
  AND2X1 U10024 ( .IN1(n9037), .IN2(g2844), .Q(n10022) );
  OR2X1 U10025 ( .IN1(n10024), .IN2(n10025), .Q(g34608) );
  AND2X1 U10026 ( .IN1(n9159), .IN2(g2697), .Q(n10025) );
  AND2X1 U10027 ( .IN1(n9037), .IN2(g2704), .Q(n10024) );
  OR2X1 U10028 ( .IN1(n10026), .IN2(n10027), .Q(g34607) );
  AND2X1 U10029 ( .IN1(n9159), .IN2(g2689), .Q(n10027) );
  AND2X1 U10030 ( .IN1(n9038), .IN2(g2697), .Q(n10026) );
  AND2X1 U10031 ( .IN1(n9038), .IN2(g2689), .Q(g34606) );
  OR2X1 U10032 ( .IN1(n10028), .IN2(n10029), .Q(g34605) );
  AND2X1 U10033 ( .IN1(n9159), .IN2(g2138), .Q(n10029) );
  AND2X1 U10034 ( .IN1(n9038), .IN2(g2145), .Q(n10028) );
  OR2X1 U10035 ( .IN1(n10030), .IN2(n10031), .Q(g34604) );
  AND2X1 U10036 ( .IN1(n9159), .IN2(g2130), .Q(n10031) );
  AND2X1 U10037 ( .IN1(n9038), .IN2(g2138), .Q(n10030) );
  AND2X1 U10038 ( .IN1(n9038), .IN2(g2130), .Q(g34603) );
  AND2X1 U10039 ( .IN1(n9038), .IN2(g1291), .Q(g34602) );
  AND2X1 U10040 ( .IN1(n9038), .IN2(g947), .Q(g34601) );
  OR3X1 U10041 ( .IN1(n10032), .IN2(n10033), .IN3(n10034), .Q(g34600) );
  AND2X1 U10042 ( .IN1(n9159), .IN2(g776), .Q(n10034) );
  AND2X1 U10043 ( .IN1(n2507), .IN2(n5551), .Q(n10033) );
  AND3X1 U10044 ( .IN1(n2404), .IN2(n10035), .IN3(g781), .Q(n10032) );
  INVX0 U10045 ( .INP(n2507), .ZN(n10035) );
  OR3X1 U10046 ( .IN1(n10036), .IN2(n10037), .IN3(n10038), .Q(g34599) );
  AND2X1 U10047 ( .IN1(n9159), .IN2(g608), .Q(n10038) );
  AND2X1 U10048 ( .IN1(n2509), .IN2(n5474), .Q(n10037) );
  AND3X1 U10049 ( .IN1(n2421), .IN2(n10039), .IN3(g613), .Q(n10036) );
  INVX0 U10050 ( .INP(n2509), .ZN(n10039) );
  OR2X1 U10051 ( .IN1(n10040), .IN2(n10041), .Q(g34598) );
  AND2X1 U10052 ( .IN1(g29221), .IN2(n9016), .Q(n10041) );
  AND2X1 U10053 ( .IN1(n9159), .IN2(g550), .Q(n10040) );
  OR3X1 U10054 ( .IN1(n10042), .IN2(n10043), .IN3(n10044), .Q(g34468) );
  AND2X1 U10055 ( .IN1(n9159), .IN2(g4854), .Q(n10044) );
  AND2X1 U10056 ( .IN1(n10045), .IN2(g4859), .Q(n10043) );
  AND2X1 U10057 ( .IN1(n10046), .IN2(n10047), .Q(n10042) );
  OR2X1 U10058 ( .IN1(n10048), .IN2(n10049), .Q(g34467) );
  AND2X1 U10059 ( .IN1(n9159), .IN2(g4849), .Q(n10049) );
  AND3X1 U10060 ( .IN1(n10050), .IN2(n10051), .IN3(n10045), .Q(n10048) );
  INVX0 U10061 ( .INP(n10047), .ZN(n10051) );
  AND3X1 U10062 ( .IN1(g4849), .IN2(g4854), .IN3(n2563), .Q(n10047) );
  OR2X1 U10063 ( .IN1(n10052), .IN2(g4854), .Q(n10050) );
  AND2X1 U10064 ( .IN1(n2563), .IN2(g4849), .Q(n10052) );
  OR2X1 U10065 ( .IN1(n10053), .IN2(n10054), .Q(g34466) );
  AND3X1 U10066 ( .IN1(n10045), .IN2(g4843), .IN3(n5283), .Q(n10054) );
  AND2X1 U10067 ( .IN1(n10055), .IN2(g4878), .Q(n10053) );
  OR2X1 U10068 ( .IN1(n9135), .IN2(n10056), .Q(n10055) );
  AND2X1 U10069 ( .IN1(n8689), .IN2(n10046), .Q(n10056) );
  OR3X1 U10070 ( .IN1(n10057), .IN2(n10058), .IN3(n10059), .Q(g34465) );
  AND2X1 U10071 ( .IN1(n9159), .IN2(g4843), .Q(n10059) );
  AND2X1 U10072 ( .IN1(n2567), .IN2(n10045), .Q(n10058) );
  AND3X1 U10073 ( .IN1(n10046), .IN2(n2563), .IN3(n8766), .Q(n10057) );
  OR3X1 U10074 ( .IN1(n10060), .IN2(n10061), .IN3(n10062), .Q(g34464) );
  AND2X1 U10075 ( .IN1(n9160), .IN2(g4664), .Q(n10062) );
  AND2X1 U10076 ( .IN1(n10063), .IN2(g4669), .Q(n10061) );
  AND2X1 U10077 ( .IN1(n10064), .IN2(n10065), .Q(n10060) );
  OR2X1 U10078 ( .IN1(n10066), .IN2(n10067), .Q(g34463) );
  AND2X1 U10079 ( .IN1(n9160), .IN2(g4659), .Q(n10067) );
  AND3X1 U10080 ( .IN1(n10068), .IN2(n10069), .IN3(n10063), .Q(n10066) );
  INVX0 U10081 ( .INP(n10065), .ZN(n10069) );
  AND3X1 U10082 ( .IN1(g4659), .IN2(g4664), .IN3(n2573), .Q(n10065) );
  OR2X1 U10083 ( .IN1(n10070), .IN2(g4664), .Q(n10068) );
  AND2X1 U10084 ( .IN1(n2573), .IN2(g4659), .Q(n10070) );
  OR2X1 U10085 ( .IN1(n10071), .IN2(n10072), .Q(g34462) );
  AND3X1 U10086 ( .IN1(n10063), .IN2(test_so19), .IN3(n5656), .Q(n10072) );
  AND2X1 U10087 ( .IN1(n10073), .IN2(g4688), .Q(n10071) );
  OR2X1 U10088 ( .IN1(n9135), .IN2(n10074), .Q(n10073) );
  AND2X1 U10089 ( .IN1(n10064), .IN2(n8854), .Q(n10074) );
  OR3X1 U10090 ( .IN1(n10075), .IN2(n10076), .IN3(n10077), .Q(g34461) );
  AND2X1 U10091 ( .IN1(test_so19), .IN2(n9137), .Q(n10077) );
  AND2X1 U10092 ( .IN1(n2577), .IN2(n10063), .Q(n10076) );
  AND3X1 U10093 ( .IN1(n10064), .IN2(n2573), .IN3(n8769), .Q(n10075) );
  OR2X1 U10094 ( .IN1(n10078), .IN2(n10079), .Q(g34460) );
  AND2X1 U10095 ( .IN1(g34025), .IN2(test_so3), .Q(n10079) );
  AND2X1 U10096 ( .IN1(n10080), .IN2(g4639), .Q(n10078) );
  OR2X1 U10097 ( .IN1(n9135), .IN2(n10081), .Q(n10080) );
  AND3X1 U10098 ( .IN1(n10082), .IN2(n8842), .IN3(n5382), .Q(n10081) );
  OR2X1 U10099 ( .IN1(n10083), .IN2(n10084), .Q(g34459) );
  AND2X1 U10100 ( .IN1(n10085), .IN2(n9016), .Q(n10084) );
  OR2X1 U10101 ( .IN1(n10086), .IN2(n10087), .Q(n10085) );
  INVX0 U10102 ( .INP(n10082), .ZN(n10087) );
  AND2X1 U10103 ( .IN1(n10088), .IN2(n10089), .Q(n10086) );
  OR2X1 U10104 ( .IN1(n10090), .IN2(g4340), .Q(n10088) );
  AND2X1 U10105 ( .IN1(n9160), .IN2(g4643), .Q(n10083) );
  OR2X1 U10106 ( .IN1(n10091), .IN2(n10092), .Q(g34458) );
  AND2X1 U10107 ( .IN1(test_so99), .IN2(n10093), .Q(n10092) );
  OR2X1 U10108 ( .IN1(n9135), .IN2(n10094), .Q(n10093) );
  AND3X1 U10109 ( .IN1(n10095), .IN2(g4639), .IN3(n5844), .Q(n10094) );
  AND2X1 U10110 ( .IN1(n10096), .IN2(g4633), .Q(n10091) );
  OR2X1 U10111 ( .IN1(n10097), .IN2(n10098), .Q(n10096) );
  AND2X1 U10112 ( .IN1(n10099), .IN2(n8843), .Q(n10097) );
  OR3X1 U10113 ( .IN1(n10100), .IN2(n10101), .IN3(n10102), .Q(g34457) );
  AND2X1 U10114 ( .IN1(test_so3), .IN2(n9139), .Q(n10102) );
  AND3X1 U10115 ( .IN1(n10095), .IN2(g4639), .IN3(n8843), .Q(n10101) );
  AND2X1 U10116 ( .IN1(test_so99), .IN2(n10098), .Q(n10100) );
  OR2X1 U10117 ( .IN1(n10103), .IN2(g34025), .Q(n10098) );
  AND2X1 U10118 ( .IN1(n10099), .IN2(n8842), .Q(n10103) );
  OR2X1 U10119 ( .IN1(n10104), .IN2(n10105), .Q(g34456) );
  AND2X1 U10120 ( .IN1(n10106), .IN2(g4616), .Q(n10105) );
  AND2X1 U10121 ( .IN1(n10107), .IN2(g4608), .Q(n10104) );
  OR2X1 U10122 ( .IN1(n9135), .IN2(n10108), .Q(n10107) );
  AND2X1 U10123 ( .IN1(n2590), .IN2(n10109), .Q(n10108) );
  OR2X1 U10124 ( .IN1(n10110), .IN2(n10111), .Q(g34455) );
  AND2X1 U10125 ( .IN1(n2595), .IN2(g4332), .Q(n10111) );
  AND2X1 U10126 ( .IN1(n10112), .IN2(g4322), .Q(n10110) );
  OR2X1 U10127 ( .IN1(n9135), .IN2(n10113), .Q(n10112) );
  AND3X1 U10128 ( .IN1(n10082), .IN2(n10114), .IN3(n2594), .Q(n10113) );
  OR2X1 U10129 ( .IN1(n10115), .IN2(n10116), .Q(g34454) );
  AND2X1 U10130 ( .IN1(n9160), .IN2(g4601), .Q(n10116) );
  AND3X1 U10131 ( .IN1(n10117), .IN2(n10118), .IN3(n10106), .Q(n10115) );
  OR2X1 U10132 ( .IN1(n2590), .IN2(g4608), .Q(n10118) );
  OR2X1 U10133 ( .IN1(n5274), .IN2(n10119), .Q(n10117) );
  INVX0 U10134 ( .INP(n2590), .ZN(n10119) );
  OR3X1 U10135 ( .IN1(n10120), .IN2(n10121), .IN3(n10122), .Q(g34453) );
  AND2X1 U10136 ( .IN1(n9160), .IN2(g4593), .Q(n10122) );
  AND3X1 U10137 ( .IN1(n2598), .IN2(n10109), .IN3(n5365), .Q(n10121) );
  AND3X1 U10138 ( .IN1(n10106), .IN2(n10123), .IN3(g4601), .Q(n10120) );
  INVX0 U10139 ( .INP(n2598), .ZN(n10123) );
  OR2X1 U10140 ( .IN1(n10124), .IN2(n10125), .Q(g34452) );
  AND2X1 U10141 ( .IN1(n9160), .IN2(g4584), .Q(n10125) );
  AND3X1 U10142 ( .IN1(n10126), .IN2(n10127), .IN3(n10106), .Q(n10124) );
  OR2X1 U10143 ( .IN1(n141), .IN2(g4593), .Q(n10127) );
  INVX0 U10144 ( .INP(n10128), .ZN(n141) );
  OR2X1 U10145 ( .IN1(n5303), .IN2(n10128), .Q(n10126) );
  OR2X1 U10146 ( .IN1(n10129), .IN2(n10130), .Q(g34451) );
  AND2X1 U10147 ( .IN1(n9160), .IN2(g4332), .Q(n10130) );
  AND3X1 U10148 ( .IN1(n10131), .IN2(n10128), .IN3(n10106), .Q(n10129) );
  AND2X1 U10149 ( .IN1(n9038), .IN2(n10109), .Q(n10106) );
  AND2X1 U10150 ( .IN1(n10082), .IN2(n10132), .Q(n10109) );
  OR2X1 U10151 ( .IN1(n10128), .IN2(n5608), .Q(n10132) );
  OR2X1 U10152 ( .IN1(n5539), .IN2(n10114), .Q(n10128) );
  OR2X1 U10153 ( .IN1(n10133), .IN2(g4584), .Q(n10131) );
  OR3X1 U10154 ( .IN1(n10134), .IN2(n10135), .IN3(n10136), .Q(g34450) );
  AND2X1 U10155 ( .IN1(n9160), .IN2(g4311), .Q(n10136) );
  AND3X1 U10156 ( .IN1(n2594), .IN2(n10082), .IN3(n5506), .Q(n10135) );
  AND3X1 U10157 ( .IN1(n2595), .IN2(n10137), .IN3(g4322), .Q(n10134) );
  INVX0 U10158 ( .INP(n2594), .ZN(n10137) );
  AND2X1 U10159 ( .IN1(n10114), .IN2(n10138), .Q(n2595) );
  INVX0 U10160 ( .INP(n10133), .ZN(n10114) );
  AND3X1 U10161 ( .IN1(g4332), .IN2(g4322), .IN3(n2607), .Q(n10133) );
  AND2X1 U10162 ( .IN1(g4358), .IN2(n10139), .Q(n2607) );
  OR3X1 U10163 ( .IN1(n10140), .IN2(n10141), .IN3(n10142), .Q(g34448) );
  AND3X1 U10164 ( .IN1(n10143), .IN2(n10144), .IN3(n10145), .Q(n10142) );
  OR2X1 U10165 ( .IN1(n10146), .IN2(n10147), .Q(n10143) );
  AND2X1 U10166 ( .IN1(n8296), .IN2(n9017), .Q(n10146) );
  AND2X1 U10167 ( .IN1(n9160), .IN2(g2827), .Q(n10141) );
  AND3X1 U10168 ( .IN1(n10148), .IN2(g2819), .IN3(n9065), .Q(n10140) );
  OR3X1 U10169 ( .IN1(n10149), .IN2(n10150), .IN3(n10151), .Q(g34447) );
  AND3X1 U10170 ( .IN1(n10152), .IN2(n10144), .IN3(n10153), .Q(n10151) );
  OR2X1 U10171 ( .IN1(n10154), .IN2(n10147), .Q(n10152) );
  AND2X1 U10172 ( .IN1(n8295), .IN2(n9016), .Q(n10154) );
  AND2X1 U10173 ( .IN1(n9160), .IN2(g2815), .Q(n10150) );
  AND3X1 U10174 ( .IN1(n10155), .IN2(g2807), .IN3(n9065), .Q(n10149) );
  OR3X1 U10175 ( .IN1(n10156), .IN2(n10157), .IN3(n10158), .Q(g34446) );
  AND3X1 U10176 ( .IN1(n10159), .IN2(n10144), .IN3(n10160), .Q(n10158) );
  INVX0 U10177 ( .INP(n10161), .ZN(n10159) );
  AND2X1 U10178 ( .IN1(n10162), .IN2(n10163), .Q(n10161) );
  OR2X1 U10179 ( .IN1(n9136), .IN2(test_so37), .Q(n10162) );
  AND2X1 U10180 ( .IN1(n9160), .IN2(g2819), .Q(n10157) );
  AND3X1 U10181 ( .IN1(n10164), .IN2(g2815), .IN3(n9065), .Q(n10156) );
  OR3X1 U10182 ( .IN1(n10165), .IN2(n10166), .IN3(n10167), .Q(g34445) );
  AND3X1 U10183 ( .IN1(n10168), .IN2(n10144), .IN3(n10169), .Q(n10167) );
  OR2X1 U10184 ( .IN1(n1795), .IN2(n6005), .Q(n10144) );
  OR2X1 U10185 ( .IN1(n10170), .IN2(n10147), .Q(n10168) );
  AND2X1 U10186 ( .IN1(n8292), .IN2(n9017), .Q(n10170) );
  AND2X1 U10187 ( .IN1(n9160), .IN2(g2807), .Q(n10166) );
  AND3X1 U10188 ( .IN1(n10171), .IN2(g2803), .IN3(n9064), .Q(n10165) );
  OR3X1 U10189 ( .IN1(n10172), .IN2(n10173), .IN3(n10174), .Q(g34444) );
  AND3X1 U10190 ( .IN1(n10175), .IN2(n10176), .IN3(n10145), .Q(n10174) );
  INVX0 U10191 ( .INP(n10148), .ZN(n10145) );
  OR2X1 U10192 ( .IN1(n10177), .IN2(n10147), .Q(n10175) );
  AND2X1 U10193 ( .IN1(n8293), .IN2(n9017), .Q(n10177) );
  AND2X1 U10194 ( .IN1(n9160), .IN2(g2795), .Q(n10173) );
  AND3X1 U10195 ( .IN1(n10148), .IN2(g2787), .IN3(n9064), .Q(n10172) );
  OR2X1 U10196 ( .IN1(n10178), .IN2(n10179), .Q(n10148) );
  OR3X1 U10197 ( .IN1(n10180), .IN2(n10181), .IN3(n10182), .Q(g34443) );
  AND3X1 U10198 ( .IN1(n10183), .IN2(n10176), .IN3(n10153), .Q(n10182) );
  OR2X1 U10199 ( .IN1(n10184), .IN2(n10147), .Q(n10183) );
  AND2X1 U10200 ( .IN1(n8291), .IN2(n9017), .Q(n10184) );
  AND2X1 U10201 ( .IN1(n9160), .IN2(g2783), .Q(n10181) );
  AND3X1 U10202 ( .IN1(n10155), .IN2(g2775), .IN3(n9064), .Q(n10180) );
  INVX0 U10203 ( .INP(n10153), .ZN(n10155) );
  AND3X1 U10204 ( .IN1(g2724), .IN2(n8676), .IN3(n10185), .Q(n10153) );
  OR3X1 U10205 ( .IN1(n10186), .IN2(n10187), .IN3(n10188), .Q(g34442) );
  AND3X1 U10206 ( .IN1(n10189), .IN2(n10176), .IN3(n10160), .Q(n10188) );
  INVX0 U10207 ( .INP(n10164), .ZN(n10160) );
  OR2X1 U10208 ( .IN1(n10190), .IN2(n10147), .Q(n10189) );
  AND2X1 U10209 ( .IN1(n8294), .IN2(n9017), .Q(n10190) );
  AND2X1 U10210 ( .IN1(n9160), .IN2(g2787), .Q(n10187) );
  AND3X1 U10211 ( .IN1(n10164), .IN2(g2783), .IN3(n9064), .Q(n10186) );
  OR2X1 U10212 ( .IN1(n10179), .IN2(n10191), .Q(n10164) );
  OR3X1 U10213 ( .IN1(n10192), .IN2(n10193), .IN3(n10194), .Q(g34441) );
  AND3X1 U10214 ( .IN1(n10195), .IN2(n10176), .IN3(n10169), .Q(n10194) );
  OR2X1 U10215 ( .IN1(n1795), .IN2(n6006), .Q(n10176) );
  OR2X1 U10216 ( .IN1(n10196), .IN2(n10147), .Q(n10195) );
  AND2X1 U10217 ( .IN1(n8297), .IN2(n9017), .Q(n10196) );
  AND2X1 U10218 ( .IN1(n9160), .IN2(g2775), .Q(n10193) );
  AND3X1 U10219 ( .IN1(n10171), .IN2(g2771), .IN3(n9063), .Q(n10192) );
  INVX0 U10220 ( .INP(n10169), .ZN(n10171) );
  AND2X1 U10221 ( .IN1(n10197), .IN2(n10185), .Q(n10169) );
  OR2X1 U10222 ( .IN1(n10198), .IN2(n10199), .Q(g34440) );
  AND2X1 U10223 ( .IN1(n10200), .IN2(n9017), .Q(n10199) );
  OR2X1 U10224 ( .IN1(n10201), .IN2(n10202), .Q(n10200) );
  AND2X1 U10225 ( .IN1(g890), .IN2(g896), .Q(n10202) );
  AND2X1 U10226 ( .IN1(n10203), .IN2(g862), .Q(n10201) );
  OR2X1 U10227 ( .IN1(n10204), .IN2(n5431), .Q(n10203) );
  AND2X1 U10228 ( .IN1(n10205), .IN2(n10206), .Q(n10204) );
  OR3X1 U10229 ( .IN1(n2644), .IN2(n10207), .IN3(g703), .Q(n10205) );
  AND2X1 U10230 ( .IN1(n9160), .IN2(g446), .Q(n10198) );
  OR3X1 U10231 ( .IN1(n10208), .IN2(n10209), .IN3(n10210), .Q(g34439) );
  AND2X1 U10232 ( .IN1(n9160), .IN2(g772), .Q(n10210) );
  AND2X1 U10233 ( .IN1(n2554), .IN2(n5330), .Q(n10209) );
  AND3X1 U10234 ( .IN1(n2404), .IN2(n10211), .IN3(g776), .Q(n10208) );
  INVX0 U10235 ( .INP(n2554), .ZN(n10211) );
  OR3X1 U10236 ( .IN1(n10212), .IN2(n10213), .IN3(n10214), .Q(g34438) );
  AND2X1 U10237 ( .IN1(n9160), .IN2(g604), .Q(n10214) );
  AND2X1 U10238 ( .IN1(n2556), .IN2(n5475), .Q(n10213) );
  AND3X1 U10239 ( .IN1(n2421), .IN2(n10215), .IN3(g608), .Q(n10212) );
  INVX0 U10240 ( .INP(n2556), .ZN(n10215) );
  AND4X1 U10241 ( .IN1(n8555), .IN2(n5711), .IN3(n5416), .IN4(n10216), .Q(
        g34435) );
  OR3X1 U10242 ( .IN1(n10217), .IN2(g4141), .IN3(g4082), .Q(n10216) );
  AND4X1 U10243 ( .IN1(test_so11), .IN2(n5350), .IN3(n10218), .IN4(g4112), .Q(
        n10217) );
  OR2X1 U10244 ( .IN1(n8806), .IN2(n9468), .Q(g34425) );
  OR2X1 U10245 ( .IN1(n10219), .IN2(n10220), .Q(n9468) );
  AND2X1 U10246 ( .IN1(n10221), .IN2(n10222), .Q(n10219) );
  OR2X1 U10247 ( .IN1(n10223), .IN2(n10224), .Q(n8806) );
  AND2X1 U10248 ( .IN1(n10225), .IN2(test_so81), .Q(n10224) );
  OR2X1 U10249 ( .IN1(n10226), .IN2(n10227), .Q(n10225) );
  AND2X1 U10250 ( .IN1(n10228), .IN2(g4358), .Q(n10227) );
  OR2X1 U10251 ( .IN1(n10229), .IN2(n10230), .Q(n10228) );
  AND2X1 U10252 ( .IN1(n10231), .IN2(n9915), .Q(n10230) );
  AND2X1 U10253 ( .IN1(n10232), .IN2(n9918), .Q(n10229) );
  AND2X1 U10254 ( .IN1(n5348), .IN2(n10233), .Q(n10226) );
  OR2X1 U10255 ( .IN1(n10234), .IN2(n10235), .Q(n10233) );
  AND2X1 U10256 ( .IN1(n10236), .IN2(n9915), .Q(n10235) );
  AND2X1 U10257 ( .IN1(n10237), .IN2(n9918), .Q(n10234) );
  AND2X1 U10258 ( .IN1(n10238), .IN2(n8822), .Q(n10223) );
  OR2X1 U10259 ( .IN1(n10239), .IN2(n10240), .Q(n10238) );
  AND2X1 U10260 ( .IN1(n10241), .IN2(g4358), .Q(n10240) );
  OR2X1 U10261 ( .IN1(n10242), .IN2(n10243), .Q(n10241) );
  AND2X1 U10262 ( .IN1(n10244), .IN2(n9915), .Q(n10243) );
  AND2X1 U10263 ( .IN1(n10245), .IN2(n9918), .Q(n10242) );
  AND2X1 U10264 ( .IN1(n5348), .IN2(n10246), .Q(n10239) );
  OR2X1 U10265 ( .IN1(n10247), .IN2(n10248), .Q(n10246) );
  AND2X1 U10266 ( .IN1(n9366), .IN2(n9915), .Q(n10248) );
  AND2X1 U10267 ( .IN1(g31860), .IN2(n9918), .Q(n10247) );
  OR3X1 U10268 ( .IN1(g34843), .IN2(n10249), .IN3(n10220), .Q(g34383) );
  AND2X1 U10269 ( .IN1(n10250), .IN2(n10251), .Q(n10249) );
  AND4X1 U10270 ( .IN1(n10252), .IN2(n10253), .IN3(n10254), .IN4(n10255), .Q(
        n10251) );
  AND4X1 U10271 ( .IN1(n985), .IN2(n998), .IN3(n997), .IN4(n987), .Q(n10250)
         );
  OR2X1 U10272 ( .IN1(n10256), .IN2(n10257), .Q(g34843) );
  OR4X1 U10273 ( .IN1(n10258), .IN2(n10259), .IN3(n10260), .IN4(n10261), .Q(
        n10257) );
  AND3X1 U10274 ( .IN1(n10262), .IN2(g2495), .IN3(n5523), .Q(n10261) );
  AND3X1 U10275 ( .IN1(n10263), .IN2(g2629), .IN3(n5524), .Q(n10260) );
  AND2X1 U10276 ( .IN1(g31862), .IN2(n10264), .Q(n10259) );
  AND3X1 U10277 ( .IN1(n5505), .IN2(g2070), .IN3(n10265), .Q(n10258) );
  OR4X1 U10278 ( .IN1(n10266), .IN2(n10267), .IN3(n10268), .IN4(n10269), .Q(
        n10256) );
  INVX0 U10279 ( .INP(n10270), .ZN(n10269) );
  INVX0 U10280 ( .INP(n10271), .ZN(n10268) );
  OR3X1 U10281 ( .IN1(n10272), .IN2(n10273), .IN3(n10274), .Q(g34269) );
  AND3X1 U10282 ( .IN1(n10275), .IN2(n10276), .IN3(n10277), .Q(n10274) );
  OR2X1 U10283 ( .IN1(n10278), .IN2(g4961), .Q(n10276) );
  AND2X1 U10284 ( .IN1(n9160), .IN2(g4961), .Q(n10273) );
  AND3X1 U10285 ( .IN1(n10279), .IN2(g4955), .IN3(n9063), .Q(n10272) );
  INVX0 U10286 ( .INP(n10275), .ZN(n10279) );
  OR2X1 U10287 ( .IN1(n10280), .IN2(n10281), .Q(n10275) );
  OR3X1 U10288 ( .IN1(n10282), .IN2(n10283), .IN3(n10284), .Q(g34268) );
  AND3X1 U10289 ( .IN1(n10285), .IN2(n10286), .IN3(n10277), .Q(n10284) );
  OR2X1 U10290 ( .IN1(n10278), .IN2(g4950), .Q(n10286) );
  AND2X1 U10291 ( .IN1(n9160), .IN2(g4950), .Q(n10283) );
  AND3X1 U10292 ( .IN1(n10287), .IN2(g4944), .IN3(n9063), .Q(n10282) );
  INVX0 U10293 ( .INP(n10285), .ZN(n10287) );
  OR2X1 U10294 ( .IN1(n10288), .IN2(n10281), .Q(n10285) );
  OR3X1 U10295 ( .IN1(n10289), .IN2(n10290), .IN3(n10291), .Q(g34267) );
  AND3X1 U10296 ( .IN1(n10292), .IN2(n10293), .IN3(n10277), .Q(n10291) );
  OR2X1 U10297 ( .IN1(n10278), .IN2(g4939), .Q(n10293) );
  AND2X1 U10298 ( .IN1(n9160), .IN2(g4939), .Q(n10290) );
  AND3X1 U10299 ( .IN1(n10294), .IN2(g4933), .IN3(n9063), .Q(n10289) );
  INVX0 U10300 ( .INP(n10292), .ZN(n10294) );
  OR2X1 U10301 ( .IN1(n10295), .IN2(n10281), .Q(n10292) );
  OR3X1 U10302 ( .IN1(n10296), .IN2(n10297), .IN3(n10298), .Q(g34266) );
  AND3X1 U10303 ( .IN1(n10299), .IN2(n10300), .IN3(n10277), .Q(n10298) );
  AND2X1 U10304 ( .IN1(n9032), .IN2(n10301), .Q(n10277) );
  OR2X1 U10305 ( .IN1(n10302), .IN2(n10278), .Q(n10301) );
  OR2X1 U10306 ( .IN1(n10278), .IN2(g4894), .Q(n10300) );
  INVX0 U10307 ( .INP(n10303), .ZN(n10278) );
  OR2X1 U10308 ( .IN1(n8618), .IN2(n10302), .Q(n10303) );
  AND2X1 U10309 ( .IN1(n9161), .IN2(g4894), .Q(n10297) );
  AND3X1 U10310 ( .IN1(n10304), .IN2(g4888), .IN3(n9062), .Q(n10296) );
  INVX0 U10311 ( .INP(n10299), .ZN(n10304) );
  OR2X1 U10312 ( .IN1(n9914), .IN2(n10281), .Q(n10299) );
  INVX0 U10313 ( .INP(n10302), .ZN(n10281) );
  OR3X1 U10315 ( .IN1(test_so46), .IN2(n10305), .IN3(g5008), .Q(n10302) );
  AND2X1 U10316 ( .IN1(n10045), .IN2(n9425), .Q(g34265) );
  AND3X1 U10317 ( .IN1(n5318), .IN2(n5443), .IN3(n5713), .Q(n9425) );
  AND2X1 U10319 ( .IN1(n9040), .IN2(n10046), .Q(n10045) );
  AND2X1 U10320 ( .IN1(n10306), .IN2(n10307), .Q(n10046) );
  OR3X1 U10321 ( .IN1(n10308), .IN2(n10309), .IN3(n10310), .Q(g34264) );
  AND3X1 U10322 ( .IN1(n10311), .IN2(n10312), .IN3(n10313), .Q(n10310) );
  OR2X1 U10323 ( .IN1(n10314), .IN2(g4771), .Q(n10312) );
  AND2X1 U10324 ( .IN1(n9161), .IN2(g4771), .Q(n10309) );
  AND3X1 U10325 ( .IN1(n10315), .IN2(g4765), .IN3(n9062), .Q(n10308) );
  INVX0 U10326 ( .INP(n10311), .ZN(n10315) );
  OR2X1 U10327 ( .IN1(n10316), .IN2(n10317), .Q(n10311) );
  OR3X1 U10328 ( .IN1(n10318), .IN2(n10319), .IN3(n10320), .Q(g34263) );
  AND3X1 U10329 ( .IN1(n10321), .IN2(n10322), .IN3(n10313), .Q(n10320) );
  OR2X1 U10330 ( .IN1(n10314), .IN2(g4760), .Q(n10322) );
  AND2X1 U10331 ( .IN1(n9161), .IN2(g4760), .Q(n10319) );
  AND3X1 U10332 ( .IN1(n10323), .IN2(g4754), .IN3(n9062), .Q(n10318) );
  INVX0 U10333 ( .INP(n10321), .ZN(n10323) );
  OR2X1 U10334 ( .IN1(n10324), .IN2(n10317), .Q(n10321) );
  OR3X1 U10335 ( .IN1(n10325), .IN2(n10326), .IN3(n10327), .Q(g34262) );
  AND3X1 U10336 ( .IN1(n10328), .IN2(n10329), .IN3(n10313), .Q(n10327) );
  OR2X1 U10337 ( .IN1(n10314), .IN2(test_so18), .Q(n10329) );
  AND2X1 U10338 ( .IN1(test_so18), .IN2(n9138), .Q(n10326) );
  AND3X1 U10339 ( .IN1(n10330), .IN2(g4743), .IN3(n9062), .Q(n10325) );
  INVX0 U10340 ( .INP(n10328), .ZN(n10330) );
  OR2X1 U10341 ( .IN1(n10331), .IN2(n10317), .Q(n10328) );
  OR3X1 U10342 ( .IN1(n10332), .IN2(n10333), .IN3(n10334), .Q(g34261) );
  AND3X1 U10343 ( .IN1(n10335), .IN2(n10336), .IN3(n10313), .Q(n10334) );
  AND2X1 U10344 ( .IN1(n9039), .IN2(n10337), .Q(n10313) );
  OR2X1 U10345 ( .IN1(n10338), .IN2(n10314), .Q(n10337) );
  OR2X1 U10346 ( .IN1(n10314), .IN2(g4704), .Q(n10336) );
  INVX0 U10347 ( .INP(n10339), .ZN(n10314) );
  OR2X1 U10348 ( .IN1(n8619), .IN2(n10338), .Q(n10339) );
  AND2X1 U10349 ( .IN1(n9161), .IN2(g4704), .Q(n10333) );
  AND3X1 U10350 ( .IN1(n10340), .IN2(g4698), .IN3(n9061), .Q(n10332) );
  INVX0 U10351 ( .INP(n10335), .ZN(n10340) );
  OR2X1 U10352 ( .IN1(n9917), .IN2(n10317), .Q(n10335) );
  INVX0 U10353 ( .INP(n10338), .ZN(n10317) );
  OR3X1 U10354 ( .IN1(n10305), .IN2(g4818), .IN3(g8132), .Q(n10338) );
  AND2X1 U10355 ( .IN1(n10063), .IN2(n9395), .Q(g34260) );
  AND3X1 U10356 ( .IN1(n5440), .IN2(n5712), .IN3(n8553), .Q(n9395) );
  AND2X1 U10357 ( .IN1(n9039), .IN2(n10064), .Q(n10063) );
  AND2X1 U10358 ( .IN1(n10341), .IN2(n10342), .Q(n10064) );
  AND2X1 U10359 ( .IN1(n10343), .IN2(g4633), .Q(g34259) );
  OR2X1 U10360 ( .IN1(n9124), .IN2(n10344), .Q(n10343) );
  AND2X1 U10361 ( .IN1(n10095), .IN2(n5727), .Q(n10344) );
  AND3X1 U10362 ( .IN1(n10082), .IN2(test_so3), .IN3(n5382), .Q(n10095) );
  OR3X1 U10363 ( .IN1(n10345), .IN2(n10346), .IN3(n10347), .Q(g34258) );
  AND2X1 U10364 ( .IN1(test_so81), .IN2(n9138), .Q(n10347) );
  AND3X1 U10365 ( .IN1(n10139), .IN2(n10082), .IN3(n5348), .Q(n10346) );
  INVX0 U10366 ( .INP(n10348), .ZN(n10139) );
  AND3X1 U10367 ( .IN1(n10138), .IN2(n10348), .IN3(g4358), .Q(n10345) );
  OR2X1 U10368 ( .IN1(n8822), .IN2(n10089), .Q(n10348) );
  OR3X1 U10369 ( .IN1(n10349), .IN2(n10350), .IN3(n10351), .Q(g34257) );
  AND2X1 U10370 ( .IN1(n9161), .IN2(g4340), .Q(n10351) );
  AND3X1 U10371 ( .IN1(n10082), .IN2(n8822), .IN3(n10352), .Q(n10350) );
  AND3X1 U10372 ( .IN1(n10138), .IN2(test_so81), .IN3(n10089), .Q(n10349) );
  INVX0 U10373 ( .INP(n10352), .ZN(n10089) );
  AND2X1 U10374 ( .IN1(g4340), .IN2(n10090), .Q(n10352) );
  AND3X1 U10375 ( .IN1(n5727), .IN2(test_so3), .IN3(test_so99), .Q(n10090) );
  OR2X1 U10376 ( .IN1(n10353), .IN2(n10354), .Q(g34256) );
  AND2X1 U10377 ( .IN1(n10355), .IN2(n9017), .Q(n10354) );
  OR3X1 U10378 ( .IN1(n10356), .IN2(n10357), .IN3(g4459), .Q(n10355) );
  AND2X1 U10379 ( .IN1(n5671), .IN2(g4473), .Q(n10357) );
  AND2X1 U10380 ( .IN1(n9161), .IN2(g4369), .Q(n10353) );
  OR4X1 U10381 ( .IN1(n10358), .IN2(g4462), .IN3(n9121), .IN4(n10356), .Q(
        g34255) );
  AND2X1 U10382 ( .IN1(test_so38), .IN2(g4473), .Q(n10358) );
  OR2X1 U10383 ( .IN1(n10359), .IN2(n10360), .Q(g34254) );
  AND2X1 U10384 ( .IN1(n10356), .IN2(n9017), .Q(n10360) );
  AND2X1 U10385 ( .IN1(n10361), .IN2(g4473), .Q(n10359) );
  OR4X1 U10386 ( .IN1(n5382), .IN2(n9122), .IN3(test_so38), .IN4(n5671), .Q(
        n10361) );
  AND2X1 U10387 ( .IN1(n10362), .IN2(n9018), .Q(g34253) );
  OR3X1 U10388 ( .IN1(n5671), .IN2(n10356), .IN3(n8838), .Q(n10362) );
  AND3X1 U10389 ( .IN1(g26960), .IN2(n10363), .IN3(n5849), .Q(n10356) );
  OR2X1 U10390 ( .IN1(n9802), .IN2(n10364), .Q(n10363) );
  AND2X1 U10391 ( .IN1(n2668), .IN2(n5846), .Q(n10364) );
  OR3X1 U10392 ( .IN1(n10365), .IN2(n10366), .IN3(n10367), .Q(g34252) );
  AND2X1 U10393 ( .IN1(n9161), .IN2(g767), .Q(n10367) );
  AND2X1 U10394 ( .IN1(n2647), .IN2(n5334), .Q(n10366) );
  AND3X1 U10395 ( .IN1(n2404), .IN2(n10368), .IN3(g772), .Q(n10365) );
  INVX0 U10396 ( .INP(n2647), .ZN(n10368) );
  OR3X1 U10397 ( .IN1(n10369), .IN2(n10370), .IN3(n10371), .Q(g34251) );
  AND2X1 U10398 ( .IN1(n9161), .IN2(g599), .Q(n10371) );
  AND2X1 U10399 ( .IN1(n2649), .IN2(n5473), .Q(n10370) );
  AND3X1 U10400 ( .IN1(n2421), .IN2(n10372), .IN3(g604), .Q(n10369) );
  INVX0 U10401 ( .INP(n2649), .ZN(n10372) );
  OR3X1 U10402 ( .IN1(n10373), .IN2(n10374), .IN3(n10375), .Q(g34250) );
  AND2X1 U10403 ( .IN1(n9161), .IN2(g298), .Q(n10375) );
  AND2X1 U10404 ( .IN1(n5724), .IN2(n2707), .Q(n10374) );
  AND3X1 U10405 ( .IN1(n8803), .IN2(n10376), .IN3(g142), .Q(n10373) );
  INVX0 U10406 ( .INP(n2707), .ZN(n10376) );
  OR3X1 U10407 ( .IN1(n10377), .IN2(n10378), .IN3(n10379), .Q(g34249) );
  AND2X1 U10408 ( .IN1(n9161), .IN2(g157), .Q(n10379) );
  AND2X1 U10409 ( .IN1(n2710), .IN2(n5843), .Q(n10378) );
  AND3X1 U10410 ( .IN1(n10380), .IN2(n10381), .IN3(g160), .Q(n10377) );
  INVX0 U10411 ( .INP(n2710), .ZN(n10381) );
  OR3X1 U10412 ( .IN1(g34781), .IN2(n10382), .IN3(n10220), .Q(g34201) );
  AND4X1 U10413 ( .IN1(n790), .IN2(n788), .IN3(n10383), .IN4(n10384), .Q(
        n10382) );
  AND4X1 U10414 ( .IN1(n1370), .IN2(n1372), .IN3(n1366), .IN4(n1368), .Q(
        n10384) );
  AND2X1 U10415 ( .IN1(n794), .IN2(n1733), .Q(n10383) );
  OR2X1 U10416 ( .IN1(n10385), .IN2(n10386), .Q(g34781) );
  OR4X1 U10417 ( .IN1(n10387), .IN2(n10388), .IN3(n10389), .IN4(n10390), .Q(
        n10386) );
  AND2X1 U10418 ( .IN1(n10391), .IN2(n10392), .Q(n10390) );
  AND3X1 U10419 ( .IN1(n3005), .IN2(g1783), .IN3(n5359), .Q(n10389) );
  AND2X1 U10420 ( .IN1(g25167), .IN2(n10393), .Q(n10388) );
  AND2X1 U10421 ( .IN1(n10394), .IN2(n10395), .Q(n10387) );
  OR4X1 U10422 ( .IN1(n10396), .IN2(n10397), .IN3(n10398), .IN4(n10399), .Q(
        n10385) );
  AND3X1 U10423 ( .IN1(test_so21), .IN2(n10400), .IN3(n5511), .Q(n10399) );
  AND3X1 U10424 ( .IN1(n10401), .IN2(g2476), .IN3(n5509), .Q(n10398) );
  AND3X1 U10425 ( .IN1(n10402), .IN2(g1917), .IN3(n5510), .Q(n10397) );
  AND3X1 U10426 ( .IN1(n10403), .IN2(g2208), .IN3(n5512), .Q(n10396) );
  OR2X1 U10427 ( .IN1(n10404), .IN2(n10405), .Q(g34041) );
  AND2X1 U10428 ( .IN1(n9161), .IN2(g5008), .Q(n10405) );
  AND3X1 U10429 ( .IN1(n10406), .IN2(n10407), .IN3(n10408), .Q(n10404) );
  OR2X1 U10430 ( .IN1(n9916), .IN2(g4983), .Q(n10407) );
  OR4X1 U10431 ( .IN1(n10409), .IN2(n10410), .IN3(n10411), .IN4(n10412), .Q(
        g34040) );
  AND3X1 U10432 ( .IN1(n9435), .IN2(n10307), .IN3(n9061), .Q(n10412) );
  AND2X1 U10433 ( .IN1(n9154), .IN2(g4975), .Q(n10411) );
  AND2X1 U10434 ( .IN1(n10408), .IN2(g4899), .Q(n10410) );
  AND2X1 U10435 ( .IN1(n10413), .IN2(n9434), .Q(n10409) );
  OR2X1 U10436 ( .IN1(n10414), .IN2(n10415), .Q(g34039) );
  AND2X1 U10437 ( .IN1(n10408), .IN2(g4966), .Q(n10415) );
  AND2X1 U10438 ( .IN1(test_so58), .IN2(n10416), .Q(n10414) );
  OR2X1 U10439 ( .IN1(n9125), .IN2(n10417), .Q(n10416) );
  AND2X1 U10440 ( .IN1(n10418), .IN2(n10419), .Q(n10417) );
  OR3X1 U10441 ( .IN1(n10420), .IN2(n10421), .IN3(n10422), .Q(g34038) );
  AND2X1 U10442 ( .IN1(n9152), .IN2(g4983), .Q(n10422) );
  AND3X1 U10443 ( .IN1(n10418), .IN2(n8837), .IN3(n10419), .Q(n10421) );
  AND3X1 U10444 ( .IN1(test_so58), .IN2(n10408), .IN3(n10406), .Q(n10420) );
  OR3X1 U10445 ( .IN1(n10423), .IN2(n10424), .IN3(n10425), .Q(g34037) );
  AND2X1 U10446 ( .IN1(n9152), .IN2(g4966), .Q(n10425) );
  AND2X1 U10447 ( .IN1(n10413), .IN2(n5360), .Q(n10424) );
  AND3X1 U10448 ( .IN1(g4966), .IN2(n10307), .IN3(n10419), .Q(n10413) );
  INVX0 U10449 ( .INP(n10406), .ZN(n10419) );
  AND2X1 U10450 ( .IN1(n10408), .IN2(g4975), .Q(n10423) );
  AND2X1 U10451 ( .IN1(n9039), .IN2(n10418), .Q(n10408) );
  AND2X1 U10452 ( .IN1(n10307), .IN2(n10426), .Q(n10418) );
  OR2X1 U10453 ( .IN1(n10406), .IN2(n5706), .Q(n10426) );
  OR2X1 U10454 ( .IN1(n5367), .IN2(n10306), .Q(n10406) );
  INVX0 U10455 ( .INP(n9916), .ZN(n10306) );
  AND2X1 U10456 ( .IN1(g4878), .IN2(n10427), .Q(n9916) );
  AND2X1 U10457 ( .IN1(n10428), .IN2(g4871), .Q(g34036) );
  AND2X1 U10458 ( .IN1(n10428), .IN2(g4864), .Q(g34035) );
  AND2X1 U10459 ( .IN1(n10428), .IN2(g4836), .Q(g34034) );
  OR2X1 U10460 ( .IN1(n9125), .IN2(n10307), .Q(n10428) );
  OR3X1 U10461 ( .IN1(n8675), .IN2(n1795), .IN3(n10221), .Q(n10307) );
  OR2X1 U10462 ( .IN1(n10429), .IN2(n10430), .Q(g34033) );
  AND2X1 U10463 ( .IN1(n9152), .IN2(g4818), .Q(n10430) );
  AND3X1 U10464 ( .IN1(n10431), .IN2(n10432), .IN3(n10433), .Q(n10429) );
  OR2X1 U10465 ( .IN1(n9919), .IN2(g4793), .Q(n10432) );
  OR4X1 U10466 ( .IN1(n10434), .IN2(n10435), .IN3(n10436), .IN4(n10437), .Q(
        g34032) );
  AND3X1 U10467 ( .IN1(n9405), .IN2(n10342), .IN3(n9060), .Q(n10437) );
  AND2X1 U10468 ( .IN1(n9152), .IN2(g4785), .Q(n10436) );
  AND2X1 U10469 ( .IN1(n10433), .IN2(g4709), .Q(n10435) );
  AND2X1 U10470 ( .IN1(n10438), .IN2(n9404), .Q(n10434) );
  OR2X1 U10471 ( .IN1(n10439), .IN2(n10440), .Q(g34031) );
  AND2X1 U10472 ( .IN1(n10433), .IN2(g4776), .Q(n10440) );
  AND2X1 U10473 ( .IN1(test_so29), .IN2(n10441), .Q(n10439) );
  OR2X1 U10474 ( .IN1(n9125), .IN2(n10442), .Q(n10441) );
  AND2X1 U10475 ( .IN1(n10443), .IN2(n10444), .Q(n10442) );
  OR3X1 U10476 ( .IN1(n10445), .IN2(n10446), .IN3(n10447), .Q(g34030) );
  AND2X1 U10477 ( .IN1(n9152), .IN2(g4793), .Q(n10447) );
  AND3X1 U10478 ( .IN1(n10443), .IN2(n8836), .IN3(n10444), .Q(n10446) );
  AND3X1 U10479 ( .IN1(test_so29), .IN2(n10433), .IN3(n10431), .Q(n10445) );
  OR3X1 U10480 ( .IN1(n10448), .IN2(n10449), .IN3(n10450), .Q(g34029) );
  AND2X1 U10481 ( .IN1(n9152), .IN2(g4776), .Q(n10450) );
  AND2X1 U10482 ( .IN1(n10438), .IN2(n5361), .Q(n10449) );
  AND3X1 U10483 ( .IN1(g4776), .IN2(n10342), .IN3(n10444), .Q(n10438) );
  INVX0 U10484 ( .INP(n10431), .ZN(n10444) );
  AND2X1 U10485 ( .IN1(n10433), .IN2(g4785), .Q(n10448) );
  AND2X1 U10486 ( .IN1(n9039), .IN2(n10443), .Q(n10433) );
  AND2X1 U10487 ( .IN1(n10342), .IN2(n10451), .Q(n10443) );
  OR2X1 U10488 ( .IN1(n10431), .IN2(n5707), .Q(n10451) );
  OR2X1 U10489 ( .IN1(n5368), .IN2(n10341), .Q(n10431) );
  INVX0 U10490 ( .INP(n9919), .ZN(n10341) );
  AND2X1 U10491 ( .IN1(g4688), .IN2(n10452), .Q(n9919) );
  AND2X1 U10492 ( .IN1(n9467), .IN2(g4674), .Q(g34027) );
  AND2X1 U10493 ( .IN1(n9467), .IN2(g4646), .Q(g34026) );
  OR2X1 U10494 ( .IN1(n9126), .IN2(n10342), .Q(n9467) );
  OR3X1 U10495 ( .IN1(n8675), .IN2(n1795), .IN3(n10222), .Q(n10342) );
  AND2X1 U10496 ( .IN1(n5727), .IN2(n10099), .Q(g34025) );
  AND2X1 U10497 ( .IN1(n10138), .IN2(n5382), .Q(n10099) );
  AND2X1 U10498 ( .IN1(n9039), .IN2(n10082), .Q(n10138) );
  OR2X1 U10499 ( .IN1(n10453), .IN2(DFF_961_n1), .Q(n10082) );
  AND2X1 U10500 ( .IN1(n10454), .IN2(n1795), .Q(n10453) );
  OR2X1 U10501 ( .IN1(n10455), .IN2(n10456), .Q(g34024) );
  AND3X1 U10502 ( .IN1(n10457), .IN2(n10458), .IN3(n9060), .Q(n10456) );
  OR2X1 U10503 ( .IN1(n10459), .IN2(n10460), .Q(n10458) );
  OR2X1 U10504 ( .IN1(n10454), .IN2(n10461), .Q(n10457) );
  AND2X1 U10505 ( .IN1(n9152), .IN2(g4492), .Q(n10455) );
  OR2X1 U10506 ( .IN1(n10462), .IN2(n10463), .Q(g34023) );
  AND2X1 U10507 ( .IN1(n10464), .IN2(n9325), .Q(n10463) );
  OR2X1 U10508 ( .IN1(n9126), .IN2(n10465), .Q(n10464) );
  AND4X1 U10509 ( .IN1(n10466), .IN2(g4555), .IN3(g4558), .IN4(g4561), .Q(
        n10465) );
  AND3X1 U10510 ( .IN1(n10460), .IN2(n9051), .IN3(n10466), .Q(n10462) );
  OR2X1 U10511 ( .IN1(n10454), .IN2(n10467), .Q(n10466) );
  INVX0 U10512 ( .INP(n9802), .ZN(n10454) );
  OR2X1 U10513 ( .IN1(n9802), .IN2(g2988), .Q(n10460) );
  OR4X1 U10514 ( .IN1(n2787), .IN2(n10468), .IN3(n10469), .IN4(n10470), .Q(
        g34022) );
  AND2X1 U10515 ( .IN1(n9152), .IN2(g2759), .Q(n10470) );
  AND3X1 U10516 ( .IN1(n10471), .IN2(g2763), .IN3(n9060), .Q(n10469) );
  INVX0 U10517 ( .INP(n10472), .ZN(n10468) );
  OR2X1 U10518 ( .IN1(n10471), .IN2(g2763), .Q(n10472) );
  OR2X1 U10519 ( .IN1(n8793), .IN2(n10473), .Q(n10471) );
  OR3X1 U10520 ( .IN1(n10474), .IN2(n10475), .IN3(n10476), .Q(g34021) );
  AND2X1 U10521 ( .IN1(n9152), .IN2(g2648), .Q(n10476) );
  AND2X1 U10522 ( .IN1(n10477), .IN2(g2567), .Q(n10475) );
  AND2X1 U10523 ( .IN1(n10478), .IN2(n10479), .Q(n10474) );
  OR2X1 U10524 ( .IN1(n10480), .IN2(n10481), .Q(g34020) );
  AND2X1 U10525 ( .IN1(n10482), .IN2(n9018), .Q(n10481) );
  OR2X1 U10526 ( .IN1(n10483), .IN2(n10484), .Q(n10482) );
  AND2X1 U10527 ( .IN1(n10485), .IN2(g2643), .Q(n10484) );
  OR2X1 U10528 ( .IN1(n10486), .IN2(n10487), .Q(n10485) );
  AND2X1 U10529 ( .IN1(n10488), .IN2(g2555), .Q(n10486) );
  AND2X1 U10530 ( .IN1(n10489), .IN2(n10490), .Q(n10483) );
  INVX0 U10531 ( .INP(n10488), .ZN(n10490) );
  OR2X1 U10532 ( .IN1(n10491), .IN2(n10478), .Q(n10489) );
  AND2X1 U10533 ( .IN1(n8348), .IN2(n10492), .Q(n10491) );
  AND2X1 U10534 ( .IN1(n10493), .IN2(g2629), .Q(n10480) );
  OR2X1 U10535 ( .IN1(n9126), .IN2(n10494), .Q(n10493) );
  AND2X1 U10536 ( .IN1(n10488), .IN2(g2643), .Q(n10494) );
  AND2X1 U10537 ( .IN1(n10495), .IN2(n10496), .Q(n10488) );
  OR2X1 U10538 ( .IN1(g1589), .IN2(n10497), .Q(n10496) );
  OR3X1 U10539 ( .IN1(n10498), .IN2(n10499), .IN3(n10500), .Q(g34019) );
  AND2X1 U10540 ( .IN1(n10501), .IN2(n10479), .Q(n10500) );
  AND2X1 U10541 ( .IN1(n9152), .IN2(g2571), .Q(n10499) );
  AND3X1 U10542 ( .IN1(n10502), .IN2(g2583), .IN3(n9059), .Q(n10498) );
  INVX0 U10543 ( .INP(n10501), .ZN(n10502) );
  AND2X1 U10544 ( .IN1(g2629), .IN2(n10503), .Q(n10501) );
  OR3X1 U10545 ( .IN1(n10504), .IN2(n10505), .IN3(n10506), .Q(g34018) );
  AND2X1 U10546 ( .IN1(n10507), .IN2(n10479), .Q(n10506) );
  INVX0 U10547 ( .INP(n10508), .ZN(n10507) );
  AND2X1 U10548 ( .IN1(n9152), .IN2(g2583), .Q(n10505) );
  AND3X1 U10549 ( .IN1(test_so61), .IN2(n10508), .IN3(n9059), .Q(n10504) );
  OR2X1 U10550 ( .IN1(n10487), .IN2(n10509), .Q(n10508) );
  OR3X1 U10551 ( .IN1(n10510), .IN2(n10511), .IN3(n10512), .Q(g34017) );
  AND2X1 U10552 ( .IN1(n10513), .IN2(n10479), .Q(n10512) );
  AND2X1 U10553 ( .IN1(test_so61), .IN2(n9139), .Q(n10511) );
  AND3X1 U10554 ( .IN1(test_so66), .IN2(n10514), .IN3(n9060), .Q(n10510) );
  INVX0 U10555 ( .INP(n10513), .ZN(n10514) );
  AND3X1 U10556 ( .IN1(g2629), .IN2(g2555), .IN3(n10492), .Q(n10513) );
  OR3X1 U10557 ( .IN1(n10515), .IN2(n10516), .IN3(n10517), .Q(g34016) );
  AND2X1 U10558 ( .IN1(n10518), .IN2(n10479), .Q(n10517) );
  AND2X1 U10559 ( .IN1(n9152), .IN2(g2563), .Q(n10516) );
  AND3X1 U10560 ( .IN1(n10519), .IN2(g2571), .IN3(n9058), .Q(n10515) );
  INVX0 U10561 ( .INP(n10518), .ZN(n10519) );
  AND3X1 U10562 ( .IN1(g2599), .IN2(n10492), .IN3(n5521), .Q(n10518) );
  OR3X1 U10563 ( .IN1(n10520), .IN2(n10521), .IN3(n10522), .Q(g34015) );
  AND2X1 U10564 ( .IN1(n10523), .IN2(n10479), .Q(n10522) );
  AND2X1 U10565 ( .IN1(n9039), .IN2(n10524), .Q(n10479) );
  INVX0 U10566 ( .INP(n10525), .ZN(n10524) );
  AND2X1 U10567 ( .IN1(n10495), .IN2(n10526), .Q(n10525) );
  OR2X1 U10568 ( .IN1(n10497), .IN2(g1585), .Q(n10526) );
  OR3X1 U10569 ( .IN1(n10527), .IN2(n10528), .IN3(n10529), .Q(n10495) );
  AND2X1 U10570 ( .IN1(n5483), .IN2(n10530), .Q(n10529) );
  INVX0 U10571 ( .INP(n10497), .ZN(n10528) );
  AND2X1 U10572 ( .IN1(n9152), .IN2(g2567), .Q(n10521) );
  AND3X1 U10573 ( .IN1(n10531), .IN2(g2563), .IN3(n9058), .Q(n10520) );
  INVX0 U10574 ( .INP(n10523), .ZN(n10531) );
  AND2X1 U10575 ( .IN1(g2555), .IN2(n10503), .Q(n10523) );
  OR3X1 U10576 ( .IN1(n10532), .IN2(n10533), .IN3(n10534), .Q(g34014) );
  AND2X1 U10577 ( .IN1(n9152), .IN2(g2514), .Q(n10534) );
  AND2X1 U10578 ( .IN1(n10535), .IN2(g2433), .Q(n10533) );
  AND2X1 U10579 ( .IN1(n10536), .IN2(n10537), .Q(n10532) );
  OR2X1 U10580 ( .IN1(n10538), .IN2(n10539), .Q(g34013) );
  AND2X1 U10581 ( .IN1(n10540), .IN2(n9018), .Q(n10539) );
  OR2X1 U10582 ( .IN1(n10541), .IN2(n10542), .Q(n10540) );
  AND2X1 U10583 ( .IN1(n10543), .IN2(g2509), .Q(n10542) );
  OR2X1 U10584 ( .IN1(n10544), .IN2(n10545), .Q(n10543) );
  AND2X1 U10585 ( .IN1(test_so79), .IN2(n10546), .Q(n10544) );
  AND2X1 U10586 ( .IN1(n10547), .IN2(n10548), .Q(n10541) );
  INVX0 U10587 ( .INP(n10546), .ZN(n10548) );
  OR2X1 U10588 ( .IN1(n10549), .IN2(n10536), .Q(n10547) );
  AND2X1 U10589 ( .IN1(n8347), .IN2(n10550), .Q(n10549) );
  AND2X1 U10590 ( .IN1(n10551), .IN2(g2495), .Q(n10538) );
  OR2X1 U10591 ( .IN1(n9126), .IN2(n10552), .Q(n10551) );
  AND2X1 U10592 ( .IN1(n10546), .IN2(g2509), .Q(n10552) );
  AND2X1 U10593 ( .IN1(n10553), .IN2(n10554), .Q(n10546) );
  OR2X1 U10594 ( .IN1(n10555), .IN2(n5755), .Q(n10554) );
  OR3X1 U10595 ( .IN1(n10556), .IN2(n10557), .IN3(n10558), .Q(g34012) );
  AND2X1 U10596 ( .IN1(n10559), .IN2(n10537), .Q(n10558) );
  AND2X1 U10597 ( .IN1(n9152), .IN2(g2437), .Q(n10557) );
  AND3X1 U10598 ( .IN1(n10560), .IN2(g2449), .IN3(n9058), .Q(n10556) );
  INVX0 U10599 ( .INP(n10559), .ZN(n10560) );
  AND2X1 U10600 ( .IN1(g2495), .IN2(n10561), .Q(n10559) );
  OR3X1 U10601 ( .IN1(n10562), .IN2(n10563), .IN3(n10564), .Q(g34011) );
  AND2X1 U10602 ( .IN1(n10565), .IN2(n10537), .Q(n10564) );
  AND2X1 U10603 ( .IN1(n9152), .IN2(g2449), .Q(n10563) );
  AND3X1 U10604 ( .IN1(n10566), .IN2(n9274), .IN3(n9060), .Q(n10562) );
  INVX0 U10605 ( .INP(n10565), .ZN(n10566) );
  AND2X1 U10606 ( .IN1(n8826), .IN2(n10567), .Q(n10565) );
  OR3X1 U10607 ( .IN1(n10568), .IN2(n10569), .IN3(n10570), .Q(g34010) );
  AND2X1 U10608 ( .IN1(n10571), .IN2(n10537), .Q(n10570) );
  AND2X1 U10609 ( .IN1(n9152), .IN2(n9274), .Q(n10569) );
  AND3X1 U10610 ( .IN1(n10572), .IN2(g2441), .IN3(n9059), .Q(n10568) );
  INVX0 U10611 ( .INP(n10571), .ZN(n10572) );
  AND3X1 U10612 ( .IN1(g2495), .IN2(n10550), .IN3(test_so79), .Q(n10571) );
  OR3X1 U10613 ( .IN1(n10573), .IN2(n10574), .IN3(n10575), .Q(g34009) );
  AND2X1 U10614 ( .IN1(n10576), .IN2(n10537), .Q(n10575) );
  AND2X1 U10615 ( .IN1(n9152), .IN2(g2429), .Q(n10574) );
  AND3X1 U10616 ( .IN1(n10577), .IN2(g2437), .IN3(n9058), .Q(n10573) );
  INVX0 U10617 ( .INP(n10576), .ZN(n10577) );
  AND2X1 U10618 ( .IN1(n5522), .IN2(n10567), .Q(n10576) );
  OR3X1 U10619 ( .IN1(n10578), .IN2(n10579), .IN3(n10580), .Q(g34008) );
  AND2X1 U10620 ( .IN1(n10581), .IN2(n10537), .Q(n10580) );
  INVX0 U10621 ( .INP(n10582), .ZN(n10537) );
  OR2X1 U10622 ( .IN1(n9127), .IN2(n10583), .Q(n10582) );
  AND2X1 U10623 ( .IN1(n10553), .IN2(n10584), .Q(n10583) );
  OR2X1 U10624 ( .IN1(n5757), .IN2(n10555), .Q(n10584) );
  OR3X1 U10625 ( .IN1(n10527), .IN2(n10585), .IN3(n10586), .Q(n10553) );
  AND2X1 U10626 ( .IN1(n5290), .IN2(n10530), .Q(n10586) );
  INVX0 U10627 ( .INP(n10555), .ZN(n10585) );
  AND2X1 U10628 ( .IN1(n9152), .IN2(g2433), .Q(n10579) );
  AND3X1 U10629 ( .IN1(n10587), .IN2(g2429), .IN3(n9059), .Q(n10578) );
  INVX0 U10630 ( .INP(n10581), .ZN(n10587) );
  AND2X1 U10631 ( .IN1(test_so79), .IN2(n10561), .Q(n10581) );
  OR3X1 U10632 ( .IN1(n10588), .IN2(n10589), .IN3(n10590), .Q(g34007) );
  AND2X1 U10633 ( .IN1(n9152), .IN2(g2380), .Q(n10590) );
  AND2X1 U10634 ( .IN1(n10591), .IN2(g2299), .Q(n10589) );
  AND2X1 U10635 ( .IN1(n10592), .IN2(n10593), .Q(n10588) );
  OR2X1 U10636 ( .IN1(n10594), .IN2(n10595), .Q(g34006) );
  AND2X1 U10637 ( .IN1(n10596), .IN2(n9018), .Q(n10595) );
  OR2X1 U10638 ( .IN1(n10597), .IN2(n10598), .Q(n10596) );
  AND2X1 U10639 ( .IN1(n10599), .IN2(g2375), .Q(n10598) );
  OR2X1 U10640 ( .IN1(n10600), .IN2(n10601), .Q(n10599) );
  AND2X1 U10641 ( .IN1(n10602), .IN2(g2287), .Q(n10600) );
  AND2X1 U10642 ( .IN1(n10603), .IN2(n10604), .Q(n10597) );
  INVX0 U10643 ( .INP(n10602), .ZN(n10604) );
  OR2X1 U10644 ( .IN1(n10605), .IN2(n10592), .Q(n10603) );
  AND2X1 U10645 ( .IN1(n8349), .IN2(n10606), .Q(n10605) );
  AND2X1 U10646 ( .IN1(n10607), .IN2(g2361), .Q(n10594) );
  OR2X1 U10647 ( .IN1(n9127), .IN2(n10608), .Q(n10607) );
  AND2X1 U10648 ( .IN1(n10602), .IN2(g2375), .Q(n10608) );
  AND2X1 U10649 ( .IN1(n10609), .IN2(n10610), .Q(n10602) );
  OR2X1 U10650 ( .IN1(n10611), .IN2(g1589), .Q(n10610) );
  OR3X1 U10651 ( .IN1(n10612), .IN2(n10613), .IN3(n10614), .Q(g34005) );
  AND2X1 U10652 ( .IN1(n10615), .IN2(n10593), .Q(n10614) );
  INVX0 U10653 ( .INP(n10616), .ZN(n10615) );
  AND2X1 U10654 ( .IN1(n9152), .IN2(g2303), .Q(n10613) );
  AND3X1 U10655 ( .IN1(n10616), .IN2(g2315), .IN3(n9060), .Q(n10612) );
  OR2X1 U10656 ( .IN1(g2331), .IN2(n10617), .Q(n10616) );
  OR3X1 U10657 ( .IN1(n10618), .IN2(n10619), .IN3(n10620), .Q(g34004) );
  AND2X1 U10658 ( .IN1(n10621), .IN2(n10593), .Q(n10620) );
  AND2X1 U10659 ( .IN1(n9152), .IN2(g2315), .Q(n10619) );
  AND3X1 U10660 ( .IN1(n10622), .IN2(n9314), .IN3(n9058), .Q(n10618) );
  INVX0 U10661 ( .INP(n10621), .ZN(n10622) );
  AND2X1 U10662 ( .IN1(n5353), .IN2(n10623), .Q(n10621) );
  OR3X1 U10663 ( .IN1(n10624), .IN2(n10625), .IN3(n10626), .Q(g34003) );
  AND2X1 U10664 ( .IN1(n10627), .IN2(n10593), .Q(n10626) );
  INVX0 U10665 ( .INP(n10628), .ZN(n10627) );
  AND2X1 U10666 ( .IN1(n9153), .IN2(n9314), .Q(n10625) );
  AND3X1 U10667 ( .IN1(n10628), .IN2(g2307), .IN3(n9058), .Q(n10624) );
  OR2X1 U10668 ( .IN1(n5353), .IN2(n10617), .Q(n10628) );
  OR2X1 U10669 ( .IN1(n10601), .IN2(n5537), .Q(n10617) );
  OR3X1 U10670 ( .IN1(n10629), .IN2(n10630), .IN3(n10631), .Q(g34002) );
  AND2X1 U10671 ( .IN1(n10632), .IN2(n10593), .Q(n10631) );
  AND2X1 U10672 ( .IN1(n9153), .IN2(g2295), .Q(n10630) );
  AND3X1 U10673 ( .IN1(n10633), .IN2(g2303), .IN3(n9059), .Q(n10629) );
  INVX0 U10674 ( .INP(n10632), .ZN(n10633) );
  AND2X1 U10675 ( .IN1(n5537), .IN2(n10623), .Q(n10632) );
  OR3X1 U10676 ( .IN1(n10634), .IN2(n10635), .IN3(n10636), .Q(g34001) );
  AND2X1 U10677 ( .IN1(n10637), .IN2(n10593), .Q(n10636) );
  AND2X1 U10678 ( .IN1(n9039), .IN2(n10638), .Q(n10593) );
  INVX0 U10679 ( .INP(n10639), .ZN(n10638) );
  AND2X1 U10680 ( .IN1(n10640), .IN2(n10609), .Q(n10639) );
  OR3X1 U10681 ( .IN1(n10527), .IN2(n10641), .IN3(n10642), .Q(n10609) );
  AND2X1 U10682 ( .IN1(n5343), .IN2(n10530), .Q(n10642) );
  INVX0 U10683 ( .INP(n10611), .ZN(n10641) );
  OR2X1 U10684 ( .IN1(g1585), .IN2(n10611), .Q(n10640) );
  AND2X1 U10685 ( .IN1(n9153), .IN2(g2299), .Q(n10635) );
  AND3X1 U10686 ( .IN1(n10643), .IN2(g2295), .IN3(n9059), .Q(n10634) );
  INVX0 U10687 ( .INP(n10637), .ZN(n10643) );
  AND3X1 U10688 ( .IN1(g2287), .IN2(n10606), .IN3(n5513), .Q(n10637) );
  OR3X1 U10689 ( .IN1(n10644), .IN2(n10645), .IN3(n10646), .Q(g34000) );
  AND2X1 U10690 ( .IN1(n9153), .IN2(g2246), .Q(n10646) );
  AND2X1 U10691 ( .IN1(n10647), .IN2(g2165), .Q(n10645) );
  AND2X1 U10692 ( .IN1(n10648), .IN2(n10649), .Q(n10644) );
  OR2X1 U10693 ( .IN1(n10650), .IN2(n10651), .Q(g33999) );
  AND2X1 U10694 ( .IN1(n10652), .IN2(n9018), .Q(n10651) );
  OR2X1 U10695 ( .IN1(n10653), .IN2(n10654), .Q(n10652) );
  AND2X1 U10696 ( .IN1(n10655), .IN2(g2241), .Q(n10654) );
  OR2X1 U10697 ( .IN1(n10656), .IN2(n10657), .Q(n10655) );
  AND2X1 U10698 ( .IN1(n10658), .IN2(g2153), .Q(n10656) );
  AND2X1 U10699 ( .IN1(n10659), .IN2(n10660), .Q(n10653) );
  INVX0 U10700 ( .INP(n10658), .ZN(n10660) );
  OR2X1 U10701 ( .IN1(n10661), .IN2(n10648), .Q(n10659) );
  AND2X1 U10702 ( .IN1(n8351), .IN2(n10662), .Q(n10661) );
  AND2X1 U10703 ( .IN1(n10663), .IN2(g2227), .Q(n10650) );
  OR2X1 U10704 ( .IN1(n9127), .IN2(n10664), .Q(n10663) );
  AND2X1 U10705 ( .IN1(n10658), .IN2(g2241), .Q(n10664) );
  AND2X1 U10706 ( .IN1(n10665), .IN2(n10666), .Q(n10658) );
  OR2X1 U10707 ( .IN1(n10667), .IN2(n5755), .Q(n10666) );
  OR3X1 U10708 ( .IN1(n10668), .IN2(n10669), .IN3(n10670), .Q(g33998) );
  AND2X1 U10709 ( .IN1(n10671), .IN2(n10649), .Q(n10670) );
  INVX0 U10710 ( .INP(n10672), .ZN(n10671) );
  AND2X1 U10711 ( .IN1(n9153), .IN2(g2169), .Q(n10669) );
  AND3X1 U10712 ( .IN1(n10672), .IN2(g2181), .IN3(n9061), .Q(n10668) );
  OR2X1 U10713 ( .IN1(g2197), .IN2(n10673), .Q(n10672) );
  OR3X1 U10714 ( .IN1(n10674), .IN2(n10675), .IN3(n10676), .Q(g33997) );
  AND2X1 U10715 ( .IN1(n10677), .IN2(n10649), .Q(n10676) );
  AND2X1 U10716 ( .IN1(n9153), .IN2(g2181), .Q(n10675) );
  AND3X1 U10717 ( .IN1(n10678), .IN2(n9352), .IN3(n9058), .Q(n10674) );
  INVX0 U10718 ( .INP(n10677), .ZN(n10678) );
  AND2X1 U10719 ( .IN1(n5356), .IN2(n10679), .Q(n10677) );
  OR3X1 U10720 ( .IN1(n10680), .IN2(n10681), .IN3(n10682), .Q(g33996) );
  AND2X1 U10721 ( .IN1(n10683), .IN2(n10649), .Q(n10682) );
  INVX0 U10722 ( .INP(n10684), .ZN(n10683) );
  AND2X1 U10723 ( .IN1(n9153), .IN2(n9352), .Q(n10681) );
  AND3X1 U10724 ( .IN1(n10684), .IN2(g2173), .IN3(n9059), .Q(n10680) );
  OR2X1 U10725 ( .IN1(n5356), .IN2(n10673), .Q(n10684) );
  OR2X1 U10726 ( .IN1(n10657), .IN2(n5538), .Q(n10673) );
  OR3X1 U10727 ( .IN1(n10685), .IN2(n10686), .IN3(n10687), .Q(g33995) );
  AND2X1 U10728 ( .IN1(n10688), .IN2(n10649), .Q(n10687) );
  AND2X1 U10729 ( .IN1(n9153), .IN2(g2161), .Q(n10686) );
  AND3X1 U10730 ( .IN1(n10689), .IN2(g2169), .IN3(n9058), .Q(n10685) );
  INVX0 U10731 ( .INP(n10688), .ZN(n10689) );
  AND2X1 U10732 ( .IN1(n5538), .IN2(n10679), .Q(n10688) );
  OR3X1 U10733 ( .IN1(n10690), .IN2(n10691), .IN3(n10692), .Q(g33994) );
  AND2X1 U10734 ( .IN1(n10693), .IN2(n10649), .Q(n10692) );
  AND2X1 U10735 ( .IN1(n9039), .IN2(n10694), .Q(n10649) );
  INVX0 U10736 ( .INP(n10695), .ZN(n10694) );
  AND2X1 U10737 ( .IN1(n10696), .IN2(n10665), .Q(n10695) );
  OR3X1 U10738 ( .IN1(n10527), .IN2(n10697), .IN3(n10698), .Q(n10665) );
  AND2X1 U10739 ( .IN1(n5289), .IN2(n10530), .Q(n10698) );
  INVX0 U10740 ( .INP(n10667), .ZN(n10697) );
  AND2X1 U10741 ( .IN1(g1291), .IN2(n10530), .Q(n10527) );
  AND2X1 U10742 ( .IN1(g4180), .IN2(n10699), .Q(n10530) );
  OR2X1 U10743 ( .IN1(n5757), .IN2(n10667), .Q(n10696) );
  AND2X1 U10744 ( .IN1(n9153), .IN2(g2165), .Q(n10691) );
  AND3X1 U10745 ( .IN1(n10700), .IN2(g2161), .IN3(n9062), .Q(n10690) );
  INVX0 U10746 ( .INP(n10693), .ZN(n10700) );
  AND3X1 U10747 ( .IN1(g2153), .IN2(n10662), .IN3(n5514), .Q(n10693) );
  OR3X1 U10748 ( .IN1(n10701), .IN2(n10702), .IN3(n10703), .Q(g33993) );
  AND2X1 U10749 ( .IN1(n9153), .IN2(g2089), .Q(n10703) );
  AND2X1 U10750 ( .IN1(n10704), .IN2(g2008), .Q(n10702) );
  AND2X1 U10751 ( .IN1(n10705), .IN2(n10706), .Q(n10701) );
  OR2X1 U10752 ( .IN1(n10707), .IN2(n10708), .Q(g33992) );
  AND2X1 U10753 ( .IN1(n10709), .IN2(n9018), .Q(n10708) );
  OR2X1 U10754 ( .IN1(n10710), .IN2(n10711), .Q(n10709) );
  AND2X1 U10755 ( .IN1(n10712), .IN2(g2084), .Q(n10711) );
  OR2X1 U10756 ( .IN1(n10713), .IN2(n10714), .Q(n10712) );
  AND2X1 U10757 ( .IN1(n10715), .IN2(g1996), .Q(n10713) );
  AND2X1 U10758 ( .IN1(n10716), .IN2(n10717), .Q(n10710) );
  INVX0 U10759 ( .INP(n10715), .ZN(n10717) );
  OR2X1 U10760 ( .IN1(n10718), .IN2(n10705), .Q(n10716) );
  AND2X1 U10761 ( .IN1(n8346), .IN2(n10719), .Q(n10718) );
  AND2X1 U10762 ( .IN1(n10720), .IN2(g2070), .Q(n10707) );
  OR2X1 U10763 ( .IN1(n9128), .IN2(n10721), .Q(n10720) );
  AND2X1 U10764 ( .IN1(n10715), .IN2(g2084), .Q(n10721) );
  AND2X1 U10765 ( .IN1(n10722), .IN2(n10723), .Q(n10715) );
  OR2X1 U10766 ( .IN1(g1246), .IN2(n10724), .Q(n10723) );
  OR3X1 U10767 ( .IN1(n10725), .IN2(n10726), .IN3(n10727), .Q(g33991) );
  AND2X1 U10768 ( .IN1(n10728), .IN2(n10706), .Q(n10727) );
  INVX0 U10769 ( .INP(n10729), .ZN(n10728) );
  AND2X1 U10770 ( .IN1(n9153), .IN2(g2012), .Q(n10726) );
  AND3X1 U10771 ( .IN1(n10729), .IN2(g2024), .IN3(n9074), .Q(n10725) );
  OR2X1 U10772 ( .IN1(g2040), .IN2(n10730), .Q(n10729) );
  OR3X1 U10773 ( .IN1(n10731), .IN2(n10732), .IN3(n10733), .Q(g33990) );
  AND2X1 U10774 ( .IN1(n10734), .IN2(n10706), .Q(n10733) );
  INVX0 U10775 ( .INP(n10735), .ZN(n10734) );
  AND2X1 U10776 ( .IN1(n9153), .IN2(g2024), .Q(n10732) );
  AND3X1 U10777 ( .IN1(n10735), .IN2(n9312), .IN3(n9074), .Q(n10731) );
  OR2X1 U10778 ( .IN1(n10714), .IN2(n10736), .Q(n10735) );
  OR3X1 U10779 ( .IN1(n10737), .IN2(n10738), .IN3(n10739), .Q(g33989) );
  AND2X1 U10780 ( .IN1(n10740), .IN2(n10706), .Q(n10739) );
  INVX0 U10781 ( .INP(n10741), .ZN(n10740) );
  AND2X1 U10782 ( .IN1(n9153), .IN2(n9312), .Q(n10738) );
  AND3X1 U10783 ( .IN1(n10741), .IN2(g2016), .IN3(n9074), .Q(n10737) );
  OR2X1 U10784 ( .IN1(n5355), .IN2(n10730), .Q(n10741) );
  OR2X1 U10785 ( .IN1(n10714), .IN2(n5535), .Q(n10730) );
  OR3X1 U10786 ( .IN1(n10742), .IN2(n10743), .IN3(n10744), .Q(g33988) );
  AND2X1 U10787 ( .IN1(n10745), .IN2(n10706), .Q(n10744) );
  AND2X1 U10788 ( .IN1(n9153), .IN2(g2004), .Q(n10743) );
  AND3X1 U10789 ( .IN1(n10746), .IN2(g2012), .IN3(n9074), .Q(n10742) );
  INVX0 U10790 ( .INP(n10745), .ZN(n10746) );
  AND3X1 U10791 ( .IN1(g2040), .IN2(n10719), .IN3(n5535), .Q(n10745) );
  OR3X1 U10792 ( .IN1(n10747), .IN2(n10748), .IN3(n10749), .Q(g33987) );
  AND2X1 U10793 ( .IN1(n10750), .IN2(n10706), .Q(n10749) );
  AND2X1 U10794 ( .IN1(n9039), .IN2(n10751), .Q(n10706) );
  INVX0 U10795 ( .INP(n10752), .ZN(n10751) );
  AND2X1 U10796 ( .IN1(n10753), .IN2(n10722), .Q(n10752) );
  OR3X1 U10797 ( .IN1(n10754), .IN2(n10755), .IN3(n10756), .Q(n10722) );
  AND2X1 U10798 ( .IN1(n5341), .IN2(n10757), .Q(n10756) );
  OR2X1 U10799 ( .IN1(n10724), .IN2(g30332), .Q(n10753) );
  AND2X1 U10800 ( .IN1(n9153), .IN2(g2008), .Q(n10748) );
  AND3X1 U10801 ( .IN1(n10758), .IN2(g2004), .IN3(n9074), .Q(n10747) );
  INVX0 U10802 ( .INP(n10750), .ZN(n10758) );
  AND3X1 U10803 ( .IN1(g1996), .IN2(n10719), .IN3(n5505), .Q(n10750) );
  OR3X1 U10804 ( .IN1(n10759), .IN2(n10760), .IN3(n10761), .Q(g33986) );
  AND2X1 U10805 ( .IN1(n9153), .IN2(g1955), .Q(n10761) );
  AND2X1 U10806 ( .IN1(n10762), .IN2(g1874), .Q(n10760) );
  AND2X1 U10807 ( .IN1(n10763), .IN2(n10764), .Q(n10759) );
  OR2X1 U10808 ( .IN1(n10765), .IN2(n10766), .Q(g33985) );
  AND2X1 U10809 ( .IN1(n10767), .IN2(n9018), .Q(n10766) );
  OR2X1 U10810 ( .IN1(n10768), .IN2(n10769), .Q(n10767) );
  AND2X1 U10811 ( .IN1(n10770), .IN2(g1950), .Q(n10769) );
  OR2X1 U10812 ( .IN1(n10771), .IN2(n10772), .Q(n10770) );
  AND2X1 U10813 ( .IN1(test_so8), .IN2(n10773), .Q(n10771) );
  AND2X1 U10814 ( .IN1(n10774), .IN2(n10775), .Q(n10768) );
  INVX0 U10815 ( .INP(n10773), .ZN(n10775) );
  OR2X1 U10816 ( .IN1(n10776), .IN2(n10763), .Q(n10774) );
  AND2X1 U10817 ( .IN1(n8350), .IN2(n10777), .Q(n10776) );
  AND2X1 U10818 ( .IN1(n10778), .IN2(g1936), .Q(n10765) );
  OR2X1 U10819 ( .IN1(n9128), .IN2(n10779), .Q(n10778) );
  AND2X1 U10820 ( .IN1(n10773), .IN2(g1950), .Q(n10779) );
  AND2X1 U10821 ( .IN1(n10780), .IN2(n10781), .Q(n10773) );
  OR2X1 U10822 ( .IN1(n10782), .IN2(n5756), .Q(n10781) );
  OR3X1 U10823 ( .IN1(n10783), .IN2(n10784), .IN3(n10785), .Q(g33984) );
  AND2X1 U10824 ( .IN1(n10786), .IN2(n10764), .Q(n10785) );
  INVX0 U10825 ( .INP(n10787), .ZN(n10786) );
  AND2X1 U10826 ( .IN1(n9153), .IN2(g1878), .Q(n10784) );
  AND3X1 U10827 ( .IN1(n10787), .IN2(g1890), .IN3(n9074), .Q(n10783) );
  OR2X1 U10828 ( .IN1(g1906), .IN2(n10788), .Q(n10787) );
  OR3X1 U10829 ( .IN1(n10789), .IN2(n10790), .IN3(n10791), .Q(g33983) );
  AND2X1 U10830 ( .IN1(n10792), .IN2(n10764), .Q(n10791) );
  AND2X1 U10831 ( .IN1(n9153), .IN2(g1890), .Q(n10790) );
  AND3X1 U10832 ( .IN1(n10793), .IN2(n9280), .IN3(n9074), .Q(n10789) );
  INVX0 U10833 ( .INP(n10792), .ZN(n10793) );
  AND2X1 U10834 ( .IN1(n8827), .IN2(n10794), .Q(n10792) );
  OR3X1 U10835 ( .IN1(n10795), .IN2(n10796), .IN3(n10797), .Q(g33982) );
  AND2X1 U10836 ( .IN1(n10798), .IN2(n10764), .Q(n10797) );
  INVX0 U10837 ( .INP(n10799), .ZN(n10798) );
  AND2X1 U10838 ( .IN1(n9153), .IN2(n9280), .Q(n10796) );
  AND3X1 U10839 ( .IN1(n10799), .IN2(g1882), .IN3(n9074), .Q(n10795) );
  OR2X1 U10840 ( .IN1(n8827), .IN2(n10788), .Q(n10799) );
  OR2X1 U10841 ( .IN1(n10772), .IN2(n5534), .Q(n10788) );
  OR3X1 U10842 ( .IN1(n10800), .IN2(n10801), .IN3(n10802), .Q(g33981) );
  AND2X1 U10843 ( .IN1(n10803), .IN2(n10764), .Q(n10802) );
  AND2X1 U10844 ( .IN1(n9153), .IN2(g1870), .Q(n10801) );
  AND3X1 U10845 ( .IN1(n10804), .IN2(g1878), .IN3(n9074), .Q(n10800) );
  INVX0 U10846 ( .INP(n10803), .ZN(n10804) );
  AND2X1 U10847 ( .IN1(n5534), .IN2(n10794), .Q(n10803) );
  OR3X1 U10848 ( .IN1(n10805), .IN2(n10806), .IN3(n10807), .Q(g33980) );
  AND2X1 U10849 ( .IN1(n10808), .IN2(n10764), .Q(n10807) );
  AND2X1 U10850 ( .IN1(n9038), .IN2(n10809), .Q(n10764) );
  INVX0 U10851 ( .INP(n10810), .ZN(n10809) );
  AND2X1 U10852 ( .IN1(n10811), .IN2(n10780), .Q(n10810) );
  OR3X1 U10853 ( .IN1(n10754), .IN2(n10812), .IN3(n10813), .Q(n10780) );
  AND2X1 U10854 ( .IN1(n5329), .IN2(n10757), .Q(n10813) );
  INVX0 U10855 ( .INP(n10782), .ZN(n10812) );
  OR2X1 U10856 ( .IN1(n5526), .IN2(n10782), .Q(n10811) );
  AND2X1 U10857 ( .IN1(n9153), .IN2(g1874), .Q(n10806) );
  AND3X1 U10858 ( .IN1(n10814), .IN2(g1870), .IN3(n9074), .Q(n10805) );
  INVX0 U10859 ( .INP(n10808), .ZN(n10814) );
  AND3X1 U10860 ( .IN1(n10777), .IN2(n5503), .IN3(test_so8), .Q(n10808) );
  OR3X1 U10861 ( .IN1(n10815), .IN2(n10816), .IN3(n10817), .Q(g33979) );
  AND2X1 U10862 ( .IN1(n9153), .IN2(g1821), .Q(n10817) );
  AND2X1 U10863 ( .IN1(n10818), .IN2(g1740), .Q(n10816) );
  AND2X1 U10864 ( .IN1(n10819), .IN2(n10820), .Q(n10815) );
  OR2X1 U10865 ( .IN1(n10821), .IN2(n10822), .Q(g33978) );
  AND2X1 U10866 ( .IN1(n10823), .IN2(n9018), .Q(n10822) );
  OR2X1 U10867 ( .IN1(n10824), .IN2(n10825), .Q(n10823) );
  AND2X1 U10868 ( .IN1(n10826), .IN2(g1816), .Q(n10825) );
  OR2X1 U10869 ( .IN1(n10827), .IN2(n10828), .Q(n10826) );
  AND2X1 U10870 ( .IN1(n10829), .IN2(g1728), .Q(n10827) );
  AND2X1 U10871 ( .IN1(n10830), .IN2(n10831), .Q(n10824) );
  INVX0 U10872 ( .INP(n10829), .ZN(n10831) );
  OR2X1 U10873 ( .IN1(n10832), .IN2(n10819), .Q(n10830) );
  AND2X1 U10874 ( .IN1(n8300), .IN2(n10833), .Q(n10832) );
  AND2X1 U10875 ( .IN1(n10834), .IN2(g1802), .Q(n10821) );
  OR2X1 U10876 ( .IN1(n9128), .IN2(n10835), .Q(n10834) );
  AND2X1 U10877 ( .IN1(n10829), .IN2(g1816), .Q(n10835) );
  AND2X1 U10878 ( .IN1(n10836), .IN2(n10837), .Q(n10829) );
  OR2X1 U10879 ( .IN1(n10838), .IN2(g1246), .Q(n10837) );
  OR3X1 U10880 ( .IN1(n10839), .IN2(n10840), .IN3(n10841), .Q(g33977) );
  AND2X1 U10881 ( .IN1(n10842), .IN2(n10820), .Q(n10841) );
  INVX0 U10882 ( .INP(n10843), .ZN(n10842) );
  AND2X1 U10883 ( .IN1(n9154), .IN2(g1744), .Q(n10840) );
  AND3X1 U10884 ( .IN1(n10843), .IN2(g1756), .IN3(n9075), .Q(n10839) );
  OR2X1 U10885 ( .IN1(g1772), .IN2(n10844), .Q(n10843) );
  OR3X1 U10886 ( .IN1(n10845), .IN2(n10846), .IN3(n10847), .Q(g33976) );
  AND2X1 U10887 ( .IN1(n10848), .IN2(n10820), .Q(n10847) );
  AND2X1 U10888 ( .IN1(n9154), .IN2(g1756), .Q(n10846) );
  AND3X1 U10889 ( .IN1(n10849), .IN2(g1752), .IN3(n9075), .Q(n10845) );
  INVX0 U10890 ( .INP(n10848), .ZN(n10849) );
  AND2X1 U10891 ( .IN1(n5352), .IN2(n10850), .Q(n10848) );
  OR3X1 U10892 ( .IN1(n10851), .IN2(n10852), .IN3(n10853), .Q(g33975) );
  AND2X1 U10893 ( .IN1(n10854), .IN2(n10820), .Q(n10853) );
  INVX0 U10894 ( .INP(n10855), .ZN(n10854) );
  AND2X1 U10895 ( .IN1(n9154), .IN2(g1752), .Q(n10852) );
  AND3X1 U10896 ( .IN1(n10855), .IN2(g1748), .IN3(n9075), .Q(n10851) );
  OR2X1 U10897 ( .IN1(n5352), .IN2(n10844), .Q(n10855) );
  OR2X1 U10898 ( .IN1(n10828), .IN2(n5536), .Q(n10844) );
  OR3X1 U10899 ( .IN1(n10856), .IN2(n10857), .IN3(n10858), .Q(g33974) );
  AND2X1 U10900 ( .IN1(n10859), .IN2(n10820), .Q(n10858) );
  AND2X1 U10901 ( .IN1(n9154), .IN2(g1736), .Q(n10857) );
  AND3X1 U10902 ( .IN1(n10860), .IN2(g1744), .IN3(n9075), .Q(n10856) );
  INVX0 U10903 ( .INP(n10859), .ZN(n10860) );
  AND2X1 U10904 ( .IN1(n5536), .IN2(n10850), .Q(n10859) );
  OR3X1 U10905 ( .IN1(n10861), .IN2(n10862), .IN3(n10863), .Q(g33973) );
  AND2X1 U10906 ( .IN1(n10864), .IN2(n10820), .Q(n10863) );
  AND2X1 U10907 ( .IN1(n9038), .IN2(n10865), .Q(n10820) );
  INVX0 U10908 ( .INP(n10866), .ZN(n10865) );
  AND2X1 U10909 ( .IN1(n10867), .IN2(n10836), .Q(n10866) );
  OR3X1 U10910 ( .IN1(n10754), .IN2(n10868), .IN3(n10869), .Q(n10836) );
  AND2X1 U10911 ( .IN1(n5478), .IN2(n10757), .Q(n10869) );
  INVX0 U10912 ( .INP(n10838), .ZN(n10868) );
  OR2X1 U10913 ( .IN1(g30332), .IN2(n10838), .Q(n10867) );
  AND2X1 U10914 ( .IN1(n9154), .IN2(g1740), .Q(n10862) );
  AND3X1 U10915 ( .IN1(n10870), .IN2(g1736), .IN3(n9075), .Q(n10861) );
  INVX0 U10916 ( .INP(n10864), .ZN(n10870) );
  AND3X1 U10917 ( .IN1(g1728), .IN2(n10833), .IN3(n5504), .Q(n10864) );
  OR3X1 U10918 ( .IN1(n10871), .IN2(n10872), .IN3(n10873), .Q(g33972) );
  AND2X1 U10919 ( .IN1(n9154), .IN2(g1687), .Q(n10873) );
  AND2X1 U10920 ( .IN1(n10874), .IN2(g1604), .Q(n10872) );
  AND2X1 U10921 ( .IN1(n10875), .IN2(n10876), .Q(n10871) );
  OR2X1 U10922 ( .IN1(n10877), .IN2(n10878), .Q(g33971) );
  AND2X1 U10923 ( .IN1(n10879), .IN2(n9019), .Q(n10878) );
  OR2X1 U10924 ( .IN1(n10880), .IN2(n10881), .Q(n10879) );
  AND2X1 U10925 ( .IN1(n10882), .IN2(g1682), .Q(n10881) );
  OR2X1 U10926 ( .IN1(n10883), .IN2(n10884), .Q(n10882) );
  AND2X1 U10927 ( .IN1(n10885), .IN2(g1592), .Q(n10883) );
  AND2X1 U10928 ( .IN1(n10886), .IN2(n10887), .Q(n10880) );
  INVX0 U10929 ( .INP(n10885), .ZN(n10887) );
  OR2X1 U10930 ( .IN1(n10888), .IN2(n10875), .Q(n10886) );
  AND2X1 U10931 ( .IN1(n8352), .IN2(n10889), .Q(n10888) );
  AND2X1 U10932 ( .IN1(n10890), .IN2(g1668), .Q(n10877) );
  OR2X1 U10933 ( .IN1(n9129), .IN2(n10891), .Q(n10890) );
  AND2X1 U10934 ( .IN1(n10885), .IN2(g1682), .Q(n10891) );
  AND2X1 U10935 ( .IN1(n10892), .IN2(n10893), .Q(n10885) );
  OR2X1 U10936 ( .IN1(n10894), .IN2(n5756), .Q(n10893) );
  OR3X1 U10937 ( .IN1(n10895), .IN2(n10896), .IN3(n10897), .Q(g33970) );
  AND2X1 U10938 ( .IN1(n10898), .IN2(n10876), .Q(n10897) );
  AND2X1 U10939 ( .IN1(n9154), .IN2(g1608), .Q(n10896) );
  AND3X1 U10940 ( .IN1(n10899), .IN2(g1620), .IN3(n9075), .Q(n10895) );
  INVX0 U10941 ( .INP(n10898), .ZN(n10899) );
  AND2X1 U10942 ( .IN1(n10889), .IN2(g31862), .Q(n10898) );
  OR3X1 U10943 ( .IN1(n10900), .IN2(n10901), .IN3(n10902), .Q(g33969) );
  AND2X1 U10944 ( .IN1(n10903), .IN2(n10876), .Q(n10902) );
  AND2X1 U10945 ( .IN1(n9154), .IN2(g1620), .Q(n10901) );
  AND3X1 U10946 ( .IN1(n10904), .IN2(n9303), .IN3(n9075), .Q(n10900) );
  INVX0 U10947 ( .INP(n10903), .ZN(n10904) );
  AND2X1 U10948 ( .IN1(n5362), .IN2(n10905), .Q(n10903) );
  OR3X1 U10949 ( .IN1(n10906), .IN2(n10907), .IN3(n10908), .Q(g33968) );
  AND2X1 U10950 ( .IN1(n10909), .IN2(n10876), .Q(n10908) );
  AND2X1 U10951 ( .IN1(n9154), .IN2(n9303), .Q(n10907) );
  AND3X1 U10952 ( .IN1(n10910), .IN2(g1612), .IN3(n9075), .Q(n10906) );
  INVX0 U10953 ( .INP(n10909), .ZN(n10910) );
  AND2X1 U10954 ( .IN1(g1668), .IN2(n10911), .Q(n10909) );
  OR3X1 U10955 ( .IN1(n10912), .IN2(n10913), .IN3(n10914), .Q(g33967) );
  AND2X1 U10956 ( .IN1(n10915), .IN2(n10876), .Q(n10914) );
  AND2X1 U10957 ( .IN1(n9154), .IN2(g1600), .Q(n10913) );
  AND3X1 U10958 ( .IN1(n10916), .IN2(g1608), .IN3(n9075), .Q(n10912) );
  INVX0 U10959 ( .INP(n10915), .ZN(n10916) );
  AND2X1 U10960 ( .IN1(n5598), .IN2(n10905), .Q(n10915) );
  OR3X1 U10961 ( .IN1(n10917), .IN2(n10918), .IN3(n10919), .Q(g33966) );
  AND2X1 U10962 ( .IN1(n10920), .IN2(n10876), .Q(n10919) );
  INVX0 U10963 ( .INP(n10921), .ZN(n10876) );
  OR2X1 U10964 ( .IN1(n9129), .IN2(n10922), .Q(n10921) );
  AND2X1 U10965 ( .IN1(n10923), .IN2(n10892), .Q(n10922) );
  OR3X1 U10966 ( .IN1(n10754), .IN2(n10924), .IN3(n10925), .Q(n10892) );
  AND2X1 U10967 ( .IN1(n5328), .IN2(n10757), .Q(n10925) );
  INVX0 U10968 ( .INP(n10894), .ZN(n10924) );
  AND2X1 U10969 ( .IN1(g947), .IN2(n10757), .Q(n10754) );
  AND2X1 U10970 ( .IN1(g4180), .IN2(n10926), .Q(n10757) );
  OR2X1 U10971 ( .IN1(n5526), .IN2(n10894), .Q(n10923) );
  AND2X1 U10972 ( .IN1(n9154), .IN2(g1604), .Q(n10918) );
  AND3X1 U10973 ( .IN1(n10927), .IN2(g1600), .IN3(n9075), .Q(n10917) );
  INVX0 U10974 ( .INP(n10920), .ZN(n10927) );
  AND2X1 U10975 ( .IN1(n5549), .IN2(n10911), .Q(n10920) );
  OR3X1 U10976 ( .IN1(n10928), .IN2(n10929), .IN3(n10930), .Q(g33965) );
  AND2X1 U10977 ( .IN1(n9154), .IN2(g763), .Q(n10930) );
  AND2X1 U10978 ( .IN1(n2704), .IN2(n5333), .Q(n10929) );
  AND3X1 U10979 ( .IN1(n2404), .IN2(n10931), .IN3(g767), .Q(n10928) );
  INVX0 U10980 ( .INP(n2704), .ZN(n10931) );
  OR3X1 U10981 ( .IN1(n10932), .IN2(n10933), .IN3(n10934), .Q(g33964) );
  AND2X1 U10982 ( .IN1(n9154), .IN2(g595), .Q(n10934) );
  AND2X1 U10983 ( .IN1(n2706), .IN2(n5550), .Q(n10933) );
  AND3X1 U10984 ( .IN1(n2421), .IN2(n10935), .IN3(g599), .Q(n10932) );
  INVX0 U10985 ( .INP(n2706), .ZN(n10935) );
  OR2X1 U10986 ( .IN1(n10936), .IN2(n10937), .Q(g33963) );
  AND3X1 U10987 ( .IN1(n10938), .IN2(n10939), .IN3(n9075), .Q(n10937) );
  OR3X1 U10988 ( .IN1(g73), .IN2(n10940), .IN3(n10941), .Q(n10939) );
  AND2X1 U10989 ( .IN1(g72), .IN2(g262), .Q(n10941) );
  AND2X1 U10990 ( .IN1(n10942), .IN2(g269), .Q(n10940) );
  OR2X1 U10991 ( .IN1(n10943), .IN2(n9824), .Q(n10938) );
  AND2X1 U10992 ( .IN1(n10942), .IN2(g255), .Q(n10943) );
  AND2X1 U10993 ( .IN1(n9154), .IN2(g29215), .Q(n10936) );
  OR2X1 U10994 ( .IN1(n10944), .IN2(n10945), .Q(g33962) );
  AND3X1 U10995 ( .IN1(n10946), .IN2(n10947), .IN3(n9075), .Q(n10945) );
  OR2X1 U10996 ( .IN1(n10948), .IN2(n9824), .Q(n10947) );
  INVX0 U10997 ( .INP(g73), .ZN(n9824) );
  AND2X1 U10998 ( .IN1(n10949), .IN2(n10950), .Q(n10948) );
  OR2X1 U10999 ( .IN1(g72), .IN2(g232), .Q(n10950) );
  OR2X1 U11000 ( .IN1(n10942), .IN2(g225), .Q(n10949) );
  OR3X1 U11001 ( .IN1(g73), .IN2(n10951), .IN3(n10952), .Q(n10946) );
  AND2X1 U11002 ( .IN1(g72), .IN2(g239), .Q(n10952) );
  AND2X1 U11003 ( .IN1(n10942), .IN2(g246), .Q(n10951) );
  AND2X1 U11004 ( .IN1(n9154), .IN2(g479), .Q(n10944) );
  OR3X1 U11005 ( .IN1(n10953), .IN2(n10954), .IN3(n10955), .Q(g33961) );
  AND2X1 U11006 ( .IN1(n9154), .IN2(g294), .Q(n10955) );
  AND2X1 U11007 ( .IN1(n2989), .IN2(n5675), .Q(n10954) );
  AND3X1 U11008 ( .IN1(n8803), .IN2(n10956), .IN3(g298), .Q(n10953) );
  INVX0 U11009 ( .INP(n2989), .ZN(n10956) );
  OR3X1 U11010 ( .IN1(n10957), .IN2(n10958), .IN3(n10959), .Q(g33960) );
  AND2X1 U11011 ( .IN1(n9154), .IN2(g153), .Q(n10959) );
  AND2X1 U11012 ( .IN1(n2991), .IN2(n5678), .Q(n10958) );
  AND3X1 U11013 ( .IN1(n10380), .IN2(n10960), .IN3(g157), .Q(n10957) );
  INVX0 U11014 ( .INP(n2991), .ZN(n10960) );
  OR4X1 U11015 ( .IN1(g34649), .IN2(n10305), .IN3(n8684), .IN4(n8683), .Q(
        g33935) );
  OR4X1 U11016 ( .IN1(n10961), .IN2(n10962), .IN3(n10963), .IN4(n10964), .Q(
        g34649) );
  AND2X1 U11017 ( .IN1(n9437), .IN2(g4955), .Q(n10964) );
  AND2X1 U11018 ( .IN1(n9434), .IN2(g4933), .Q(n10962) );
  AND2X1 U11019 ( .IN1(n9435), .IN2(g4944), .Q(n10961) );
  OR3X1 U11020 ( .IN1(n5846), .IN2(n10305), .IN3(g18881), .Q(g33874) );
  OR4X1 U11021 ( .IN1(n10220), .IN2(n9339), .IN3(n10965), .IN4(n10966), .Q(
        g33659) );
  INVX0 U11022 ( .INP(n9337), .ZN(n10966) );
  OR2X1 U11023 ( .IN1(n10967), .IN2(n10968), .Q(n9337) );
  AND2X1 U11024 ( .IN1(n5715), .IN2(n9476), .Q(n10968) );
  AND2X1 U11025 ( .IN1(g72), .IN2(g4108), .Q(n10967) );
  INVX0 U11026 ( .INP(n9338), .ZN(n10965) );
  OR2X1 U11027 ( .IN1(n10969), .IN2(n10970), .Q(n9338) );
  AND2X1 U11028 ( .IN1(g73), .IN2(g4104), .Q(n10970) );
  AND2X1 U11029 ( .IN1(n8693), .IN2(n9473), .Q(n10969) );
  OR2X1 U11030 ( .IN1(n10971), .IN2(n10972), .Q(n9339) );
  AND2X1 U11031 ( .IN1(n10973), .IN2(g4098), .Q(n10972) );
  OR3X1 U11032 ( .IN1(n10974), .IN2(n10975), .IN3(n10976), .Q(n10973) );
  AND2X1 U11033 ( .IN1(n10977), .IN2(n10978), .Q(n10976) );
  AND2X1 U11034 ( .IN1(n10979), .IN2(n10218), .Q(n10975) );
  AND3X1 U11035 ( .IN1(n10980), .IN2(n10981), .IN3(g4093), .Q(n10974) );
  OR2X1 U11036 ( .IN1(n10982), .IN2(g4087), .Q(n10981) );
  OR2X1 U11037 ( .IN1(n5480), .IN2(n9376), .Q(n10980) );
  AND2X1 U11038 ( .IN1(n5350), .IN2(n10983), .Q(n10971) );
  OR3X1 U11039 ( .IN1(n10984), .IN2(n10985), .IN3(n10986), .Q(n10983) );
  AND2X1 U11040 ( .IN1(n10987), .IN2(n10978), .Q(n10986) );
  AND2X1 U11041 ( .IN1(g32975), .IN2(n10218), .Q(n10985) );
  AND3X1 U11042 ( .IN1(n10988), .IN2(n10989), .IN3(g4093), .Q(n10984) );
  OR2X1 U11043 ( .IN1(n10990), .IN2(g4087), .Q(n10989) );
  OR2X1 U11044 ( .IN1(n5480), .IN2(n10991), .Q(n10988) );
  OR2X1 U11045 ( .IN1(n10305), .IN2(n10992), .Q(n10220) );
  OR4X1 U11046 ( .IN1(g34657), .IN2(n10305), .IN3(n8682), .IN4(n8681), .Q(
        g33636) );
  INVX0 U11047 ( .INP(n2668), .ZN(n10305) );
  OR2X1 U11048 ( .IN1(n10993), .IN2(g134), .Q(n2668) );
  AND2X1 U11049 ( .IN1(g99), .IN2(g37), .Q(n10993) );
  OR4X1 U11050 ( .IN1(n10994), .IN2(n10995), .IN3(n10996), .IN4(n10997), .Q(
        g34657) );
  AND2X1 U11051 ( .IN1(n9407), .IN2(g4765), .Q(n10997) );
  AND2X1 U11052 ( .IN1(n9404), .IN2(g4743), .Q(n10995) );
  AND2X1 U11053 ( .IN1(n9405), .IN2(g4754), .Q(n10994) );
  OR2X1 U11054 ( .IN1(n10998), .IN2(n10999), .Q(g33627) );
  AND2X1 U11055 ( .IN1(n9154), .IN2(g6741), .Q(n10999) );
  AND2X1 U11056 ( .IN1(n11000), .IN2(n11001), .Q(n10998) );
  OR2X1 U11057 ( .IN1(n11002), .IN2(n11003), .Q(n11000) );
  AND2X1 U11058 ( .IN1(n9365), .IN2(n11004), .Q(n11003) );
  AND2X1 U11059 ( .IN1(n11005), .IN2(n9019), .Q(n11002) );
  OR2X1 U11060 ( .IN1(n11006), .IN2(n9369), .Q(n11005) );
  AND2X1 U11061 ( .IN1(n8809), .IN2(g6682), .Q(n11006) );
  OR3X1 U11062 ( .IN1(n11007), .IN2(n11008), .IN3(n11009), .Q(g33626) );
  AND2X1 U11063 ( .IN1(n11010), .IN2(g6741), .Q(n11009) );
  AND2X1 U11064 ( .IN1(n9154), .IN2(g6736), .Q(n11008) );
  AND4X1 U11065 ( .IN1(n11001), .IN2(n11004), .IN3(n5398), .IN4(n9050), .Q(
        n11007) );
  OR4X1 U11066 ( .IN1(n10221), .IN2(n11011), .IN3(test_so81), .IN4(n8809), .Q(
        n11001) );
  OR2X1 U11067 ( .IN1(n11012), .IN2(n11013), .Q(g33625) );
  AND2X1 U11068 ( .IN1(n9154), .IN2(g6395), .Q(n11013) );
  AND2X1 U11069 ( .IN1(n11014), .IN2(n11015), .Q(n11012) );
  OR2X1 U11070 ( .IN1(n11016), .IN2(n11017), .Q(n11014) );
  AND2X1 U11071 ( .IN1(n11018), .IN2(n11019), .Q(n11017) );
  AND2X1 U11072 ( .IN1(n11020), .IN2(n9019), .Q(n11016) );
  OR2X1 U11073 ( .IN1(n11021), .IN2(n11022), .Q(n11020) );
  AND2X1 U11074 ( .IN1(n11023), .IN2(g6336), .Q(n11021) );
  OR3X1 U11075 ( .IN1(n11024), .IN2(n11025), .IN3(n11026), .Q(g33624) );
  AND2X1 U11076 ( .IN1(n11027), .IN2(g6395), .Q(n11026) );
  AND2X1 U11077 ( .IN1(n9154), .IN2(g6390), .Q(n11025) );
  AND4X1 U11078 ( .IN1(n11019), .IN2(n11015), .IN3(n5396), .IN4(n9050), .Q(
        n11024) );
  OR4X1 U11079 ( .IN1(n11023), .IN2(n11028), .IN3(n10222), .IN4(n8822), .Q(
        n11015) );
  OR2X1 U11080 ( .IN1(n11029), .IN2(n11030), .Q(g33623) );
  AND2X1 U11081 ( .IN1(test_so57), .IN2(n9139), .Q(n11030) );
  AND2X1 U11082 ( .IN1(n11031), .IN2(n11032), .Q(n11029) );
  OR2X1 U11083 ( .IN1(n11033), .IN2(n11034), .Q(n11031) );
  AND2X1 U11084 ( .IN1(n11035), .IN2(n11036), .Q(n11034) );
  AND2X1 U11085 ( .IN1(n11037), .IN2(n9019), .Q(n11033) );
  OR2X1 U11086 ( .IN1(n11038), .IN2(n11039), .Q(n11037) );
  AND2X1 U11087 ( .IN1(n11040), .IN2(g5990), .Q(n11038) );
  OR3X1 U11088 ( .IN1(n11041), .IN2(n11042), .IN3(n11043), .Q(g33622) );
  AND2X1 U11089 ( .IN1(n11044), .IN2(test_so57), .Q(n11043) );
  AND2X1 U11090 ( .IN1(test_so50), .IN2(n9140), .Q(n11042) );
  AND4X1 U11091 ( .IN1(n11032), .IN2(n8835), .IN3(n11036), .IN4(n9049), .Q(
        n11041) );
  OR4X1 U11092 ( .IN1(n11028), .IN2(n11040), .IN3(test_so81), .IN4(n10222), 
        .Q(n11032) );
  OR2X1 U11093 ( .IN1(n11045), .IN2(n11046), .Q(g33621) );
  AND2X1 U11094 ( .IN1(n9155), .IN2(g5703), .Q(n11046) );
  AND2X1 U11095 ( .IN1(n11047), .IN2(n11048), .Q(n11045) );
  OR2X1 U11096 ( .IN1(n11049), .IN2(n11050), .Q(n11047) );
  AND2X1 U11097 ( .IN1(n11051), .IN2(n11052), .Q(n11050) );
  AND2X1 U11098 ( .IN1(n11053), .IN2(n9019), .Q(n11049) );
  OR2X1 U11099 ( .IN1(n11054), .IN2(n11055), .Q(n11053) );
  AND2X1 U11100 ( .IN1(n11056), .IN2(g5644), .Q(n11054) );
  OR3X1 U11101 ( .IN1(n11057), .IN2(n11058), .IN3(n11059), .Q(g33620) );
  AND2X1 U11102 ( .IN1(n11060), .IN2(g5703), .Q(n11059) );
  AND2X1 U11103 ( .IN1(n9155), .IN2(g5698), .Q(n11058) );
  AND4X1 U11104 ( .IN1(n11052), .IN2(n11048), .IN3(n5397), .IN4(n9049), .Q(
        n11057) );
  OR4X1 U11105 ( .IN1(n11011), .IN2(n11056), .IN3(n10222), .IN4(n8822), .Q(
        n11048) );
  OR2X1 U11106 ( .IN1(n11061), .IN2(n11062), .Q(g33619) );
  AND2X1 U11107 ( .IN1(n9155), .IN2(g5357), .Q(n11062) );
  AND2X1 U11108 ( .IN1(n11063), .IN2(n11064), .Q(n11061) );
  OR2X1 U11109 ( .IN1(n11065), .IN2(n11066), .Q(n11063) );
  AND2X1 U11110 ( .IN1(n9360), .IN2(g33959), .Q(n11066) );
  AND2X1 U11111 ( .IN1(n11067), .IN2(n9019), .Q(n11065) );
  OR2X1 U11112 ( .IN1(n11068), .IN2(n9359), .Q(n11067) );
  AND2X1 U11113 ( .IN1(n8804), .IN2(g5297), .Q(n11068) );
  OR3X1 U11114 ( .IN1(n11069), .IN2(n11070), .IN3(n11071), .Q(g33618) );
  AND2X1 U11115 ( .IN1(n11072), .IN2(g5357), .Q(n11071) );
  AND2X1 U11116 ( .IN1(n9155), .IN2(g5352), .Q(n11070) );
  AND4X1 U11117 ( .IN1(n11064), .IN2(g33959), .IN3(n5393), .IN4(n9049), .Q(
        n11069) );
  OR4X1 U11118 ( .IN1(n10222), .IN2(n11011), .IN3(test_so81), .IN4(n8804), .Q(
        n11064) );
  INVX0 U11119 ( .INP(n9918), .ZN(n10222) );
  AND3X1 U11120 ( .IN1(n9826), .IN2(n11073), .IN3(n5323), .Q(n9918) );
  OR2X1 U11121 ( .IN1(n11074), .IN2(n11075), .Q(g33617) );
  AND2X1 U11122 ( .IN1(n10467), .IN2(n9019), .Q(n11075) );
  OR2X1 U11123 ( .IN1(n11076), .IN2(n11077), .Q(n10467) );
  AND2X1 U11124 ( .IN1(n11078), .IN2(g4581), .Q(n11077) );
  OR2X1 U11125 ( .IN1(n9802), .IN2(g4575), .Q(n11078) );
  AND2X1 U11126 ( .IN1(n5670), .IN2(g4552), .Q(n11076) );
  AND2X1 U11127 ( .IN1(n9155), .IN2(g4552), .Q(n11074) );
  OR2X1 U11128 ( .IN1(n11079), .IN2(n11080), .Q(g33616) );
  AND2X1 U11129 ( .IN1(n10461), .IN2(n9019), .Q(n11080) );
  OR2X1 U11130 ( .IN1(n11081), .IN2(n11082), .Q(n10461) );
  AND2X1 U11131 ( .IN1(n11083), .IN2(g4581), .Q(n11082) );
  OR2X1 U11132 ( .IN1(test_so100), .IN2(n9802), .Q(n11083) );
  AND2X1 U11133 ( .IN1(n5670), .IN2(g4512), .Q(n11081) );
  AND2X1 U11134 ( .IN1(n9155), .IN2(g4515), .Q(n11079) );
  OR2X1 U11135 ( .IN1(n11084), .IN2(n11085), .Q(g33614) );
  AND2X1 U11136 ( .IN1(n9155), .IN2(g4054), .Q(n11085) );
  AND2X1 U11137 ( .IN1(n11086), .IN2(n11087), .Q(n11084) );
  OR2X1 U11138 ( .IN1(n11088), .IN2(n11089), .Q(n11086) );
  AND2X1 U11139 ( .IN1(n11090), .IN2(n11091), .Q(n11089) );
  AND2X1 U11140 ( .IN1(n11092), .IN2(n9019), .Q(n11088) );
  OR2X1 U11141 ( .IN1(n11093), .IN2(n11094), .Q(n11092) );
  AND2X1 U11142 ( .IN1(n11095), .IN2(g3990), .Q(n11093) );
  OR3X1 U11143 ( .IN1(n11096), .IN2(n11097), .IN3(n11098), .Q(g33613) );
  AND2X1 U11144 ( .IN1(n11099), .IN2(g4054), .Q(n11098) );
  AND2X1 U11145 ( .IN1(n9155), .IN2(g4049), .Q(n11097) );
  AND4X1 U11146 ( .IN1(n11091), .IN2(n11087), .IN3(n5395), .IN4(n9049), .Q(
        n11096) );
  OR4X1 U11147 ( .IN1(n11028), .IN2(n11095), .IN3(n10221), .IN4(n8822), .Q(
        n11087) );
  OR2X1 U11148 ( .IN1(n11100), .IN2(n11101), .Q(g33612) );
  AND2X1 U11149 ( .IN1(n9151), .IN2(g3703), .Q(n11101) );
  AND2X1 U11150 ( .IN1(n11102), .IN2(n11103), .Q(n11100) );
  OR2X1 U11151 ( .IN1(n11104), .IN2(n11105), .Q(n11102) );
  AND2X1 U11152 ( .IN1(n11106), .IN2(n11107), .Q(n11105) );
  AND2X1 U11153 ( .IN1(n11108), .IN2(n9019), .Q(n11104) );
  OR2X1 U11154 ( .IN1(n11109), .IN2(n11110), .Q(n11108) );
  AND2X1 U11155 ( .IN1(n11111), .IN2(g3639), .Q(n11109) );
  OR3X1 U11156 ( .IN1(n11112), .IN2(n11113), .IN3(n11114), .Q(g33611) );
  AND2X1 U11157 ( .IN1(n11115), .IN2(g3703), .Q(n11114) );
  AND2X1 U11158 ( .IN1(n9155), .IN2(g3698), .Q(n11113) );
  AND4X1 U11159 ( .IN1(n11107), .IN2(n11103), .IN3(n5399), .IN4(n9049), .Q(
        n11112) );
  OR4X1 U11160 ( .IN1(n11111), .IN2(n11028), .IN3(test_so81), .IN4(n10221), 
        .Q(n11103) );
  INVX0 U11161 ( .INP(n3033), .ZN(n11028) );
  OR2X1 U11162 ( .IN1(n11116), .IN2(n11117), .Q(g33610) );
  AND3X1 U11163 ( .IN1(n11118), .IN2(n11119), .IN3(n9076), .Q(n11117) );
  OR3X1 U11164 ( .IN1(n11120), .IN2(n11121), .IN3(n11122), .Q(n11118) );
  AND2X1 U11165 ( .IN1(n11123), .IN2(g3288), .Q(n11121) );
  AND2X1 U11166 ( .IN1(n11124), .IN2(n11125), .Q(n11120) );
  AND2X1 U11167 ( .IN1(n9155), .IN2(g3352), .Q(n11116) );
  OR3X1 U11168 ( .IN1(n11126), .IN2(n11127), .IN3(n11128), .Q(g33609) );
  AND2X1 U11169 ( .IN1(n11129), .IN2(g3352), .Q(n11128) );
  AND2X1 U11170 ( .IN1(n9155), .IN2(g3347), .Q(n11127) );
  AND4X1 U11171 ( .IN1(n11125), .IN2(n11119), .IN3(n5604), .IN4(n9049), .Q(
        n11126) );
  OR4X1 U11172 ( .IN1(n11011), .IN2(n11123), .IN3(n10221), .IN4(n8822), .Q(
        n11119) );
  INVX0 U11173 ( .INP(n9915), .ZN(n10221) );
  AND3X1 U11174 ( .IN1(g4311), .IN2(n9826), .IN3(n11073), .Q(n9915) );
  OR2X1 U11175 ( .IN1(n11130), .IN2(n11131), .Q(n11073) );
  AND2X1 U11176 ( .IN1(g73), .IN2(g4332), .Q(n11131) );
  AND2X1 U11177 ( .IN1(n5540), .IN2(n9473), .Q(n11130) );
  OR2X1 U11178 ( .IN1(n11132), .IN2(n11133), .Q(n9826) );
  AND2X1 U11179 ( .IN1(g72), .IN2(g4322), .Q(n11133) );
  AND2X1 U11180 ( .IN1(n5506), .IN2(n10942), .Q(n11132) );
  INVX0 U11181 ( .INP(g72), .ZN(n10942) );
  INVX0 U11182 ( .INP(n3023), .ZN(n11011) );
  OR4X1 U11183 ( .IN1(n2787), .IN2(n11134), .IN3(n11135), .IN4(n11136), .Q(
        g33608) );
  AND2X1 U11184 ( .IN1(test_so30), .IN2(n9139), .Q(n11136) );
  AND3X1 U11185 ( .IN1(n10473), .IN2(g2759), .IN3(n9076), .Q(n11135) );
  INVX0 U11186 ( .INP(n11137), .ZN(n10473) );
  AND2X1 U11187 ( .IN1(n11137), .IN2(n8793), .Q(n11134) );
  AND2X1 U11188 ( .IN1(test_so30), .IN2(n2790), .Q(n11137) );
  INVX0 U11189 ( .INP(n11138), .ZN(g33607) );
  AND3X1 U11190 ( .IN1(n11139), .IN2(n11140), .IN3(n11141), .Q(n11138) );
  OR2X1 U11191 ( .IN1(n5351), .IN2(n9007), .Q(n11141) );
  OR3X1 U11192 ( .IN1(n11142), .IN2(n11143), .IN3(n11144), .Q(n11140) );
  AND2X1 U11193 ( .IN1(n11145), .IN2(n11146), .Q(n11143) );
  OR4X1 U11194 ( .IN1(n10163), .IN2(g2599), .IN3(n5521), .IN4(n985), .Q(n11146) );
  INVX0 U11195 ( .INP(n10263), .ZN(n985) );
  AND3X1 U11196 ( .IN1(g518), .IN2(n3116), .IN3(n5519), .Q(n10263) );
  OR2X1 U11197 ( .IN1(n9129), .IN2(n11147), .Q(n11145) );
  AND3X1 U11198 ( .IN1(g2629), .IN2(g112), .IN3(n5524), .Q(n11142) );
  OR2X1 U11199 ( .IN1(n5311), .IN2(n11148), .Q(n11139) );
  AND2X1 U11200 ( .IN1(n11149), .IN2(n11150), .Q(n11148) );
  OR2X1 U11201 ( .IN1(n3105), .IN2(n9122), .Q(n11150) );
  OR3X1 U11202 ( .IN1(n11151), .IN2(n11152), .IN3(n11153), .Q(g33606) );
  AND2X1 U11203 ( .IN1(n10477), .IN2(g2675), .Q(n11153) );
  AND2X1 U11204 ( .IN1(n9155), .IN2(g2671), .Q(n11152) );
  AND3X1 U11205 ( .IN1(n5457), .IN2(n10478), .IN3(n9076), .Q(n11151) );
  OR3X1 U11206 ( .IN1(n11154), .IN2(n11155), .IN3(n11156), .Q(g33605) );
  AND2X1 U11207 ( .IN1(n10477), .IN2(g2671), .Q(n11156) );
  AND4X1 U11208 ( .IN1(n10478), .IN2(n9081), .IN3(n5418), .IN4(n8860), .Q(
        n11155) );
  AND2X1 U11209 ( .IN1(test_so48), .IN2(n11157), .Q(n11154) );
  OR2X1 U11210 ( .IN1(n9129), .IN2(n11158), .Q(n11157) );
  AND2X1 U11211 ( .IN1(n10478), .IN2(g2661), .Q(n11158) );
  OR2X1 U11212 ( .IN1(n11159), .IN2(n11160), .Q(g33604) );
  AND2X1 U11213 ( .IN1(n11161), .IN2(g2661), .Q(n11160) );
  AND2X1 U11214 ( .IN1(test_so48), .IN2(n10477), .Q(n11159) );
  OR2X1 U11215 ( .IN1(n11162), .IN2(n11163), .Q(g33603) );
  AND2X1 U11216 ( .IN1(n11161), .IN2(g2643), .Q(n11163) );
  AND2X1 U11217 ( .IN1(n10477), .IN2(g2648), .Q(n11162) );
  INVX0 U11218 ( .INP(n11161), .ZN(n10477) );
  OR2X1 U11219 ( .IN1(n9129), .IN2(n10478), .Q(n11161) );
  AND3X1 U11220 ( .IN1(n10492), .IN2(n5351), .IN3(n5521), .Q(n10478) );
  OR2X1 U11221 ( .IN1(n11164), .IN2(n11165), .Q(g33602) );
  AND2X1 U11222 ( .IN1(n11166), .IN2(g2629), .Q(n11165) );
  AND2X1 U11223 ( .IN1(n11167), .IN2(g2599), .Q(n11164) );
  OR2X1 U11224 ( .IN1(n9129), .IN2(n11168), .Q(n11167) );
  AND2X1 U11225 ( .IN1(n10492), .IN2(n11147), .Q(n11168) );
  OR3X1 U11226 ( .IN1(n11169), .IN2(n11170), .IN3(n11171), .Q(g33601) );
  AND2X1 U11227 ( .IN1(n11166), .IN2(g2599), .Q(n11171) );
  AND4X1 U11228 ( .IN1(n11147), .IN2(g2555), .IN3(n10492), .IN4(n9048), .Q(
        n11170) );
  AND2X1 U11229 ( .IN1(n9155), .IN2(g2606), .Q(n11169) );
  OR2X1 U11230 ( .IN1(n11172), .IN2(n11173), .Q(g33600) );
  AND2X1 U11231 ( .IN1(n11166), .IN2(g2555), .Q(n11173) );
  AND2X1 U11232 ( .IN1(n9037), .IN2(n10487), .Q(n11166) );
  INVX0 U11233 ( .INP(n10492), .ZN(n10487) );
  AND4X1 U11234 ( .IN1(n5521), .IN2(n11174), .IN3(n9048), .IN4(n11147), .Q(
        n11172) );
  INVX0 U11235 ( .INP(n3111), .ZN(n11147) );
  OR2X1 U11236 ( .IN1(n10503), .IN2(g2555), .Q(n11174) );
  AND2X1 U11237 ( .IN1(n10492), .IN2(n5524), .Q(n10503) );
  OR2X1 U11238 ( .IN1(n705), .IN2(n10497), .Q(n10492) );
  OR3X1 U11239 ( .IN1(n11175), .IN2(n11176), .IN3(n11177), .Q(n10497) );
  AND2X1 U11240 ( .IN1(n2549), .IN2(g1300), .Q(n11177) );
  AND3X1 U11241 ( .IN1(g2689), .IN2(g2704), .IN3(g2697), .Q(n11176) );
  INVX0 U11242 ( .INP(n11144), .ZN(n705) );
  OR2X1 U11243 ( .IN1(n11178), .IN2(n8544), .Q(n11144) );
  AND3X1 U11244 ( .IN1(n11179), .IN2(n8819), .IN3(n5364), .Q(n11178) );
  INVX0 U11245 ( .INP(n11180), .ZN(g33599) );
  AND4X1 U11246 ( .IN1(n549), .IN2(n11181), .IN3(n11182), .IN4(n11183), .Q(
        n11180) );
  OR4X1 U11247 ( .IN1(n11184), .IN2(n11185), .IN3(n11186), .IN4(n9121), .Q(
        n11183) );
  OR2X1 U11248 ( .IN1(n8826), .IN2(n9007), .Q(n11182) );
  OR2X1 U11249 ( .IN1(n11187), .IN2(n5619), .Q(n11181) );
  AND2X1 U11250 ( .IN1(n11188), .IN2(n11149), .Q(n11187) );
  OR2X1 U11251 ( .IN1(n9128), .IN2(n3125), .Q(n11188) );
  OR4X1 U11252 ( .IN1(g2465), .IN2(n11184), .IN3(n10163), .IN4(n11189), .Q(
        n549) );
  OR3X1 U11253 ( .IN1(n5522), .IN2(n998), .IN3(n11185), .Q(n11189) );
  AND3X1 U11254 ( .IN1(g112), .IN2(g2495), .IN3(n5523), .Q(n11185) );
  INVX0 U11255 ( .INP(n10262), .ZN(n998) );
  AND3X1 U11256 ( .IN1(g504), .IN2(g518), .IN3(n3116), .Q(n10262) );
  OR3X1 U11257 ( .IN1(n11190), .IN2(n11191), .IN3(n11192), .Q(g33598) );
  AND2X1 U11258 ( .IN1(n10535), .IN2(g2541), .Q(n11192) );
  AND2X1 U11259 ( .IN1(n9155), .IN2(g2537), .Q(n11191) );
  AND3X1 U11260 ( .IN1(n5461), .IN2(n10536), .IN3(n9076), .Q(n11190) );
  OR3X1 U11261 ( .IN1(n11193), .IN2(n11194), .IN3(n11195), .Q(g33597) );
  AND2X1 U11262 ( .IN1(n10535), .IN2(g2537), .Q(n11195) );
  AND4X1 U11263 ( .IN1(n10536), .IN2(n9081), .IN3(n5420), .IN4(n5761), .Q(
        n11194) );
  AND2X1 U11264 ( .IN1(n11196), .IN2(g2533), .Q(n11193) );
  OR2X1 U11265 ( .IN1(n9128), .IN2(n11197), .Q(n11196) );
  AND2X1 U11266 ( .IN1(n10536), .IN2(g2527), .Q(n11197) );
  OR2X1 U11267 ( .IN1(n11198), .IN2(n11199), .Q(g33596) );
  AND2X1 U11268 ( .IN1(n11200), .IN2(g2527), .Q(n11199) );
  AND2X1 U11269 ( .IN1(n10535), .IN2(g2533), .Q(n11198) );
  OR2X1 U11270 ( .IN1(n11201), .IN2(n11202), .Q(g33595) );
  AND2X1 U11271 ( .IN1(n11200), .IN2(g2509), .Q(n11202) );
  AND2X1 U11272 ( .IN1(n10535), .IN2(g2514), .Q(n11201) );
  INVX0 U11273 ( .INP(n11200), .ZN(n10535) );
  OR2X1 U11274 ( .IN1(n9128), .IN2(n10536), .Q(n11200) );
  AND3X1 U11275 ( .IN1(n8826), .IN2(n10550), .IN3(n5522), .Q(n10536) );
  OR3X1 U11276 ( .IN1(n11203), .IN2(n11204), .IN3(n11205), .Q(g33594) );
  AND2X1 U11277 ( .IN1(n9155), .IN2(g2465), .Q(n11205) );
  AND2X1 U11278 ( .IN1(n10567), .IN2(n11186), .Q(n11204) );
  AND2X1 U11279 ( .IN1(n10550), .IN2(g2465), .Q(n10567) );
  AND2X1 U11280 ( .IN1(n11206), .IN2(g2495), .Q(n11203) );
  OR3X1 U11281 ( .IN1(n11207), .IN2(n11208), .IN3(n11209), .Q(g33593) );
  AND2X1 U11282 ( .IN1(n11206), .IN2(g2465), .Q(n11209) );
  AND4X1 U11283 ( .IN1(n10550), .IN2(n11186), .IN3(test_so79), .IN4(n9048), 
        .Q(n11208) );
  AND2X1 U11284 ( .IN1(n9155), .IN2(g2472), .Q(n11207) );
  OR2X1 U11285 ( .IN1(n11210), .IN2(n11211), .Q(g33592) );
  AND2X1 U11286 ( .IN1(n11206), .IN2(test_so79), .Q(n11211) );
  AND2X1 U11287 ( .IN1(n9037), .IN2(n10545), .Q(n11206) );
  INVX0 U11288 ( .INP(n10550), .ZN(n10545) );
  AND4X1 U11289 ( .IN1(n5522), .IN2(n11212), .IN3(n9047), .IN4(n11186), .Q(
        n11210) );
  INVX0 U11290 ( .INP(n3131), .ZN(n11186) );
  OR2X1 U11291 ( .IN1(n10561), .IN2(test_so79), .Q(n11212) );
  AND2X1 U11292 ( .IN1(n10550), .IN2(n5523), .Q(n10561) );
  OR2X1 U11293 ( .IN1(n724), .IN2(n10555), .Q(n10550) );
  OR3X1 U11294 ( .IN1(n11175), .IN2(n11213), .IN3(n11214), .Q(n10555) );
  AND2X1 U11295 ( .IN1(n2549), .IN2(g1472), .Q(n11214) );
  AND3X1 U11296 ( .IN1(g2697), .IN2(g2689), .IN3(n5377), .Q(n11213) );
  INVX0 U11297 ( .INP(n11184), .ZN(n724) );
  OR2X1 U11298 ( .IN1(n11215), .IN2(n8734), .Q(n11184) );
  AND2X1 U11299 ( .IN1(n11179), .IN2(n11216), .Q(n11215) );
  INVX0 U11300 ( .INP(n11217), .ZN(g33591) );
  AND3X1 U11301 ( .IN1(n11218), .IN2(n11219), .IN3(n11220), .Q(n11217) );
  OR2X1 U11302 ( .IN1(n5353), .IN2(n9007), .Q(n11220) );
  OR3X1 U11303 ( .IN1(n11221), .IN2(n11222), .IN3(n11223), .Q(n11219) );
  AND2X1 U11304 ( .IN1(n11224), .IN2(n11225), .Q(n11222) );
  OR2X1 U11305 ( .IN1(n10163), .IN2(n10270), .Q(n11225) );
  OR3X1 U11306 ( .IN1(n5537), .IN2(n997), .IN3(g2331), .Q(n10270) );
  OR2X1 U11307 ( .IN1(n9128), .IN2(n11226), .Q(n11224) );
  AND3X1 U11308 ( .IN1(g2361), .IN2(g112), .IN3(n5513), .Q(n11221) );
  OR2X1 U11309 ( .IN1(n5310), .IN2(n11227), .Q(n11218) );
  AND2X1 U11310 ( .IN1(n11149), .IN2(n11228), .Q(n11227) );
  OR2X1 U11311 ( .IN1(n3145), .IN2(n9122), .Q(n11228) );
  OR3X1 U11312 ( .IN1(n11229), .IN2(n11230), .IN3(n11231), .Q(g33590) );
  AND2X1 U11313 ( .IN1(n10591), .IN2(g2407), .Q(n11231) );
  AND2X1 U11314 ( .IN1(test_so31), .IN2(n9139), .Q(n11230) );
  AND3X1 U11315 ( .IN1(n5459), .IN2(n10592), .IN3(n9076), .Q(n11229) );
  OR3X1 U11316 ( .IN1(n11232), .IN2(n11233), .IN3(n11234), .Q(g33589) );
  AND2X1 U11317 ( .IN1(test_so31), .IN2(n10591), .Q(n11234) );
  AND4X1 U11318 ( .IN1(n10592), .IN2(n9081), .IN3(n5421), .IN4(n5762), .Q(
        n11233) );
  AND2X1 U11319 ( .IN1(n11235), .IN2(g2399), .Q(n11232) );
  OR2X1 U11320 ( .IN1(n9128), .IN2(n11236), .Q(n11235) );
  AND2X1 U11321 ( .IN1(n10592), .IN2(g2393), .Q(n11236) );
  OR2X1 U11322 ( .IN1(n11237), .IN2(n11238), .Q(g33588) );
  AND2X1 U11323 ( .IN1(n11239), .IN2(g2393), .Q(n11238) );
  AND2X1 U11324 ( .IN1(n10591), .IN2(g2399), .Q(n11237) );
  OR2X1 U11325 ( .IN1(n11240), .IN2(n11241), .Q(g33587) );
  AND2X1 U11326 ( .IN1(n11239), .IN2(g2375), .Q(n11241) );
  AND2X1 U11327 ( .IN1(n10591), .IN2(g2380), .Q(n11240) );
  INVX0 U11328 ( .INP(n11239), .ZN(n10591) );
  OR2X1 U11329 ( .IN1(n9128), .IN2(n10592), .Q(n11239) );
  AND3X1 U11330 ( .IN1(n10606), .IN2(n5353), .IN3(n5537), .Q(n10592) );
  OR3X1 U11331 ( .IN1(n11242), .IN2(n11243), .IN3(n11244), .Q(g33586) );
  AND2X1 U11332 ( .IN1(n9155), .IN2(g2331), .Q(n11244) );
  AND2X1 U11333 ( .IN1(n10623), .IN2(n11226), .Q(n11243) );
  AND2X1 U11334 ( .IN1(n10606), .IN2(g2331), .Q(n10623) );
  AND2X1 U11335 ( .IN1(n11245), .IN2(g2361), .Q(n11242) );
  OR3X1 U11336 ( .IN1(n11246), .IN2(n11247), .IN3(n11248), .Q(g33585) );
  AND2X1 U11337 ( .IN1(n11245), .IN2(g2331), .Q(n11248) );
  AND4X1 U11338 ( .IN1(n10606), .IN2(g2287), .IN3(n11226), .IN4(n9048), .Q(
        n11247) );
  AND2X1 U11339 ( .IN1(n9155), .IN2(g2338), .Q(n11246) );
  OR2X1 U11340 ( .IN1(n11249), .IN2(n11250), .Q(g33584) );
  AND2X1 U11341 ( .IN1(n11245), .IN2(g2287), .Q(n11250) );
  AND2X1 U11342 ( .IN1(n9037), .IN2(n10601), .Q(n11245) );
  INVX0 U11343 ( .INP(n10606), .ZN(n10601) );
  AND4X1 U11344 ( .IN1(n5537), .IN2(n11251), .IN3(n11226), .IN4(n9048), .Q(
        n11249) );
  OR2X1 U11345 ( .IN1(n997), .IN2(n11252), .Q(n11226) );
  OR3X1 U11346 ( .IN1(n5519), .IN2(n11253), .IN3(g518), .Q(n997) );
  OR2X1 U11347 ( .IN1(n11254), .IN2(g2287), .Q(n11251) );
  AND2X1 U11348 ( .IN1(n5513), .IN2(n10606), .Q(n11254) );
  OR2X1 U11349 ( .IN1(n388), .IN2(n10611), .Q(n10606) );
  OR3X1 U11350 ( .IN1(n11175), .IN2(n11255), .IN3(n11256), .Q(n10611) );
  AND2X1 U11351 ( .IN1(n2549), .IN2(g1448), .Q(n11256) );
  AND3X1 U11352 ( .IN1(g2689), .IN2(g2704), .IN3(n5308), .Q(n11255) );
  INVX0 U11353 ( .INP(n11223), .ZN(n388) );
  OR2X1 U11354 ( .IN1(n11257), .IN2(n8733), .Q(n11223) );
  AND2X1 U11355 ( .IN1(n11258), .IN2(n11179), .Q(n11257) );
  INVX0 U11356 ( .INP(n11259), .ZN(g33583) );
  AND3X1 U11357 ( .IN1(n11260), .IN2(n11261), .IN3(n11262), .Q(n11259) );
  OR2X1 U11358 ( .IN1(n5356), .IN2(n9007), .Q(n11262) );
  OR3X1 U11359 ( .IN1(n11263), .IN2(n11264), .IN3(n11265), .Q(n11261) );
  AND2X1 U11360 ( .IN1(n11266), .IN2(n11267), .Q(n11264) );
  OR2X1 U11361 ( .IN1(n10163), .IN2(n10271), .Q(n11267) );
  OR3X1 U11362 ( .IN1(n5538), .IN2(n987), .IN3(g2197), .Q(n10271) );
  OR2X1 U11363 ( .IN1(n9128), .IN2(n11268), .Q(n11266) );
  AND3X1 U11364 ( .IN1(g2227), .IN2(g112), .IN3(n5514), .Q(n11263) );
  OR2X1 U11365 ( .IN1(n5620), .IN2(n11269), .Q(n11260) );
  AND2X1 U11366 ( .IN1(n11149), .IN2(n11270), .Q(n11269) );
  OR2X1 U11367 ( .IN1(n3164), .IN2(n9123), .Q(n11270) );
  OR3X1 U11368 ( .IN1(n11271), .IN2(n11272), .IN3(n11273), .Q(g33582) );
  AND2X1 U11369 ( .IN1(n10647), .IN2(g2273), .Q(n11273) );
  AND2X1 U11370 ( .IN1(n9155), .IN2(g2269), .Q(n11272) );
  AND3X1 U11371 ( .IN1(n5458), .IN2(n10648), .IN3(n9076), .Q(n11271) );
  OR3X1 U11372 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .Q(g33581) );
  AND2X1 U11373 ( .IN1(n10647), .IN2(g2269), .Q(n11276) );
  AND4X1 U11374 ( .IN1(n10648), .IN2(n9081), .IN3(n5419), .IN4(n8861), .Q(
        n11275) );
  AND2X1 U11375 ( .IN1(test_so62), .IN2(n11277), .Q(n11274) );
  OR2X1 U11376 ( .IN1(n9127), .IN2(n11278), .Q(n11277) );
  AND2X1 U11377 ( .IN1(n10648), .IN2(g2259), .Q(n11278) );
  OR2X1 U11378 ( .IN1(n11279), .IN2(n11280), .Q(g33580) );
  AND2X1 U11379 ( .IN1(n11281), .IN2(g2259), .Q(n11280) );
  AND2X1 U11380 ( .IN1(test_so62), .IN2(n10647), .Q(n11279) );
  OR2X1 U11381 ( .IN1(n11282), .IN2(n11283), .Q(g33579) );
  AND2X1 U11382 ( .IN1(n11281), .IN2(g2241), .Q(n11283) );
  AND2X1 U11383 ( .IN1(n10647), .IN2(g2246), .Q(n11282) );
  INVX0 U11384 ( .INP(n11281), .ZN(n10647) );
  OR2X1 U11385 ( .IN1(n9127), .IN2(n10648), .Q(n11281) );
  AND3X1 U11386 ( .IN1(n10662), .IN2(n5356), .IN3(n5538), .Q(n10648) );
  OR3X1 U11387 ( .IN1(n11284), .IN2(n11285), .IN3(n11286), .Q(g33578) );
  AND2X1 U11388 ( .IN1(n9155), .IN2(g2197), .Q(n11286) );
  AND2X1 U11389 ( .IN1(n10679), .IN2(n11268), .Q(n11285) );
  AND2X1 U11390 ( .IN1(n10662), .IN2(g2197), .Q(n10679) );
  AND2X1 U11391 ( .IN1(n11287), .IN2(g2227), .Q(n11284) );
  OR3X1 U11392 ( .IN1(n11288), .IN2(n11289), .IN3(n11290), .Q(g33577) );
  AND2X1 U11393 ( .IN1(n11287), .IN2(g2197), .Q(n11290) );
  AND4X1 U11394 ( .IN1(n10662), .IN2(g2153), .IN3(n11268), .IN4(n9049), .Q(
        n11289) );
  AND2X1 U11395 ( .IN1(n9155), .IN2(g2204), .Q(n11288) );
  OR2X1 U11396 ( .IN1(n11291), .IN2(n11292), .Q(g33576) );
  AND2X1 U11397 ( .IN1(n11287), .IN2(g2153), .Q(n11292) );
  AND2X1 U11398 ( .IN1(n9037), .IN2(n10657), .Q(n11287) );
  INVX0 U11399 ( .INP(n10662), .ZN(n10657) );
  AND4X1 U11400 ( .IN1(n5538), .IN2(n11293), .IN3(n11268), .IN4(n9048), .Q(
        n11291) );
  OR2X1 U11401 ( .IN1(n987), .IN2(n11252), .Q(n11268) );
  OR3X1 U11402 ( .IN1(n11253), .IN2(g518), .IN3(g504), .Q(n987) );
  INVX0 U11403 ( .INP(n3116), .ZN(n11253) );
  OR2X1 U11404 ( .IN1(n11294), .IN2(g2153), .Q(n11293) );
  AND2X1 U11405 ( .IN1(n5514), .IN2(n10662), .Q(n11294) );
  OR2X1 U11406 ( .IN1(n719), .IN2(n10667), .Q(n10662) );
  OR3X1 U11407 ( .IN1(n11175), .IN2(n11295), .IN3(n11296), .Q(n10667) );
  AND2X1 U11408 ( .IN1(n2549), .IN2(g1478), .Q(n11296) );
  AND3X1 U11409 ( .IN1(n5377), .IN2(g2689), .IN3(n5308), .Q(n11295) );
  INVX0 U11410 ( .INP(n10699), .ZN(n11175) );
  OR2X1 U11411 ( .IN1(n11297), .IN2(g134), .Q(n10699) );
  AND3X1 U11412 ( .IN1(n11298), .IN2(g691), .IN3(n5595), .Q(n11297) );
  INVX0 U11413 ( .INP(n11265), .ZN(n719) );
  OR2X1 U11414 ( .IN1(n11299), .IN2(n8735), .Q(n11265) );
  AND2X1 U11415 ( .IN1(n11300), .IN2(n11179), .Q(n11299) );
  AND4X1 U11416 ( .IN1(n5768), .IN2(n8729), .IN3(test_so68), .IN4(n11301), .Q(
        n11179) );
  AND3X1 U11417 ( .IN1(g1404), .IN2(n5441), .IN3(n5546), .Q(n11301) );
  OR4X1 U11418 ( .IN1(n11302), .IN2(n11303), .IN3(n11304), .IN4(n11305), .Q(
        g33575) );
  INVX0 U11419 ( .INP(n11306), .ZN(n11305) );
  OR4X1 U11420 ( .IN1(n11307), .IN2(n11308), .IN3(n11309), .IN4(n9121), .Q(
        n11306) );
  AND2X1 U11421 ( .IN1(n9156), .IN2(g1996), .Q(n11304) );
  AND2X1 U11422 ( .IN1(n11310), .IN2(g2047), .Q(n11303) );
  OR2X1 U11423 ( .IN1(n11311), .IN2(n11312), .Q(n11310) );
  AND2X1 U11424 ( .IN1(n11313), .IN2(n9020), .Q(n11311) );
  INVX0 U11425 ( .INP(n282), .ZN(n11302) );
  OR4X1 U11426 ( .IN1(g2040), .IN2(n11313), .IN3(n10163), .IN4(n11314), .Q(
        n282) );
  OR2X1 U11427 ( .IN1(n5535), .IN2(n11308), .Q(n11314) );
  AND3X1 U11428 ( .IN1(g112), .IN2(g2070), .IN3(n5505), .Q(n11308) );
  OR2X1 U11429 ( .IN1(n11307), .IN2(n10252), .Q(n11313) );
  OR3X1 U11430 ( .IN1(n11315), .IN2(n11316), .IN3(n11317), .Q(g33574) );
  AND2X1 U11431 ( .IN1(n10704), .IN2(g2116), .Q(n11317) );
  AND2X1 U11432 ( .IN1(n9156), .IN2(g2112), .Q(n11316) );
  AND3X1 U11433 ( .IN1(n5463), .IN2(n10705), .IN3(n9076), .Q(n11315) );
  OR3X1 U11434 ( .IN1(n11318), .IN2(n11319), .IN3(n11320), .Q(g33573) );
  AND2X1 U11435 ( .IN1(n10704), .IN2(g2112), .Q(n11320) );
  AND4X1 U11436 ( .IN1(n10705), .IN2(n9082), .IN3(n5666), .IN4(n5452), .Q(
        n11319) );
  AND2X1 U11437 ( .IN1(n11321), .IN2(g2108), .Q(n11318) );
  OR2X1 U11438 ( .IN1(n9127), .IN2(n11322), .Q(n11321) );
  AND2X1 U11439 ( .IN1(n10705), .IN2(g2102), .Q(n11322) );
  OR2X1 U11440 ( .IN1(n11323), .IN2(n11324), .Q(g33572) );
  AND2X1 U11441 ( .IN1(n11325), .IN2(g2102), .Q(n11324) );
  AND2X1 U11442 ( .IN1(n10704), .IN2(g2108), .Q(n11323) );
  OR2X1 U11443 ( .IN1(n11326), .IN2(n11327), .Q(g33571) );
  AND2X1 U11444 ( .IN1(n11325), .IN2(g2084), .Q(n11327) );
  AND2X1 U11445 ( .IN1(n10704), .IN2(g2089), .Q(n11326) );
  INVX0 U11446 ( .INP(n11325), .ZN(n10704) );
  OR2X1 U11447 ( .IN1(n9127), .IN2(n10705), .Q(n11325) );
  AND3X1 U11448 ( .IN1(n10719), .IN2(n5355), .IN3(n5535), .Q(n10705) );
  OR2X1 U11449 ( .IN1(n11328), .IN2(n11329), .Q(g33570) );
  AND2X1 U11450 ( .IN1(n11330), .IN2(g2070), .Q(n11329) );
  AND2X1 U11451 ( .IN1(n11331), .IN2(g2040), .Q(n11328) );
  OR2X1 U11452 ( .IN1(n9127), .IN2(n11332), .Q(n11331) );
  AND2X1 U11453 ( .IN1(n11309), .IN2(n10719), .Q(n11332) );
  OR3X1 U11454 ( .IN1(n11333), .IN2(n11334), .IN3(n11335), .Q(g33569) );
  AND2X1 U11455 ( .IN1(n11330), .IN2(g2040), .Q(n11335) );
  AND4X1 U11456 ( .IN1(n10719), .IN2(g1996), .IN3(n11309), .IN4(n9048), .Q(
        n11334) );
  AND2X1 U11457 ( .IN1(n9156), .IN2(g2047), .Q(n11333) );
  OR2X1 U11458 ( .IN1(n11336), .IN2(n11337), .Q(g33568) );
  AND2X1 U11459 ( .IN1(n11330), .IN2(g1996), .Q(n11337) );
  AND2X1 U11460 ( .IN1(n9037), .IN2(n10714), .Q(n11330) );
  AND4X1 U11461 ( .IN1(n5535), .IN2(n11338), .IN3(n11309), .IN4(n9050), .Q(
        n11336) );
  OR2X1 U11462 ( .IN1(n10252), .IN2(n11252), .Q(n11309) );
  INVX0 U11463 ( .INP(n10265), .ZN(n10252) );
  AND3X1 U11464 ( .IN1(g518), .IN2(n5519), .IN3(n3195), .Q(n10265) );
  OR2X1 U11465 ( .IN1(n11339), .IN2(g1996), .Q(n11338) );
  AND2X1 U11466 ( .IN1(n5505), .IN2(n10719), .Q(n11339) );
  INVX0 U11467 ( .INP(n10714), .ZN(n10719) );
  AND2X1 U11468 ( .IN1(n11307), .IN2(n10755), .Q(n10714) );
  INVX0 U11469 ( .INP(n10724), .ZN(n10755) );
  OR3X1 U11470 ( .IN1(n11340), .IN2(n11341), .IN3(n11342), .Q(n10724) );
  AND2X1 U11471 ( .IN1(n5286), .IN2(g956), .Q(n11342) );
  AND3X1 U11472 ( .IN1(g2145), .IN2(g2130), .IN3(g2138), .Q(n11341) );
  OR2X1 U11473 ( .IN1(n11343), .IN2(n8543), .Q(n11307) );
  AND3X1 U11474 ( .IN1(n5363), .IN2(n11344), .IN3(n5599), .Q(n11343) );
  OR3X1 U11475 ( .IN1(n11345), .IN2(n11346), .IN3(n11347), .Q(g33567) );
  AND2X1 U11476 ( .IN1(test_so8), .IN2(n9139), .Q(n11347) );
  AND2X1 U11477 ( .IN1(n11348), .IN2(g1913), .Q(n11346) );
  OR2X1 U11478 ( .IN1(n11349), .IN2(n11312), .Q(n11348) );
  AND2X1 U11479 ( .IN1(n11350), .IN2(n9020), .Q(n11349) );
  OR2X1 U11480 ( .IN1(n10253), .IN2(n11351), .Q(n11350) );
  INVX0 U11481 ( .INP(n11352), .ZN(n10253) );
  AND3X1 U11482 ( .IN1(n11353), .IN2(n11354), .IN3(n11355), .Q(n11345) );
  OR3X1 U11483 ( .IN1(n8671), .IN2(n5534), .IN3(g1906), .Q(n11354) );
  OR2X1 U11484 ( .IN1(n11356), .IN2(n11357), .Q(n11353) );
  AND2X1 U11485 ( .IN1(n11358), .IN2(n9020), .Q(n11357) );
  AND2X1 U11486 ( .IN1(n10267), .IN2(n10147), .Q(n11356) );
  AND3X1 U11487 ( .IN1(g1936), .IN2(n11352), .IN3(n5503), .Q(n10267) );
  OR3X1 U11488 ( .IN1(n11359), .IN2(n11360), .IN3(n11361), .Q(g33566) );
  AND2X1 U11489 ( .IN1(n10762), .IN2(g1982), .Q(n11361) );
  AND2X1 U11490 ( .IN1(n9156), .IN2(g1978), .Q(n11360) );
  AND3X1 U11491 ( .IN1(n5462), .IN2(n10763), .IN3(n9077), .Q(n11359) );
  OR3X1 U11492 ( .IN1(n11362), .IN2(n11363), .IN3(n11364), .Q(g33565) );
  AND2X1 U11493 ( .IN1(n10762), .IN2(g1978), .Q(n11364) );
  AND4X1 U11494 ( .IN1(n10763), .IN2(n9081), .IN3(n5664), .IN4(n5450), .Q(
        n11363) );
  AND2X1 U11495 ( .IN1(n11365), .IN2(g1974), .Q(n11362) );
  OR2X1 U11496 ( .IN1(n9127), .IN2(n11366), .Q(n11365) );
  AND2X1 U11497 ( .IN1(n10763), .IN2(g1968), .Q(n11366) );
  OR2X1 U11498 ( .IN1(n11367), .IN2(n11368), .Q(g33564) );
  AND2X1 U11499 ( .IN1(n11369), .IN2(g1968), .Q(n11368) );
  AND2X1 U11500 ( .IN1(n10762), .IN2(g1974), .Q(n11367) );
  OR2X1 U11501 ( .IN1(n11370), .IN2(n11371), .Q(g33563) );
  AND2X1 U11502 ( .IN1(n11369), .IN2(g1950), .Q(n11371) );
  AND2X1 U11503 ( .IN1(n10762), .IN2(g1955), .Q(n11370) );
  INVX0 U11504 ( .INP(n11369), .ZN(n10762) );
  OR2X1 U11505 ( .IN1(n9127), .IN2(n10763), .Q(n11369) );
  AND3X1 U11506 ( .IN1(n8827), .IN2(n10777), .IN3(n5534), .Q(n10763) );
  OR3X1 U11507 ( .IN1(n11372), .IN2(n11373), .IN3(n11374), .Q(g33562) );
  AND2X1 U11508 ( .IN1(n9156), .IN2(g1906), .Q(n11374) );
  AND2X1 U11509 ( .IN1(n10794), .IN2(n11375), .Q(n11373) );
  AND2X1 U11510 ( .IN1(n10777), .IN2(g1906), .Q(n10794) );
  AND2X1 U11511 ( .IN1(n11376), .IN2(g1936), .Q(n11372) );
  OR3X1 U11512 ( .IN1(n11377), .IN2(n11378), .IN3(n11379), .Q(g33561) );
  AND2X1 U11513 ( .IN1(n11376), .IN2(g1906), .Q(n11379) );
  AND4X1 U11514 ( .IN1(n11375), .IN2(n10777), .IN3(test_so8), .IN4(n9048), .Q(
        n11378) );
  AND2X1 U11515 ( .IN1(n9156), .IN2(g1913), .Q(n11377) );
  OR2X1 U11516 ( .IN1(n11380), .IN2(n11381), .Q(g33560) );
  AND2X1 U11517 ( .IN1(n11376), .IN2(test_so8), .Q(n11381) );
  AND2X1 U11518 ( .IN1(n9036), .IN2(n10772), .Q(n11376) );
  INVX0 U11519 ( .INP(n10777), .ZN(n10772) );
  AND4X1 U11520 ( .IN1(n5534), .IN2(n11382), .IN3(n11375), .IN4(n9048), .Q(
        n11380) );
  INVX0 U11521 ( .INP(n11358), .ZN(n11375) );
  AND2X1 U11522 ( .IN1(n11352), .IN2(n3115), .Q(n11358) );
  AND3X1 U11523 ( .IN1(g504), .IN2(g518), .IN3(n3195), .Q(n11352) );
  OR2X1 U11524 ( .IN1(n11383), .IN2(test_so8), .Q(n11382) );
  AND2X1 U11525 ( .IN1(n5503), .IN2(n10777), .Q(n11383) );
  OR2X1 U11526 ( .IN1(n11355), .IN2(n10782), .Q(n10777) );
  OR3X1 U11527 ( .IN1(n11340), .IN2(n11384), .IN3(n11385), .Q(n10782) );
  AND2X1 U11528 ( .IN1(n5286), .IN2(g1129), .Q(n11385) );
  AND3X1 U11529 ( .IN1(g2138), .IN2(g2130), .IN3(n5307), .Q(n11384) );
  INVX0 U11530 ( .INP(n11351), .ZN(n11355) );
  OR2X1 U11531 ( .IN1(n11386), .IN2(n8698), .Q(n11351) );
  AND2X1 U11532 ( .IN1(n11387), .IN2(n11344), .Q(n11386) );
  OR3X1 U11533 ( .IN1(n11388), .IN2(n11389), .IN3(n11390), .Q(g33559) );
  AND2X1 U11534 ( .IN1(n9156), .IN2(g1728), .Q(n11390) );
  AND2X1 U11535 ( .IN1(n11391), .IN2(g1779), .Q(n11389) );
  OR2X1 U11536 ( .IN1(n11392), .IN2(n11312), .Q(n11391) );
  AND2X1 U11537 ( .IN1(n11393), .IN2(n9020), .Q(n11392) );
  OR2X1 U11538 ( .IN1(n10254), .IN2(n11394), .Q(n11393) );
  INVX0 U11539 ( .INP(n11395), .ZN(n10254) );
  AND3X1 U11540 ( .IN1(n11396), .IN2(n11397), .IN3(n11398), .Q(n11388) );
  OR3X1 U11541 ( .IN1(n8671), .IN2(n5536), .IN3(g1772), .Q(n11397) );
  OR2X1 U11542 ( .IN1(n11399), .IN2(n11400), .Q(n11396) );
  AND2X1 U11543 ( .IN1(n11401), .IN2(n9021), .Q(n11400) );
  AND2X1 U11544 ( .IN1(n10266), .IN2(n10147), .Q(n11399) );
  AND3X1 U11545 ( .IN1(g1802), .IN2(n11395), .IN3(n5504), .Q(n10266) );
  OR3X1 U11546 ( .IN1(n11402), .IN2(n11403), .IN3(n11404), .Q(g33558) );
  AND2X1 U11547 ( .IN1(n10818), .IN2(g1848), .Q(n11404) );
  AND2X1 U11548 ( .IN1(n9156), .IN2(g1844), .Q(n11403) );
  AND3X1 U11549 ( .IN1(n5464), .IN2(n10819), .IN3(n9077), .Q(n11402) );
  OR3X1 U11550 ( .IN1(n11405), .IN2(n11406), .IN3(n11407), .Q(g33557) );
  AND2X1 U11551 ( .IN1(n10818), .IN2(g1844), .Q(n11407) );
  AND4X1 U11552 ( .IN1(n10819), .IN2(n9081), .IN3(n5665), .IN4(n5451), .Q(
        n11406) );
  AND2X1 U11553 ( .IN1(n11408), .IN2(g1840), .Q(n11405) );
  OR2X1 U11554 ( .IN1(n9127), .IN2(n11409), .Q(n11408) );
  AND2X1 U11555 ( .IN1(n10819), .IN2(g1834), .Q(n11409) );
  OR2X1 U11556 ( .IN1(n11410), .IN2(n11411), .Q(g33556) );
  AND2X1 U11557 ( .IN1(n11412), .IN2(g1834), .Q(n11411) );
  AND2X1 U11558 ( .IN1(n10818), .IN2(g1840), .Q(n11410) );
  OR2X1 U11559 ( .IN1(n11413), .IN2(n11414), .Q(g33555) );
  AND2X1 U11560 ( .IN1(n11412), .IN2(g1816), .Q(n11414) );
  AND2X1 U11561 ( .IN1(n10818), .IN2(g1821), .Q(n11413) );
  INVX0 U11562 ( .INP(n11412), .ZN(n10818) );
  OR2X1 U11563 ( .IN1(n9127), .IN2(n10819), .Q(n11412) );
  AND3X1 U11564 ( .IN1(n10833), .IN2(n5352), .IN3(n5536), .Q(n10819) );
  OR3X1 U11565 ( .IN1(n11415), .IN2(n11416), .IN3(n11417), .Q(g33554) );
  AND2X1 U11566 ( .IN1(n9156), .IN2(g1772), .Q(n11417) );
  AND2X1 U11567 ( .IN1(n10850), .IN2(n11418), .Q(n11416) );
  AND2X1 U11568 ( .IN1(n10833), .IN2(g1772), .Q(n10850) );
  AND2X1 U11569 ( .IN1(n11419), .IN2(g1802), .Q(n11415) );
  OR3X1 U11570 ( .IN1(n11420), .IN2(n11421), .IN3(n11422), .Q(g33553) );
  AND2X1 U11571 ( .IN1(n11419), .IN2(g1772), .Q(n11422) );
  AND4X1 U11572 ( .IN1(n10833), .IN2(g1728), .IN3(n11418), .IN4(n9050), .Q(
        n11421) );
  AND2X1 U11573 ( .IN1(n9156), .IN2(g1779), .Q(n11420) );
  OR2X1 U11574 ( .IN1(n11423), .IN2(n11424), .Q(g33552) );
  AND2X1 U11575 ( .IN1(n11419), .IN2(g1728), .Q(n11424) );
  AND2X1 U11576 ( .IN1(n9036), .IN2(n10828), .Q(n11419) );
  INVX0 U11577 ( .INP(n10833), .ZN(n10828) );
  AND4X1 U11578 ( .IN1(n5536), .IN2(n11425), .IN3(n11418), .IN4(n9048), .Q(
        n11423) );
  INVX0 U11579 ( .INP(n11401), .ZN(n11418) );
  AND2X1 U11580 ( .IN1(n11395), .IN2(n3115), .Q(n11401) );
  AND3X1 U11581 ( .IN1(g504), .IN2(n5287), .IN3(n3195), .Q(n11395) );
  OR2X1 U11582 ( .IN1(n11426), .IN2(g1728), .Q(n11425) );
  AND2X1 U11583 ( .IN1(n5504), .IN2(n10833), .Q(n11426) );
  OR2X1 U11584 ( .IN1(n11398), .IN2(n10838), .Q(n10833) );
  OR3X1 U11585 ( .IN1(n11340), .IN2(n11427), .IN3(n11428), .Q(n10838) );
  AND2X1 U11586 ( .IN1(n5286), .IN2(g1105), .Q(n11428) );
  AND3X1 U11587 ( .IN1(g2145), .IN2(g2130), .IN3(n5275), .Q(n11427) );
  INVX0 U11588 ( .INP(n11394), .ZN(n11398) );
  OR2X1 U11589 ( .IN1(n11429), .IN2(n8841), .Q(n11394) );
  AND2X1 U11590 ( .IN1(n11430), .IN2(n11344), .Q(n11429) );
  OR4X1 U11591 ( .IN1(n11431), .IN2(n11432), .IN3(n11433), .IN4(n11434), .Q(
        g33551) );
  AND2X1 U11592 ( .IN1(n11435), .IN2(n9021), .Q(n11434) );
  OR2X1 U11593 ( .IN1(n11436), .IN2(n11437), .Q(n11435) );
  AND2X1 U11594 ( .IN1(test_so75), .IN2(n11438), .Q(n11437) );
  OR2X1 U11595 ( .IN1(n10255), .IN2(n11439), .Q(n11438) );
  INVX0 U11596 ( .INP(n11440), .ZN(n11436) );
  OR3X1 U11597 ( .IN1(n11439), .IN2(n11441), .IN3(n11442), .Q(n11440) );
  AND2X1 U11598 ( .IN1(g112), .IN2(g31862), .Q(n11441) );
  AND2X1 U11599 ( .IN1(n9156), .IN2(g1592), .Q(n11433) );
  AND2X1 U11600 ( .IN1(test_so75), .IN2(n11312), .Q(n11432) );
  AND3X1 U11601 ( .IN1(n8671), .IN2(g33533), .IN3(n11443), .Q(n11431) );
  AND3X1 U11602 ( .IN1(n10264), .IN2(n10147), .IN3(g31862), .Q(n11443) );
  OR3X1 U11603 ( .IN1(n11444), .IN2(n11445), .IN3(n11446), .Q(g33550) );
  AND2X1 U11604 ( .IN1(n10874), .IN2(g1714), .Q(n11446) );
  AND2X1 U11605 ( .IN1(n9156), .IN2(g1710), .Q(n11445) );
  AND3X1 U11606 ( .IN1(n5460), .IN2(n10875), .IN3(n9077), .Q(n11444) );
  OR3X1 U11607 ( .IN1(n11447), .IN2(n11448), .IN3(n11449), .Q(g33549) );
  AND2X1 U11608 ( .IN1(n10874), .IN2(g1710), .Q(n11449) );
  AND4X1 U11609 ( .IN1(n10875), .IN2(n9081), .IN3(n5417), .IN4(n8862), .Q(
        n11448) );
  AND2X1 U11610 ( .IN1(test_so15), .IN2(n11450), .Q(n11447) );
  OR2X1 U11611 ( .IN1(n9126), .IN2(n11451), .Q(n11450) );
  AND2X1 U11612 ( .IN1(n10875), .IN2(g1700), .Q(n11451) );
  OR2X1 U11613 ( .IN1(n11452), .IN2(n11453), .Q(g33548) );
  AND2X1 U11614 ( .IN1(n11454), .IN2(g1700), .Q(n11453) );
  AND2X1 U11615 ( .IN1(test_so15), .IN2(n10874), .Q(n11452) );
  OR2X1 U11616 ( .IN1(n11455), .IN2(n11456), .Q(g33547) );
  AND2X1 U11617 ( .IN1(n11454), .IN2(g1682), .Q(n11456) );
  AND2X1 U11618 ( .IN1(n10874), .IN2(g1687), .Q(n11455) );
  INVX0 U11619 ( .INP(n11454), .ZN(n10874) );
  OR2X1 U11620 ( .IN1(n9126), .IN2(n10875), .Q(n11454) );
  AND3X1 U11621 ( .IN1(n10889), .IN2(n5362), .IN3(n5598), .Q(n10875) );
  OR3X1 U11622 ( .IN1(n11457), .IN2(n11458), .IN3(n11459), .Q(g33546) );
  AND2X1 U11623 ( .IN1(n9156), .IN2(g1636), .Q(n11459) );
  AND2X1 U11624 ( .IN1(n10905), .IN2(n11442), .Q(n11458) );
  AND2X1 U11625 ( .IN1(n10889), .IN2(g1636), .Q(n10905) );
  AND2X1 U11626 ( .IN1(n11460), .IN2(g1668), .Q(n11457) );
  OR3X1 U11627 ( .IN1(n11461), .IN2(n11462), .IN3(n11463), .Q(g33545) );
  AND2X1 U11628 ( .IN1(n11460), .IN2(g1636), .Q(n11463) );
  AND3X1 U11629 ( .IN1(n10911), .IN2(n11442), .IN3(n9077), .Q(n11462) );
  AND2X1 U11630 ( .IN1(n10889), .IN2(g1592), .Q(n10911) );
  AND2X1 U11631 ( .IN1(test_so75), .IN2(n9138), .Q(n11461) );
  OR2X1 U11632 ( .IN1(n11464), .IN2(n11465), .Q(g33544) );
  AND2X1 U11633 ( .IN1(n11460), .IN2(g1592), .Q(n11465) );
  AND2X1 U11634 ( .IN1(n9036), .IN2(n10884), .Q(n11460) );
  INVX0 U11635 ( .INP(n10889), .ZN(n10884) );
  AND4X1 U11636 ( .IN1(n5598), .IN2(n11466), .IN3(n11442), .IN4(n9048), .Q(
        n11464) );
  OR2X1 U11637 ( .IN1(n10255), .IN2(n11252), .Q(n11442) );
  INVX0 U11638 ( .INP(n3115), .ZN(n11252) );
  INVX0 U11639 ( .INP(n10264), .ZN(n10255) );
  AND3X1 U11640 ( .IN1(n5287), .IN2(n5519), .IN3(n3195), .Q(n10264) );
  OR2X1 U11641 ( .IN1(n11467), .IN2(g1592), .Q(n11466) );
  AND2X1 U11642 ( .IN1(n5549), .IN2(n10889), .Q(n11467) );
  OR2X1 U11643 ( .IN1(g33533), .IN2(n10894), .Q(n10889) );
  OR3X1 U11644 ( .IN1(n11340), .IN2(n11468), .IN3(n11469), .Q(n10894) );
  AND2X1 U11645 ( .IN1(n5286), .IN2(g1135), .Q(n11469) );
  AND3X1 U11646 ( .IN1(n5307), .IN2(g2130), .IN3(n5275), .Q(n11468) );
  INVX0 U11647 ( .INP(n10926), .ZN(n11340) );
  OR2X1 U11648 ( .IN1(n11470), .IN2(g134), .Q(n10926) );
  AND3X1 U11649 ( .IN1(n11471), .IN2(g691), .IN3(n5595), .Q(n11470) );
  OR2X1 U11650 ( .IN1(n11472), .IN2(n11473), .Q(g33543) );
  AND2X1 U11651 ( .IN1(n11474), .IN2(g1373), .Q(n11473) );
  OR2X1 U11652 ( .IN1(n9126), .IN2(n11475), .Q(n11474) );
  AND3X1 U11653 ( .IN1(n11476), .IN2(n11477), .IN3(n8797), .Q(n11475) );
  AND3X1 U11654 ( .IN1(n9054), .IN2(g1379), .IN3(n11478), .Q(n11472) );
  OR2X1 U11655 ( .IN1(n11479), .IN2(n11480), .Q(n11478) );
  AND2X1 U11656 ( .IN1(n8657), .IN2(n11477), .Q(n11479) );
  OR3X1 U11657 ( .IN1(n11481), .IN2(n11482), .IN3(n11483), .Q(g33542) );
  AND2X1 U11658 ( .IN1(n9156), .IN2(g1270), .Q(n11483) );
  AND2X1 U11659 ( .IN1(n5730), .IN2(n11484), .Q(n11482) );
  AND3X1 U11660 ( .IN1(n11485), .IN2(n11486), .IN3(g1274), .Q(n11481) );
  OR2X1 U11661 ( .IN1(n11487), .IN2(n11488), .Q(g33541) );
  AND2X1 U11662 ( .IN1(n11489), .IN2(g1030), .Q(n11488) );
  OR2X1 U11663 ( .IN1(n9126), .IN2(n11490), .Q(n11489) );
  AND3X1 U11664 ( .IN1(n11491), .IN2(n11492), .IN3(n8794), .Q(n11490) );
  AND3X1 U11665 ( .IN1(n9054), .IN2(g1036), .IN3(n11493), .Q(n11487) );
  OR2X1 U11666 ( .IN1(n11494), .IN2(n11495), .Q(n11493) );
  AND2X1 U11667 ( .IN1(n8656), .IN2(n11492), .Q(n11494) );
  OR3X1 U11668 ( .IN1(n11496), .IN2(n11497), .IN3(n11498), .Q(g33540) );
  AND2X1 U11669 ( .IN1(n9156), .IN2(g925), .Q(n11498) );
  AND2X1 U11670 ( .IN1(n5731), .IN2(n11499), .Q(n11497) );
  AND3X1 U11671 ( .IN1(n11500), .IN2(n11501), .IN3(g930), .Q(n11496) );
  OR3X1 U11672 ( .IN1(n11502), .IN2(n11503), .IN3(n11504), .Q(g33539) );
  AND2X1 U11673 ( .IN1(n9156), .IN2(g758), .Q(n11504) );
  AND2X1 U11674 ( .IN1(n2980), .IN2(n5332), .Q(n11503) );
  AND3X1 U11675 ( .IN1(n2404), .IN2(n11505), .IN3(g763), .Q(n11502) );
  INVX0 U11676 ( .INP(n2980), .ZN(n11505) );
  OR3X1 U11677 ( .IN1(n11506), .IN2(n11507), .IN3(n11508), .Q(g33538) );
  AND2X1 U11678 ( .IN1(n9156), .IN2(g590), .Q(n11508) );
  AND2X1 U11679 ( .IN1(n2982), .IN2(n5476), .Q(n11507) );
  AND3X1 U11680 ( .IN1(n2421), .IN2(n11509), .IN3(g595), .Q(n11506) );
  INVX0 U11681 ( .INP(n2982), .ZN(n11509) );
  OR2X1 U11682 ( .IN1(n11510), .IN2(n11511), .Q(g33537) );
  AND3X1 U11683 ( .IN1(n2707), .IN2(g142), .IN3(n9077), .Q(n11511) );
  AND2X1 U11684 ( .IN1(n9168), .IN2(g301), .Q(n11510) );
  AND2X1 U11685 ( .IN1(n11512), .IN2(g160), .Q(g33536) );
  OR2X1 U11686 ( .IN1(n2710), .IN2(n9123), .Q(n11512) );
  OR3X1 U11687 ( .IN1(n11513), .IN2(n11514), .IN3(n11515), .Q(g33535) );
  AND2X1 U11688 ( .IN1(n9166), .IN2(g291), .Q(n11515) );
  AND2X1 U11689 ( .IN1(n3276), .IN2(n5680), .Q(n11514) );
  AND3X1 U11690 ( .IN1(n8803), .IN2(n11516), .IN3(g294), .Q(n11513) );
  INVX0 U11691 ( .INP(n3276), .ZN(n11516) );
  OR3X1 U11692 ( .IN1(n11517), .IN2(n11518), .IN3(n11519), .Q(g33534) );
  AND2X1 U11693 ( .IN1(n9166), .IN2(g150), .Q(n11519) );
  AND2X1 U11694 ( .IN1(n3277), .IN2(n5677), .Q(n11518) );
  AND3X1 U11695 ( .IN1(n10380), .IN2(n11520), .IN3(g153), .Q(n11517) );
  INVX0 U11696 ( .INP(n3277), .ZN(n11520) );
  INVX0 U11697 ( .INP(n11439), .ZN(g33533) );
  OR2X1 U11698 ( .IN1(n11521), .IN2(n8699), .Q(n11439) );
  AND3X1 U11699 ( .IN1(n11344), .IN2(g1171), .IN3(n5599), .Q(n11521) );
  AND4X1 U11700 ( .IN1(n8730), .IN2(n5442), .IN3(n5547), .IN4(n11522), .Q(
        n11344) );
  AND3X1 U11701 ( .IN1(n8839), .IN2(g1061), .IN3(g979), .Q(n11522) );
  AND3X1 U11702 ( .IN1(n11523), .IN2(n11524), .IN3(n11525), .Q(g33435) );
  OR2X1 U11703 ( .IN1(n5610), .IN2(n10178), .Q(n11525) );
  OR3X1 U11704 ( .IN1(n11526), .IN2(n11527), .IN3(g2729), .Q(n11524) );
  AND2X1 U11705 ( .IN1(n5544), .IN2(n5301), .Q(n11527) );
  AND2X1 U11706 ( .IN1(n5378), .IN2(g2724), .Q(n11526) );
  OR2X1 U11707 ( .IN1(n5403), .IN2(n10191), .Q(n11523) );
  AND3X1 U11708 ( .IN1(n11528), .IN2(n11529), .IN3(n11530), .Q(g33079) );
  OR2X1 U11709 ( .IN1(n5609), .IN2(n10178), .Q(n11530) );
  OR3X1 U11710 ( .IN1(n11531), .IN2(n11532), .IN3(g2729), .Q(n11529) );
  AND2X1 U11711 ( .IN1(n5545), .IN2(n5301), .Q(n11532) );
  AND2X1 U11712 ( .IN1(n5379), .IN2(g2724), .Q(n11531) );
  OR2X1 U11713 ( .IN1(n5404), .IN2(n10191), .Q(n11528) );
  OR2X1 U11714 ( .IN1(n8676), .IN2(g2724), .Q(n10191) );
  OR2X1 U11715 ( .IN1(n11533), .IN2(n11534), .Q(g33070) );
  AND2X1 U11716 ( .IN1(n9166), .IN2(g6565), .Q(n11534) );
  AND2X1 U11717 ( .IN1(n11535), .IN2(n11536), .Q(n11533) );
  OR3X1 U11718 ( .IN1(n11537), .IN2(n11538), .IN3(n11539), .Q(n11535) );
  AND2X1 U11719 ( .IN1(g25756), .IN2(n5646), .Q(n11539) );
  AND2X1 U11720 ( .IN1(n11540), .IN2(n9021), .Q(n11538) );
  OR2X1 U11721 ( .IN1(n11541), .IN2(n11542), .Q(g33069) );
  AND2X1 U11722 ( .IN1(n11543), .IN2(g6565), .Q(n11542) );
  AND2X1 U11723 ( .IN1(n11544), .IN2(g6561), .Q(n11541) );
  OR2X1 U11724 ( .IN1(n9125), .IN2(n11545), .Q(n11544) );
  AND2X1 U11725 ( .IN1(n5386), .IN2(n11536), .Q(n11545) );
  OR2X1 U11726 ( .IN1(n11546), .IN2(n11547), .Q(g33068) );
  AND2X1 U11727 ( .IN1(n9166), .IN2(g6555), .Q(n11547) );
  AND3X1 U11728 ( .IN1(n11536), .IN2(n11548), .IN3(n5646), .Q(n11546) );
  INVX0 U11729 ( .INP(n769), .ZN(n11548) );
  OR2X1 U11730 ( .IN1(n11549), .IN2(n11550), .Q(g33067) );
  AND2X1 U11731 ( .IN1(n9166), .IN2(g6549), .Q(n11550) );
  AND2X1 U11732 ( .IN1(n11551), .IN2(n11536), .Q(n11549) );
  INVX0 U11733 ( .INP(n11552), .ZN(n11551) );
  AND2X1 U11734 ( .IN1(n11553), .IN2(n3407), .Q(n11552) );
  OR2X1 U11735 ( .IN1(n9124), .IN2(n3406), .Q(n11553) );
  OR2X1 U11736 ( .IN1(n11554), .IN2(n11555), .Q(g33065) );
  AND2X1 U11737 ( .IN1(n9166), .IN2(g6219), .Q(n11555) );
  AND2X1 U11738 ( .IN1(n11556), .IN2(n11557), .Q(n11554) );
  OR3X1 U11739 ( .IN1(n11558), .IN2(n11559), .IN3(n11560), .Q(n11556) );
  AND2X1 U11740 ( .IN1(g25742), .IN2(n5651), .Q(n11560) );
  AND2X1 U11741 ( .IN1(n9036), .IN2(n11561), .Q(n11559) );
  OR2X1 U11742 ( .IN1(n11562), .IN2(n11563), .Q(g33064) );
  AND2X1 U11743 ( .IN1(n11564), .IN2(g6219), .Q(n11563) );
  AND2X1 U11744 ( .IN1(n11565), .IN2(g6215), .Q(n11562) );
  OR2X1 U11745 ( .IN1(n9125), .IN2(n11566), .Q(n11565) );
  AND2X1 U11746 ( .IN1(n5385), .IN2(n11557), .Q(n11566) );
  OR2X1 U11747 ( .IN1(n11567), .IN2(n11568), .Q(g33063) );
  AND2X1 U11748 ( .IN1(n9166), .IN2(g6209), .Q(n11568) );
  AND3X1 U11749 ( .IN1(n11557), .IN2(n11569), .IN3(n5651), .Q(n11567) );
  INVX0 U11750 ( .INP(n1022), .ZN(n11569) );
  OR2X1 U11751 ( .IN1(n11570), .IN2(n11571), .Q(g33062) );
  AND2X1 U11752 ( .IN1(n9166), .IN2(g6203), .Q(n11571) );
  AND2X1 U11753 ( .IN1(n11572), .IN2(n11557), .Q(n11570) );
  INVX0 U11754 ( .INP(n11573), .ZN(n11572) );
  AND2X1 U11755 ( .IN1(n11574), .IN2(n3417), .Q(n11573) );
  OR2X1 U11756 ( .IN1(n9125), .IN2(n3416), .Q(n11574) );
  OR2X1 U11757 ( .IN1(n11575), .IN2(n11576), .Q(g33060) );
  AND2X1 U11758 ( .IN1(n9166), .IN2(g5873), .Q(n11576) );
  AND2X1 U11759 ( .IN1(n11577), .IN2(n11578), .Q(n11575) );
  OR3X1 U11760 ( .IN1(n11579), .IN2(n11580), .IN3(n11581), .Q(n11577) );
  AND2X1 U11761 ( .IN1(g25728), .IN2(n5649), .Q(n11581) );
  AND2X1 U11762 ( .IN1(n9036), .IN2(n11582), .Q(n11580) );
  OR2X1 U11763 ( .IN1(n11583), .IN2(n11584), .Q(g33059) );
  AND2X1 U11764 ( .IN1(n11585), .IN2(g5873), .Q(n11584) );
  AND2X1 U11765 ( .IN1(n11586), .IN2(g5869), .Q(n11583) );
  OR2X1 U11766 ( .IN1(n9125), .IN2(n11587), .Q(n11586) );
  AND2X1 U11767 ( .IN1(n5388), .IN2(n11578), .Q(n11587) );
  OR2X1 U11768 ( .IN1(n11588), .IN2(n11589), .Q(g33058) );
  AND2X1 U11769 ( .IN1(n9166), .IN2(g5863), .Q(n11589) );
  AND3X1 U11770 ( .IN1(n11578), .IN2(n11590), .IN3(n5649), .Q(n11588) );
  INVX0 U11771 ( .INP(n1084), .ZN(n11590) );
  OR2X1 U11772 ( .IN1(n11591), .IN2(n11592), .Q(g33057) );
  AND2X1 U11773 ( .IN1(n9166), .IN2(g5857), .Q(n11592) );
  AND2X1 U11774 ( .IN1(n11593), .IN2(n11578), .Q(n11591) );
  INVX0 U11775 ( .INP(n11594), .ZN(n11593) );
  AND2X1 U11776 ( .IN1(n11595), .IN2(n3427), .Q(n11594) );
  OR2X1 U11777 ( .IN1(n9124), .IN2(n3426), .Q(n11595) );
  OR2X1 U11778 ( .IN1(n11596), .IN2(n11597), .Q(g33055) );
  AND2X1 U11779 ( .IN1(n9166), .IN2(g5527), .Q(n11597) );
  AND2X1 U11780 ( .IN1(n11598), .IN2(n11599), .Q(n11596) );
  OR3X1 U11781 ( .IN1(n11600), .IN2(n11601), .IN3(n11602), .Q(n11598) );
  AND2X1 U11782 ( .IN1(g25714), .IN2(n5647), .Q(n11602) );
  AND2X1 U11783 ( .IN1(n9035), .IN2(n11603), .Q(n11601) );
  OR2X1 U11784 ( .IN1(n11604), .IN2(n11605), .Q(g33054) );
  AND2X1 U11785 ( .IN1(n11606), .IN2(g5527), .Q(n11605) );
  AND2X1 U11786 ( .IN1(n11607), .IN2(g5523), .Q(n11604) );
  OR2X1 U11787 ( .IN1(n9125), .IN2(n11608), .Q(n11607) );
  AND2X1 U11788 ( .IN1(n5389), .IN2(n11599), .Q(n11608) );
  OR2X1 U11789 ( .IN1(n11609), .IN2(n11610), .Q(g33053) );
  AND2X1 U11790 ( .IN1(n9166), .IN2(g5517), .Q(n11610) );
  AND3X1 U11791 ( .IN1(n11599), .IN2(n11611), .IN3(n5647), .Q(n11609) );
  INVX0 U11792 ( .INP(n528), .ZN(n11611) );
  OR2X1 U11793 ( .IN1(n11612), .IN2(n11613), .Q(g33052) );
  AND2X1 U11794 ( .IN1(n9166), .IN2(g5511), .Q(n11613) );
  AND2X1 U11795 ( .IN1(n11614), .IN2(n11599), .Q(n11612) );
  INVX0 U11796 ( .INP(n11615), .ZN(n11614) );
  AND2X1 U11797 ( .IN1(n11616), .IN2(n3437), .Q(n11615) );
  OR2X1 U11798 ( .IN1(n9124), .IN2(n3436), .Q(n11616) );
  OR2X1 U11799 ( .IN1(n11617), .IN2(n11618), .Q(g33050) );
  AND2X1 U11800 ( .IN1(n9166), .IN2(g5180), .Q(n11618) );
  AND2X1 U11801 ( .IN1(n11619), .IN2(n11620), .Q(n11617) );
  OR3X1 U11802 ( .IN1(n11621), .IN2(n11622), .IN3(n11623), .Q(n11619) );
  AND2X1 U11803 ( .IN1(g25700), .IN2(n5650), .Q(n11623) );
  AND2X1 U11804 ( .IN1(n9035), .IN2(n11624), .Q(n11622) );
  OR2X1 U11805 ( .IN1(n11625), .IN2(n11626), .Q(g33049) );
  AND2X1 U11806 ( .IN1(n11627), .IN2(g5180), .Q(n11626) );
  AND2X1 U11807 ( .IN1(n11628), .IN2(g5176), .Q(n11625) );
  OR2X1 U11808 ( .IN1(n9124), .IN2(n11629), .Q(n11628) );
  AND2X1 U11809 ( .IN1(n5384), .IN2(n11620), .Q(n11629) );
  OR2X1 U11810 ( .IN1(n11630), .IN2(n11631), .Q(g33048) );
  AND2X1 U11811 ( .IN1(n9167), .IN2(g5170), .Q(n11631) );
  AND3X1 U11812 ( .IN1(n11620), .IN2(n11632), .IN3(n5650), .Q(n11630) );
  INVX0 U11813 ( .INP(n764), .ZN(n11632) );
  OR2X1 U11814 ( .IN1(n11633), .IN2(n11634), .Q(g33047) );
  AND2X1 U11815 ( .IN1(n9167), .IN2(g5164), .Q(n11634) );
  AND2X1 U11816 ( .IN1(n11635), .IN2(n11620), .Q(n11633) );
  INVX0 U11817 ( .INP(n11636), .ZN(n11635) );
  AND2X1 U11818 ( .IN1(n11637), .IN2(n3447), .Q(n11636) );
  OR2X1 U11819 ( .IN1(n9124), .IN2(n3446), .Q(n11637) );
  OR3X1 U11820 ( .IN1(n11638), .IN2(n11639), .IN3(n11640), .Q(g33046) );
  AND2X1 U11821 ( .IN1(n9167), .IN2(g5052), .Q(n11640) );
  AND3X1 U11822 ( .IN1(n11641), .IN2(n11642), .IN3(g5057), .Q(n11639) );
  INVX0 U11823 ( .INP(n11643), .ZN(n11642) );
  AND2X1 U11824 ( .IN1(n5615), .IN2(n11644), .Q(n11638) );
  OR2X1 U11825 ( .IN1(n11643), .IN2(n11645), .Q(n11644) );
  AND2X1 U11826 ( .IN1(g5052), .IN2(n11646), .Q(n11643) );
  OR3X1 U11827 ( .IN1(n11647), .IN2(n11648), .IN3(n11649), .Q(g33045) );
  AND2X1 U11828 ( .IN1(n11650), .IN2(g4567), .Q(n11649) );
  OR3X1 U11829 ( .IN1(n11651), .IN2(n11652), .IN3(n11648), .Q(g33044) );
  AND2X1 U11830 ( .IN1(test_so93), .IN2(n11650), .Q(n11651) );
  OR3X1 U11831 ( .IN1(n11653), .IN2(n11654), .IN3(n11655), .Q(g33043) );
  AND2X1 U11832 ( .IN1(test_so16), .IN2(n11650), .Q(n11655) );
  OR3X1 U11833 ( .IN1(n11653), .IN2(n11648), .IN3(n11656), .Q(g33042) );
  AND2X1 U11834 ( .IN1(n11650), .IN2(g4540), .Q(n11656) );
  INVX0 U11835 ( .INP(n11657), .ZN(n11648) );
  OR2X1 U11836 ( .IN1(n8775), .IN2(n11650), .Q(n11657) );
  OR3X1 U11837 ( .IN1(n11647), .IN2(n11654), .IN3(n11658), .Q(g33041) );
  AND2X1 U11838 ( .IN1(test_so56), .IN2(n11650), .Q(n11658) );
  OR3X1 U11839 ( .IN1(n11659), .IN2(n11652), .IN3(n11660), .Q(g33040) );
  AND2X1 U11840 ( .IN1(n11661), .IN2(n9802), .Q(n11652) );
  OR2X1 U11841 ( .IN1(g72), .IN2(g73), .Q(n9802) );
  AND2X1 U11842 ( .IN1(n11650), .IN2(g4504), .Q(n11659) );
  OR3X1 U11843 ( .IN1(n11647), .IN2(n11662), .IN3(n11663), .Q(g33039) );
  AND2X1 U11844 ( .IN1(n11650), .IN2(g4501), .Q(n11663) );
  OR3X1 U11845 ( .IN1(n11647), .IN2(n11660), .IN3(n11664), .Q(g33038) );
  AND2X1 U11846 ( .IN1(n11650), .IN2(g4498), .Q(n11664) );
  AND2X1 U11847 ( .IN1(n11665), .IN2(n11661), .Q(n11647) );
  OR2X1 U11848 ( .IN1(n9476), .IN2(g73), .Q(n11665) );
  OR3X1 U11849 ( .IN1(n11653), .IN2(n11662), .IN3(n11666), .Q(g33037) );
  AND2X1 U11850 ( .IN1(n11650), .IN2(g4495), .Q(n11666) );
  OR3X1 U11851 ( .IN1(n11653), .IN2(n11660), .IN3(n11667), .Q(g33036) );
  AND2X1 U11852 ( .IN1(n11650), .IN2(g4480), .Q(n11667) );
  AND2X1 U11853 ( .IN1(g4572), .IN2(n11661), .Q(n11660) );
  AND2X1 U11854 ( .IN1(n11668), .IN2(n11661), .Q(n11653) );
  OR2X1 U11855 ( .IN1(n9473), .IN2(g72), .Q(n11668) );
  OR4X1 U11856 ( .IN1(n8811), .IN2(n11669), .IN3(n11670), .IN4(n11671), .Q(
        g33035) );
  AND2X1 U11857 ( .IN1(n9167), .IN2(g4098), .Q(n11671) );
  AND3X1 U11858 ( .IN1(n9454), .IN2(g4108), .IN3(n9077), .Q(n11670) );
  AND2X1 U11859 ( .IN1(n9478), .IN2(n5715), .Q(n11669) );
  OR2X1 U11860 ( .IN1(n11672), .IN2(n11673), .Q(g33034) );
  AND2X1 U11861 ( .IN1(n9167), .IN2(g3873), .Q(n11673) );
  AND2X1 U11862 ( .IN1(n11674), .IN2(n11675), .Q(n11672) );
  OR3X1 U11863 ( .IN1(n11676), .IN2(n11677), .IN3(n11678), .Q(n11674) );
  AND2X1 U11864 ( .IN1(g25676), .IN2(n8823), .Q(n11678) );
  AND2X1 U11865 ( .IN1(n9035), .IN2(n11679), .Q(n11677) );
  OR2X1 U11866 ( .IN1(n11680), .IN2(n11681), .Q(g33033) );
  AND2X1 U11867 ( .IN1(n11682), .IN2(g3873), .Q(n11681) );
  AND2X1 U11868 ( .IN1(test_so33), .IN2(n11683), .Q(n11680) );
  OR2X1 U11869 ( .IN1(n9136), .IN2(n11684), .Q(n11683) );
  AND2X1 U11870 ( .IN1(n5387), .IN2(n11675), .Q(n11684) );
  OR2X1 U11871 ( .IN1(n11685), .IN2(n11686), .Q(g33032) );
  AND2X1 U11872 ( .IN1(n9167), .IN2(g3863), .Q(n11686) );
  AND3X1 U11873 ( .IN1(n11687), .IN2(n8823), .IN3(n11675), .Q(n11685) );
  INVX0 U11874 ( .INP(n1151), .ZN(n11687) );
  OR2X1 U11875 ( .IN1(n11688), .IN2(n11689), .Q(g33031) );
  AND2X1 U11876 ( .IN1(n9167), .IN2(g3857), .Q(n11689) );
  AND2X1 U11877 ( .IN1(n11690), .IN2(n11675), .Q(n11688) );
  INVX0 U11878 ( .INP(n11691), .ZN(n11690) );
  AND2X1 U11879 ( .IN1(n11692), .IN2(n3482), .Q(n11691) );
  OR2X1 U11880 ( .IN1(n9135), .IN2(n3481), .Q(n11692) );
  OR2X1 U11881 ( .IN1(n11693), .IN2(n11694), .Q(g33029) );
  AND2X1 U11882 ( .IN1(n9167), .IN2(g3522), .Q(n11694) );
  AND2X1 U11883 ( .IN1(n11695), .IN2(n11696), .Q(n11693) );
  OR3X1 U11884 ( .IN1(n11697), .IN2(n11698), .IN3(n11699), .Q(n11695) );
  AND2X1 U11885 ( .IN1(g25662), .IN2(n5645), .Q(n11699) );
  AND2X1 U11886 ( .IN1(n9035), .IN2(n11700), .Q(n11698) );
  OR2X1 U11887 ( .IN1(n11701), .IN2(n11702), .Q(g33028) );
  AND2X1 U11888 ( .IN1(n11703), .IN2(g3522), .Q(n11702) );
  AND2X1 U11889 ( .IN1(n11704), .IN2(g3518), .Q(n11701) );
  OR2X1 U11890 ( .IN1(n9135), .IN2(n11705), .Q(n11704) );
  AND2X1 U11891 ( .IN1(n5383), .IN2(n11696), .Q(n11705) );
  OR2X1 U11892 ( .IN1(n11706), .IN2(n11707), .Q(g33027) );
  AND2X1 U11893 ( .IN1(n9167), .IN2(g3512), .Q(n11707) );
  AND3X1 U11894 ( .IN1(n11696), .IN2(n11708), .IN3(n5645), .Q(n11706) );
  INVX0 U11895 ( .INP(n115), .ZN(n11708) );
  OR2X1 U11896 ( .IN1(n11709), .IN2(n11710), .Q(g33026) );
  AND2X1 U11897 ( .IN1(n9167), .IN2(g3506), .Q(n11710) );
  AND2X1 U11898 ( .IN1(n11711), .IN2(n11696), .Q(n11709) );
  INVX0 U11899 ( .INP(n11712), .ZN(n11711) );
  AND2X1 U11900 ( .IN1(n11713), .IN2(n3492), .Q(n11712) );
  OR2X1 U11901 ( .IN1(n9135), .IN2(n3491), .Q(n11713) );
  OR3X1 U11902 ( .IN1(n11714), .IN2(n11715), .IN3(n11716), .Q(g33024) );
  AND2X1 U11903 ( .IN1(g25648), .IN2(n11717), .Q(n11716) );
  AND3X1 U11904 ( .IN1(n11718), .IN2(n11719), .IN3(n9077), .Q(n11715) );
  OR2X1 U11905 ( .IN1(n11720), .IN2(n11721), .Q(n11718) );
  AND2X1 U11906 ( .IN1(n9167), .IN2(g3171), .Q(n11714) );
  OR2X1 U11907 ( .IN1(n11722), .IN2(n11723), .Q(g33023) );
  AND2X1 U11908 ( .IN1(n11724), .IN2(g3167), .Q(n11723) );
  OR2X1 U11909 ( .IN1(n9135), .IN2(n11725), .Q(n11724) );
  AND2X1 U11910 ( .IN1(n5603), .IN2(n11719), .Q(n11725) );
  AND3X1 U11911 ( .IN1(n9054), .IN2(g3171), .IN3(n11717), .Q(n11722) );
  OR2X1 U11912 ( .IN1(n11726), .IN2(n11727), .Q(g33022) );
  AND2X1 U11913 ( .IN1(n9167), .IN2(g3161), .Q(n11727) );
  AND2X1 U11914 ( .IN1(n11717), .IN2(n11728), .Q(n11726) );
  INVX0 U11915 ( .INP(n130), .ZN(n11728) );
  OR2X1 U11916 ( .IN1(n11729), .IN2(n11730), .Q(g33021) );
  AND2X1 U11917 ( .IN1(n9167), .IN2(g3155), .Q(n11730) );
  AND2X1 U11918 ( .IN1(n11731), .IN2(n11719), .Q(n11729) );
  INVX0 U11919 ( .INP(n11732), .ZN(n11731) );
  AND2X1 U11920 ( .IN1(n11733), .IN2(n3501), .Q(n11732) );
  OR2X1 U11921 ( .IN1(n9134), .IN2(n3502), .Q(n11733) );
  OR3X1 U11922 ( .IN1(n11734), .IN2(n11735), .IN3(n2787), .Q(g33019) );
  AND2X1 U11923 ( .IN1(n11736), .IN2(n9021), .Q(n11735) );
  OR2X1 U11924 ( .IN1(n11737), .IN2(n11738), .Q(n11736) );
  AND2X1 U11925 ( .IN1(n2790), .IN2(n5300), .Q(n11738) );
  AND2X1 U11926 ( .IN1(test_so30), .IN2(n11739), .Q(n11737) );
  INVX0 U11927 ( .INP(n2790), .ZN(n11739) );
  AND2X1 U11928 ( .IN1(n9167), .IN2(g2748), .Q(n11734) );
  OR4X1 U11929 ( .IN1(n11740), .IN2(n11741), .IN3(n11742), .IN4(n11743), .Q(
        g33018) );
  AND4X1 U11930 ( .IN1(n3511), .IN2(n11744), .IN3(n11745), .IN4(n8772), .Q(
        n11743) );
  AND2X1 U11931 ( .IN1(n10147), .IN2(g2619), .Q(n11745) );
  AND2X1 U11932 ( .IN1(n9167), .IN2(g2610), .Q(n11742) );
  AND2X1 U11933 ( .IN1(test_so40), .IN2(n11746), .Q(n11741) );
  OR3X1 U11934 ( .IN1(n11312), .IN2(n11747), .IN3(n11748), .Q(n11746) );
  AND2X1 U11935 ( .IN1(n1370), .IN2(n9022), .Q(n11748) );
  INVX0 U11936 ( .INP(n10392), .ZN(n1370) );
  AND3X1 U11937 ( .IN1(n3512), .IN2(n9507), .IN3(n3517), .Q(n11740) );
  AND2X1 U11938 ( .IN1(n10392), .IN2(n3524), .Q(n9507) );
  AND2X1 U11939 ( .IN1(n3505), .IN2(n3525), .Q(n10392) );
  OR3X1 U11940 ( .IN1(n8800), .IN2(n5508), .IN3(g2610), .Q(n3512) );
  OR4X1 U11941 ( .IN1(n11749), .IN2(n11750), .IN3(n3519), .IN4(n11751), .Q(
        g33017) );
  AND2X1 U11942 ( .IN1(n11747), .IN2(g2619), .Q(n11751) );
  AND2X1 U11943 ( .IN1(test_so40), .IN2(n9137), .Q(n11750) );
  AND2X1 U11944 ( .IN1(n3517), .IN2(g2610), .Q(n11749) );
  OR3X1 U11945 ( .IN1(n11752), .IN2(n11753), .IN3(n3519), .Q(g33016) );
  INVX0 U11946 ( .INP(n11754), .ZN(n11753) );
  OR2X1 U11947 ( .IN1(n11747), .IN2(n5372), .Q(n11754) );
  AND2X1 U11948 ( .IN1(n11747), .IN2(g2610), .Q(n11752) );
  OR4X1 U11949 ( .IN1(n11755), .IN2(n11756), .IN3(n3519), .IN4(n11757), .Q(
        g33015) );
  AND3X1 U11950 ( .IN1(n5508), .IN2(n11758), .IN3(n3517), .Q(n11757) );
  AND2X1 U11951 ( .IN1(test_so34), .IN2(n9138), .Q(n11756) );
  AND2X1 U11952 ( .IN1(n11747), .IN2(g2587), .Q(n11755) );
  OR4X1 U11953 ( .IN1(n11759), .IN2(n11760), .IN3(n11761), .IN4(n11762), .Q(
        g33014) );
  AND4X1 U11954 ( .IN1(n3530), .IN2(n11763), .IN3(n11764), .IN4(n8773), .Q(
        n11762) );
  AND2X1 U11955 ( .IN1(n10147), .IN2(g2485), .Q(n11764) );
  AND2X1 U11956 ( .IN1(n9167), .IN2(g2476), .Q(n11761) );
  AND2X1 U11957 ( .IN1(n11765), .IN2(g2491), .Q(n11760) );
  OR3X1 U11958 ( .IN1(n11312), .IN2(n11766), .IN3(n11767), .Q(n11765) );
  AND2X1 U11959 ( .IN1(n1372), .IN2(n9022), .Q(n11767) );
  INVX0 U11960 ( .INP(n10401), .ZN(n1372) );
  AND3X1 U11961 ( .IN1(n3531), .IN2(n9506), .IN3(n3536), .Q(n11759) );
  AND2X1 U11962 ( .IN1(n10401), .IN2(n3524), .Q(n9506) );
  AND3X1 U11963 ( .IN1(g2748), .IN2(n5349), .IN3(n3525), .Q(n10401) );
  OR3X1 U11964 ( .IN1(n8800), .IN2(n5509), .IN3(g2476), .Q(n3531) );
  OR4X1 U11965 ( .IN1(n11768), .IN2(n11769), .IN3(n3538), .IN4(n11770), .Q(
        g33013) );
  AND2X1 U11966 ( .IN1(n11766), .IN2(g2485), .Q(n11770) );
  AND2X1 U11967 ( .IN1(n9167), .IN2(g2491), .Q(n11769) );
  AND2X1 U11968 ( .IN1(n3536), .IN2(g2476), .Q(n11768) );
  OR3X1 U11969 ( .IN1(n11771), .IN2(n11772), .IN3(n3538), .Q(g33012) );
  INVX0 U11970 ( .INP(n11773), .ZN(n11772) );
  OR2X1 U11971 ( .IN1(n11766), .IN2(n5373), .Q(n11773) );
  AND2X1 U11972 ( .IN1(n11766), .IN2(g2476), .Q(n11771) );
  OR4X1 U11973 ( .IN1(n11774), .IN2(n11775), .IN3(n3538), .IN4(n11776), .Q(
        g33011) );
  AND3X1 U11974 ( .IN1(n5509), .IN2(n11777), .IN3(n3536), .Q(n11776) );
  AND2X1 U11975 ( .IN1(n9167), .IN2(g2461), .Q(n11775) );
  AND2X1 U11976 ( .IN1(n11766), .IN2(g2453), .Q(n11774) );
  OR4X1 U11977 ( .IN1(n11778), .IN2(n11779), .IN3(n11780), .IN4(n11781), .Q(
        g33010) );
  AND4X1 U11978 ( .IN1(n3548), .IN2(n11782), .IN3(n11783), .IN4(n8830), .Q(
        n11781) );
  AND2X1 U11979 ( .IN1(n10147), .IN2(g2351), .Q(n11783) );
  AND2X1 U11980 ( .IN1(test_so21), .IN2(n9137), .Q(n11780) );
  AND2X1 U11981 ( .IN1(n11784), .IN2(g2357), .Q(n11779) );
  OR3X1 U11982 ( .IN1(n11312), .IN2(n11785), .IN3(n11786), .Q(n11784) );
  AND2X1 U11983 ( .IN1(n1366), .IN2(n9022), .Q(n11786) );
  INVX0 U11984 ( .INP(n10400), .ZN(n1366) );
  AND3X1 U11985 ( .IN1(n3549), .IN2(n9509), .IN3(n3555), .Q(n11778) );
  AND2X1 U11986 ( .IN1(n10400), .IN2(n3524), .Q(n9509) );
  AND3X1 U11987 ( .IN1(g2741), .IN2(n5516), .IN3(n3525), .Q(n10400) );
  OR3X1 U11988 ( .IN1(test_so21), .IN2(n8800), .IN3(n5511), .Q(n3549) );
  OR4X1 U11989 ( .IN1(n11787), .IN2(n11788), .IN3(n3557), .IN4(n11789), .Q(
        g33009) );
  AND2X1 U11990 ( .IN1(n11785), .IN2(g2351), .Q(n11789) );
  AND2X1 U11991 ( .IN1(n9167), .IN2(g2357), .Q(n11788) );
  AND2X1 U11992 ( .IN1(n3555), .IN2(test_so21), .Q(n11787) );
  OR3X1 U11993 ( .IN1(n11790), .IN2(n11791), .IN3(n3557), .Q(g33008) );
  INVX0 U11994 ( .INP(n11792), .ZN(n11791) );
  OR2X1 U11995 ( .IN1(n11785), .IN2(n5375), .Q(n11792) );
  AND2X1 U11996 ( .IN1(n11785), .IN2(test_so21), .Q(n11790) );
  OR4X1 U11997 ( .IN1(n11793), .IN2(n11794), .IN3(n3557), .IN4(n11795), .Q(
        g33007) );
  AND3X1 U11998 ( .IN1(n5511), .IN2(n11796), .IN3(n3555), .Q(n11795) );
  AND2X1 U11999 ( .IN1(n9167), .IN2(g2327), .Q(n11794) );
  AND2X1 U12000 ( .IN1(n11785), .IN2(g2319), .Q(n11793) );
  OR4X1 U12001 ( .IN1(n11797), .IN2(n11798), .IN3(n11799), .IN4(n11800), .Q(
        g33006) );
  AND4X1 U12002 ( .IN1(n3567), .IN2(n11801), .IN3(n11802), .IN4(n8721), .Q(
        n11800) );
  AND2X1 U12003 ( .IN1(n10147), .IN2(g2217), .Q(n11802) );
  AND2X1 U12004 ( .IN1(n9167), .IN2(g2208), .Q(n11799) );
  AND2X1 U12005 ( .IN1(n11803), .IN2(g2223), .Q(n11798) );
  OR3X1 U12006 ( .IN1(n11312), .IN2(n11804), .IN3(n11805), .Q(n11803) );
  AND2X1 U12007 ( .IN1(n1368), .IN2(n9023), .Q(n11805) );
  INVX0 U12008 ( .INP(n10403), .ZN(n1368) );
  AND3X1 U12009 ( .IN1(n3568), .IN2(n9508), .IN3(n3574), .Q(n11797) );
  AND2X1 U12010 ( .IN1(n10403), .IN2(n3524), .Q(n9508) );
  AND3X1 U12011 ( .IN1(n5516), .IN2(n5349), .IN3(n3525), .Q(n10403) );
  OR3X1 U12012 ( .IN1(n8800), .IN2(n5512), .IN3(g2208), .Q(n3568) );
  OR4X1 U12013 ( .IN1(n11806), .IN2(n11807), .IN3(n3576), .IN4(n11808), .Q(
        g33005) );
  AND2X1 U12014 ( .IN1(n11804), .IN2(g2217), .Q(n11808) );
  AND2X1 U12015 ( .IN1(n9167), .IN2(g2223), .Q(n11807) );
  AND2X1 U12016 ( .IN1(n3574), .IN2(g2208), .Q(n11806) );
  OR3X1 U12017 ( .IN1(n11809), .IN2(n11810), .IN3(n3576), .Q(g33004) );
  INVX0 U12018 ( .INP(n11811), .ZN(n11810) );
  OR2X1 U12019 ( .IN1(n11804), .IN2(n5376), .Q(n11811) );
  AND2X1 U12020 ( .IN1(n11804), .IN2(g2208), .Q(n11809) );
  OR4X1 U12021 ( .IN1(n11812), .IN2(n11813), .IN3(n3576), .IN4(n11814), .Q(
        g33003) );
  AND3X1 U12022 ( .IN1(n5512), .IN2(n11815), .IN3(n3574), .Q(n11814) );
  AND2X1 U12023 ( .IN1(n9168), .IN2(g2193), .Q(n11813) );
  AND2X1 U12024 ( .IN1(n11804), .IN2(g2185), .Q(n11812) );
  OR4X1 U12025 ( .IN1(n11816), .IN2(n11817), .IN3(n11818), .IN4(n11819), .Q(
        g33002) );
  AND4X1 U12026 ( .IN1(n3586), .IN2(n11820), .IN3(n11821), .IN4(n8778), .Q(
        n11819) );
  AND2X1 U12027 ( .IN1(n10147), .IN2(g2060), .Q(n11821) );
  AND2X1 U12028 ( .IN1(n9168), .IN2(g2051), .Q(n11818) );
  AND2X1 U12029 ( .IN1(n11822), .IN2(g2066), .Q(n11817) );
  OR3X1 U12030 ( .IN1(n11312), .IN2(n11823), .IN3(n11824), .Q(n11822) );
  AND2X1 U12031 ( .IN1(n790), .IN2(n9023), .Q(n11824) );
  INVX0 U12032 ( .INP(n10395), .ZN(n790) );
  AND3X1 U12033 ( .IN1(n3587), .IN2(n9343), .IN3(n3593), .Q(n11816) );
  AND2X1 U12034 ( .IN1(n10395), .IN2(n3524), .Q(n9343) );
  AND3X1 U12035 ( .IN1(n5300), .IN2(n822), .IN3(n3505), .Q(n10395) );
  OR3X1 U12036 ( .IN1(n8800), .IN2(n5507), .IN3(g2051), .Q(n3587) );
  OR4X1 U12037 ( .IN1(n11825), .IN2(n11826), .IN3(n3595), .IN4(n11827), .Q(
        g33001) );
  AND2X1 U12038 ( .IN1(n11823), .IN2(g2060), .Q(n11827) );
  AND2X1 U12039 ( .IN1(n9168), .IN2(g2066), .Q(n11826) );
  AND2X1 U12040 ( .IN1(n3593), .IN2(g2051), .Q(n11825) );
  OR3X1 U12041 ( .IN1(n11828), .IN2(n11829), .IN3(n3595), .Q(g33000) );
  INVX0 U12042 ( .INP(n11830), .ZN(n11829) );
  OR2X1 U12043 ( .IN1(n11823), .IN2(n5371), .Q(n11830) );
  AND2X1 U12044 ( .IN1(n11823), .IN2(g2051), .Q(n11828) );
  OR4X1 U12045 ( .IN1(n11831), .IN2(n11832), .IN3(n3595), .IN4(n11833), .Q(
        g32999) );
  AND3X1 U12046 ( .IN1(n5507), .IN2(n11834), .IN3(n3593), .Q(n11833) );
  AND2X1 U12047 ( .IN1(test_so59), .IN2(n9138), .Q(n11832) );
  AND2X1 U12048 ( .IN1(n11823), .IN2(g2028), .Q(n11831) );
  OR4X1 U12049 ( .IN1(n11835), .IN2(n11836), .IN3(n11837), .IN4(n11838), .Q(
        g32998) );
  AND4X1 U12050 ( .IN1(n3604), .IN2(n11839), .IN3(n11840), .IN4(n8779), .Q(
        n11838) );
  AND2X1 U12051 ( .IN1(n10147), .IN2(g1926), .Q(n11840) );
  AND2X1 U12052 ( .IN1(n9168), .IN2(g1917), .Q(n11837) );
  AND2X1 U12053 ( .IN1(n11841), .IN2(g1932), .Q(n11836) );
  OR3X1 U12054 ( .IN1(n11312), .IN2(n11842), .IN3(n11843), .Q(n11841) );
  AND2X1 U12055 ( .IN1(n788), .IN2(n9023), .Q(n11843) );
  AND3X1 U12056 ( .IN1(n3605), .IN2(n9344), .IN3(n3611), .Q(n11835) );
  AND2X1 U12057 ( .IN1(n10402), .IN2(n3524), .Q(n9344) );
  INVX0 U12058 ( .INP(n788), .ZN(n10402) );
  OR4X1 U12059 ( .IN1(g2741), .IN2(n11844), .IN3(test_so30), .IN4(n5516), .Q(
        n788) );
  OR3X1 U12060 ( .IN1(n8800), .IN2(n5510), .IN3(g1917), .Q(n3605) );
  OR4X1 U12061 ( .IN1(n11845), .IN2(n11846), .IN3(n3613), .IN4(n11847), .Q(
        g32997) );
  AND2X1 U12062 ( .IN1(n11842), .IN2(g1926), .Q(n11847) );
  AND2X1 U12063 ( .IN1(n9168), .IN2(g1932), .Q(n11846) );
  AND2X1 U12064 ( .IN1(n3611), .IN2(g1917), .Q(n11845) );
  OR3X1 U12065 ( .IN1(n11848), .IN2(n11849), .IN3(n3613), .Q(g32996) );
  INVX0 U12066 ( .INP(n11850), .ZN(n11849) );
  OR2X1 U12067 ( .IN1(n11842), .IN2(n5374), .Q(n11850) );
  AND2X1 U12068 ( .IN1(n11842), .IN2(g1917), .Q(n11848) );
  OR4X1 U12069 ( .IN1(n11851), .IN2(n11852), .IN3(n3613), .IN4(n11853), .Q(
        g32995) );
  AND3X1 U12070 ( .IN1(n5510), .IN2(n11854), .IN3(n3611), .Q(n11853) );
  AND2X1 U12071 ( .IN1(n9168), .IN2(g1902), .Q(n11852) );
  AND2X1 U12072 ( .IN1(n11842), .IN2(g1894), .Q(n11851) );
  OR4X1 U12073 ( .IN1(n11855), .IN2(n11856), .IN3(n11857), .IN4(n11858), .Q(
        g32994) );
  AND4X1 U12074 ( .IN1(n3622), .IN2(n11859), .IN3(n11860), .IN4(n5596), .Q(
        n11858) );
  AND2X1 U12075 ( .IN1(n10147), .IN2(g1792), .Q(n11860) );
  AND2X1 U12076 ( .IN1(n9168), .IN2(g1783), .Q(n11857) );
  AND2X1 U12077 ( .IN1(n11861), .IN2(g1798), .Q(n11856) );
  OR3X1 U12078 ( .IN1(n11312), .IN2(n11862), .IN3(n11863), .Q(n11861) );
  AND2X1 U12079 ( .IN1(n9033), .IN2(n1733), .Q(n11863) );
  INVX0 U12080 ( .INP(n3005), .ZN(n1733) );
  AND3X1 U12081 ( .IN1(n3623), .IN2(n9505), .IN3(n3628), .Q(n11855) );
  AND2X1 U12082 ( .IN1(n3005), .IN2(n3524), .Q(n9505) );
  OR3X1 U12083 ( .IN1(n8800), .IN2(n5359), .IN3(g1783), .Q(n3623) );
  OR4X1 U12084 ( .IN1(n11864), .IN2(n11865), .IN3(n3630), .IN4(n11866), .Q(
        g32993) );
  AND2X1 U12085 ( .IN1(n11862), .IN2(g1792), .Q(n11866) );
  AND2X1 U12086 ( .IN1(n9168), .IN2(g1798), .Q(n11865) );
  AND2X1 U12087 ( .IN1(n3628), .IN2(g1783), .Q(n11864) );
  OR3X1 U12088 ( .IN1(n11867), .IN2(n11868), .IN3(n3630), .Q(g32992) );
  INVX0 U12089 ( .INP(n11869), .ZN(n11868) );
  OR2X1 U12090 ( .IN1(n11862), .IN2(n5602), .Q(n11869) );
  AND2X1 U12091 ( .IN1(n11862), .IN2(g1783), .Q(n11867) );
  OR4X1 U12092 ( .IN1(n11870), .IN2(n11871), .IN3(n3630), .IN4(n11872), .Q(
        g32991) );
  AND3X1 U12093 ( .IN1(n5359), .IN2(n11873), .IN3(n3628), .Q(n11872) );
  AND2X1 U12094 ( .IN1(n9168), .IN2(g1768), .Q(n11871) );
  AND2X1 U12095 ( .IN1(n11862), .IN2(g1760), .Q(n11870) );
  OR4X1 U12096 ( .IN1(n11874), .IN2(n11875), .IN3(n11876), .IN4(n11877), .Q(
        g32990) );
  AND4X1 U12097 ( .IN1(n3640), .IN2(n11878), .IN3(n11879), .IN4(n8831), .Q(
        n11877) );
  AND2X1 U12098 ( .IN1(n10147), .IN2(g1657), .Q(n11879) );
  AND2X1 U12099 ( .IN1(test_so94), .IN2(n9138), .Q(n11876) );
  AND2X1 U12100 ( .IN1(n11880), .IN2(g1664), .Q(n11875) );
  OR3X1 U12101 ( .IN1(n11312), .IN2(n11881), .IN3(n11882), .Q(n11880) );
  AND2X1 U12102 ( .IN1(n794), .IN2(n9023), .Q(n11882) );
  INVX0 U12103 ( .INP(n10393), .ZN(n794) );
  INVX0 U12104 ( .INP(n11149), .ZN(n11312) );
  OR2X1 U12105 ( .IN1(n2760), .IN2(n9122), .Q(n11149) );
  AND3X1 U12106 ( .IN1(n3641), .IN2(n9342), .IN3(n3646), .Q(n11874) );
  AND2X1 U12107 ( .IN1(n10393), .IN2(n3524), .Q(n9342) );
  AND2X1 U12108 ( .IN1(n822), .IN2(n797), .Q(n10393) );
  INVX0 U12109 ( .INP(n11844), .ZN(n822) );
  OR2X1 U12110 ( .IN1(n11883), .IN2(n11884), .Q(n11844) );
  AND2X1 U12111 ( .IN1(n11885), .IN2(n11886), .Q(n11884) );
  OR2X1 U12112 ( .IN1(g72), .IN2(g2759), .Q(n11886) );
  OR2X1 U12113 ( .IN1(n8793), .IN2(n9476), .Q(n11885) );
  AND2X1 U12114 ( .IN1(n11887), .IN2(n11888), .Q(n11883) );
  OR2X1 U12115 ( .IN1(g73), .IN2(g2763), .Q(n11888) );
  OR2X1 U12116 ( .IN1(n8284), .IN2(n9473), .Q(n11887) );
  OR3X1 U12117 ( .IN1(test_so94), .IN2(n8800), .IN3(n5525), .Q(n3641) );
  OR4X1 U12118 ( .IN1(n11889), .IN2(n11890), .IN3(n3648), .IN4(n11891), .Q(
        g32989) );
  AND2X1 U12119 ( .IN1(n11881), .IN2(g1657), .Q(n11891) );
  AND2X1 U12120 ( .IN1(n9168), .IN2(g1664), .Q(n11890) );
  AND2X1 U12121 ( .IN1(n3646), .IN2(test_so94), .Q(n11889) );
  OR3X1 U12122 ( .IN1(n11892), .IN2(n11893), .IN3(n3648), .Q(g32988) );
  INVX0 U12123 ( .INP(n11894), .ZN(n11893) );
  OR2X1 U12124 ( .IN1(n11881), .IN2(n5370), .Q(n11894) );
  AND2X1 U12125 ( .IN1(n11881), .IN2(test_so94), .Q(n11892) );
  OR4X1 U12126 ( .IN1(n11895), .IN2(n11896), .IN3(n3648), .IN4(n11897), .Q(
        g32987) );
  AND3X1 U12127 ( .IN1(n5525), .IN2(n11898), .IN3(n3646), .Q(n11897) );
  AND2X1 U12128 ( .IN1(n9168), .IN2(g1632), .Q(n11896) );
  AND2X1 U12129 ( .IN1(n11881), .IN2(g1624), .Q(n11895) );
  OR3X1 U12130 ( .IN1(n11899), .IN2(n11900), .IN3(n11901), .Q(g32986) );
  AND3X1 U12131 ( .IN1(n11476), .IN2(n8657), .IN3(n11902), .Q(n11901) );
  INVX0 U12132 ( .INP(n11480), .ZN(n11476) );
  AND2X1 U12133 ( .IN1(n9168), .IN2(g1367), .Q(n11900) );
  AND3X1 U12134 ( .IN1(n11480), .IN2(g1373), .IN3(n9078), .Q(n11899) );
  OR2X1 U12135 ( .IN1(n11903), .IN2(n9494), .Q(n11480) );
  AND2X1 U12136 ( .IN1(n8798), .IN2(n11477), .Q(n11903) );
  AND2X1 U12137 ( .IN1(n11904), .IN2(g1274), .Q(g32985) );
  OR2X1 U12138 ( .IN1(n9134), .IN2(n11905), .Q(n11904) );
  AND2X1 U12139 ( .IN1(n11484), .IN2(n9854), .Q(n11905) );
  INVX0 U12140 ( .INP(n11486), .ZN(n11484) );
  OR2X1 U12141 ( .IN1(n5716), .IN2(n11906), .Q(n11486) );
  OR3X1 U12142 ( .IN1(n11907), .IN2(n11908), .IN3(n11909), .Q(g32984) );
  AND2X1 U12143 ( .IN1(n9168), .IN2(g1263), .Q(n11909) );
  AND2X1 U12144 ( .IN1(n5716), .IN2(n3662), .Q(n11908) );
  AND3X1 U12145 ( .IN1(n11485), .IN2(n11906), .IN3(g1270), .Q(n11907) );
  INVX0 U12146 ( .INP(n3662), .ZN(n11906) );
  OR3X1 U12147 ( .IN1(n11910), .IN2(n11911), .IN3(n11912), .Q(g32983) );
  AND3X1 U12148 ( .IN1(n11491), .IN2(n8656), .IN3(n11913), .Q(n11912) );
  INVX0 U12149 ( .INP(n11495), .ZN(n11491) );
  AND2X1 U12150 ( .IN1(n9168), .IN2(g1024), .Q(n11911) );
  AND3X1 U12151 ( .IN1(n11495), .IN2(g1030), .IN3(n9078), .Q(n11910) );
  OR2X1 U12152 ( .IN1(n11914), .IN2(n9371), .Q(n11495) );
  AND2X1 U12153 ( .IN1(n8795), .IN2(n11492), .Q(n11914) );
  AND2X1 U12154 ( .IN1(n11915), .IN2(g930), .Q(g32982) );
  OR2X1 U12155 ( .IN1(n9134), .IN2(n11916), .Q(n11915) );
  AND2X1 U12156 ( .IN1(n11499), .IN2(n9855), .Q(n11916) );
  INVX0 U12157 ( .INP(n11501), .ZN(n11499) );
  OR2X1 U12158 ( .IN1(n5725), .IN2(n11917), .Q(n11501) );
  OR3X1 U12159 ( .IN1(n11918), .IN2(n11919), .IN3(n11920), .Q(g32981) );
  AND2X1 U12160 ( .IN1(n9168), .IN2(g918), .Q(n11920) );
  AND2X1 U12161 ( .IN1(n5725), .IN2(n3671), .Q(n11919) );
  AND3X1 U12162 ( .IN1(n11500), .IN2(n11917), .IN3(g925), .Q(n11918) );
  INVX0 U12163 ( .INP(n3671), .ZN(n11917) );
  AND3X1 U12164 ( .IN1(n11921), .IN2(n11922), .IN3(n9078), .Q(g32980) );
  OR2X1 U12165 ( .IN1(n11923), .IN2(g854), .Q(n11922) );
  INVX0 U12166 ( .INP(n11924), .ZN(n11921) );
  AND2X1 U12167 ( .IN1(n11923), .IN2(n2644), .Q(n11924) );
  INVX0 U12168 ( .INP(n10207), .ZN(n11923) );
  OR4X1 U12169 ( .IN1(n5633), .IN2(g385), .IN3(n8690), .IN4(n8636), .Q(n10207)
         );
  OR3X1 U12170 ( .IN1(n11925), .IN2(n11926), .IN3(n11927), .Q(g32979) );
  AND2X1 U12171 ( .IN1(test_so2), .IN2(n9139), .Q(n11927) );
  AND2X1 U12172 ( .IN1(n3272), .IN2(n5331), .Q(n11926) );
  AND3X1 U12173 ( .IN1(n2404), .IN2(n11928), .IN3(g758), .Q(n11925) );
  INVX0 U12174 ( .INP(n3272), .ZN(n11928) );
  OR3X1 U12175 ( .IN1(n11929), .IN2(n11930), .IN3(n11931), .Q(g32978) );
  AND2X1 U12176 ( .IN1(n9168), .IN2(g582), .Q(n11931) );
  AND2X1 U12177 ( .IN1(n3274), .IN2(n5472), .Q(n11930) );
  AND3X1 U12178 ( .IN1(n2421), .IN2(n11932), .IN3(g590), .Q(n11929) );
  INVX0 U12179 ( .INP(n3274), .ZN(n11932) );
  OR3X1 U12180 ( .IN1(n11933), .IN2(n11934), .IN3(n11935), .Q(g32977) );
  AND2X1 U12181 ( .IN1(test_so51), .IN2(n9139), .Q(n11935) );
  AND2X1 U12182 ( .IN1(n3279), .IN2(n5679), .Q(n11934) );
  AND3X1 U12183 ( .IN1(n8803), .IN2(n11936), .IN3(g291), .Q(n11933) );
  INVX0 U12184 ( .INP(n3279), .ZN(n11936) );
  AND3X1 U12185 ( .IN1(n11937), .IN2(test_so51), .IN3(test_so55), .Q(n3279) );
  OR3X1 U12186 ( .IN1(n11938), .IN2(n11939), .IN3(n11940), .Q(g32976) );
  AND2X1 U12187 ( .IN1(n9168), .IN2(g164), .Q(n11940) );
  AND2X1 U12188 ( .IN1(n3281), .IN2(n5676), .Q(n11939) );
  AND3X1 U12189 ( .IN1(n10380), .IN2(n11941), .IN3(g150), .Q(n11938) );
  INVX0 U12190 ( .INP(n3281), .ZN(n11941) );
  AND4X1 U12191 ( .IN1(n11942), .IN2(n11943), .IN3(n11944), .IN4(n11945), .Q(
        g32185) );
  AND4X1 U12192 ( .IN1(n11946), .IN2(n11947), .IN3(n11948), .IN4(n11949), .Q(
        n11945) );
  OR2X1 U12193 ( .IN1(n8366), .IN2(n8850), .Q(n11949) );
  OR2X1 U12194 ( .IN1(n5750), .IN2(n8521), .Q(n11948) );
  OR2X1 U12195 ( .IN1(n8364), .IN2(n8522), .Q(n11947) );
  OR2X1 U12196 ( .IN1(n8363), .IN2(n8523), .Q(n11946) );
  OR2X1 U12197 ( .IN1(n8365), .IN2(n8851), .Q(n11944) );
  OR2X1 U12198 ( .IN1(n8525), .IN2(n8526), .Q(n11943) );
  OR2X1 U12199 ( .IN1(n8367), .IN2(n8524), .Q(n11942) );
  OR4X1 U12200 ( .IN1(n11950), .IN2(n11951), .IN3(n11952), .IN4(n11953), .Q(
        g31904) );
  AND2X1 U12201 ( .IN1(n8739), .IN2(n11954), .Q(n11953) );
  INVX0 U12202 ( .INP(n11955), .ZN(n11952) );
  OR4X1 U12203 ( .IN1(n11956), .IN2(n11954), .IN3(n11957), .IN4(n8739), .Q(
        n11955) );
  AND2X1 U12204 ( .IN1(n11958), .IN2(n9023), .Q(n11951) );
  AND2X1 U12205 ( .IN1(n9168), .IN2(g5029), .Q(n11950) );
  OR4X1 U12206 ( .IN1(n11645), .IN2(n11959), .IN3(n11960), .IN4(n11961), .Q(
        g31903) );
  AND2X1 U12207 ( .IN1(n11646), .IN2(n5607), .Q(n11961) );
  INVX0 U12208 ( .INP(n11962), .ZN(n11960) );
  OR4X1 U12209 ( .IN1(n11646), .IN2(n11963), .IN3(n11957), .IN4(n5607), .Q(
        n11962) );
  AND2X1 U12210 ( .IN1(g5046), .IN2(n11964), .Q(n11646) );
  AND2X1 U12211 ( .IN1(n9168), .IN2(g5046), .Q(n11959) );
  AND3X1 U12212 ( .IN1(n9055), .IN2(n5607), .IN3(n11963), .Q(n11645) );
  OR3X1 U12213 ( .IN1(n11965), .IN2(n11966), .IN3(n11967), .Q(g31902) );
  AND2X1 U12214 ( .IN1(n11956), .IN2(n9022), .Q(n11967) );
  AND2X1 U12215 ( .IN1(n11968), .IN2(g5016), .Q(n11966) );
  OR2X1 U12216 ( .IN1(n9134), .IN2(n11969), .Q(n11968) );
  AND2X1 U12217 ( .IN1(n5601), .IN2(g5062), .Q(n11969) );
  AND4X1 U12218 ( .IN1(n11641), .IN2(g5029), .IN3(n11970), .IN4(n11971), .Q(
        n11965) );
  OR2X1 U12219 ( .IN1(n8767), .IN2(g5016), .Q(n11971) );
  OR2X1 U12220 ( .IN1(n8768), .IN2(n5369), .Q(n11970) );
  OR4X1 U12221 ( .IN1(n11972), .IN2(n11973), .IN3(n11974), .IN4(n11975), .Q(
        g31901) );
  AND2X1 U12222 ( .IN1(n11964), .IN2(n5578), .Q(n11975) );
  INVX0 U12223 ( .INP(n11976), .ZN(n11974) );
  OR4X1 U12224 ( .IN1(n11977), .IN2(n11964), .IN3(n11957), .IN4(n5578), .Q(
        n11976) );
  INVX0 U12225 ( .INP(n11641), .ZN(n11957) );
  AND3X1 U12226 ( .IN1(g5037), .IN2(g5041), .IN3(n11978), .Q(n11964) );
  AND2X1 U12227 ( .IN1(n11963), .IN2(n9022), .Q(n11973) );
  AND2X1 U12228 ( .IN1(n5578), .IN2(n11977), .Q(n11963) );
  AND3X1 U12229 ( .IN1(n5605), .IN2(n11958), .IN3(n5611), .Q(n11977) );
  AND2X1 U12230 ( .IN1(n9168), .IN2(g5041), .Q(n11972) );
  OR3X1 U12231 ( .IN1(n11979), .IN2(n11980), .IN3(n11981), .Q(g31900) );
  AND2X1 U12232 ( .IN1(n11982), .IN2(n5605), .Q(n11981) );
  AND2X1 U12233 ( .IN1(n11983), .IN2(g5037), .Q(n11980) );
  OR3X1 U12234 ( .IN1(n11984), .IN2(n11985), .IN3(n9122), .Q(n11983) );
  AND2X1 U12235 ( .IN1(n11978), .IN2(n5605), .Q(n11985) );
  AND3X1 U12236 ( .IN1(n11641), .IN2(n11986), .IN3(g5041), .Q(n11984) );
  AND4X1 U12237 ( .IN1(n11987), .IN2(g5041), .IN3(n11641), .IN4(n5611), .Q(
        n11979) );
  OR4X1 U12238 ( .IN1(n11982), .IN2(n11988), .IN3(n11989), .IN4(n11990), .Q(
        g31899) );
  AND2X1 U12239 ( .IN1(n5611), .IN2(n11978), .Q(n11990) );
  AND4X1 U12240 ( .IN1(n11986), .IN2(n11987), .IN3(n11641), .IN4(g5037), .Q(
        n11989) );
  INVX0 U12241 ( .INP(n11958), .ZN(n11987) );
  INVX0 U12242 ( .INP(n11978), .ZN(n11986) );
  AND2X1 U12243 ( .IN1(g5033), .IN2(n11954), .Q(n11978) );
  AND3X1 U12244 ( .IN1(g5062), .IN2(g5029), .IN3(g5016), .Q(n11954) );
  AND2X1 U12245 ( .IN1(n9168), .IN2(g5033), .Q(n11988) );
  AND3X1 U12246 ( .IN1(n9055), .IN2(n11958), .IN3(n5611), .Q(n11982) );
  AND2X1 U12247 ( .IN1(n11956), .IN2(n8739), .Q(n11958) );
  AND3X1 U12248 ( .IN1(g5022), .IN2(n5369), .IN3(n5601), .Q(n11956) );
  OR3X1 U12249 ( .IN1(n11991), .IN2(n11992), .IN3(n11993), .Q(g31898) );
  AND3X1 U12250 ( .IN1(n11641), .IN2(n11994), .IN3(n5369), .Q(n11993) );
  AND4X1 U12251 ( .IN1(n11995), .IN2(n11996), .IN3(n11997), .IN4(n11998), .Q(
        n11641) );
  AND2X1 U12252 ( .IN1(n9033), .IN2(n11999), .Q(n11998) );
  AND2X1 U12253 ( .IN1(n9169), .IN2(g5022), .Q(n11992) );
  AND3X1 U12254 ( .IN1(n12000), .IN2(g5016), .IN3(n9078), .Q(n11991) );
  INVX0 U12255 ( .INP(n11994), .ZN(n12000) );
  OR2X1 U12256 ( .IN1(g5022), .IN2(g5062), .Q(n11994) );
  OR3X1 U12257 ( .IN1(n11654), .IN2(n12001), .IN3(n12002), .Q(g31897) );
  AND2X1 U12258 ( .IN1(n9169), .IN2(g4423), .Q(n12001) );
  AND2X1 U12259 ( .IN1(g4575), .IN2(n11661), .Q(n11654) );
  OR3X1 U12260 ( .IN1(n11662), .IN2(n12003), .IN3(n12002), .Q(g31896) );
  OR2X1 U12261 ( .IN1(n12004), .IN2(n12005), .Q(n12002) );
  AND2X1 U12262 ( .IN1(n11661), .IN2(n12006), .Q(n12005) );
  OR2X1 U12263 ( .IN1(n9473), .IN2(n9476), .Q(n12006) );
  INVX0 U12264 ( .INP(g72), .ZN(n9476) );
  INVX0 U12265 ( .INP(g73), .ZN(n9473) );
  AND3X1 U12266 ( .IN1(n9055), .IN2(g4372), .IN3(n5670), .Q(n12004) );
  INVX0 U12267 ( .INP(n12007), .ZN(n12003) );
  OR2X1 U12268 ( .IN1(n9008), .IN2(n5849), .Q(n12007) );
  AND2X1 U12269 ( .IN1(n11661), .IN2(test_so100), .Q(n11662) );
  INVX0 U12270 ( .INP(n11650), .ZN(n11661) );
  OR2X1 U12271 ( .IN1(n5670), .IN2(n9123), .Q(n11650) );
  OR2X1 U12272 ( .IN1(n12008), .IN2(n10147), .Q(g31895) );
  INVX0 U12273 ( .INP(n10163), .ZN(n10147) );
  OR2X1 U12274 ( .IN1(n9134), .IN2(n1795), .Q(n10163) );
  INVX0 U12275 ( .INP(n2760), .ZN(n1795) );
  AND2X1 U12276 ( .IN1(n9169), .IN2(g4382), .Q(n12008) );
  OR3X1 U12277 ( .IN1(n8811), .IN2(n12009), .IN3(n12010), .Q(g31894) );
  AND2X1 U12278 ( .IN1(n12011), .IN2(g4093), .Q(n12010) );
  OR2X1 U12279 ( .IN1(n9134), .IN2(n12012), .Q(n12011) );
  AND2X1 U12280 ( .IN1(n9454), .IN2(n12013), .Q(n12012) );
  AND3X1 U12281 ( .IN1(n9055), .IN2(g4098), .IN3(n9454), .Q(n12009) );
  INVX0 U12282 ( .INP(n9478), .ZN(n9454) );
  AND3X1 U12283 ( .IN1(g4098), .IN2(g4093), .IN3(n12013), .Q(n9478) );
  OR2X1 U12284 ( .IN1(n12014), .IN2(n12015), .Q(g31872) );
  AND2X1 U12285 ( .IN1(n9169), .IN2(g2741), .Q(n12015) );
  AND3X1 U12286 ( .IN1(n12016), .IN2(n12017), .IN3(n3730), .Q(n12014) );
  OR2X1 U12287 ( .IN1(n12018), .IN2(g2748), .Q(n12017) );
  OR2X1 U12288 ( .IN1(n5516), .IN2(n12019), .Q(n12016) );
  OR3X1 U12289 ( .IN1(n12020), .IN2(n12021), .IN3(n12022), .Q(g31871) );
  AND2X1 U12290 ( .IN1(n3733), .IN2(n11902), .Q(n12022) );
  AND3X1 U12291 ( .IN1(n9494), .IN2(g1367), .IN3(n9079), .Q(n12021) );
  OR2X1 U12292 ( .IN1(n12023), .IN2(n9493), .Q(n9494) );
  AND2X1 U12293 ( .IN1(n8654), .IN2(n11477), .Q(n12023) );
  AND2X1 U12294 ( .IN1(n9169), .IN2(g1361), .Q(n12020) );
  OR3X1 U12295 ( .IN1(n12024), .IN2(n12025), .IN3(n12026), .Q(g31870) );
  AND2X1 U12296 ( .IN1(n9169), .IN2(g1259), .Q(n12026) );
  AND2X1 U12297 ( .IN1(n3664), .IN2(n5674), .Q(n12025) );
  AND3X1 U12298 ( .IN1(n11485), .IN2(n12027), .IN3(g1263), .Q(n12024) );
  INVX0 U12299 ( .INP(n3664), .ZN(n12027) );
  OR3X1 U12300 ( .IN1(n12028), .IN2(n12029), .IN3(n12030), .Q(g31869) );
  AND2X1 U12301 ( .IN1(n3738), .IN2(n11913), .Q(n12030) );
  AND3X1 U12302 ( .IN1(n9371), .IN2(g1024), .IN3(n9078), .Q(n12029) );
  OR2X1 U12303 ( .IN1(n12031), .IN2(n9370), .Q(n9371) );
  AND2X1 U12304 ( .IN1(n8653), .IN2(n11492), .Q(n12031) );
  AND2X1 U12305 ( .IN1(n9169), .IN2(g1018), .Q(n12028) );
  OR3X1 U12306 ( .IN1(n12032), .IN2(n12033), .IN3(n12034), .Q(g31868) );
  AND2X1 U12307 ( .IN1(n9169), .IN2(g914), .Q(n12034) );
  AND2X1 U12308 ( .IN1(n3673), .IN2(n5673), .Q(n12033) );
  AND3X1 U12309 ( .IN1(n11500), .IN2(n12035), .IN3(g918), .Q(n12032) );
  INVX0 U12310 ( .INP(n3673), .ZN(n12035) );
  OR3X1 U12311 ( .IN1(n12036), .IN2(n12037), .IN3(n12038), .Q(g31867) );
  AND2X1 U12312 ( .IN1(n9169), .IN2(g744), .Q(n12038) );
  AND2X1 U12313 ( .IN1(n3682), .IN2(n5471), .Q(n12037) );
  AND3X1 U12314 ( .IN1(n2404), .IN2(test_so2), .IN3(n12039), .Q(n12036) );
  INVX0 U12315 ( .INP(n3682), .ZN(n12039) );
  OR3X1 U12316 ( .IN1(n12040), .IN2(n12041), .IN3(n12042), .Q(g31866) );
  AND2X1 U12317 ( .IN1(n9169), .IN2(g577), .Q(n12042) );
  AND2X1 U12318 ( .IN1(n3684), .IN2(n5552), .Q(n12041) );
  AND3X1 U12319 ( .IN1(n2421), .IN2(n12043), .IN3(g582), .Q(n12040) );
  INVX0 U12320 ( .INP(n3684), .ZN(n12043) );
  OR2X1 U12321 ( .IN1(n12044), .IN2(n12045), .Q(g31865) );
  AND3X1 U12322 ( .IN1(n8803), .IN2(test_so51), .IN3(n8847), .Q(n12045) );
  AND2X1 U12323 ( .IN1(test_so55), .IN2(n12046), .Q(n12044) );
  OR2X1 U12324 ( .IN1(n9134), .IN2(n12047), .Q(n12046) );
  AND2X1 U12325 ( .IN1(n11937), .IN2(n8855), .Q(n12047) );
  OR3X1 U12326 ( .IN1(n12048), .IN2(n12049), .IN3(n12050), .Q(g31864) );
  AND2X1 U12327 ( .IN1(test_so73), .IN2(n9137), .Q(n12050) );
  AND2X1 U12328 ( .IN1(n3687), .IN2(n5561), .Q(n12049) );
  AND3X1 U12329 ( .IN1(n10380), .IN2(n12051), .IN3(g164), .Q(n12048) );
  INVX0 U12330 ( .INP(n3687), .ZN(n12051) );
  AND3X1 U12331 ( .IN1(n12052), .IN2(n12053), .IN3(test_so73), .Q(n3687) );
  AND2X1 U12332 ( .IN1(g1668), .IN2(n5549), .Q(g31862) );
  OR2X1 U12333 ( .IN1(n12054), .IN2(n12055), .Q(g31793) );
  AND3X1 U12334 ( .IN1(n12056), .IN2(n9888), .IN3(n9890), .Q(n12055) );
  OR2X1 U12335 ( .IN1(n12057), .IN2(n12058), .Q(n12056) );
  AND2X1 U12336 ( .IN1(n12059), .IN2(n12060), .Q(n12058) );
  AND3X1 U12337 ( .IN1(n8647), .IN2(n12061), .IN3(n8648), .Q(n12057) );
  OR2X1 U12338 ( .IN1(n12062), .IN2(n12059), .Q(n12061) );
  AND2X1 U12339 ( .IN1(n12063), .IN2(n12060), .Q(n12062) );
  OR2X1 U12340 ( .IN1(n12064), .IN2(n12065), .Q(n12063) );
  AND3X1 U12341 ( .IN1(n12066), .IN2(n12067), .IN3(n12068), .Q(n12064) );
  OR2X1 U12342 ( .IN1(n12069), .IN2(n12070), .Q(n12068) );
  AND2X1 U12343 ( .IN1(n12071), .IN2(n12072), .Q(n12069) );
  OR2X1 U12344 ( .IN1(n12071), .IN2(n12072), .Q(n12066) );
  AND2X1 U12345 ( .IN1(n9889), .IN2(n12073), .Q(n12054) );
  OR2X1 U12346 ( .IN1(n12074), .IN2(n9890), .Q(n12073) );
  AND2X1 U12347 ( .IN1(n9500), .IN2(n12075), .Q(n9890) );
  AND2X1 U12348 ( .IN1(n12076), .IN2(n9888), .Q(n12074) );
  OR2X1 U12349 ( .IN1(n9500), .IN2(n12075), .Q(n12076) );
  OR2X1 U12350 ( .IN1(n8760), .IN2(n9123), .Q(n9500) );
  AND4X1 U12351 ( .IN1(n8647), .IN2(n8648), .IN3(n12060), .IN4(n12059), .Q(
        n9889) );
  AND2X1 U12352 ( .IN1(n12067), .IN2(n12065), .Q(n12059) );
  AND3X1 U12353 ( .IN1(n12070), .IN2(n12072), .IN3(n12071), .Q(n12065) );
  OR2X1 U12354 ( .IN1(n8680), .IN2(n10992), .Q(g31665) );
  OR2X1 U12355 ( .IN1(n5488), .IN2(n10992), .Q(g31656) );
  INVX0 U12356 ( .INP(g113), .ZN(n10992) );
  OR3X1 U12357 ( .IN1(n12077), .IN2(n12078), .IN3(n12079), .Q(g30563) );
  AND2X1 U12358 ( .IN1(n9169), .IN2(g6653), .Q(n12079) );
  AND2X1 U12359 ( .IN1(n3765), .IN2(n10979), .Q(n12078) );
  AND2X1 U12360 ( .IN1(n12080), .IN2(g6657), .Q(n12077) );
  OR3X1 U12361 ( .IN1(n12081), .IN2(n12082), .IN3(n12083), .Q(g30562) );
  AND2X1 U12362 ( .IN1(n12084), .IN2(n3765), .Q(n12083) );
  INVX0 U12363 ( .INP(n12085), .ZN(n12084) );
  AND2X1 U12364 ( .IN1(n9169), .IN2(g6649), .Q(n12082) );
  AND3X1 U12365 ( .IN1(n12085), .IN2(g6605), .IN3(n9079), .Q(n12081) );
  OR2X1 U12366 ( .IN1(n5646), .IN2(n1423), .Q(n12085) );
  OR3X1 U12367 ( .IN1(n12086), .IN2(n12087), .IN3(n12088), .Q(g30561) );
  AND2X1 U12368 ( .IN1(n11537), .IN2(n3765), .Q(n12088) );
  INVX0 U12369 ( .INP(n12089), .ZN(n11537) );
  AND2X1 U12370 ( .IN1(n9169), .IN2(g6645), .Q(n12087) );
  AND3X1 U12371 ( .IN1(n12089), .IN2(g6597), .IN3(n9078), .Q(n12086) );
  OR2X1 U12372 ( .IN1(n5646), .IN2(n1416), .Q(n12089) );
  OR3X1 U12373 ( .IN1(n12090), .IN2(n12091), .IN3(n12092), .Q(g30560) );
  AND2X1 U12374 ( .IN1(n12093), .IN2(n3765), .Q(n12092) );
  INVX0 U12375 ( .INP(n12094), .ZN(n12093) );
  AND2X1 U12376 ( .IN1(n9169), .IN2(g6641), .Q(n12091) );
  AND3X1 U12377 ( .IN1(n12094), .IN2(g6589), .IN3(n9079), .Q(n12090) );
  OR2X1 U12378 ( .IN1(n5646), .IN2(n1418), .Q(n12094) );
  OR3X1 U12379 ( .IN1(n12095), .IN2(n12096), .IN3(n12097), .Q(g30559) );
  AND2X1 U12380 ( .IN1(n3774), .IN2(n12098), .Q(n12097) );
  AND3X1 U12381 ( .IN1(n12099), .IN2(g6653), .IN3(n9078), .Q(n12096) );
  OR2X1 U12382 ( .IN1(n769), .IN2(n1422), .Q(n12099) );
  AND2X1 U12383 ( .IN1(n9169), .IN2(g6637), .Q(n12095) );
  OR3X1 U12384 ( .IN1(n12100), .IN2(n12101), .IN3(n12102), .Q(g30558) );
  AND2X1 U12385 ( .IN1(n3774), .IN2(n11540), .Q(n12102) );
  AND3X1 U12386 ( .IN1(n12103), .IN2(g6649), .IN3(n9079), .Q(n12101) );
  OR2X1 U12387 ( .IN1(n769), .IN2(n1423), .Q(n12103) );
  AND2X1 U12388 ( .IN1(n9169), .IN2(g6633), .Q(n12100) );
  OR3X1 U12389 ( .IN1(n12104), .IN2(n12105), .IN3(n12106), .Q(g30557) );
  AND2X1 U12390 ( .IN1(n3774), .IN2(n12107), .Q(n12106) );
  AND3X1 U12391 ( .IN1(n12108), .IN2(g6645), .IN3(n9078), .Q(n12105) );
  OR2X1 U12392 ( .IN1(n769), .IN2(n1416), .Q(n12108) );
  AND2X1 U12393 ( .IN1(n9169), .IN2(g6629), .Q(n12104) );
  OR3X1 U12394 ( .IN1(n12109), .IN2(n12110), .IN3(n12111), .Q(g30556) );
  AND2X1 U12395 ( .IN1(n3774), .IN2(n12112), .Q(n12111) );
  AND3X1 U12396 ( .IN1(n12113), .IN2(g6641), .IN3(n9080), .Q(n12110) );
  OR2X1 U12397 ( .IN1(n769), .IN2(n1418), .Q(n12113) );
  OR2X1 U12398 ( .IN1(n8643), .IN2(n5571), .Q(n769) );
  AND2X1 U12399 ( .IN1(n9169), .IN2(g6625), .Q(n12109) );
  OR3X1 U12400 ( .IN1(n12114), .IN2(n12115), .IN3(n12116), .Q(g30555) );
  AND2X1 U12401 ( .IN1(n3780), .IN2(n12098), .Q(n12116) );
  AND3X1 U12402 ( .IN1(n12117), .IN2(g6637), .IN3(n9079), .Q(n12115) );
  OR2X1 U12403 ( .IN1(n3406), .IN2(n1422), .Q(n12117) );
  AND2X1 U12404 ( .IN1(n9169), .IN2(g6621), .Q(n12114) );
  OR3X1 U12405 ( .IN1(n12118), .IN2(n12119), .IN3(n12120), .Q(g30554) );
  AND2X1 U12406 ( .IN1(n3780), .IN2(n11540), .Q(n12120) );
  AND3X1 U12407 ( .IN1(n12121), .IN2(g6633), .IN3(n9080), .Q(n12119) );
  OR2X1 U12408 ( .IN1(n3406), .IN2(n1423), .Q(n12121) );
  AND2X1 U12409 ( .IN1(n9169), .IN2(g6617), .Q(n12118) );
  OR3X1 U12410 ( .IN1(n12122), .IN2(n12123), .IN3(n12124), .Q(g30553) );
  AND2X1 U12411 ( .IN1(n3780), .IN2(n12107), .Q(n12124) );
  AND3X1 U12412 ( .IN1(n12125), .IN2(g6629), .IN3(n9079), .Q(n12123) );
  OR2X1 U12413 ( .IN1(n3406), .IN2(n1416), .Q(n12125) );
  AND2X1 U12414 ( .IN1(n9169), .IN2(g6613), .Q(n12122) );
  OR3X1 U12415 ( .IN1(n12126), .IN2(n12127), .IN3(n12128), .Q(g30552) );
  AND2X1 U12416 ( .IN1(n3780), .IN2(n12112), .Q(n12128) );
  AND3X1 U12417 ( .IN1(n12129), .IN2(g6625), .IN3(n9079), .Q(n12127) );
  OR2X1 U12418 ( .IN1(n3406), .IN2(n1418), .Q(n12129) );
  OR2X1 U12419 ( .IN1(n8643), .IN2(g6549), .Q(n3406) );
  AND2X1 U12420 ( .IN1(n9169), .IN2(g6609), .Q(n12126) );
  OR3X1 U12421 ( .IN1(n12130), .IN2(n12131), .IN3(n12132), .Q(g30551) );
  AND2X1 U12422 ( .IN1(n3785), .IN2(n12098), .Q(n12132) );
  AND3X1 U12423 ( .IN1(n12133), .IN2(g6621), .IN3(n9080), .Q(n12131) );
  OR2X1 U12424 ( .IN1(n3407), .IN2(n1422), .Q(n12133) );
  AND2X1 U12425 ( .IN1(n9170), .IN2(g6601), .Q(n12130) );
  OR3X1 U12426 ( .IN1(n12134), .IN2(n12135), .IN3(n12136), .Q(g30550) );
  AND2X1 U12427 ( .IN1(n3785), .IN2(n11540), .Q(n12136) );
  INVX0 U12428 ( .INP(n1423), .ZN(n11540) );
  AND3X1 U12429 ( .IN1(n12137), .IN2(g6617), .IN3(n9078), .Q(n12135) );
  OR2X1 U12430 ( .IN1(n3407), .IN2(n1423), .Q(n12137) );
  OR2X1 U12431 ( .IN1(n5563), .IN2(g6565), .Q(n1423) );
  AND2X1 U12432 ( .IN1(n9170), .IN2(g6593), .Q(n12134) );
  OR3X1 U12433 ( .IN1(n12138), .IN2(n12139), .IN3(n12140), .Q(g30549) );
  AND2X1 U12434 ( .IN1(n3785), .IN2(n12107), .Q(n12140) );
  INVX0 U12435 ( .INP(n1416), .ZN(n12107) );
  AND3X1 U12436 ( .IN1(n12141), .IN2(g6613), .IN3(n9079), .Q(n12139) );
  OR2X1 U12437 ( .IN1(n3407), .IN2(n1416), .Q(n12141) );
  OR2X1 U12438 ( .IN1(n5386), .IN2(g6573), .Q(n1416) );
  AND2X1 U12439 ( .IN1(test_so71), .IN2(n9139), .Q(n12138) );
  OR3X1 U12440 ( .IN1(n12142), .IN2(n12143), .IN3(n12144), .Q(g30548) );
  AND2X1 U12441 ( .IN1(n3785), .IN2(n12112), .Q(n12144) );
  INVX0 U12442 ( .INP(n1418), .ZN(n12112) );
  AND3X1 U12443 ( .IN1(n12145), .IN2(g6609), .IN3(n9080), .Q(n12143) );
  OR2X1 U12444 ( .IN1(n3407), .IN2(n1418), .Q(n12145) );
  OR2X1 U12445 ( .IN1(g6565), .IN2(g6573), .Q(n1418) );
  OR2X1 U12446 ( .IN1(n5571), .IN2(g6555), .Q(n3407) );
  AND2X1 U12447 ( .IN1(n9170), .IN2(g6581), .Q(n12142) );
  OR3X1 U12448 ( .IN1(n12146), .IN2(n12147), .IN3(n12148), .Q(g30547) );
  AND2X1 U12449 ( .IN1(n9170), .IN2(g6605), .Q(n12148) );
  AND2X1 U12450 ( .IN1(n3790), .IN2(n3765), .Q(n12147) );
  AND3X1 U12451 ( .IN1(n9055), .IN2(g6601), .IN3(n12149), .Q(n12146) );
  INVX0 U12452 ( .INP(n3790), .ZN(n12149) );
  OR3X1 U12453 ( .IN1(n12150), .IN2(n12151), .IN3(n12152), .Q(g30546) );
  AND2X1 U12454 ( .IN1(n9170), .IN2(g6597), .Q(n12152) );
  AND2X1 U12455 ( .IN1(n3793), .IN2(n3765), .Q(n12151) );
  AND3X1 U12456 ( .IN1(n9055), .IN2(g6593), .IN3(n12153), .Q(n12150) );
  INVX0 U12457 ( .INP(n3793), .ZN(n12153) );
  OR3X1 U12458 ( .IN1(n12154), .IN2(n12155), .IN3(n12156), .Q(g30545) );
  AND2X1 U12459 ( .IN1(n9170), .IN2(g6589), .Q(n12156) );
  AND2X1 U12460 ( .IN1(n3795), .IN2(n3765), .Q(n12155) );
  AND3X1 U12461 ( .IN1(test_so71), .IN2(n9052), .IN3(n12157), .Q(n12154) );
  INVX0 U12462 ( .INP(n3795), .ZN(n12157) );
  OR3X1 U12463 ( .IN1(n12158), .IN2(n12159), .IN3(n12160), .Q(g30544) );
  AND2X1 U12464 ( .IN1(n9170), .IN2(g6573), .Q(n12160) );
  AND2X1 U12465 ( .IN1(n3797), .IN2(n3765), .Q(n12159) );
  AND3X1 U12466 ( .IN1(n9056), .IN2(g6581), .IN3(n12161), .Q(n12158) );
  INVX0 U12467 ( .INP(n3797), .ZN(n12161) );
  AND2X1 U12468 ( .IN1(n11543), .IN2(n5571), .Q(g30543) );
  AND3X1 U12469 ( .IN1(n9057), .IN2(n11536), .IN3(n5646), .Q(n11543) );
  OR2X1 U12470 ( .IN1(n12162), .IN2(n12163), .Q(n11536) );
  OR3X1 U12471 ( .IN1(n12164), .IN2(n12165), .IN3(n12166), .Q(g30542) );
  AND2X1 U12472 ( .IN1(n9170), .IN2(g6307), .Q(n12166) );
  AND2X1 U12473 ( .IN1(n10991), .IN2(n3765), .Q(n12165) );
  AND2X1 U12474 ( .IN1(n12167), .IN2(g6311), .Q(n12164) );
  OR3X1 U12475 ( .IN1(n12168), .IN2(n12169), .IN3(n12170), .Q(g30541) );
  AND2X1 U12476 ( .IN1(n12171), .IN2(n3765), .Q(n12170) );
  INVX0 U12477 ( .INP(n12172), .ZN(n12171) );
  AND2X1 U12478 ( .IN1(n9170), .IN2(g6303), .Q(n12169) );
  AND3X1 U12479 ( .IN1(n12172), .IN2(g6259), .IN3(n9080), .Q(n12168) );
  OR2X1 U12480 ( .IN1(n5651), .IN2(n55), .Q(n12172) );
  OR3X1 U12481 ( .IN1(n12173), .IN2(n12174), .IN3(n12175), .Q(g30540) );
  AND2X1 U12482 ( .IN1(n11558), .IN2(n3765), .Q(n12175) );
  INVX0 U12483 ( .INP(n12176), .ZN(n11558) );
  AND2X1 U12484 ( .IN1(n9170), .IN2(g6299), .Q(n12174) );
  AND3X1 U12485 ( .IN1(n12176), .IN2(g6251), .IN3(n9080), .Q(n12173) );
  OR2X1 U12486 ( .IN1(n5651), .IN2(n93), .Q(n12176) );
  OR3X1 U12487 ( .IN1(n12177), .IN2(n12178), .IN3(n12179), .Q(g30539) );
  AND2X1 U12488 ( .IN1(n12180), .IN2(n3765), .Q(n12179) );
  INVX0 U12489 ( .INP(n12181), .ZN(n12180) );
  AND2X1 U12490 ( .IN1(n9170), .IN2(g6295), .Q(n12178) );
  AND3X1 U12491 ( .IN1(n12181), .IN2(g6243), .IN3(n9080), .Q(n12177) );
  OR2X1 U12492 ( .IN1(n5651), .IN2(n57), .Q(n12181) );
  OR3X1 U12493 ( .IN1(n12182), .IN2(n12183), .IN3(n12184), .Q(g30538) );
  AND2X1 U12494 ( .IN1(n3808), .IN2(n12185), .Q(n12184) );
  AND3X1 U12495 ( .IN1(n12186), .IN2(g6307), .IN3(n9079), .Q(n12183) );
  OR2X1 U12496 ( .IN1(n92), .IN2(n1022), .Q(n12186) );
  AND2X1 U12497 ( .IN1(n9170), .IN2(g6291), .Q(n12182) );
  OR3X1 U12498 ( .IN1(n12187), .IN2(n12188), .IN3(n12189), .Q(g30537) );
  AND2X1 U12499 ( .IN1(n3808), .IN2(n11561), .Q(n12189) );
  AND3X1 U12500 ( .IN1(n12190), .IN2(g6303), .IN3(n9080), .Q(n12188) );
  OR2X1 U12501 ( .IN1(n55), .IN2(n1022), .Q(n12190) );
  AND2X1 U12502 ( .IN1(n9170), .IN2(g6287), .Q(n12187) );
  OR3X1 U12503 ( .IN1(n12191), .IN2(n12192), .IN3(n12193), .Q(g30536) );
  AND2X1 U12504 ( .IN1(n3808), .IN2(n12194), .Q(n12193) );
  AND3X1 U12505 ( .IN1(n12195), .IN2(g6299), .IN3(n9079), .Q(n12192) );
  OR2X1 U12506 ( .IN1(n93), .IN2(n1022), .Q(n12195) );
  AND2X1 U12507 ( .IN1(n9170), .IN2(g6283), .Q(n12191) );
  OR3X1 U12508 ( .IN1(n12196), .IN2(n12197), .IN3(n12198), .Q(g30535) );
  AND2X1 U12509 ( .IN1(n3808), .IN2(n12199), .Q(n12198) );
  AND3X1 U12510 ( .IN1(n12200), .IN2(g6295), .IN3(n9079), .Q(n12197) );
  OR2X1 U12511 ( .IN1(n57), .IN2(n1022), .Q(n12200) );
  OR2X1 U12512 ( .IN1(n8641), .IN2(n5574), .Q(n1022) );
  AND2X1 U12513 ( .IN1(n9170), .IN2(g6279), .Q(n12196) );
  OR3X1 U12514 ( .IN1(n12201), .IN2(n12202), .IN3(n12203), .Q(g30534) );
  AND2X1 U12515 ( .IN1(n3814), .IN2(n12185), .Q(n12203) );
  AND3X1 U12516 ( .IN1(n12204), .IN2(g6291), .IN3(n9080), .Q(n12202) );
  OR2X1 U12517 ( .IN1(n92), .IN2(n3416), .Q(n12204) );
  AND2X1 U12518 ( .IN1(n9170), .IN2(g6275), .Q(n12201) );
  OR3X1 U12519 ( .IN1(n12205), .IN2(n12206), .IN3(n12207), .Q(g30533) );
  AND2X1 U12520 ( .IN1(n3814), .IN2(n11561), .Q(n12207) );
  AND3X1 U12521 ( .IN1(n12208), .IN2(g6287), .IN3(n9080), .Q(n12206) );
  OR2X1 U12522 ( .IN1(n55), .IN2(n3416), .Q(n12208) );
  AND2X1 U12523 ( .IN1(n9170), .IN2(g6271), .Q(n12205) );
  OR3X1 U12524 ( .IN1(n12209), .IN2(n12210), .IN3(n12211), .Q(g30532) );
  AND2X1 U12525 ( .IN1(n3814), .IN2(n12194), .Q(n12211) );
  AND3X1 U12526 ( .IN1(n12212), .IN2(g6283), .IN3(n9080), .Q(n12210) );
  OR2X1 U12527 ( .IN1(n93), .IN2(n3416), .Q(n12212) );
  AND2X1 U12528 ( .IN1(n9170), .IN2(g6267), .Q(n12209) );
  OR3X1 U12529 ( .IN1(n12213), .IN2(n12214), .IN3(n12215), .Q(g30531) );
  AND2X1 U12530 ( .IN1(n3814), .IN2(n12199), .Q(n12215) );
  AND3X1 U12531 ( .IN1(n12216), .IN2(g6279), .IN3(n9080), .Q(n12214) );
  OR2X1 U12532 ( .IN1(n57), .IN2(n3416), .Q(n12216) );
  OR2X1 U12533 ( .IN1(n8641), .IN2(g6203), .Q(n3416) );
  AND2X1 U12534 ( .IN1(n9170), .IN2(g6263), .Q(n12213) );
  OR3X1 U12535 ( .IN1(n12217), .IN2(n12218), .IN3(n12219), .Q(g30530) );
  AND2X1 U12536 ( .IN1(n3819), .IN2(n12185), .Q(n12219) );
  AND3X1 U12537 ( .IN1(n12220), .IN2(g6275), .IN3(n9079), .Q(n12218) );
  OR2X1 U12538 ( .IN1(n92), .IN2(n3417), .Q(n12220) );
  AND2X1 U12539 ( .IN1(n9170), .IN2(g6255), .Q(n12217) );
  OR3X1 U12540 ( .IN1(n12221), .IN2(n12222), .IN3(n12223), .Q(g30529) );
  AND2X1 U12541 ( .IN1(n3819), .IN2(n11561), .Q(n12223) );
  INVX0 U12542 ( .INP(n55), .ZN(n11561) );
  AND3X1 U12543 ( .IN1(n12224), .IN2(g6271), .IN3(n9073), .Q(n12222) );
  OR2X1 U12544 ( .IN1(n55), .IN2(n3417), .Q(n12224) );
  OR2X1 U12545 ( .IN1(n5568), .IN2(g6219), .Q(n55) );
  AND2X1 U12546 ( .IN1(n9170), .IN2(g6247), .Q(n12221) );
  OR3X1 U12547 ( .IN1(n12225), .IN2(n12226), .IN3(n12227), .Q(g30528) );
  AND2X1 U12548 ( .IN1(n3819), .IN2(n12194), .Q(n12227) );
  INVX0 U12549 ( .INP(n93), .ZN(n12194) );
  AND3X1 U12550 ( .IN1(n12228), .IN2(g6267), .IN3(n9073), .Q(n12226) );
  OR2X1 U12551 ( .IN1(n93), .IN2(n3417), .Q(n12228) );
  OR2X1 U12552 ( .IN1(n5385), .IN2(g6227), .Q(n93) );
  AND2X1 U12553 ( .IN1(n9170), .IN2(g6239), .Q(n12225) );
  OR3X1 U12554 ( .IN1(n12229), .IN2(n12230), .IN3(n12231), .Q(g30527) );
  AND2X1 U12555 ( .IN1(n3819), .IN2(n12199), .Q(n12231) );
  INVX0 U12556 ( .INP(n57), .ZN(n12199) );
  AND3X1 U12557 ( .IN1(n12232), .IN2(g6263), .IN3(n9073), .Q(n12230) );
  OR2X1 U12558 ( .IN1(n57), .IN2(n3417), .Q(n12232) );
  OR2X1 U12559 ( .IN1(n5574), .IN2(g6209), .Q(n3417) );
  OR2X1 U12560 ( .IN1(g6227), .IN2(g6219), .Q(n57) );
  AND2X1 U12561 ( .IN1(n9136), .IN2(g6235), .Q(n12229) );
  OR3X1 U12562 ( .IN1(n12233), .IN2(n12234), .IN3(n12235), .Q(g30526) );
  AND2X1 U12563 ( .IN1(n9136), .IN2(g6259), .Q(n12235) );
  AND2X1 U12564 ( .IN1(n3824), .IN2(n3765), .Q(n12234) );
  AND3X1 U12565 ( .IN1(n9057), .IN2(g6255), .IN3(n12236), .Q(n12233) );
  INVX0 U12566 ( .INP(n3824), .ZN(n12236) );
  OR3X1 U12567 ( .IN1(n12237), .IN2(n12238), .IN3(n12239), .Q(g30525) );
  AND2X1 U12568 ( .IN1(n9163), .IN2(g6251), .Q(n12239) );
  AND2X1 U12569 ( .IN1(n3827), .IN2(n3765), .Q(n12238) );
  AND3X1 U12570 ( .IN1(n9057), .IN2(g6247), .IN3(n12240), .Q(n12237) );
  INVX0 U12571 ( .INP(n3827), .ZN(n12240) );
  OR3X1 U12572 ( .IN1(n12241), .IN2(n12242), .IN3(n12243), .Q(g30524) );
  AND2X1 U12573 ( .IN1(n9161), .IN2(g6243), .Q(n12243) );
  AND2X1 U12574 ( .IN1(n3829), .IN2(n3765), .Q(n12242) );
  AND3X1 U12575 ( .IN1(n9056), .IN2(g6239), .IN3(n12244), .Q(n12241) );
  INVX0 U12576 ( .INP(n3829), .ZN(n12244) );
  OR3X1 U12577 ( .IN1(n12245), .IN2(n12246), .IN3(n12247), .Q(g30523) );
  AND2X1 U12578 ( .IN1(n9161), .IN2(g6227), .Q(n12247) );
  AND2X1 U12579 ( .IN1(n3831), .IN2(n3765), .Q(n12246) );
  AND3X1 U12580 ( .IN1(n9057), .IN2(g6235), .IN3(n12248), .Q(n12245) );
  INVX0 U12581 ( .INP(n3831), .ZN(n12248) );
  AND2X1 U12582 ( .IN1(n11564), .IN2(n5574), .Q(g30522) );
  AND3X1 U12583 ( .IN1(n9056), .IN2(n11557), .IN3(n5651), .Q(n11564) );
  OR3X1 U12584 ( .IN1(n5480), .IN2(n5340), .IN3(n12249), .Q(n11557) );
  OR3X1 U12585 ( .IN1(n12250), .IN2(n12251), .IN3(n12252), .Q(g30521) );
  AND2X1 U12586 ( .IN1(n9161), .IN2(g5961), .Q(n12252) );
  AND2X1 U12587 ( .IN1(n10990), .IN2(n3765), .Q(n12251) );
  AND2X1 U12588 ( .IN1(test_so13), .IN2(n12253), .Q(n12250) );
  OR3X1 U12589 ( .IN1(n12254), .IN2(n12255), .IN3(n12256), .Q(g30520) );
  AND2X1 U12590 ( .IN1(n12257), .IN2(n3765), .Q(n12256) );
  INVX0 U12591 ( .INP(n12258), .ZN(n12257) );
  AND2X1 U12592 ( .IN1(n9161), .IN2(g5957), .Q(n12255) );
  AND3X1 U12593 ( .IN1(n12258), .IN2(g5913), .IN3(n9073), .Q(n12254) );
  OR2X1 U12594 ( .IN1(n5649), .IN2(n729), .Q(n12258) );
  OR3X1 U12595 ( .IN1(n12259), .IN2(n12260), .IN3(n12261), .Q(g30519) );
  AND2X1 U12596 ( .IN1(n11579), .IN2(n3765), .Q(n12261) );
  INVX0 U12597 ( .INP(n12262), .ZN(n11579) );
  AND2X1 U12598 ( .IN1(n9161), .IN2(g5953), .Q(n12260) );
  AND3X1 U12599 ( .IN1(n12262), .IN2(g5905), .IN3(n9073), .Q(n12259) );
  OR2X1 U12600 ( .IN1(n5649), .IN2(n736), .Q(n12262) );
  OR3X1 U12601 ( .IN1(n12263), .IN2(n12264), .IN3(n12265), .Q(g30518) );
  AND2X1 U12602 ( .IN1(n12266), .IN2(n3765), .Q(n12265) );
  INVX0 U12603 ( .INP(n12267), .ZN(n12266) );
  AND2X1 U12604 ( .IN1(n9161), .IN2(g5949), .Q(n12264) );
  AND3X1 U12605 ( .IN1(n12267), .IN2(g5897), .IN3(n9073), .Q(n12263) );
  OR2X1 U12606 ( .IN1(n5649), .IN2(n731), .Q(n12267) );
  OR3X1 U12607 ( .IN1(n12268), .IN2(n12269), .IN3(n12270), .Q(g30517) );
  AND2X1 U12608 ( .IN1(n3842), .IN2(n12271), .Q(n12270) );
  AND3X1 U12609 ( .IN1(n12272), .IN2(g5961), .IN3(n9073), .Q(n12269) );
  OR2X1 U12610 ( .IN1(n735), .IN2(n1084), .Q(n12272) );
  AND2X1 U12611 ( .IN1(n9161), .IN2(g5945), .Q(n12268) );
  OR3X1 U12612 ( .IN1(n12273), .IN2(n12274), .IN3(n12275), .Q(g30516) );
  AND2X1 U12613 ( .IN1(n3842), .IN2(n11582), .Q(n12275) );
  AND3X1 U12614 ( .IN1(n12276), .IN2(g5957), .IN3(n9073), .Q(n12274) );
  OR2X1 U12615 ( .IN1(n729), .IN2(n1084), .Q(n12276) );
  AND2X1 U12616 ( .IN1(n9161), .IN2(g5941), .Q(n12273) );
  OR3X1 U12617 ( .IN1(n12277), .IN2(n12278), .IN3(n12279), .Q(g30515) );
  AND2X1 U12618 ( .IN1(n3842), .IN2(n12280), .Q(n12279) );
  AND3X1 U12619 ( .IN1(n12281), .IN2(g5953), .IN3(n9073), .Q(n12278) );
  OR2X1 U12620 ( .IN1(n736), .IN2(n1084), .Q(n12281) );
  AND2X1 U12621 ( .IN1(n9161), .IN2(g5937), .Q(n12277) );
  OR3X1 U12622 ( .IN1(n12282), .IN2(n12283), .IN3(n12284), .Q(g30514) );
  AND2X1 U12623 ( .IN1(n3842), .IN2(n12285), .Q(n12284) );
  AND3X1 U12624 ( .IN1(n12286), .IN2(g5949), .IN3(n9073), .Q(n12283) );
  OR2X1 U12625 ( .IN1(n731), .IN2(n1084), .Q(n12286) );
  OR2X1 U12626 ( .IN1(n8638), .IN2(n5573), .Q(n1084) );
  AND2X1 U12627 ( .IN1(n9161), .IN2(g5933), .Q(n12282) );
  OR3X1 U12628 ( .IN1(n12287), .IN2(n12288), .IN3(n12289), .Q(g30513) );
  AND2X1 U12629 ( .IN1(n3848), .IN2(n12271), .Q(n12289) );
  AND3X1 U12630 ( .IN1(n12290), .IN2(g5945), .IN3(n9073), .Q(n12288) );
  OR2X1 U12631 ( .IN1(n735), .IN2(n3426), .Q(n12290) );
  AND2X1 U12632 ( .IN1(n9162), .IN2(g5929), .Q(n12287) );
  OR3X1 U12633 ( .IN1(n12291), .IN2(n12292), .IN3(n12293), .Q(g30512) );
  AND2X1 U12634 ( .IN1(n3848), .IN2(n11582), .Q(n12293) );
  AND3X1 U12635 ( .IN1(n12294), .IN2(g5941), .IN3(n9073), .Q(n12292) );
  OR2X1 U12636 ( .IN1(n729), .IN2(n3426), .Q(n12294) );
  AND2X1 U12637 ( .IN1(n9162), .IN2(g5925), .Q(n12291) );
  OR3X1 U12638 ( .IN1(n12295), .IN2(n12296), .IN3(n12297), .Q(g30511) );
  AND2X1 U12639 ( .IN1(n3848), .IN2(n12280), .Q(n12297) );
  AND3X1 U12640 ( .IN1(n12298), .IN2(g5937), .IN3(n9072), .Q(n12296) );
  OR2X1 U12641 ( .IN1(n736), .IN2(n3426), .Q(n12298) );
  AND2X1 U12642 ( .IN1(n9162), .IN2(g5921), .Q(n12295) );
  OR3X1 U12643 ( .IN1(n12299), .IN2(n12300), .IN3(n12301), .Q(g30510) );
  AND2X1 U12644 ( .IN1(n3848), .IN2(n12285), .Q(n12301) );
  AND3X1 U12645 ( .IN1(n12302), .IN2(g5933), .IN3(n9072), .Q(n12300) );
  OR2X1 U12646 ( .IN1(n731), .IN2(n3426), .Q(n12302) );
  OR2X1 U12647 ( .IN1(n8638), .IN2(g5857), .Q(n3426) );
  AND2X1 U12648 ( .IN1(test_so28), .IN2(n9138), .Q(n12299) );
  OR3X1 U12649 ( .IN1(n12303), .IN2(n12304), .IN3(n12305), .Q(g30509) );
  AND2X1 U12650 ( .IN1(n3853), .IN2(n12271), .Q(n12305) );
  AND3X1 U12651 ( .IN1(n12306), .IN2(g5929), .IN3(n9072), .Q(n12304) );
  OR2X1 U12652 ( .IN1(n735), .IN2(n3427), .Q(n12306) );
  AND2X1 U12653 ( .IN1(n9162), .IN2(g5909), .Q(n12303) );
  OR3X1 U12654 ( .IN1(n12307), .IN2(n12308), .IN3(n12309), .Q(g30508) );
  AND2X1 U12655 ( .IN1(n3853), .IN2(n11582), .Q(n12309) );
  INVX0 U12656 ( .INP(n729), .ZN(n11582) );
  AND3X1 U12657 ( .IN1(n12310), .IN2(g5925), .IN3(n9072), .Q(n12308) );
  OR2X1 U12658 ( .IN1(n729), .IN2(n3427), .Q(n12310) );
  OR2X1 U12659 ( .IN1(n8832), .IN2(g5873), .Q(n729) );
  AND2X1 U12660 ( .IN1(n9162), .IN2(g5901), .Q(n12307) );
  OR3X1 U12661 ( .IN1(n12311), .IN2(n12312), .IN3(n12313), .Q(g30507) );
  AND2X1 U12662 ( .IN1(n3853), .IN2(n12280), .Q(n12313) );
  INVX0 U12663 ( .INP(n736), .ZN(n12280) );
  AND3X1 U12664 ( .IN1(n12314), .IN2(g5921), .IN3(n9072), .Q(n12312) );
  OR2X1 U12665 ( .IN1(n736), .IN2(n3427), .Q(n12314) );
  OR2X1 U12666 ( .IN1(test_so36), .IN2(n5388), .Q(n736) );
  AND2X1 U12667 ( .IN1(n9162), .IN2(g5893), .Q(n12311) );
  OR3X1 U12668 ( .IN1(n12315), .IN2(n12316), .IN3(n12317), .Q(g30506) );
  AND2X1 U12669 ( .IN1(n3853), .IN2(n12285), .Q(n12317) );
  INVX0 U12670 ( .INP(n731), .ZN(n12285) );
  AND3X1 U12671 ( .IN1(test_so28), .IN2(n12318), .IN3(n9072), .Q(n12316) );
  OR2X1 U12672 ( .IN1(n731), .IN2(n3427), .Q(n12318) );
  OR2X1 U12673 ( .IN1(n5573), .IN2(g5863), .Q(n3427) );
  OR2X1 U12674 ( .IN1(test_so36), .IN2(g5873), .Q(n731) );
  AND2X1 U12675 ( .IN1(n9162), .IN2(g5889), .Q(n12315) );
  OR3X1 U12676 ( .IN1(n12319), .IN2(n12320), .IN3(n12321), .Q(g30505) );
  AND2X1 U12677 ( .IN1(n9162), .IN2(g5913), .Q(n12321) );
  AND2X1 U12678 ( .IN1(n3858), .IN2(n3765), .Q(n12320) );
  AND3X1 U12679 ( .IN1(n9057), .IN2(g5909), .IN3(n12322), .Q(n12319) );
  INVX0 U12680 ( .INP(n3858), .ZN(n12322) );
  OR3X1 U12681 ( .IN1(n12323), .IN2(n12324), .IN3(n12325), .Q(g30504) );
  AND2X1 U12682 ( .IN1(n9162), .IN2(g5905), .Q(n12325) );
  AND2X1 U12683 ( .IN1(n3861), .IN2(n3765), .Q(n12324) );
  AND3X1 U12684 ( .IN1(n9055), .IN2(g5901), .IN3(n12326), .Q(n12323) );
  INVX0 U12685 ( .INP(n3861), .ZN(n12326) );
  OR3X1 U12686 ( .IN1(n12327), .IN2(n12328), .IN3(n12329), .Q(g30503) );
  AND2X1 U12687 ( .IN1(n9162), .IN2(g5897), .Q(n12329) );
  AND2X1 U12688 ( .IN1(n3863), .IN2(n3765), .Q(n12328) );
  AND3X1 U12689 ( .IN1(n9056), .IN2(g5893), .IN3(n12330), .Q(n12327) );
  INVX0 U12690 ( .INP(n3863), .ZN(n12330) );
  OR3X1 U12691 ( .IN1(n12331), .IN2(n12332), .IN3(n12333), .Q(g30502) );
  AND2X1 U12692 ( .IN1(test_so36), .IN2(n9137), .Q(n12333) );
  AND2X1 U12693 ( .IN1(n3865), .IN2(n3765), .Q(n12332) );
  AND3X1 U12694 ( .IN1(n9057), .IN2(g5889), .IN3(n12334), .Q(n12331) );
  INVX0 U12695 ( .INP(n3865), .ZN(n12334) );
  AND2X1 U12696 ( .IN1(n11585), .IN2(n5573), .Q(g30501) );
  AND3X1 U12697 ( .IN1(n9056), .IN2(n11578), .IN3(n5649), .Q(n11585) );
  OR3X1 U12698 ( .IN1(n5340), .IN2(g4087), .IN3(n12249), .Q(n11578) );
  OR3X1 U12699 ( .IN1(n12335), .IN2(n12336), .IN3(n12337), .Q(g30500) );
  AND2X1 U12700 ( .IN1(n9162), .IN2(g5615), .Q(n12337) );
  AND2X1 U12701 ( .IN1(n3765), .IN2(n10987), .Q(n12336) );
  AND2X1 U12702 ( .IN1(n12338), .IN2(g5619), .Q(n12335) );
  OR3X1 U12703 ( .IN1(n12339), .IN2(n12340), .IN3(n12341), .Q(g30499) );
  AND2X1 U12704 ( .IN1(n12342), .IN2(n3765), .Q(n12341) );
  INVX0 U12705 ( .INP(n12343), .ZN(n12342) );
  AND2X1 U12706 ( .IN1(n9162), .IN2(g5611), .Q(n12340) );
  AND3X1 U12707 ( .IN1(n12343), .IN2(g5567), .IN3(n9072), .Q(n12339) );
  OR2X1 U12708 ( .IN1(n5647), .IN2(n946), .Q(n12343) );
  OR3X1 U12709 ( .IN1(n12344), .IN2(n12345), .IN3(n12346), .Q(g30498) );
  AND2X1 U12710 ( .IN1(n11600), .IN2(n3765), .Q(n12346) );
  INVX0 U12711 ( .INP(n12347), .ZN(n11600) );
  AND2X1 U12712 ( .IN1(n9162), .IN2(g5607), .Q(n12345) );
  AND3X1 U12713 ( .IN1(test_so6), .IN2(n12347), .IN3(n9072), .Q(n12344) );
  OR2X1 U12714 ( .IN1(n5647), .IN2(n943), .Q(n12347) );
  OR3X1 U12715 ( .IN1(n12348), .IN2(n12349), .IN3(n12350), .Q(g30497) );
  AND2X1 U12716 ( .IN1(n12351), .IN2(n3765), .Q(n12350) );
  INVX0 U12717 ( .INP(n12352), .ZN(n12351) );
  AND2X1 U12718 ( .IN1(n9162), .IN2(g5603), .Q(n12349) );
  AND3X1 U12719 ( .IN1(n12352), .IN2(g5551), .IN3(n9072), .Q(n12348) );
  OR2X1 U12720 ( .IN1(n5647), .IN2(n944), .Q(n12352) );
  OR3X1 U12721 ( .IN1(n12353), .IN2(n12354), .IN3(n12355), .Q(g30496) );
  AND2X1 U12722 ( .IN1(n3875), .IN2(n12356), .Q(n12355) );
  AND3X1 U12723 ( .IN1(n12357), .IN2(g5615), .IN3(n9072), .Q(n12354) );
  OR2X1 U12724 ( .IN1(n945), .IN2(n528), .Q(n12357) );
  AND2X1 U12725 ( .IN1(n9162), .IN2(g5599), .Q(n12353) );
  OR3X1 U12726 ( .IN1(n12358), .IN2(n12359), .IN3(n12360), .Q(g30495) );
  AND2X1 U12727 ( .IN1(n3875), .IN2(n11603), .Q(n12360) );
  AND3X1 U12728 ( .IN1(n12361), .IN2(g5611), .IN3(n9072), .Q(n12359) );
  OR2X1 U12729 ( .IN1(n946), .IN2(n528), .Q(n12361) );
  AND2X1 U12730 ( .IN1(n9162), .IN2(g5595), .Q(n12358) );
  OR3X1 U12731 ( .IN1(n12362), .IN2(n12363), .IN3(n12364), .Q(g30494) );
  AND2X1 U12732 ( .IN1(n3875), .IN2(n12365), .Q(n12364) );
  AND3X1 U12733 ( .IN1(n12366), .IN2(g5607), .IN3(n9072), .Q(n12363) );
  OR2X1 U12734 ( .IN1(n943), .IN2(n528), .Q(n12366) );
  AND2X1 U12735 ( .IN1(test_so5), .IN2(n9137), .Q(n12362) );
  OR3X1 U12736 ( .IN1(n12367), .IN2(n12368), .IN3(n12369), .Q(g30493) );
  AND2X1 U12737 ( .IN1(n3875), .IN2(n12370), .Q(n12369) );
  AND3X1 U12738 ( .IN1(n12371), .IN2(g5603), .IN3(n9072), .Q(n12368) );
  OR2X1 U12739 ( .IN1(n944), .IN2(n528), .Q(n12371) );
  OR2X1 U12740 ( .IN1(n8640), .IN2(n5575), .Q(n528) );
  AND2X1 U12741 ( .IN1(n9162), .IN2(g5587), .Q(n12367) );
  OR3X1 U12742 ( .IN1(n12372), .IN2(n12373), .IN3(n12374), .Q(g30492) );
  AND2X1 U12743 ( .IN1(n3881), .IN2(n12356), .Q(n12374) );
  AND3X1 U12744 ( .IN1(n12375), .IN2(g5599), .IN3(n9071), .Q(n12373) );
  OR2X1 U12745 ( .IN1(n945), .IN2(n3436), .Q(n12375) );
  AND2X1 U12746 ( .IN1(n9162), .IN2(g5583), .Q(n12372) );
  OR3X1 U12747 ( .IN1(n12376), .IN2(n12377), .IN3(n12378), .Q(g30491) );
  AND2X1 U12748 ( .IN1(n3881), .IN2(n11603), .Q(n12378) );
  AND3X1 U12749 ( .IN1(n12379), .IN2(g5595), .IN3(n9071), .Q(n12377) );
  OR2X1 U12750 ( .IN1(n946), .IN2(n3436), .Q(n12379) );
  AND2X1 U12751 ( .IN1(n9162), .IN2(g5579), .Q(n12376) );
  OR3X1 U12752 ( .IN1(n12380), .IN2(n12381), .IN3(n12382), .Q(g30490) );
  AND2X1 U12753 ( .IN1(n3881), .IN2(n12365), .Q(n12382) );
  AND3X1 U12754 ( .IN1(test_so5), .IN2(n12383), .IN3(n9071), .Q(n12381) );
  OR2X1 U12755 ( .IN1(n943), .IN2(n3436), .Q(n12383) );
  AND2X1 U12756 ( .IN1(n9162), .IN2(g5575), .Q(n12380) );
  OR3X1 U12757 ( .IN1(n12384), .IN2(n12385), .IN3(n12386), .Q(g30489) );
  AND2X1 U12758 ( .IN1(n3881), .IN2(n12370), .Q(n12386) );
  AND3X1 U12759 ( .IN1(n12387), .IN2(g5587), .IN3(n9071), .Q(n12385) );
  OR2X1 U12760 ( .IN1(n944), .IN2(n3436), .Q(n12387) );
  OR2X1 U12761 ( .IN1(n8640), .IN2(g5511), .Q(n3436) );
  AND2X1 U12762 ( .IN1(n9162), .IN2(g5571), .Q(n12384) );
  OR3X1 U12763 ( .IN1(n12388), .IN2(n12389), .IN3(n12390), .Q(g30488) );
  AND2X1 U12764 ( .IN1(n3886), .IN2(n12356), .Q(n12390) );
  AND3X1 U12765 ( .IN1(n12391), .IN2(g5583), .IN3(n9071), .Q(n12389) );
  OR2X1 U12766 ( .IN1(n945), .IN2(n3437), .Q(n12391) );
  AND2X1 U12767 ( .IN1(n9162), .IN2(g5563), .Q(n12388) );
  OR3X1 U12768 ( .IN1(n12392), .IN2(n12393), .IN3(n12394), .Q(g30487) );
  AND2X1 U12769 ( .IN1(n3886), .IN2(n11603), .Q(n12394) );
  INVX0 U12770 ( .INP(n946), .ZN(n11603) );
  AND3X1 U12771 ( .IN1(n12395), .IN2(g5579), .IN3(n9071), .Q(n12393) );
  OR2X1 U12772 ( .IN1(n946), .IN2(n3437), .Q(n12395) );
  OR2X1 U12773 ( .IN1(n5566), .IN2(g5527), .Q(n946) );
  AND2X1 U12774 ( .IN1(n9163), .IN2(g5555), .Q(n12392) );
  OR3X1 U12775 ( .IN1(n12396), .IN2(n12397), .IN3(n12398), .Q(g30486) );
  AND2X1 U12776 ( .IN1(n3886), .IN2(n12365), .Q(n12398) );
  INVX0 U12777 ( .INP(n943), .ZN(n12365) );
  AND3X1 U12778 ( .IN1(n12399), .IN2(g5575), .IN3(n9071), .Q(n12397) );
  OR2X1 U12779 ( .IN1(n943), .IN2(n3437), .Q(n12399) );
  OR2X1 U12780 ( .IN1(n5389), .IN2(g5535), .Q(n943) );
  AND2X1 U12781 ( .IN1(n9163), .IN2(g5547), .Q(n12396) );
  OR3X1 U12782 ( .IN1(n12400), .IN2(n12401), .IN3(n12402), .Q(g30485) );
  AND2X1 U12783 ( .IN1(n3886), .IN2(n12370), .Q(n12402) );
  INVX0 U12784 ( .INP(n944), .ZN(n12370) );
  AND3X1 U12785 ( .IN1(n12403), .IN2(g5571), .IN3(n9071), .Q(n12401) );
  OR2X1 U12786 ( .IN1(n944), .IN2(n3437), .Q(n12403) );
  OR2X1 U12787 ( .IN1(n5575), .IN2(g5517), .Q(n3437) );
  OR2X1 U12788 ( .IN1(g5527), .IN2(g5535), .Q(n944) );
  AND2X1 U12789 ( .IN1(n9163), .IN2(g5543), .Q(n12400) );
  OR3X1 U12790 ( .IN1(n12404), .IN2(n12405), .IN3(n12406), .Q(g30484) );
  AND2X1 U12791 ( .IN1(n9163), .IN2(g5567), .Q(n12406) );
  AND2X1 U12792 ( .IN1(n3891), .IN2(n3765), .Q(n12405) );
  AND3X1 U12793 ( .IN1(n9056), .IN2(g5563), .IN3(n12407), .Q(n12404) );
  INVX0 U12794 ( .INP(n3891), .ZN(n12407) );
  OR3X1 U12795 ( .IN1(n12408), .IN2(n12409), .IN3(n12410), .Q(g30483) );
  AND2X1 U12796 ( .IN1(test_so6), .IN2(n9138), .Q(n12410) );
  AND2X1 U12797 ( .IN1(n3894), .IN2(n3765), .Q(n12409) );
  AND3X1 U12798 ( .IN1(n9057), .IN2(g5555), .IN3(n12411), .Q(n12408) );
  INVX0 U12799 ( .INP(n3894), .ZN(n12411) );
  OR3X1 U12800 ( .IN1(n12412), .IN2(n12413), .IN3(n12414), .Q(g30482) );
  AND2X1 U12801 ( .IN1(n9163), .IN2(g5551), .Q(n12414) );
  AND2X1 U12802 ( .IN1(n3896), .IN2(n3765), .Q(n12413) );
  AND3X1 U12803 ( .IN1(n9056), .IN2(g5547), .IN3(n12415), .Q(n12412) );
  INVX0 U12804 ( .INP(n3896), .ZN(n12415) );
  OR3X1 U12805 ( .IN1(n12416), .IN2(n12417), .IN3(n12418), .Q(g30481) );
  AND2X1 U12806 ( .IN1(n9163), .IN2(g5535), .Q(n12418) );
  AND2X1 U12807 ( .IN1(n3898), .IN2(n3765), .Q(n12417) );
  AND3X1 U12808 ( .IN1(n9056), .IN2(g5543), .IN3(n12419), .Q(n12416) );
  INVX0 U12809 ( .INP(n3898), .ZN(n12419) );
  AND2X1 U12810 ( .IN1(n11606), .IN2(n5575), .Q(g30480) );
  AND3X1 U12811 ( .IN1(n9056), .IN2(n11599), .IN3(n5647), .Q(n11606) );
  OR2X1 U12812 ( .IN1(n12420), .IN2(n12249), .Q(n11599) );
  OR3X1 U12813 ( .IN1(n12421), .IN2(n12422), .IN3(n12423), .Q(g30479) );
  AND2X1 U12814 ( .IN1(n9163), .IN2(g5268), .Q(n12423) );
  AND2X1 U12815 ( .IN1(n3765), .IN2(g32975), .Q(n12422) );
  AND2X1 U12816 ( .IN1(n9490), .IN2(g5272), .Q(n12421) );
  OR3X1 U12817 ( .IN1(n12424), .IN2(n12425), .IN3(n12426), .Q(g30478) );
  AND2X1 U12818 ( .IN1(n12427), .IN2(n3765), .Q(n12426) );
  INVX0 U12819 ( .INP(n12428), .ZN(n12427) );
  AND2X1 U12820 ( .IN1(n9163), .IN2(g5264), .Q(n12425) );
  AND3X1 U12821 ( .IN1(n12428), .IN2(g5220), .IN3(n9071), .Q(n12424) );
  OR2X1 U12822 ( .IN1(n5650), .IN2(n223), .Q(n12428) );
  OR3X1 U12823 ( .IN1(n12429), .IN2(n12430), .IN3(n12431), .Q(g30477) );
  AND2X1 U12824 ( .IN1(n11621), .IN2(n3765), .Q(n12431) );
  INVX0 U12825 ( .INP(n12432), .ZN(n11621) );
  AND2X1 U12826 ( .IN1(n9163), .IN2(g5260), .Q(n12430) );
  AND3X1 U12827 ( .IN1(n12432), .IN2(g5212), .IN3(n9071), .Q(n12429) );
  OR2X1 U12828 ( .IN1(n5650), .IN2(n232), .Q(n12432) );
  OR3X1 U12829 ( .IN1(n12433), .IN2(n12434), .IN3(n12435), .Q(g30476) );
  AND2X1 U12830 ( .IN1(n12436), .IN2(n3765), .Q(n12435) );
  INVX0 U12831 ( .INP(n12437), .ZN(n12436) );
  AND2X1 U12832 ( .IN1(n9163), .IN2(g5256), .Q(n12434) );
  AND3X1 U12833 ( .IN1(n12437), .IN2(g5204), .IN3(n9071), .Q(n12433) );
  OR2X1 U12834 ( .IN1(n5650), .IN2(n225), .Q(n12437) );
  OR3X1 U12835 ( .IN1(n12438), .IN2(n12439), .IN3(n12440), .Q(g30475) );
  AND2X1 U12836 ( .IN1(n3908), .IN2(n12441), .Q(n12440) );
  AND3X1 U12837 ( .IN1(n12442), .IN2(g5268), .IN3(n9071), .Q(n12439) );
  OR2X1 U12838 ( .IN1(n764), .IN2(n231), .Q(n12442) );
  AND2X1 U12839 ( .IN1(n9163), .IN2(g5252), .Q(n12438) );
  OR3X1 U12840 ( .IN1(n12443), .IN2(n12444), .IN3(n12445), .Q(g30474) );
  AND2X1 U12841 ( .IN1(n3908), .IN2(n11624), .Q(n12445) );
  AND3X1 U12842 ( .IN1(n12446), .IN2(g5264), .IN3(n9071), .Q(n12444) );
  OR2X1 U12843 ( .IN1(n764), .IN2(n223), .Q(n12446) );
  AND2X1 U12844 ( .IN1(n9163), .IN2(g5248), .Q(n12443) );
  OR3X1 U12845 ( .IN1(n12447), .IN2(n12448), .IN3(n12449), .Q(g30473) );
  AND2X1 U12846 ( .IN1(n3908), .IN2(n12450), .Q(n12449) );
  AND3X1 U12847 ( .IN1(n12451), .IN2(g5260), .IN3(n9070), .Q(n12448) );
  OR2X1 U12848 ( .IN1(n764), .IN2(n232), .Q(n12451) );
  AND2X1 U12849 ( .IN1(n9163), .IN2(g5244), .Q(n12447) );
  OR3X1 U12850 ( .IN1(n12452), .IN2(n12453), .IN3(n12454), .Q(g30472) );
  AND2X1 U12851 ( .IN1(n3908), .IN2(n12455), .Q(n12454) );
  AND3X1 U12852 ( .IN1(n12456), .IN2(g5256), .IN3(n9070), .Q(n12453) );
  OR2X1 U12853 ( .IN1(n764), .IN2(n225), .Q(n12456) );
  OR2X1 U12854 ( .IN1(n8642), .IN2(n5570), .Q(n764) );
  AND2X1 U12855 ( .IN1(n9163), .IN2(g5240), .Q(n12452) );
  OR3X1 U12856 ( .IN1(n12457), .IN2(n12458), .IN3(n12459), .Q(g30471) );
  AND2X1 U12857 ( .IN1(n3914), .IN2(n12441), .Q(n12459) );
  AND3X1 U12858 ( .IN1(n12460), .IN2(g5252), .IN3(n9070), .Q(n12458) );
  OR2X1 U12859 ( .IN1(n3446), .IN2(n231), .Q(n12460) );
  AND2X1 U12860 ( .IN1(n9163), .IN2(g5236), .Q(n12457) );
  OR3X1 U12861 ( .IN1(n12461), .IN2(n12462), .IN3(n12463), .Q(g30470) );
  AND2X1 U12862 ( .IN1(n3914), .IN2(n11624), .Q(n12463) );
  AND3X1 U12863 ( .IN1(n12464), .IN2(g5248), .IN3(n9070), .Q(n12462) );
  OR2X1 U12864 ( .IN1(n3446), .IN2(n223), .Q(n12464) );
  AND2X1 U12865 ( .IN1(n9163), .IN2(g5232), .Q(n12461) );
  OR3X1 U12866 ( .IN1(n12465), .IN2(n12466), .IN3(n12467), .Q(g30469) );
  AND2X1 U12867 ( .IN1(n3914), .IN2(n12450), .Q(n12467) );
  AND3X1 U12868 ( .IN1(n12468), .IN2(g5244), .IN3(n9070), .Q(n12466) );
  OR2X1 U12869 ( .IN1(n3446), .IN2(n232), .Q(n12468) );
  AND2X1 U12870 ( .IN1(test_so82), .IN2(n9138), .Q(n12465) );
  OR3X1 U12871 ( .IN1(n12469), .IN2(n12470), .IN3(n12471), .Q(g30468) );
  AND2X1 U12872 ( .IN1(n3914), .IN2(n12455), .Q(n12471) );
  AND3X1 U12873 ( .IN1(n12472), .IN2(g5240), .IN3(n9070), .Q(n12470) );
  OR2X1 U12874 ( .IN1(n3446), .IN2(n225), .Q(n12472) );
  OR2X1 U12875 ( .IN1(n8642), .IN2(g5164), .Q(n3446) );
  AND2X1 U12876 ( .IN1(n9163), .IN2(g5224), .Q(n12469) );
  OR3X1 U12877 ( .IN1(n12473), .IN2(n12474), .IN3(n12475), .Q(g30467) );
  AND2X1 U12878 ( .IN1(n3919), .IN2(n12441), .Q(n12475) );
  AND3X1 U12879 ( .IN1(n12476), .IN2(g5236), .IN3(n9070), .Q(n12474) );
  OR2X1 U12880 ( .IN1(n3447), .IN2(n231), .Q(n12476) );
  AND2X1 U12881 ( .IN1(n9163), .IN2(g5216), .Q(n12473) );
  OR3X1 U12882 ( .IN1(n12477), .IN2(n12478), .IN3(n12479), .Q(g30466) );
  AND2X1 U12883 ( .IN1(n3919), .IN2(n11624), .Q(n12479) );
  INVX0 U12884 ( .INP(n223), .ZN(n11624) );
  AND3X1 U12885 ( .IN1(n12480), .IN2(g5232), .IN3(n9070), .Q(n12478) );
  OR2X1 U12886 ( .IN1(n3447), .IN2(n223), .Q(n12480) );
  OR2X1 U12887 ( .IN1(n5567), .IN2(g5180), .Q(n223) );
  AND2X1 U12888 ( .IN1(n9163), .IN2(g5208), .Q(n12477) );
  OR3X1 U12889 ( .IN1(n12481), .IN2(n12482), .IN3(n12483), .Q(g30465) );
  AND2X1 U12890 ( .IN1(n3919), .IN2(n12450), .Q(n12483) );
  INVX0 U12891 ( .INP(n232), .ZN(n12450) );
  AND3X1 U12892 ( .IN1(test_so82), .IN2(n12484), .IN3(n9070), .Q(n12482) );
  OR2X1 U12893 ( .IN1(n3447), .IN2(n232), .Q(n12484) );
  OR2X1 U12894 ( .IN1(n5384), .IN2(g5188), .Q(n232) );
  AND2X1 U12895 ( .IN1(n9163), .IN2(g5200), .Q(n12481) );
  OR3X1 U12896 ( .IN1(n12485), .IN2(n12486), .IN3(n12487), .Q(g30464) );
  AND2X1 U12897 ( .IN1(n3919), .IN2(n12455), .Q(n12487) );
  INVX0 U12898 ( .INP(n225), .ZN(n12455) );
  AND3X1 U12899 ( .IN1(n12488), .IN2(g5224), .IN3(n9070), .Q(n12486) );
  OR2X1 U12900 ( .IN1(n3447), .IN2(n225), .Q(n12488) );
  OR2X1 U12901 ( .IN1(g5188), .IN2(g5180), .Q(n225) );
  OR2X1 U12902 ( .IN1(n5570), .IN2(g5170), .Q(n3447) );
  AND2X1 U12903 ( .IN1(n9163), .IN2(g5196), .Q(n12485) );
  OR3X1 U12904 ( .IN1(n12489), .IN2(n12490), .IN3(n12491), .Q(g30463) );
  AND2X1 U12905 ( .IN1(n9164), .IN2(g5220), .Q(n12491) );
  AND2X1 U12906 ( .IN1(n3924), .IN2(n3765), .Q(n12490) );
  AND3X1 U12907 ( .IN1(n9055), .IN2(g5216), .IN3(n12492), .Q(n12489) );
  INVX0 U12908 ( .INP(n3924), .ZN(n12492) );
  OR3X1 U12909 ( .IN1(n12493), .IN2(n12494), .IN3(n12495), .Q(g30462) );
  AND2X1 U12910 ( .IN1(n9164), .IN2(g5212), .Q(n12495) );
  AND2X1 U12911 ( .IN1(n3927), .IN2(n3765), .Q(n12494) );
  AND3X1 U12912 ( .IN1(n9055), .IN2(g5208), .IN3(n12496), .Q(n12493) );
  INVX0 U12913 ( .INP(n3927), .ZN(n12496) );
  OR3X1 U12914 ( .IN1(n12497), .IN2(n12498), .IN3(n12499), .Q(g30461) );
  AND2X1 U12915 ( .IN1(n9164), .IN2(g5204), .Q(n12499) );
  AND2X1 U12916 ( .IN1(n3929), .IN2(n3765), .Q(n12498) );
  AND3X1 U12917 ( .IN1(n9055), .IN2(g5200), .IN3(n12500), .Q(n12497) );
  INVX0 U12918 ( .INP(n3929), .ZN(n12500) );
  OR3X1 U12919 ( .IN1(n12501), .IN2(n12502), .IN3(n12503), .Q(g30460) );
  AND2X1 U12920 ( .IN1(n9164), .IN2(g5188), .Q(n12503) );
  AND2X1 U12921 ( .IN1(n3931), .IN2(n3765), .Q(n12502) );
  AND3X1 U12922 ( .IN1(n9054), .IN2(g5196), .IN3(n12504), .Q(n12501) );
  INVX0 U12923 ( .INP(n3931), .ZN(n12504) );
  AND2X1 U12924 ( .IN1(n11627), .IN2(n5570), .Q(g30459) );
  AND3X1 U12925 ( .IN1(n9054), .IN2(n11620), .IN3(n5650), .Q(n11627) );
  OR2X1 U12926 ( .IN1(n12162), .IN2(n12249), .Q(n11620) );
  INVX0 U12927 ( .INP(n3833), .ZN(n12249) );
  OR3X1 U12928 ( .IN1(n12505), .IN2(n12506), .IN3(n9121), .Q(g30458) );
  INVX0 U12929 ( .INP(n12507), .ZN(n12506) );
  OR2X1 U12930 ( .IN1(n12508), .IN2(n5846), .Q(n12507) );
  AND2X1 U12931 ( .IN1(n12508), .IN2(g113), .Q(n12505) );
  AND2X1 U12932 ( .IN1(g4473), .IN2(n5765), .Q(n12508) );
  OR2X1 U12933 ( .IN1(n12509), .IN2(n12510), .Q(g30457) );
  AND2X1 U12934 ( .IN1(n12511), .IN2(n9022), .Q(n12510) );
  OR2X1 U12935 ( .IN1(n12512), .IN2(n12513), .Q(n12511) );
  AND3X1 U12936 ( .IN1(n12514), .IN2(n12515), .IN3(n5983), .Q(n12513) );
  OR2X1 U12937 ( .IN1(n12516), .IN2(n12517), .Q(n12515) );
  INVX0 U12938 ( .INP(n12518), .ZN(n12514) );
  AND2X1 U12939 ( .IN1(n12517), .IN2(n12516), .Q(n12518) );
  INVX0 U12940 ( .INP(g115), .ZN(n12517) );
  AND3X1 U12941 ( .IN1(n12519), .IN2(n12520), .IN3(n5981), .Q(n12512) );
  OR2X1 U12942 ( .IN1(n12521), .IN2(n12522), .Q(n12520) );
  INVX0 U12943 ( .INP(n12523), .ZN(n12519) );
  AND2X1 U12944 ( .IN1(n12522), .IN2(n12521), .Q(n12523) );
  INVX0 U12945 ( .INP(g126), .ZN(n12522) );
  AND2X1 U12946 ( .IN1(n9164), .IN2(g4122), .Q(n12509) );
  OR3X1 U12947 ( .IN1(n12524), .IN2(n12525), .IN3(n12526), .Q(g30456) );
  AND2X1 U12948 ( .IN1(n9164), .IN2(g4087), .Q(n12526) );
  AND2X1 U12949 ( .IN1(n3941), .IN2(n12527), .Q(n12525) );
  AND4X1 U12950 ( .IN1(test_so11), .IN2(n12528), .IN3(n10978), .IN4(g4169), 
        .Q(n12524) );
  OR3X1 U12951 ( .IN1(n12529), .IN2(n12530), .IN3(n12531), .Q(g30455) );
  AND2X1 U12952 ( .IN1(n9164), .IN2(g3961), .Q(n12531) );
  AND2X1 U12953 ( .IN1(n3765), .IN2(n9376), .Q(n12530) );
  AND2X1 U12954 ( .IN1(n9375), .IN2(g3965), .Q(n12529) );
  OR3X1 U12955 ( .IN1(n12532), .IN2(n12533), .IN3(n12534), .Q(g30454) );
  AND2X1 U12956 ( .IN1(n12535), .IN2(n3765), .Q(n12534) );
  INVX0 U12957 ( .INP(n12536), .ZN(n12535) );
  AND2X1 U12958 ( .IN1(n9164), .IN2(g3957), .Q(n12533) );
  AND3X1 U12959 ( .IN1(n12536), .IN2(g3913), .IN3(n9070), .Q(n12532) );
  OR2X1 U12960 ( .IN1(n837), .IN2(n8823), .Q(n12536) );
  OR3X1 U12961 ( .IN1(n12537), .IN2(n12538), .IN3(n12539), .Q(g30453) );
  AND2X1 U12962 ( .IN1(n11676), .IN2(n3765), .Q(n12539) );
  INVX0 U12963 ( .INP(n12540), .ZN(n11676) );
  AND2X1 U12964 ( .IN1(n9164), .IN2(g3953), .Q(n12538) );
  AND3X1 U12965 ( .IN1(n12540), .IN2(g3905), .IN3(n9073), .Q(n12537) );
  OR2X1 U12966 ( .IN1(n844), .IN2(n8823), .Q(n12540) );
  OR3X1 U12967 ( .IN1(n12541), .IN2(n12542), .IN3(n12543), .Q(g30452) );
  AND2X1 U12968 ( .IN1(n12544), .IN2(n3765), .Q(n12543) );
  INVX0 U12969 ( .INP(n12545), .ZN(n12544) );
  AND2X1 U12970 ( .IN1(test_so65), .IN2(n9139), .Q(n12542) );
  AND3X1 U12971 ( .IN1(n12545), .IN2(g3897), .IN3(n9070), .Q(n12541) );
  OR2X1 U12972 ( .IN1(n839), .IN2(n8823), .Q(n12545) );
  OR3X1 U12973 ( .IN1(n12546), .IN2(n12547), .IN3(n12548), .Q(g30451) );
  AND2X1 U12974 ( .IN1(n3951), .IN2(n12549), .Q(n12548) );
  AND3X1 U12975 ( .IN1(n12550), .IN2(g3961), .IN3(n9070), .Q(n12547) );
  OR2X1 U12976 ( .IN1(n843), .IN2(n1151), .Q(n12550) );
  AND2X1 U12977 ( .IN1(n9164), .IN2(g3945), .Q(n12546) );
  OR3X1 U12978 ( .IN1(n12551), .IN2(n12552), .IN3(n12553), .Q(g30450) );
  AND2X1 U12979 ( .IN1(n3951), .IN2(n11679), .Q(n12553) );
  AND3X1 U12980 ( .IN1(n12554), .IN2(g3957), .IN3(n9069), .Q(n12552) );
  OR2X1 U12981 ( .IN1(n837), .IN2(n1151), .Q(n12554) );
  AND2X1 U12982 ( .IN1(n9164), .IN2(g3941), .Q(n12551) );
  OR3X1 U12983 ( .IN1(n12555), .IN2(n12556), .IN3(n12557), .Q(g30449) );
  AND2X1 U12984 ( .IN1(n3951), .IN2(n12558), .Q(n12557) );
  AND3X1 U12985 ( .IN1(n12559), .IN2(g3953), .IN3(n9069), .Q(n12556) );
  OR2X1 U12986 ( .IN1(n844), .IN2(n1151), .Q(n12559) );
  AND2X1 U12987 ( .IN1(n9164), .IN2(g3937), .Q(n12555) );
  OR3X1 U12988 ( .IN1(n12560), .IN2(n12561), .IN3(n12562), .Q(g30448) );
  AND2X1 U12989 ( .IN1(n3951), .IN2(n12563), .Q(n12562) );
  AND3X1 U12990 ( .IN1(test_so65), .IN2(n12564), .IN3(n9069), .Q(n12561) );
  OR2X1 U12991 ( .IN1(n839), .IN2(n1151), .Q(n12564) );
  OR2X1 U12992 ( .IN1(n8639), .IN2(n5572), .Q(n1151) );
  AND2X1 U12993 ( .IN1(n9164), .IN2(g3933), .Q(n12560) );
  OR3X1 U12994 ( .IN1(n12565), .IN2(n12566), .IN3(n12567), .Q(g30447) );
  AND2X1 U12995 ( .IN1(n3957), .IN2(n12549), .Q(n12567) );
  AND3X1 U12996 ( .IN1(n12568), .IN2(g3945), .IN3(n9069), .Q(n12566) );
  OR2X1 U12997 ( .IN1(n843), .IN2(n3481), .Q(n12568) );
  AND2X1 U12998 ( .IN1(n9164), .IN2(g3929), .Q(n12565) );
  OR3X1 U12999 ( .IN1(n12569), .IN2(n12570), .IN3(n12571), .Q(g30446) );
  AND2X1 U13000 ( .IN1(n3957), .IN2(n11679), .Q(n12571) );
  AND3X1 U13001 ( .IN1(n12572), .IN2(g3941), .IN3(n9069), .Q(n12570) );
  OR2X1 U13002 ( .IN1(n837), .IN2(n3481), .Q(n12572) );
  AND2X1 U13003 ( .IN1(n9164), .IN2(g3925), .Q(n12569) );
  OR3X1 U13004 ( .IN1(n12573), .IN2(n12574), .IN3(n12575), .Q(g30445) );
  AND2X1 U13005 ( .IN1(n3957), .IN2(n12558), .Q(n12575) );
  AND3X1 U13006 ( .IN1(n12576), .IN2(g3937), .IN3(n9069), .Q(n12574) );
  OR2X1 U13007 ( .IN1(n844), .IN2(n3481), .Q(n12576) );
  AND2X1 U13008 ( .IN1(n9164), .IN2(g3921), .Q(n12573) );
  OR3X1 U13009 ( .IN1(n12577), .IN2(n12578), .IN3(n12579), .Q(g30444) );
  AND2X1 U13010 ( .IN1(n3957), .IN2(n12563), .Q(n12579) );
  AND3X1 U13011 ( .IN1(n12580), .IN2(g3933), .IN3(n9069), .Q(n12578) );
  OR2X1 U13012 ( .IN1(n839), .IN2(n3481), .Q(n12580) );
  OR2X1 U13013 ( .IN1(n8639), .IN2(g3857), .Q(n3481) );
  AND2X1 U13014 ( .IN1(n9164), .IN2(g3917), .Q(n12577) );
  OR3X1 U13015 ( .IN1(n12581), .IN2(n12582), .IN3(n12583), .Q(g30443) );
  AND2X1 U13016 ( .IN1(n3962), .IN2(n12549), .Q(n12583) );
  AND3X1 U13017 ( .IN1(n12584), .IN2(g3929), .IN3(n9069), .Q(n12582) );
  OR2X1 U13018 ( .IN1(n843), .IN2(n3482), .Q(n12584) );
  AND2X1 U13019 ( .IN1(n9164), .IN2(g3909), .Q(n12581) );
  OR3X1 U13020 ( .IN1(n12585), .IN2(n12586), .IN3(n12587), .Q(g30442) );
  AND2X1 U13021 ( .IN1(n3962), .IN2(n11679), .Q(n12587) );
  INVX0 U13022 ( .INP(n837), .ZN(n11679) );
  AND3X1 U13023 ( .IN1(n12588), .IN2(g3925), .IN3(n9069), .Q(n12586) );
  OR2X1 U13024 ( .IN1(n837), .IN2(n3482), .Q(n12588) );
  OR2X1 U13025 ( .IN1(n5564), .IN2(g3873), .Q(n837) );
  AND2X1 U13026 ( .IN1(n9164), .IN2(g3901), .Q(n12585) );
  OR3X1 U13027 ( .IN1(n12589), .IN2(n12590), .IN3(n12591), .Q(g30441) );
  AND2X1 U13028 ( .IN1(n3962), .IN2(n12558), .Q(n12591) );
  INVX0 U13029 ( .INP(n844), .ZN(n12558) );
  AND3X1 U13030 ( .IN1(n12592), .IN2(g3921), .IN3(n9069), .Q(n12590) );
  OR2X1 U13031 ( .IN1(n844), .IN2(n3482), .Q(n12592) );
  OR2X1 U13032 ( .IN1(n5387), .IN2(g3881), .Q(n844) );
  AND2X1 U13033 ( .IN1(n9164), .IN2(g3893), .Q(n12589) );
  OR3X1 U13034 ( .IN1(n12593), .IN2(n12594), .IN3(n12595), .Q(g30440) );
  AND2X1 U13035 ( .IN1(n3962), .IN2(n12563), .Q(n12595) );
  INVX0 U13036 ( .INP(n839), .ZN(n12563) );
  AND3X1 U13037 ( .IN1(n12596), .IN2(g3917), .IN3(n9069), .Q(n12594) );
  OR2X1 U13038 ( .IN1(n839), .IN2(n3482), .Q(n12596) );
  OR2X1 U13039 ( .IN1(n5572), .IN2(g3863), .Q(n3482) );
  OR2X1 U13040 ( .IN1(g3881), .IN2(g3873), .Q(n839) );
  AND2X1 U13041 ( .IN1(test_so24), .IN2(n9139), .Q(n12593) );
  OR3X1 U13042 ( .IN1(n12597), .IN2(n12598), .IN3(n12599), .Q(g30439) );
  AND2X1 U13043 ( .IN1(n9164), .IN2(g3913), .Q(n12599) );
  AND2X1 U13044 ( .IN1(n3967), .IN2(n3765), .Q(n12598) );
  AND3X1 U13045 ( .IN1(n9054), .IN2(g3909), .IN3(n12600), .Q(n12597) );
  INVX0 U13046 ( .INP(n3967), .ZN(n12600) );
  OR3X1 U13047 ( .IN1(n12601), .IN2(n12602), .IN3(n12603), .Q(g30438) );
  AND2X1 U13048 ( .IN1(n9164), .IN2(g3905), .Q(n12603) );
  AND2X1 U13049 ( .IN1(n3970), .IN2(n3765), .Q(n12602) );
  AND3X1 U13050 ( .IN1(n9053), .IN2(g3901), .IN3(n12604), .Q(n12601) );
  INVX0 U13051 ( .INP(n3970), .ZN(n12604) );
  OR3X1 U13052 ( .IN1(n12605), .IN2(n12606), .IN3(n12607), .Q(g30437) );
  AND2X1 U13053 ( .IN1(n9165), .IN2(g3897), .Q(n12607) );
  AND2X1 U13054 ( .IN1(n3972), .IN2(n3765), .Q(n12606) );
  AND3X1 U13055 ( .IN1(n9054), .IN2(g3893), .IN3(n12608), .Q(n12605) );
  INVX0 U13056 ( .INP(n3972), .ZN(n12608) );
  OR3X1 U13057 ( .IN1(n12609), .IN2(n12610), .IN3(n12611), .Q(g30436) );
  AND2X1 U13058 ( .IN1(n9165), .IN2(g3881), .Q(n12611) );
  AND2X1 U13059 ( .IN1(n3974), .IN2(n3765), .Q(n12610) );
  AND3X1 U13060 ( .IN1(test_so24), .IN2(n9052), .IN3(n12612), .Q(n12609) );
  INVX0 U13061 ( .INP(n3974), .ZN(n12612) );
  AND2X1 U13062 ( .IN1(n11682), .IN2(n5572), .Q(g30435) );
  AND3X1 U13063 ( .IN1(n8823), .IN2(n9052), .IN3(n11675), .Q(n11682) );
  OR3X1 U13064 ( .IN1(n5480), .IN2(n5340), .IN3(n12163), .Q(n11675) );
  OR3X1 U13065 ( .IN1(n12613), .IN2(n12614), .IN3(n12615), .Q(g30434) );
  AND2X1 U13066 ( .IN1(n9165), .IN2(g3610), .Q(n12615) );
  AND2X1 U13067 ( .IN1(n10982), .IN2(n3765), .Q(n12614) );
  AND2X1 U13068 ( .IN1(n12616), .IN2(g3614), .Q(n12613) );
  OR3X1 U13069 ( .IN1(n12617), .IN2(n12618), .IN3(n12619), .Q(g30433) );
  AND2X1 U13070 ( .IN1(n12620), .IN2(n3765), .Q(n12619) );
  INVX0 U13071 ( .INP(n12621), .ZN(n12620) );
  AND2X1 U13072 ( .IN1(n9165), .IN2(g3606), .Q(n12618) );
  AND3X1 U13073 ( .IN1(n12621), .IN2(g3562), .IN3(n9069), .Q(n12617) );
  OR2X1 U13074 ( .IN1(n5645), .IN2(n471), .Q(n12621) );
  OR3X1 U13075 ( .IN1(n12622), .IN2(n12623), .IN3(n12624), .Q(g30432) );
  AND2X1 U13076 ( .IN1(n11697), .IN2(n3765), .Q(n12624) );
  INVX0 U13077 ( .INP(n12625), .ZN(n11697) );
  AND2X1 U13078 ( .IN1(test_so43), .IN2(n9139), .Q(n12623) );
  AND3X1 U13079 ( .IN1(n12625), .IN2(g3554), .IN3(n9069), .Q(n12622) );
  OR2X1 U13080 ( .IN1(n5645), .IN2(n463), .Q(n12625) );
  OR3X1 U13081 ( .IN1(n12626), .IN2(n12627), .IN3(n12628), .Q(g30431) );
  AND2X1 U13082 ( .IN1(n12629), .IN2(n3765), .Q(n12628) );
  INVX0 U13083 ( .INP(n12630), .ZN(n12629) );
  AND2X1 U13084 ( .IN1(n9165), .IN2(g3598), .Q(n12627) );
  AND3X1 U13085 ( .IN1(n12630), .IN2(g3546), .IN3(n9068), .Q(n12626) );
  OR2X1 U13086 ( .IN1(n5645), .IN2(n465), .Q(n12630) );
  OR3X1 U13087 ( .IN1(n12631), .IN2(n12632), .IN3(n12633), .Q(g30430) );
  AND2X1 U13088 ( .IN1(n3984), .IN2(n12634), .Q(n12633) );
  AND3X1 U13089 ( .IN1(n12635), .IN2(g3610), .IN3(n9068), .Q(n12632) );
  OR2X1 U13090 ( .IN1(n470), .IN2(n115), .Q(n12635) );
  AND2X1 U13091 ( .IN1(n9165), .IN2(g3594), .Q(n12631) );
  OR3X1 U13092 ( .IN1(n12636), .IN2(n12637), .IN3(n12638), .Q(g30429) );
  AND2X1 U13093 ( .IN1(n3984), .IN2(n11700), .Q(n12638) );
  AND3X1 U13094 ( .IN1(n12639), .IN2(g3606), .IN3(n9068), .Q(n12637) );
  OR2X1 U13095 ( .IN1(n471), .IN2(n115), .Q(n12639) );
  AND2X1 U13096 ( .IN1(n9165), .IN2(g3590), .Q(n12636) );
  OR3X1 U13097 ( .IN1(n12640), .IN2(n12641), .IN3(n12642), .Q(g30428) );
  AND2X1 U13098 ( .IN1(n3984), .IN2(n12643), .Q(n12642) );
  AND3X1 U13099 ( .IN1(test_so43), .IN2(n12644), .IN3(n9068), .Q(n12641) );
  OR2X1 U13100 ( .IN1(n463), .IN2(n115), .Q(n12644) );
  AND2X1 U13101 ( .IN1(n9165), .IN2(g3586), .Q(n12640) );
  OR3X1 U13102 ( .IN1(n12645), .IN2(n12646), .IN3(n12647), .Q(g30427) );
  AND2X1 U13103 ( .IN1(n3984), .IN2(n12648), .Q(n12647) );
  AND3X1 U13104 ( .IN1(n12649), .IN2(g3598), .IN3(n9068), .Q(n12646) );
  OR2X1 U13105 ( .IN1(n465), .IN2(n115), .Q(n12649) );
  OR2X1 U13106 ( .IN1(n8637), .IN2(n5576), .Q(n115) );
  AND2X1 U13107 ( .IN1(n9165), .IN2(g3582), .Q(n12645) );
  OR3X1 U13108 ( .IN1(n12650), .IN2(n12651), .IN3(n12652), .Q(g30426) );
  AND2X1 U13109 ( .IN1(n3990), .IN2(n12634), .Q(n12652) );
  AND3X1 U13110 ( .IN1(n12653), .IN2(g3594), .IN3(n9068), .Q(n12651) );
  OR2X1 U13111 ( .IN1(n470), .IN2(n3491), .Q(n12653) );
  AND2X1 U13112 ( .IN1(n9165), .IN2(g3578), .Q(n12650) );
  OR3X1 U13113 ( .IN1(n12654), .IN2(n12655), .IN3(n12656), .Q(g30425) );
  AND2X1 U13114 ( .IN1(n3990), .IN2(n11700), .Q(n12656) );
  AND3X1 U13115 ( .IN1(n12657), .IN2(g3590), .IN3(n9068), .Q(n12655) );
  OR2X1 U13116 ( .IN1(n471), .IN2(n3491), .Q(n12657) );
  AND2X1 U13117 ( .IN1(n9165), .IN2(g3574), .Q(n12654) );
  OR3X1 U13118 ( .IN1(n12658), .IN2(n12659), .IN3(n12660), .Q(g30424) );
  AND2X1 U13119 ( .IN1(n3990), .IN2(n12643), .Q(n12660) );
  AND3X1 U13120 ( .IN1(n12661), .IN2(g3586), .IN3(n9068), .Q(n12659) );
  OR2X1 U13121 ( .IN1(n463), .IN2(n3491), .Q(n12661) );
  AND2X1 U13122 ( .IN1(n9165), .IN2(g3570), .Q(n12658) );
  OR3X1 U13123 ( .IN1(n12662), .IN2(n12663), .IN3(n12664), .Q(g30423) );
  AND2X1 U13124 ( .IN1(n3990), .IN2(n12648), .Q(n12664) );
  AND3X1 U13125 ( .IN1(n12665), .IN2(g3582), .IN3(n9068), .Q(n12663) );
  OR2X1 U13126 ( .IN1(n465), .IN2(n3491), .Q(n12665) );
  OR2X1 U13127 ( .IN1(n8637), .IN2(g3506), .Q(n3491) );
  AND2X1 U13128 ( .IN1(n9165), .IN2(g3566), .Q(n12662) );
  OR3X1 U13129 ( .IN1(n12666), .IN2(n12667), .IN3(n12668), .Q(g30422) );
  AND2X1 U13130 ( .IN1(n3995), .IN2(n12634), .Q(n12668) );
  AND3X1 U13131 ( .IN1(n12669), .IN2(g3578), .IN3(n9068), .Q(n12667) );
  OR2X1 U13132 ( .IN1(n470), .IN2(n3492), .Q(n12669) );
  AND2X1 U13133 ( .IN1(n9165), .IN2(g3558), .Q(n12666) );
  OR3X1 U13134 ( .IN1(n12670), .IN2(n12671), .IN3(n12672), .Q(g30421) );
  AND2X1 U13135 ( .IN1(n3995), .IN2(n11700), .Q(n12672) );
  INVX0 U13136 ( .INP(n471), .ZN(n11700) );
  AND3X1 U13137 ( .IN1(n12673), .IN2(g3574), .IN3(n9068), .Q(n12671) );
  OR2X1 U13138 ( .IN1(n471), .IN2(n3492), .Q(n12673) );
  OR2X1 U13139 ( .IN1(n5569), .IN2(g3522), .Q(n471) );
  AND2X1 U13140 ( .IN1(n9165), .IN2(g3550), .Q(n12670) );
  OR3X1 U13141 ( .IN1(n12674), .IN2(n12675), .IN3(n12676), .Q(g30420) );
  AND2X1 U13142 ( .IN1(n3995), .IN2(n12643), .Q(n12676) );
  INVX0 U13143 ( .INP(n463), .ZN(n12643) );
  AND3X1 U13144 ( .IN1(n12677), .IN2(g3570), .IN3(n9068), .Q(n12675) );
  OR2X1 U13145 ( .IN1(n463), .IN2(n3492), .Q(n12677) );
  OR2X1 U13146 ( .IN1(n5383), .IN2(g3530), .Q(n463) );
  AND2X1 U13147 ( .IN1(n9165), .IN2(g3542), .Q(n12674) );
  OR3X1 U13148 ( .IN1(n12678), .IN2(n12679), .IN3(n12680), .Q(g30419) );
  AND2X1 U13149 ( .IN1(n3995), .IN2(n12648), .Q(n12680) );
  INVX0 U13150 ( .INP(n465), .ZN(n12648) );
  AND3X1 U13151 ( .IN1(n12681), .IN2(g3566), .IN3(n9068), .Q(n12679) );
  OR2X1 U13152 ( .IN1(n465), .IN2(n3492), .Q(n12681) );
  OR2X1 U13153 ( .IN1(n5576), .IN2(g3512), .Q(n3492) );
  OR2X1 U13154 ( .IN1(g3522), .IN2(g3530), .Q(n465) );
  AND2X1 U13155 ( .IN1(n9165), .IN2(g3538), .Q(n12678) );
  OR3X1 U13156 ( .IN1(n12682), .IN2(n12683), .IN3(n12684), .Q(g30418) );
  AND2X1 U13157 ( .IN1(n9165), .IN2(g3562), .Q(n12684) );
  AND2X1 U13158 ( .IN1(n4000), .IN2(n3765), .Q(n12683) );
  AND3X1 U13159 ( .IN1(n9054), .IN2(g3558), .IN3(n12685), .Q(n12682) );
  INVX0 U13160 ( .INP(n4000), .ZN(n12685) );
  OR3X1 U13161 ( .IN1(n12686), .IN2(n12687), .IN3(n12688), .Q(g30417) );
  AND2X1 U13162 ( .IN1(n9165), .IN2(g3554), .Q(n12688) );
  AND2X1 U13163 ( .IN1(n4003), .IN2(n3765), .Q(n12687) );
  AND3X1 U13164 ( .IN1(n9054), .IN2(g3550), .IN3(n12689), .Q(n12686) );
  INVX0 U13165 ( .INP(n4003), .ZN(n12689) );
  OR3X1 U13166 ( .IN1(n12690), .IN2(n12691), .IN3(n12692), .Q(g30416) );
  AND2X1 U13167 ( .IN1(n9165), .IN2(g3546), .Q(n12692) );
  AND2X1 U13168 ( .IN1(n4005), .IN2(n3765), .Q(n12691) );
  AND3X1 U13169 ( .IN1(n9053), .IN2(g3542), .IN3(n12693), .Q(n12690) );
  INVX0 U13170 ( .INP(n4005), .ZN(n12693) );
  OR3X1 U13171 ( .IN1(n12694), .IN2(n12695), .IN3(n12696), .Q(g30415) );
  AND2X1 U13172 ( .IN1(n9165), .IN2(g3530), .Q(n12696) );
  AND2X1 U13173 ( .IN1(n4007), .IN2(n3765), .Q(n12695) );
  AND3X1 U13174 ( .IN1(n9054), .IN2(g3538), .IN3(n12697), .Q(n12694) );
  INVX0 U13175 ( .INP(n4007), .ZN(n12697) );
  AND2X1 U13176 ( .IN1(n11703), .IN2(n5576), .Q(g30414) );
  AND3X1 U13177 ( .IN1(n9053), .IN2(n11696), .IN3(n5645), .Q(n11703) );
  OR3X1 U13178 ( .IN1(n5340), .IN2(g4087), .IN3(n12163), .Q(n11696) );
  OR3X1 U13179 ( .IN1(n12698), .IN2(n12699), .IN3(n12700), .Q(g30413) );
  AND2X1 U13180 ( .IN1(test_so84), .IN2(n9140), .Q(n12700) );
  AND2X1 U13181 ( .IN1(n3765), .IN2(n10977), .Q(n12699) );
  AND2X1 U13182 ( .IN1(n12701), .IN2(g3263), .Q(n12698) );
  OR3X1 U13183 ( .IN1(n12702), .IN2(n12703), .IN3(n12704), .Q(g30412) );
  AND2X1 U13184 ( .IN1(n12705), .IN2(n3765), .Q(n12704) );
  INVX0 U13185 ( .INP(n12706), .ZN(n12705) );
  AND2X1 U13186 ( .IN1(n9165), .IN2(g3255), .Q(n12703) );
  AND3X1 U13187 ( .IN1(n12706), .IN2(g3211), .IN3(n9067), .Q(n12702) );
  OR2X1 U13188 ( .IN1(n5652), .IN2(n564), .Q(n12706) );
  OR3X1 U13189 ( .IN1(n12707), .IN2(n12708), .IN3(n12709), .Q(g30411) );
  AND2X1 U13190 ( .IN1(n11720), .IN2(n3765), .Q(n12709) );
  INVX0 U13191 ( .INP(n12710), .ZN(n11720) );
  AND2X1 U13192 ( .IN1(n9166), .IN2(g3251), .Q(n12708) );
  AND3X1 U13193 ( .IN1(n12710), .IN2(g3203), .IN3(n9067), .Q(n12707) );
  OR2X1 U13194 ( .IN1(n5652), .IN2(n561), .Q(n12710) );
  OR3X1 U13195 ( .IN1(n12711), .IN2(n12712), .IN3(n12713), .Q(g30410) );
  AND2X1 U13196 ( .IN1(n12714), .IN2(n3765), .Q(n12713) );
  INVX0 U13197 ( .INP(n12715), .ZN(n12714) );
  AND2X1 U13198 ( .IN1(n9166), .IN2(g3247), .Q(n12712) );
  AND3X1 U13199 ( .IN1(test_so88), .IN2(n12715), .IN3(n9067), .Q(n12711) );
  OR2X1 U13200 ( .IN1(n5652), .IN2(n562), .Q(n12715) );
  OR3X1 U13201 ( .IN1(n12716), .IN2(n12717), .IN3(n12718), .Q(g30409) );
  AND2X1 U13202 ( .IN1(n4015), .IN2(n12719), .Q(n12718) );
  AND3X1 U13203 ( .IN1(test_so84), .IN2(n12720), .IN3(n9067), .Q(n12717) );
  OR2X1 U13204 ( .IN1(n563), .IN2(n130), .Q(n12720) );
  AND2X1 U13205 ( .IN1(n9166), .IN2(g3243), .Q(n12716) );
  OR3X1 U13206 ( .IN1(n12721), .IN2(n12722), .IN3(n12723), .Q(g30408) );
  AND2X1 U13207 ( .IN1(n4015), .IN2(n11721), .Q(n12723) );
  AND3X1 U13208 ( .IN1(n12724), .IN2(g3255), .IN3(n9067), .Q(n12722) );
  OR2X1 U13209 ( .IN1(n564), .IN2(n130), .Q(n12724) );
  AND2X1 U13210 ( .IN1(n9166), .IN2(g3239), .Q(n12721) );
  OR3X1 U13211 ( .IN1(n12725), .IN2(n12726), .IN3(n12727), .Q(g30407) );
  AND2X1 U13212 ( .IN1(n4015), .IN2(n12728), .Q(n12727) );
  AND3X1 U13213 ( .IN1(n12729), .IN2(g3251), .IN3(n9067), .Q(n12726) );
  OR2X1 U13214 ( .IN1(n561), .IN2(n130), .Q(n12729) );
  AND2X1 U13215 ( .IN1(n9166), .IN2(g3235), .Q(n12725) );
  OR3X1 U13216 ( .IN1(n12730), .IN2(n12731), .IN3(n12732), .Q(g30406) );
  AND2X1 U13217 ( .IN1(n4015), .IN2(n12733), .Q(n12732) );
  AND3X1 U13218 ( .IN1(n12734), .IN2(g3247), .IN3(n9067), .Q(n12731) );
  OR2X1 U13219 ( .IN1(n562), .IN2(n130), .Q(n12734) );
  OR2X1 U13220 ( .IN1(n8644), .IN2(n5366), .Q(n130) );
  AND2X1 U13221 ( .IN1(n9166), .IN2(g3231), .Q(n12730) );
  OR3X1 U13222 ( .IN1(n12735), .IN2(n12736), .IN3(n12737), .Q(g30405) );
  AND2X1 U13223 ( .IN1(n4022), .IN2(n12719), .Q(n12737) );
  AND3X1 U13224 ( .IN1(n12738), .IN2(g3243), .IN3(n9067), .Q(n12736) );
  OR2X1 U13225 ( .IN1(n563), .IN2(n3502), .Q(n12738) );
  AND2X1 U13226 ( .IN1(n9166), .IN2(g3227), .Q(n12735) );
  OR3X1 U13227 ( .IN1(n12739), .IN2(n12740), .IN3(n12741), .Q(g30404) );
  AND2X1 U13228 ( .IN1(n4022), .IN2(n11721), .Q(n12741) );
  AND3X1 U13229 ( .IN1(n12742), .IN2(g3239), .IN3(n9067), .Q(n12740) );
  OR2X1 U13230 ( .IN1(n564), .IN2(n3502), .Q(n12742) );
  AND2X1 U13231 ( .IN1(n9148), .IN2(g3223), .Q(n12739) );
  OR3X1 U13232 ( .IN1(n12743), .IN2(n12744), .IN3(n12745), .Q(g30403) );
  AND2X1 U13233 ( .IN1(n4022), .IN2(n12728), .Q(n12745) );
  AND3X1 U13234 ( .IN1(n12746), .IN2(g3235), .IN3(n9067), .Q(n12744) );
  OR2X1 U13235 ( .IN1(n561), .IN2(n3502), .Q(n12746) );
  AND2X1 U13236 ( .IN1(n9145), .IN2(g3219), .Q(n12743) );
  OR3X1 U13237 ( .IN1(n12747), .IN2(n12748), .IN3(n12749), .Q(g30402) );
  AND2X1 U13238 ( .IN1(n4022), .IN2(n12733), .Q(n12749) );
  AND3X1 U13239 ( .IN1(n12750), .IN2(g3231), .IN3(n9067), .Q(n12748) );
  OR2X1 U13240 ( .IN1(n562), .IN2(n3502), .Q(n12750) );
  OR2X1 U13241 ( .IN1(n8644), .IN2(g3155), .Q(n3502) );
  AND2X1 U13242 ( .IN1(n9144), .IN2(g3215), .Q(n12747) );
  OR3X1 U13243 ( .IN1(n12751), .IN2(n12752), .IN3(n12753), .Q(g30401) );
  AND2X1 U13244 ( .IN1(n4027), .IN2(n12719), .Q(n12753) );
  AND3X1 U13245 ( .IN1(n12754), .IN2(g3227), .IN3(n9067), .Q(n12752) );
  OR2X1 U13246 ( .IN1(n563), .IN2(n3501), .Q(n12754) );
  AND2X1 U13247 ( .IN1(n9144), .IN2(g3207), .Q(n12751) );
  OR3X1 U13248 ( .IN1(n12755), .IN2(n12756), .IN3(n12757), .Q(g30400) );
  AND2X1 U13249 ( .IN1(n4027), .IN2(n11721), .Q(n12757) );
  INVX0 U13250 ( .INP(n564), .ZN(n11721) );
  AND3X1 U13251 ( .IN1(n12758), .IN2(g3223), .IN3(n9067), .Q(n12756) );
  OR2X1 U13252 ( .IN1(n564), .IN2(n3501), .Q(n12758) );
  OR2X1 U13253 ( .IN1(n5390), .IN2(g3171), .Q(n564) );
  AND2X1 U13254 ( .IN1(n9144), .IN2(g3199), .Q(n12755) );
  OR3X1 U13255 ( .IN1(n12759), .IN2(n12760), .IN3(n12761), .Q(g30399) );
  AND2X1 U13256 ( .IN1(n4027), .IN2(n12728), .Q(n12761) );
  INVX0 U13257 ( .INP(n561), .ZN(n12728) );
  AND3X1 U13258 ( .IN1(n12762), .IN2(g3219), .IN3(n9066), .Q(n12760) );
  OR2X1 U13259 ( .IN1(n561), .IN2(n3501), .Q(n12762) );
  OR2X1 U13260 ( .IN1(n5603), .IN2(g3179), .Q(n561) );
  AND2X1 U13261 ( .IN1(n9144), .IN2(g3191), .Q(n12759) );
  OR3X1 U13262 ( .IN1(n12763), .IN2(n12764), .IN3(n12765), .Q(g30398) );
  AND2X1 U13263 ( .IN1(n4027), .IN2(n12733), .Q(n12765) );
  INVX0 U13264 ( .INP(n562), .ZN(n12733) );
  AND3X1 U13265 ( .IN1(n12766), .IN2(g3215), .IN3(n9066), .Q(n12764) );
  OR2X1 U13266 ( .IN1(n562), .IN2(n3501), .Q(n12766) );
  OR2X1 U13267 ( .IN1(n5366), .IN2(g3161), .Q(n3501) );
  OR2X1 U13268 ( .IN1(g3171), .IN2(g3179), .Q(n562) );
  AND2X1 U13269 ( .IN1(n9144), .IN2(g3187), .Q(n12763) );
  OR3X1 U13270 ( .IN1(n12767), .IN2(n12768), .IN3(n12769), .Q(g30397) );
  AND2X1 U13271 ( .IN1(n9144), .IN2(g3211), .Q(n12769) );
  AND2X1 U13272 ( .IN1(n4032), .IN2(n3765), .Q(n12768) );
  AND3X1 U13273 ( .IN1(n9053), .IN2(g3207), .IN3(n12770), .Q(n12767) );
  INVX0 U13274 ( .INP(n4032), .ZN(n12770) );
  OR3X1 U13275 ( .IN1(n12771), .IN2(n12772), .IN3(n12773), .Q(g30396) );
  AND2X1 U13276 ( .IN1(n9144), .IN2(g3203), .Q(n12773) );
  AND2X1 U13277 ( .IN1(n4035), .IN2(n3765), .Q(n12772) );
  AND3X1 U13278 ( .IN1(n9053), .IN2(g3199), .IN3(n12774), .Q(n12771) );
  INVX0 U13279 ( .INP(n4035), .ZN(n12774) );
  OR3X1 U13280 ( .IN1(n12775), .IN2(n12776), .IN3(n12777), .Q(g30395) );
  AND2X1 U13281 ( .IN1(test_so88), .IN2(n9139), .Q(n12777) );
  AND2X1 U13282 ( .IN1(n4037), .IN2(n3765), .Q(n12776) );
  AND3X1 U13283 ( .IN1(n9053), .IN2(g3191), .IN3(n12778), .Q(n12775) );
  INVX0 U13284 ( .INP(n4037), .ZN(n12778) );
  OR3X1 U13285 ( .IN1(n12779), .IN2(n12780), .IN3(n12781), .Q(g30394) );
  AND2X1 U13286 ( .IN1(n9144), .IN2(g3179), .Q(n12781) );
  AND2X1 U13287 ( .IN1(n4039), .IN2(n3765), .Q(n12780) );
  AND3X1 U13288 ( .IN1(n9053), .IN2(g3187), .IN3(n12782), .Q(n12779) );
  INVX0 U13289 ( .INP(n4039), .ZN(n12782) );
  AND3X1 U13290 ( .IN1(n5366), .IN2(n9051), .IN3(n11717), .Q(g30393) );
  AND2X1 U13291 ( .IN1(n11719), .IN2(n5652), .Q(n11717) );
  OR2X1 U13292 ( .IN1(n12420), .IN2(n12163), .Q(n11719) );
  INVX0 U13293 ( .INP(n3799), .ZN(n12163) );
  OR2X1 U13294 ( .IN1(n12783), .IN2(n12784), .Q(g30392) );
  AND2X1 U13295 ( .IN1(n9144), .IN2(g2803), .Q(n12783) );
  OR2X1 U13296 ( .IN1(n12785), .IN2(n12786), .Q(g30391) );
  AND2X1 U13297 ( .IN1(n9144), .IN2(g2771), .Q(n12785) );
  OR2X1 U13298 ( .IN1(n12787), .IN2(n12784), .Q(g30390) );
  AND2X1 U13299 ( .IN1(n12788), .IN2(n9022), .Q(n12784) );
  OR2X1 U13300 ( .IN1(n12789), .IN2(n12790), .Q(n12788) );
  AND2X1 U13301 ( .IN1(n12791), .IN2(n12792), .Q(n12790) );
  AND4X1 U13302 ( .IN1(n12793), .IN2(n12794), .IN3(n12795), .IN4(n12796), .Q(
        n12791) );
  OR2X1 U13303 ( .IN1(n5545), .IN2(n12797), .Q(n12796) );
  OR2X1 U13304 ( .IN1(n5379), .IN2(n1256), .Q(n12795) );
  OR2X1 U13305 ( .IN1(n5609), .IN2(n12798), .Q(n12794) );
  OR2X1 U13306 ( .IN1(n5404), .IN2(n12799), .Q(n12793) );
  AND2X1 U13307 ( .IN1(n12800), .IN2(n12801), .Q(n12789) );
  AND4X1 U13308 ( .IN1(n12802), .IN2(n12803), .IN3(n12804), .IN4(n12805), .Q(
        n12800) );
  OR2X1 U13309 ( .IN1(n12797), .IN2(g2236), .Q(n12805) );
  OR2X1 U13310 ( .IN1(n1256), .IN2(g2370), .Q(n12804) );
  OR2X1 U13311 ( .IN1(n12798), .IN2(g2638), .Q(n12803) );
  OR2X1 U13312 ( .IN1(n12799), .IN2(g2504), .Q(n12802) );
  AND2X1 U13313 ( .IN1(g2834), .IN2(n9139), .Q(n12787) );
  OR2X1 U13314 ( .IN1(n12806), .IN2(n12786), .Q(g30389) );
  AND2X1 U13315 ( .IN1(n12807), .IN2(n9022), .Q(n12786) );
  OR2X1 U13316 ( .IN1(n12808), .IN2(n12809), .Q(n12807) );
  AND2X1 U13317 ( .IN1(n12810), .IN2(n12792), .Q(n12809) );
  AND4X1 U13318 ( .IN1(n12811), .IN2(n12812), .IN3(n12813), .IN4(n12814), .Q(
        n12810) );
  OR2X1 U13319 ( .IN1(n5544), .IN2(n12797), .Q(n12814) );
  OR2X1 U13320 ( .IN1(n5378), .IN2(n1256), .Q(n12813) );
  OR2X1 U13321 ( .IN1(n5610), .IN2(n12798), .Q(n12812) );
  OR2X1 U13322 ( .IN1(n5403), .IN2(n12799), .Q(n12811) );
  AND2X1 U13323 ( .IN1(n12815), .IN2(n12801), .Q(n12808) );
  INVX0 U13324 ( .INP(n12792), .ZN(n12801) );
  AND3X1 U13325 ( .IN1(n797), .IN2(n10197), .IN3(n5600), .Q(n12792) );
  AND2X1 U13326 ( .IN1(n12816), .IN2(n5349), .Q(n797) );
  INVX0 U13327 ( .INP(n9463), .ZN(n12816) );
  AND4X1 U13328 ( .IN1(n12817), .IN2(n12818), .IN3(n12819), .IN4(n12820), .Q(
        n12815) );
  OR2X1 U13329 ( .IN1(n12797), .IN2(g1677), .Q(n12820) );
  OR2X1 U13330 ( .IN1(n1256), .IN2(g1811), .Q(n12819) );
  OR2X1 U13331 ( .IN1(n12798), .IN2(g2079), .Q(n12818) );
  OR2X1 U13332 ( .IN1(test_so53), .IN2(n12799), .Q(n12817) );
  AND2X1 U13333 ( .IN1(g2831), .IN2(n9139), .Q(n12806) );
  OR2X1 U13334 ( .IN1(n12821), .IN2(n12822), .Q(g30388) );
  AND2X1 U13335 ( .IN1(n9144), .IN2(g2735), .Q(n12822) );
  AND3X1 U13336 ( .IN1(n12823), .IN2(n12019), .IN3(n3730), .Q(n12821) );
  INVX0 U13337 ( .INP(n12018), .ZN(n12019) );
  AND2X1 U13338 ( .IN1(g2741), .IN2(n9510), .Q(n12018) );
  OR2X1 U13339 ( .IN1(n9510), .IN2(g2741), .Q(n12823) );
  AND2X1 U13340 ( .IN1(g2735), .IN2(n12824), .Q(n9510) );
  OR3X1 U13341 ( .IN1(n12825), .IN2(n12826), .IN3(n12827), .Q(g30387) );
  AND2X1 U13342 ( .IN1(n12828), .IN2(n9262), .Q(n12827) );
  AND3X1 U13343 ( .IN1(n12829), .IN2(n5457), .IN3(n5777), .Q(n12826) );
  AND2X1 U13344 ( .IN1(n12830), .IN2(g2681), .Q(n12825) );
  OR2X1 U13345 ( .IN1(n9124), .IN2(n12831), .Q(n12830) );
  AND2X1 U13346 ( .IN1(n12832), .IN2(g2675), .Q(n12831) );
  OR2X1 U13347 ( .IN1(n12833), .IN2(n12834), .Q(g30386) );
  AND2X1 U13348 ( .IN1(n12835), .IN2(g2675), .Q(n12834) );
  AND2X1 U13349 ( .IN1(n12828), .IN2(g2681), .Q(n12833) );
  OR3X1 U13350 ( .IN1(n12836), .IN2(n12837), .IN3(n12838), .Q(g30385) );
  AND2X1 U13351 ( .IN1(n9144), .IN2(g2657), .Q(n12838) );
  AND2X1 U13352 ( .IN1(n12829), .IN2(n5418), .Q(n12837) );
  AND2X1 U13353 ( .IN1(n12828), .IN2(g2661), .Q(n12836) );
  INVX0 U13354 ( .INP(n12835), .ZN(n12828) );
  OR2X1 U13355 ( .IN1(n9133), .IN2(n12832), .Q(n12835) );
  OR3X1 U13356 ( .IN1(n12839), .IN2(n12840), .IN3(n12841), .Q(g30384) );
  AND2X1 U13357 ( .IN1(n9144), .IN2(g2652), .Q(n12841) );
  AND2X1 U13358 ( .IN1(n12842), .IN2(g2657), .Q(n12840) );
  OR2X1 U13359 ( .IN1(n12843), .IN2(n11747), .Q(n12842) );
  AND2X1 U13360 ( .IN1(n9033), .IN2(n11758), .Q(n12843) );
  AND3X1 U13361 ( .IN1(n3517), .IN2(n12844), .IN3(n8808), .Q(n12839) );
  OR2X1 U13362 ( .IN1(n12845), .IN2(n12846), .Q(n12844) );
  AND2X1 U13363 ( .IN1(n8333), .IN2(g2652), .Q(n12846) );
  AND2X1 U13364 ( .IN1(n8622), .IN2(g2648), .Q(n12845) );
  OR3X1 U13365 ( .IN1(n12847), .IN2(n12848), .IN3(n12849), .Q(g30383) );
  AND2X1 U13366 ( .IN1(test_so66), .IN2(n9139), .Q(n12849) );
  AND2X1 U13367 ( .IN1(test_so34), .IN2(n12850), .Q(n12848) );
  OR2X1 U13368 ( .IN1(n12851), .IN2(n11747), .Q(n12850) );
  INVX0 U13369 ( .INP(n12852), .ZN(n12851) );
  OR2X1 U13370 ( .IN1(n10391), .IN2(n9122), .Q(n12852) );
  AND3X1 U13371 ( .IN1(n10391), .IN2(n10509), .IN3(n3517), .Q(n12847) );
  OR2X1 U13372 ( .IN1(n5524), .IN2(g2555), .Q(n10509) );
  OR3X1 U13373 ( .IN1(n12853), .IN2(n12854), .IN3(n12855), .Q(g30382) );
  AND2X1 U13374 ( .IN1(n12856), .IN2(n9295), .Q(n12855) );
  AND3X1 U13375 ( .IN1(n12857), .IN2(n5461), .IN3(n5782), .Q(n12854) );
  AND2X1 U13376 ( .IN1(n12858), .IN2(g2547), .Q(n12853) );
  OR2X1 U13377 ( .IN1(n9129), .IN2(n12859), .Q(n12858) );
  AND2X1 U13378 ( .IN1(n12860), .IN2(g2541), .Q(n12859) );
  OR2X1 U13379 ( .IN1(n12861), .IN2(n12862), .Q(g30381) );
  AND2X1 U13380 ( .IN1(n12863), .IN2(g2541), .Q(n12862) );
  AND2X1 U13381 ( .IN1(n12856), .IN2(g2547), .Q(n12861) );
  OR3X1 U13382 ( .IN1(n12864), .IN2(n12865), .IN3(n12866), .Q(g30380) );
  AND2X1 U13383 ( .IN1(n9144), .IN2(g2523), .Q(n12866) );
  AND2X1 U13384 ( .IN1(n12857), .IN2(n5420), .Q(n12865) );
  AND2X1 U13385 ( .IN1(n12856), .IN2(g2527), .Q(n12864) );
  INVX0 U13386 ( .INP(n12863), .ZN(n12856) );
  OR2X1 U13387 ( .IN1(n9129), .IN2(n12860), .Q(n12863) );
  OR3X1 U13388 ( .IN1(n12867), .IN2(n12868), .IN3(n12869), .Q(g30379) );
  AND2X1 U13389 ( .IN1(n9144), .IN2(g2518), .Q(n12869) );
  AND2X1 U13390 ( .IN1(n12870), .IN2(g2523), .Q(n12868) );
  OR2X1 U13391 ( .IN1(n12871), .IN2(n11766), .Q(n12870) );
  AND2X1 U13392 ( .IN1(n9034), .IN2(n11777), .Q(n12871) );
  AND3X1 U13393 ( .IN1(n3536), .IN2(n12872), .IN3(n8815), .Q(n12867) );
  OR2X1 U13394 ( .IN1(n12873), .IN2(n12874), .Q(n12872) );
  AND2X1 U13395 ( .IN1(n8330), .IN2(g2518), .Q(n12874) );
  AND2X1 U13396 ( .IN1(n8624), .IN2(g2514), .Q(n12873) );
  OR2X1 U13397 ( .IN1(n12875), .IN2(n12876), .Q(g30378) );
  AND2X1 U13398 ( .IN1(n12877), .IN2(n9022), .Q(n12876) );
  OR2X1 U13399 ( .IN1(n12878), .IN2(n12879), .Q(n12877) );
  AND2X1 U13400 ( .IN1(n12880), .IN2(n12881), .Q(n12879) );
  OR2X1 U13401 ( .IN1(n5523), .IN2(test_so79), .Q(n12881) );
  INVX0 U13402 ( .INP(n12882), .ZN(n12878) );
  OR2X1 U13403 ( .IN1(n12880), .IN2(n5840), .Q(n12882) );
  AND2X1 U13404 ( .IN1(n9144), .IN2(g2441), .Q(n12875) );
  OR3X1 U13405 ( .IN1(n12883), .IN2(n12884), .IN3(n12885), .Q(g30377) );
  AND2X1 U13406 ( .IN1(n12886), .IN2(n9324), .Q(n12885) );
  AND3X1 U13407 ( .IN1(n12887), .IN2(n5459), .IN3(n8863), .Q(n12884) );
  AND2X1 U13408 ( .IN1(test_so89), .IN2(n12888), .Q(n12883) );
  OR2X1 U13409 ( .IN1(n9129), .IN2(n12889), .Q(n12888) );
  AND2X1 U13410 ( .IN1(n12890), .IN2(g2407), .Q(n12889) );
  OR2X1 U13411 ( .IN1(n12891), .IN2(n12892), .Q(g30376) );
  AND2X1 U13412 ( .IN1(n12893), .IN2(g2407), .Q(n12892) );
  AND2X1 U13413 ( .IN1(test_so89), .IN2(n12886), .Q(n12891) );
  OR3X1 U13414 ( .IN1(n12894), .IN2(n12895), .IN3(n12896), .Q(g30375) );
  AND2X1 U13415 ( .IN1(n9144), .IN2(g2389), .Q(n12896) );
  AND2X1 U13416 ( .IN1(n12887), .IN2(n5421), .Q(n12895) );
  AND2X1 U13417 ( .IN1(n12886), .IN2(g2393), .Q(n12894) );
  INVX0 U13418 ( .INP(n12893), .ZN(n12886) );
  OR2X1 U13419 ( .IN1(n9129), .IN2(n12890), .Q(n12893) );
  OR3X1 U13420 ( .IN1(n12897), .IN2(n12898), .IN3(n12899), .Q(g30374) );
  AND2X1 U13421 ( .IN1(n9144), .IN2(g2384), .Q(n12899) );
  AND2X1 U13422 ( .IN1(n12900), .IN2(g2389), .Q(n12898) );
  OR2X1 U13423 ( .IN1(n12901), .IN2(n11785), .Q(n12900) );
  AND2X1 U13424 ( .IN1(n9033), .IN2(n11796), .Q(n12901) );
  AND3X1 U13425 ( .IN1(n3555), .IN2(n12902), .IN3(n8810), .Q(n12897) );
  OR2X1 U13426 ( .IN1(n12903), .IN2(n12904), .Q(n12902) );
  AND2X1 U13427 ( .IN1(n8329), .IN2(g2384), .Q(n12904) );
  AND2X1 U13428 ( .IN1(n8629), .IN2(g2380), .Q(n12903) );
  OR2X1 U13429 ( .IN1(n12905), .IN2(n12906), .Q(g30373) );
  AND2X1 U13430 ( .IN1(n12907), .IN2(n9021), .Q(n12906) );
  OR2X1 U13431 ( .IN1(n12908), .IN2(n12909), .Q(n12907) );
  AND2X1 U13432 ( .IN1(n12910), .IN2(n12911), .Q(n12909) );
  OR2X1 U13433 ( .IN1(n5513), .IN2(g2287), .Q(n12911) );
  INVX0 U13434 ( .INP(n12912), .ZN(n12908) );
  OR2X1 U13435 ( .IN1(n12910), .IN2(n5841), .Q(n12912) );
  AND2X1 U13436 ( .IN1(n9144), .IN2(g2307), .Q(n12905) );
  OR3X1 U13437 ( .IN1(n12913), .IN2(n12914), .IN3(n12915), .Q(g30372) );
  AND2X1 U13438 ( .IN1(n12916), .IN2(n9273), .Q(n12915) );
  AND3X1 U13439 ( .IN1(n12917), .IN2(n5458), .IN3(n5778), .Q(n12914) );
  AND2X1 U13440 ( .IN1(n12918), .IN2(g2279), .Q(n12913) );
  OR2X1 U13441 ( .IN1(n9130), .IN2(n12919), .Q(n12918) );
  AND2X1 U13442 ( .IN1(n12920), .IN2(g2273), .Q(n12919) );
  OR2X1 U13443 ( .IN1(n12921), .IN2(n12922), .Q(g30371) );
  AND2X1 U13444 ( .IN1(n12923), .IN2(g2273), .Q(n12922) );
  AND2X1 U13445 ( .IN1(n12916), .IN2(g2279), .Q(n12921) );
  OR3X1 U13446 ( .IN1(n12924), .IN2(n12925), .IN3(n12926), .Q(g30370) );
  AND2X1 U13447 ( .IN1(n9144), .IN2(g2255), .Q(n12926) );
  AND2X1 U13448 ( .IN1(n12917), .IN2(n5419), .Q(n12925) );
  AND2X1 U13449 ( .IN1(n12916), .IN2(g2259), .Q(n12924) );
  INVX0 U13450 ( .INP(n12923), .ZN(n12916) );
  OR2X1 U13451 ( .IN1(n9130), .IN2(n12920), .Q(n12923) );
  OR3X1 U13452 ( .IN1(n12927), .IN2(n12928), .IN3(n12929), .Q(g30369) );
  AND2X1 U13453 ( .IN1(n9144), .IN2(g2250), .Q(n12929) );
  AND2X1 U13454 ( .IN1(n12930), .IN2(g2255), .Q(n12928) );
  OR2X1 U13455 ( .IN1(n12931), .IN2(n11804), .Q(n12930) );
  AND2X1 U13456 ( .IN1(n9033), .IN2(n11815), .Q(n12931) );
  AND3X1 U13457 ( .IN1(n3574), .IN2(n12932), .IN3(n8816), .Q(n12927) );
  OR2X1 U13458 ( .IN1(n12933), .IN2(n12934), .Q(n12932) );
  AND2X1 U13459 ( .IN1(n8332), .IN2(g2250), .Q(n12934) );
  AND2X1 U13460 ( .IN1(n8633), .IN2(g2246), .Q(n12933) );
  OR2X1 U13461 ( .IN1(n12935), .IN2(n12936), .Q(g30368) );
  AND2X1 U13462 ( .IN1(n12937), .IN2(n9020), .Q(n12936) );
  OR2X1 U13463 ( .IN1(n12938), .IN2(n12939), .Q(n12937) );
  AND2X1 U13464 ( .IN1(n12940), .IN2(n12941), .Q(n12939) );
  OR2X1 U13465 ( .IN1(n5514), .IN2(g2153), .Q(n12941) );
  INVX0 U13466 ( .INP(n12942), .ZN(n12938) );
  OR2X1 U13467 ( .IN1(n12940), .IN2(n5839), .Q(n12942) );
  AND2X1 U13468 ( .IN1(n9144), .IN2(g2173), .Q(n12935) );
  OR3X1 U13469 ( .IN1(n12943), .IN2(n12944), .IN3(n12945), .Q(g30367) );
  AND2X1 U13470 ( .IN1(n12946), .IN2(g2126), .Q(n12945) );
  AND3X1 U13471 ( .IN1(n12947), .IN2(n5463), .IN3(n5784), .Q(n12944) );
  AND2X1 U13472 ( .IN1(n12948), .IN2(g2122), .Q(n12943) );
  OR2X1 U13473 ( .IN1(n9130), .IN2(n12949), .Q(n12948) );
  AND2X1 U13474 ( .IN1(n12950), .IN2(g2116), .Q(n12949) );
  OR2X1 U13475 ( .IN1(n12951), .IN2(n12952), .Q(g30366) );
  AND2X1 U13476 ( .IN1(n12953), .IN2(g2116), .Q(n12952) );
  AND2X1 U13477 ( .IN1(n12946), .IN2(g2122), .Q(n12951) );
  OR3X1 U13478 ( .IN1(n12954), .IN2(n12955), .IN3(n12956), .Q(g30365) );
  AND2X1 U13479 ( .IN1(n9143), .IN2(g2098), .Q(n12956) );
  AND2X1 U13480 ( .IN1(n12947), .IN2(n5666), .Q(n12955) );
  AND2X1 U13481 ( .IN1(n12946), .IN2(g2102), .Q(n12954) );
  INVX0 U13482 ( .INP(n12953), .ZN(n12946) );
  OR2X1 U13483 ( .IN1(n9130), .IN2(n12950), .Q(n12953) );
  OR3X1 U13484 ( .IN1(n12957), .IN2(n12958), .IN3(n12959), .Q(g30364) );
  AND2X1 U13485 ( .IN1(test_so78), .IN2(n9139), .Q(n12959) );
  AND2X1 U13486 ( .IN1(n12960), .IN2(g2098), .Q(n12958) );
  OR2X1 U13487 ( .IN1(n12961), .IN2(n11823), .Q(n12960) );
  AND2X1 U13488 ( .IN1(n9034), .IN2(n11834), .Q(n12961) );
  AND4X1 U13489 ( .IN1(n8818), .IN2(n3593), .IN3(n12962), .IN4(n12963), .Q(
        n12957) );
  OR2X1 U13490 ( .IN1(n8328), .IN2(n8833), .Q(n12963) );
  OR2X1 U13491 ( .IN1(test_so78), .IN2(g2089), .Q(n12962) );
  OR3X1 U13492 ( .IN1(n12964), .IN2(n12965), .IN3(n12966), .Q(g30363) );
  AND2X1 U13493 ( .IN1(n9143), .IN2(g2016), .Q(n12966) );
  AND2X1 U13494 ( .IN1(test_so59), .IN2(n12967), .Q(n12965) );
  OR2X1 U13495 ( .IN1(n12968), .IN2(n11823), .Q(n12967) );
  INVX0 U13496 ( .INP(n12969), .ZN(n12968) );
  OR2X1 U13497 ( .IN1(n10394), .IN2(n9122), .Q(n12969) );
  AND3X1 U13498 ( .IN1(n10394), .IN2(n10736), .IN3(n3593), .Q(n12964) );
  OR2X1 U13499 ( .IN1(n5505), .IN2(g1996), .Q(n10736) );
  OR3X1 U13500 ( .IN1(n12970), .IN2(n12971), .IN3(n12972), .Q(g30362) );
  AND2X1 U13501 ( .IN1(n12973), .IN2(g1992), .Q(n12972) );
  AND3X1 U13502 ( .IN1(n12974), .IN2(n5462), .IN3(n5783), .Q(n12971) );
  AND2X1 U13503 ( .IN1(n12975), .IN2(g1988), .Q(n12970) );
  OR2X1 U13504 ( .IN1(n9130), .IN2(n12976), .Q(n12975) );
  AND2X1 U13505 ( .IN1(n12977), .IN2(g1982), .Q(n12976) );
  OR2X1 U13506 ( .IN1(n12978), .IN2(n12979), .Q(g30361) );
  AND2X1 U13507 ( .IN1(n12980), .IN2(g1982), .Q(n12979) );
  AND2X1 U13508 ( .IN1(n12973), .IN2(g1988), .Q(n12978) );
  OR3X1 U13509 ( .IN1(n12981), .IN2(n12982), .IN3(n12983), .Q(g30360) );
  AND2X1 U13510 ( .IN1(n9143), .IN2(g1964), .Q(n12983) );
  AND2X1 U13511 ( .IN1(n12974), .IN2(n5664), .Q(n12982) );
  AND2X1 U13512 ( .IN1(n12973), .IN2(g1968), .Q(n12981) );
  INVX0 U13513 ( .INP(n12980), .ZN(n12973) );
  OR2X1 U13514 ( .IN1(n9130), .IN2(n12977), .Q(n12980) );
  OR3X1 U13515 ( .IN1(n12984), .IN2(n12985), .IN3(n12986), .Q(g30359) );
  AND2X1 U13516 ( .IN1(n9143), .IN2(g1959), .Q(n12986) );
  AND2X1 U13517 ( .IN1(n12987), .IN2(g1964), .Q(n12985) );
  OR2X1 U13518 ( .IN1(n12988), .IN2(n11842), .Q(n12987) );
  AND2X1 U13519 ( .IN1(n9034), .IN2(n11854), .Q(n12988) );
  AND3X1 U13520 ( .IN1(n3611), .IN2(n12989), .IN3(n8807), .Q(n12984) );
  OR2X1 U13521 ( .IN1(n12990), .IN2(n12991), .Q(n12989) );
  AND2X1 U13522 ( .IN1(n8326), .IN2(g1959), .Q(n12991) );
  AND2X1 U13523 ( .IN1(n8625), .IN2(g1955), .Q(n12990) );
  OR2X1 U13524 ( .IN1(n12992), .IN2(n12993), .Q(g30358) );
  AND2X1 U13525 ( .IN1(n12994), .IN2(n9015), .Q(n12993) );
  OR2X1 U13526 ( .IN1(n12995), .IN2(n12996), .Q(n12994) );
  AND2X1 U13527 ( .IN1(n12997), .IN2(n12998), .Q(n12996) );
  OR2X1 U13528 ( .IN1(n5503), .IN2(test_so8), .Q(n12998) );
  INVX0 U13529 ( .INP(n12999), .ZN(n12995) );
  OR2X1 U13530 ( .IN1(n12997), .IN2(n5837), .Q(n12999) );
  AND2X1 U13531 ( .IN1(n9143), .IN2(g1882), .Q(n12992) );
  OR3X1 U13532 ( .IN1(n13000), .IN2(n13001), .IN3(n13002), .Q(g30357) );
  AND2X1 U13533 ( .IN1(n13003), .IN2(g1858), .Q(n13002) );
  AND3X1 U13534 ( .IN1(n13004), .IN2(n5464), .IN3(n5785), .Q(n13001) );
  AND2X1 U13535 ( .IN1(n13005), .IN2(g1854), .Q(n13000) );
  OR2X1 U13536 ( .IN1(n9130), .IN2(n13006), .Q(n13005) );
  AND2X1 U13537 ( .IN1(n13007), .IN2(g1848), .Q(n13006) );
  OR2X1 U13538 ( .IN1(n13008), .IN2(n13009), .Q(g30356) );
  AND2X1 U13539 ( .IN1(n13010), .IN2(g1848), .Q(n13009) );
  AND2X1 U13540 ( .IN1(n13003), .IN2(g1854), .Q(n13008) );
  OR3X1 U13541 ( .IN1(n13011), .IN2(n13012), .IN3(n13013), .Q(g30355) );
  AND2X1 U13542 ( .IN1(n9143), .IN2(g1830), .Q(n13013) );
  AND2X1 U13543 ( .IN1(n13004), .IN2(n5665), .Q(n13012) );
  AND2X1 U13544 ( .IN1(n13003), .IN2(g1834), .Q(n13011) );
  INVX0 U13545 ( .INP(n13010), .ZN(n13003) );
  OR2X1 U13546 ( .IN1(n9130), .IN2(n13007), .Q(n13010) );
  OR3X1 U13547 ( .IN1(n13014), .IN2(n13015), .IN3(n13016), .Q(g30354) );
  AND2X1 U13548 ( .IN1(n9143), .IN2(g1825), .Q(n13016) );
  AND2X1 U13549 ( .IN1(n13017), .IN2(g1830), .Q(n13015) );
  OR2X1 U13550 ( .IN1(n13018), .IN2(n11862), .Q(n13017) );
  AND2X1 U13551 ( .IN1(n9032), .IN2(n11873), .Q(n13018) );
  AND3X1 U13552 ( .IN1(n3628), .IN2(n13019), .IN3(n8813), .Q(n13014) );
  OR2X1 U13553 ( .IN1(n13020), .IN2(n13021), .Q(n13019) );
  AND2X1 U13554 ( .IN1(n8327), .IN2(g1825), .Q(n13021) );
  AND2X1 U13555 ( .IN1(n8631), .IN2(g1821), .Q(n13020) );
  OR2X1 U13556 ( .IN1(n13022), .IN2(n13023), .Q(g30353) );
  AND2X1 U13557 ( .IN1(n13024), .IN2(n9018), .Q(n13023) );
  OR2X1 U13558 ( .IN1(n13025), .IN2(n13026), .Q(n13024) );
  AND2X1 U13559 ( .IN1(n13027), .IN2(n13028), .Q(n13026) );
  OR2X1 U13560 ( .IN1(n5504), .IN2(g1728), .Q(n13028) );
  INVX0 U13561 ( .INP(n13029), .ZN(n13025) );
  OR2X1 U13562 ( .IN1(n13027), .IN2(n5834), .Q(n13029) );
  AND2X1 U13563 ( .IN1(n9143), .IN2(g1748), .Q(n13022) );
  OR3X1 U13564 ( .IN1(n13030), .IN2(n13031), .IN3(n13032), .Q(g30352) );
  AND2X1 U13565 ( .IN1(n13033), .IN2(n9236), .Q(n13032) );
  AND4X1 U13566 ( .IN1(n5460), .IN2(n9082), .IN3(n13034), .IN4(n5780), .Q(
        n13031) );
  AND2X1 U13567 ( .IN1(n13035), .IN2(g1720), .Q(n13030) );
  OR2X1 U13568 ( .IN1(n9130), .IN2(n13036), .Q(n13035) );
  AND2X1 U13569 ( .IN1(n13034), .IN2(g1714), .Q(n13036) );
  OR2X1 U13570 ( .IN1(n13037), .IN2(n13038), .Q(g30351) );
  AND2X1 U13571 ( .IN1(n13039), .IN2(g1714), .Q(n13038) );
  AND2X1 U13572 ( .IN1(n13033), .IN2(g1720), .Q(n13037) );
  OR3X1 U13573 ( .IN1(n13040), .IN2(n13041), .IN3(n13042), .Q(g30350) );
  AND2X1 U13574 ( .IN1(n13033), .IN2(g1700), .Q(n13042) );
  INVX0 U13575 ( .INP(n13039), .ZN(n13033) );
  OR2X1 U13576 ( .IN1(n9130), .IN2(n13034), .Q(n13039) );
  AND2X1 U13577 ( .IN1(n9143), .IN2(g1696), .Q(n13041) );
  AND3X1 U13578 ( .IN1(n13034), .IN2(n5417), .IN3(n9066), .Q(n13040) );
  OR3X1 U13579 ( .IN1(n13043), .IN2(n13044), .IN3(n13045), .Q(g30349) );
  AND2X1 U13580 ( .IN1(n9143), .IN2(g1691), .Q(n13045) );
  AND2X1 U13581 ( .IN1(n13046), .IN2(g1696), .Q(n13044) );
  OR2X1 U13582 ( .IN1(n13047), .IN2(n11881), .Q(n13046) );
  AND2X1 U13583 ( .IN1(n9047), .IN2(n11898), .Q(n13047) );
  AND3X1 U13584 ( .IN1(n3646), .IN2(n13048), .IN3(n8817), .Q(n13043) );
  OR2X1 U13585 ( .IN1(n13049), .IN2(n13050), .Q(n13048) );
  AND2X1 U13586 ( .IN1(n8331), .IN2(g1691), .Q(n13050) );
  AND2X1 U13587 ( .IN1(n8627), .IN2(g1687), .Q(n13049) );
  OR3X1 U13588 ( .IN1(n13051), .IN2(n13052), .IN3(n13053), .Q(g30348) );
  AND2X1 U13589 ( .IN1(n9143), .IN2(g1612), .Q(n13053) );
  AND2X1 U13590 ( .IN1(n13054), .IN2(g1632), .Q(n13052) );
  OR2X1 U13591 ( .IN1(n13055), .IN2(n11881), .Q(n13054) );
  INVX0 U13592 ( .INP(n13056), .ZN(n13055) );
  OR2X1 U13593 ( .IN1(g25167), .IN2(n9122), .Q(n13056) );
  AND3X1 U13594 ( .IN1(g25167), .IN2(n13057), .IN3(n3646), .Q(n13051) );
  OR2X1 U13595 ( .IN1(n5549), .IN2(g1592), .Q(n13057) );
  OR2X1 U13596 ( .IN1(n13058), .IN2(n13059), .Q(g30347) );
  INVX0 U13597 ( .INP(n13060), .ZN(n13059) );
  OR2X1 U13598 ( .IN1(n9007), .IN2(n8378), .Q(n13060) );
  AND3X1 U13599 ( .IN1(n13061), .IN2(n13062), .IN3(n13063), .Q(n13058) );
  INVX0 U13600 ( .INP(n13064), .ZN(n13061) );
  AND2X1 U13601 ( .IN1(n13065), .IN2(n13066), .Q(n13064) );
  OR2X1 U13602 ( .IN1(n9130), .IN2(n8791), .Q(n13066) );
  OR2X1 U13603 ( .IN1(n13067), .IN2(n13068), .Q(g30346) );
  AND4X1 U13604 ( .IN1(n13069), .IN2(n13065), .IN3(n13063), .IN4(n9050), .Q(
        n13068) );
  INVX0 U13605 ( .INP(n13070), .ZN(n13063) );
  INVX0 U13606 ( .INP(n13071), .ZN(n13069) );
  AND2X1 U13607 ( .IN1(n13072), .IN2(n8378), .Q(n13071) );
  AND2X1 U13608 ( .IN1(n9143), .IN2(g1536), .Q(n13067) );
  OR2X1 U13609 ( .IN1(n13073), .IN2(n13074), .Q(g30345) );
  AND2X1 U13610 ( .IN1(n13075), .IN2(g1514), .Q(n13074) );
  OR2X1 U13611 ( .IN1(n9130), .IN2(n13076), .Q(n13075) );
  AND2X1 U13612 ( .IN1(n13077), .IN2(n13078), .Q(n13076) );
  OR2X1 U13613 ( .IN1(n5302), .IN2(n8819), .Q(n13078) );
  OR2X1 U13614 ( .IN1(test_so49), .IN2(g7946), .Q(n13077) );
  AND2X1 U13615 ( .IN1(n13079), .IN2(n9018), .Q(n13073) );
  OR2X1 U13616 ( .IN1(n11258), .IN2(n13070), .Q(n13079) );
  AND2X1 U13617 ( .IN1(n13080), .IN2(n9020), .Q(g30344) );
  OR3X1 U13618 ( .IN1(n13081), .IN2(n13082), .IN3(n13070), .Q(n13080) );
  OR2X1 U13619 ( .IN1(n13083), .IN2(n4173), .Q(n13070) );
  AND2X1 U13620 ( .IN1(n4172), .IN2(n11258), .Q(n13083) );
  AND3X1 U13621 ( .IN1(n13084), .IN2(g7946), .IN3(n4895), .Q(n4172) );
  AND2X1 U13622 ( .IN1(n5302), .IN2(g1514), .Q(n13082) );
  AND2X1 U13623 ( .IN1(n5364), .IN2(g7946), .Q(n13081) );
  OR3X1 U13624 ( .IN1(n13085), .IN2(n13086), .IN3(n13087), .Q(g30343) );
  AND2X1 U13625 ( .IN1(n4175), .IN2(n11902), .Q(n13087) );
  AND3X1 U13626 ( .IN1(n9493), .IN2(g1361), .IN3(n9066), .Q(n13086) );
  OR2X1 U13627 ( .IN1(n13088), .IN2(n13089), .Q(n9493) );
  AND2X1 U13628 ( .IN1(n8799), .IN2(n11477), .Q(n13088) );
  AND2X1 U13629 ( .IN1(n9143), .IN2(g1345), .Q(n13085) );
  OR3X1 U13630 ( .IN1(n13090), .IN2(n13091), .IN3(n13092), .Q(g30342) );
  AND2X1 U13631 ( .IN1(n9143), .IN2(g1256), .Q(n13092) );
  AND2X1 U13632 ( .IN1(n3736), .IN2(n5553), .Q(n13091) );
  AND3X1 U13633 ( .IN1(n11485), .IN2(n13093), .IN3(g1259), .Q(n13090) );
  INVX0 U13634 ( .INP(n3736), .ZN(n13093) );
  OR2X1 U13635 ( .IN1(n13094), .IN2(n13095), .Q(g30341) );
  INVX0 U13636 ( .INP(n13096), .ZN(n13095) );
  OR2X1 U13637 ( .IN1(n9007), .IN2(n8379), .Q(n13096) );
  AND3X1 U13638 ( .IN1(n13097), .IN2(n13098), .IN3(n13099), .Q(n13094) );
  INVX0 U13639 ( .INP(n13100), .ZN(n13097) );
  AND2X1 U13640 ( .IN1(n13101), .IN2(n13102), .Q(n13100) );
  OR2X1 U13641 ( .IN1(n9130), .IN2(n8792), .Q(n13102) );
  OR2X1 U13642 ( .IN1(n13103), .IN2(n13104), .Q(g30340) );
  AND4X1 U13643 ( .IN1(n13105), .IN2(n13101), .IN3(n13099), .IN4(n9050), .Q(
        n13104) );
  INVX0 U13644 ( .INP(n13106), .ZN(n13099) );
  INVX0 U13645 ( .INP(n13107), .ZN(n13105) );
  AND2X1 U13646 ( .IN1(n13108), .IN2(n8379), .Q(n13107) );
  AND2X1 U13647 ( .IN1(n9143), .IN2(g1193), .Q(n13103) );
  OR2X1 U13648 ( .IN1(n13109), .IN2(n13110), .Q(g30339) );
  AND2X1 U13649 ( .IN1(n13111), .IN2(g1171), .Q(n13110) );
  OR3X1 U13650 ( .IN1(n13112), .IN2(n13113), .IN3(n9121), .Q(n13111) );
  AND2X1 U13651 ( .IN1(n5304), .IN2(g1183), .Q(n13113) );
  AND2X1 U13652 ( .IN1(n5599), .IN2(g7916), .Q(n13112) );
  AND2X1 U13653 ( .IN1(n13114), .IN2(n9021), .Q(n13109) );
  OR2X1 U13654 ( .IN1(n11430), .IN2(n13106), .Q(n13114) );
  AND2X1 U13655 ( .IN1(n13115), .IN2(n9021), .Q(g30338) );
  OR3X1 U13656 ( .IN1(n13116), .IN2(n13117), .IN3(n13106), .Q(n13115) );
  OR2X1 U13657 ( .IN1(n13118), .IN2(n4191), .Q(n13106) );
  AND2X1 U13658 ( .IN1(n4190), .IN2(n11430), .Q(n13118) );
  AND3X1 U13659 ( .IN1(n13119), .IN2(g7916), .IN3(n4920), .Q(n4190) );
  AND2X1 U13660 ( .IN1(n5304), .IN2(g1171), .Q(n13117) );
  AND2X1 U13661 ( .IN1(n5363), .IN2(g7916), .Q(n13116) );
  OR3X1 U13662 ( .IN1(n13120), .IN2(n13121), .IN3(n13122), .Q(g30337) );
  AND2X1 U13663 ( .IN1(n4193), .IN2(n11913), .Q(n13122) );
  AND3X1 U13664 ( .IN1(n9370), .IN2(g1018), .IN3(n9066), .Q(n13121) );
  OR2X1 U13665 ( .IN1(n13123), .IN2(n13124), .Q(n9370) );
  AND2X1 U13666 ( .IN1(n8796), .IN2(n11492), .Q(n13123) );
  AND2X1 U13667 ( .IN1(n9143), .IN2(g1002), .Q(n13120) );
  OR3X1 U13668 ( .IN1(n13125), .IN2(n13126), .IN3(n13127), .Q(g30336) );
  AND2X1 U13669 ( .IN1(n9143), .IN2(g911), .Q(n13127) );
  AND2X1 U13670 ( .IN1(n3741), .IN2(n5560), .Q(n13126) );
  AND3X1 U13671 ( .IN1(n11500), .IN2(n13128), .IN3(g914), .Q(n13125) );
  INVX0 U13672 ( .INP(n3741), .ZN(n13128) );
  OR3X1 U13673 ( .IN1(n13129), .IN2(n13130), .IN3(n13131), .Q(g30335) );
  AND2X1 U13674 ( .IN1(test_so60), .IN2(n9138), .Q(n13131) );
  AND2X1 U13675 ( .IN1(n3743), .IN2(n5470), .Q(n13130) );
  AND3X1 U13676 ( .IN1(n2404), .IN2(n13132), .IN3(g744), .Q(n13129) );
  INVX0 U13677 ( .INP(n3743), .ZN(n13132) );
  AND3X1 U13678 ( .IN1(n4198), .IN2(test_so60), .IN3(n13133), .Q(n3743) );
  OR2X1 U13679 ( .IN1(n5482), .IN2(g736), .Q(n4198) );
  OR3X1 U13680 ( .IN1(n13134), .IN2(n13135), .IN3(n13136), .Q(g30334) );
  AND2X1 U13681 ( .IN1(n9143), .IN2(g586), .Q(n13136) );
  AND2X1 U13682 ( .IN1(n3745), .IN2(n5294), .Q(n13135) );
  AND3X1 U13683 ( .IN1(n2421), .IN2(n13137), .IN3(g577), .Q(n13134) );
  INVX0 U13684 ( .INP(n3745), .ZN(n13137) );
  OR2X1 U13685 ( .IN1(n13138), .IN2(n13139), .Q(g30333) );
  AND2X1 U13686 ( .IN1(n9143), .IN2(g142), .Q(n13139) );
  AND2X1 U13687 ( .IN1(n10380), .IN2(n13140), .Q(n13138) );
  OR2X1 U13688 ( .IN1(n13141), .IN2(n13142), .Q(n13140) );
  INVX0 U13689 ( .INP(n13143), .ZN(n13142) );
  OR2X1 U13690 ( .IN1(n13144), .IN2(test_so73), .Q(n13143) );
  AND2X1 U13691 ( .IN1(test_so73), .IN2(n13144), .Q(n13141) );
  AND2X1 U13692 ( .IN1(n9047), .IN2(n12053), .Q(n10380) );
  AND3X1 U13693 ( .IN1(g691), .IN2(n13145), .IN3(n13146), .Q(n12053) );
  OR2X1 U13694 ( .IN1(n13144), .IN2(n13147), .Q(n13146) );
  AND3X1 U13695 ( .IN1(n8834), .IN2(n5402), .IN3(n5606), .Q(n13147) );
  OR3X1 U13696 ( .IN1(n13148), .IN2(n13149), .IN3(n13150), .Q(g29309) );
  AND2X1 U13697 ( .IN1(n3765), .IN2(n13151), .Q(n13150) );
  OR2X1 U13698 ( .IN1(n10979), .IN2(n5739), .Q(n13151) );
  AND3X1 U13699 ( .IN1(n9449), .IN2(g6541), .IN3(n12080), .Q(n13149) );
  OR3X1 U13700 ( .IN1(n13152), .IN2(n13153), .IN3(n13154), .Q(g29308) );
  AND2X1 U13701 ( .IN1(n9142), .IN2(g6523), .Q(n13154) );
  AND2X1 U13702 ( .IN1(n5659), .IN2(n13155), .Q(n13153) );
  AND2X1 U13703 ( .IN1(n13156), .IN2(g6527), .Q(n13152) );
  OR3X1 U13704 ( .IN1(n13157), .IN2(n13158), .IN3(n13159), .Q(g29307) );
  AND2X1 U13705 ( .IN1(n13156), .IN2(g6523), .Q(n13159) );
  AND3X1 U13706 ( .IN1(n5426), .IN2(n13155), .IN3(n5806), .Q(n13158) );
  AND2X1 U13707 ( .IN1(n13160), .IN2(g6519), .Q(n13157) );
  OR2X1 U13708 ( .IN1(n9131), .IN2(n13161), .Q(n13160) );
  AND2X1 U13709 ( .IN1(n13162), .IN2(g6513), .Q(n13161) );
  OR2X1 U13710 ( .IN1(n13163), .IN2(n13164), .Q(g29306) );
  AND2X1 U13711 ( .IN1(n13165), .IN2(g6513), .Q(n13164) );
  AND2X1 U13712 ( .IN1(n13156), .IN2(g6519), .Q(n13163) );
  INVX0 U13713 ( .INP(n13165), .ZN(n13156) );
  OR2X1 U13714 ( .IN1(n9131), .IN2(n13162), .Q(n13165) );
  OR3X1 U13715 ( .IN1(n13166), .IN2(n13167), .IN3(n13168), .Q(g29305) );
  INVX0 U13716 ( .INP(n13169), .ZN(n13168) );
  OR2X1 U13717 ( .IN1(n12060), .IN2(n13162), .Q(n13169) );
  OR2X1 U13718 ( .IN1(n8737), .IN2(n9123), .Q(n12060) );
  AND3X1 U13719 ( .IN1(n13155), .IN2(g6505), .IN3(n5748), .Q(n13167) );
  AND2X1 U13720 ( .IN1(n9046), .IN2(n13162), .Q(n13155) );
  AND2X1 U13721 ( .IN1(n13170), .IN2(g6500), .Q(n13166) );
  OR2X1 U13722 ( .IN1(n9131), .IN2(n13171), .Q(n13170) );
  AND2X1 U13723 ( .IN1(n8695), .IN2(n13162), .Q(n13171) );
  OR3X1 U13724 ( .IN1(n13172), .IN2(n13173), .IN3(n13174), .Q(g29304) );
  AND2X1 U13725 ( .IN1(n11010), .IN2(g6500), .Q(n13174) );
  AND3X1 U13726 ( .IN1(n13175), .IN2(n13176), .IN3(n9066), .Q(n13173) );
  OR2X1 U13727 ( .IN1(n13177), .IN2(n13162), .Q(n13176) );
  AND2X1 U13728 ( .IN1(n11004), .IN2(n13178), .Q(n13162) );
  INVX0 U13729 ( .INP(n13179), .ZN(n13177) );
  OR2X1 U13730 ( .IN1(n13180), .IN2(n8809), .Q(n13179) );
  AND2X1 U13731 ( .IN1(g6500), .IN2(n13181), .Q(n13180) );
  OR2X1 U13732 ( .IN1(n13182), .IN2(n13181), .Q(n13175) );
  INVX0 U13733 ( .INP(n13183), .ZN(n13182) );
  OR2X1 U13734 ( .IN1(n13178), .IN2(n5748), .Q(n13183) );
  AND3X1 U13735 ( .IN1(g17722), .IN2(g6727), .IN3(n9366), .Q(n13178) );
  AND2X1 U13736 ( .IN1(n9142), .IN2(g6505), .Q(n13172) );
  OR3X1 U13737 ( .IN1(n13148), .IN2(n13184), .IN3(n13185), .Q(g29303) );
  AND2X1 U13738 ( .IN1(n3765), .IN2(n13186), .Q(n13185) );
  OR2X1 U13739 ( .IN1(n10991), .IN2(n5741), .Q(n13186) );
  AND3X1 U13740 ( .IN1(n9449), .IN2(g6195), .IN3(n12167), .Q(n13184) );
  OR3X1 U13741 ( .IN1(n13187), .IN2(n13188), .IN3(n13189), .Q(g29302) );
  AND2X1 U13742 ( .IN1(n9142), .IN2(g6177), .Q(n13189) );
  AND2X1 U13743 ( .IN1(n5667), .IN2(n13190), .Q(n13188) );
  AND2X1 U13744 ( .IN1(n13191), .IN2(g6181), .Q(n13187) );
  OR3X1 U13745 ( .IN1(n13192), .IN2(n13193), .IN3(n13194), .Q(g29301) );
  AND2X1 U13746 ( .IN1(n13191), .IN2(g6177), .Q(n13194) );
  AND3X1 U13747 ( .IN1(n5430), .IN2(n13190), .IN3(n5810), .Q(n13193) );
  AND2X1 U13748 ( .IN1(n13195), .IN2(g6173), .Q(n13192) );
  OR2X1 U13749 ( .IN1(n9131), .IN2(n13196), .Q(n13195) );
  AND2X1 U13750 ( .IN1(n13197), .IN2(g6167), .Q(n13196) );
  OR2X1 U13751 ( .IN1(n13198), .IN2(n13199), .Q(g29300) );
  AND2X1 U13752 ( .IN1(n13200), .IN2(g6167), .Q(n13199) );
  AND2X1 U13753 ( .IN1(n13191), .IN2(g6173), .Q(n13198) );
  INVX0 U13754 ( .INP(n13200), .ZN(n13191) );
  OR2X1 U13755 ( .IN1(n9131), .IN2(n13197), .Q(n13200) );
  OR3X1 U13756 ( .IN1(n13201), .IN2(n13202), .IN3(n13203), .Q(g29299) );
  INVX0 U13757 ( .INP(n13204), .ZN(n13203) );
  OR2X1 U13758 ( .IN1(n12071), .IN2(n13197), .Q(n13204) );
  OR2X1 U13759 ( .IN1(n8781), .IN2(n9123), .Q(n12071) );
  AND3X1 U13760 ( .IN1(n13190), .IN2(g6159), .IN3(n5747), .Q(n13202) );
  AND2X1 U13761 ( .IN1(n9047), .IN2(n13197), .Q(n13190) );
  AND2X1 U13762 ( .IN1(n13205), .IN2(g6154), .Q(n13201) );
  OR2X1 U13763 ( .IN1(n9131), .IN2(n13206), .Q(n13205) );
  AND2X1 U13764 ( .IN1(n8696), .IN2(n13197), .Q(n13206) );
  OR3X1 U13765 ( .IN1(n13207), .IN2(n13208), .IN3(n13209), .Q(g29298) );
  AND2X1 U13766 ( .IN1(n11027), .IN2(g6154), .Q(n13209) );
  AND3X1 U13767 ( .IN1(n13210), .IN2(n13211), .IN3(n9066), .Q(n13208) );
  OR2X1 U13768 ( .IN1(n13212), .IN2(n13197), .Q(n13211) );
  AND2X1 U13769 ( .IN1(n11019), .IN2(n13213), .Q(n13197) );
  INVX0 U13770 ( .INP(n13214), .ZN(n13212) );
  OR2X1 U13771 ( .IN1(n11023), .IN2(n13215), .Q(n13214) );
  AND2X1 U13772 ( .IN1(g6154), .IN2(n13216), .Q(n13215) );
  OR2X1 U13773 ( .IN1(n13217), .IN2(n13216), .Q(n13210) );
  INVX0 U13774 ( .INP(n13218), .ZN(n13217) );
  OR2X1 U13775 ( .IN1(n13213), .IN2(n5747), .Q(n13218) );
  AND3X1 U13776 ( .IN1(g17685), .IN2(n10232), .IN3(test_so69), .Q(n13213) );
  AND2X1 U13777 ( .IN1(n9142), .IN2(g6159), .Q(n13207) );
  OR3X1 U13778 ( .IN1(n13148), .IN2(n13219), .IN3(n13220), .Q(g29297) );
  AND2X1 U13779 ( .IN1(n3765), .IN2(n13221), .Q(n13220) );
  OR2X1 U13780 ( .IN1(n10990), .IN2(n5736), .Q(n13221) );
  AND3X1 U13781 ( .IN1(n9449), .IN2(g5849), .IN3(n12253), .Q(n13219) );
  OR3X1 U13782 ( .IN1(n13222), .IN2(n13223), .IN3(n13224), .Q(g29296) );
  AND2X1 U13783 ( .IN1(n9142), .IN2(g5831), .Q(n13224) );
  AND2X1 U13784 ( .IN1(n5663), .IN2(n13225), .Q(n13223) );
  AND2X1 U13785 ( .IN1(n13226), .IN2(g5835), .Q(n13222) );
  OR3X1 U13786 ( .IN1(n13227), .IN2(n13228), .IN3(n13229), .Q(g29295) );
  AND2X1 U13787 ( .IN1(n13226), .IN2(g5831), .Q(n13229) );
  AND3X1 U13788 ( .IN1(n5429), .IN2(n13225), .IN3(n5809), .Q(n13228) );
  AND2X1 U13789 ( .IN1(n13230), .IN2(g5827), .Q(n13227) );
  OR2X1 U13790 ( .IN1(n9131), .IN2(n13231), .Q(n13230) );
  AND2X1 U13791 ( .IN1(n13232), .IN2(g5821), .Q(n13231) );
  OR2X1 U13792 ( .IN1(n13233), .IN2(n13234), .Q(g29294) );
  AND2X1 U13793 ( .IN1(n13235), .IN2(g5821), .Q(n13234) );
  AND2X1 U13794 ( .IN1(n13226), .IN2(g5827), .Q(n13233) );
  INVX0 U13795 ( .INP(n13235), .ZN(n13226) );
  OR2X1 U13796 ( .IN1(n9131), .IN2(n13232), .Q(n13235) );
  OR3X1 U13797 ( .IN1(n13236), .IN2(n13237), .IN3(n13238), .Q(g29293) );
  INVX0 U13798 ( .INP(n13239), .ZN(n13238) );
  OR2X1 U13799 ( .IN1(n12072), .IN2(n13232), .Q(n13239) );
  OR2X1 U13800 ( .IN1(n8782), .IN2(n9123), .Q(n12072) );
  AND3X1 U13801 ( .IN1(n13225), .IN2(g5813), .IN3(n5749), .Q(n13237) );
  AND2X1 U13802 ( .IN1(n9043), .IN2(n13232), .Q(n13225) );
  AND2X1 U13803 ( .IN1(n13240), .IN2(g5808), .Q(n13236) );
  OR2X1 U13804 ( .IN1(n9131), .IN2(n13241), .Q(n13240) );
  AND2X1 U13805 ( .IN1(n8694), .IN2(n13232), .Q(n13241) );
  OR3X1 U13806 ( .IN1(n13242), .IN2(n13243), .IN3(n13244), .Q(g29292) );
  AND2X1 U13807 ( .IN1(n11044), .IN2(g5808), .Q(n13244) );
  AND3X1 U13808 ( .IN1(n13245), .IN2(n13246), .IN3(n9078), .Q(n13243) );
  OR2X1 U13809 ( .IN1(n13247), .IN2(n13232), .Q(n13246) );
  AND2X1 U13810 ( .IN1(n11036), .IN2(n13248), .Q(n13232) );
  INVX0 U13811 ( .INP(n13249), .ZN(n13247) );
  OR2X1 U13812 ( .IN1(n11040), .IN2(n13250), .Q(n13249) );
  AND2X1 U13813 ( .IN1(g5808), .IN2(n13251), .Q(n13250) );
  OR2X1 U13814 ( .IN1(n13252), .IN2(n13251), .Q(n13245) );
  INVX0 U13815 ( .INP(n13253), .ZN(n13252) );
  OR2X1 U13816 ( .IN1(n13248), .IN2(n5749), .Q(n13253) );
  AND3X1 U13817 ( .IN1(g17646), .IN2(g6035), .IN3(n10245), .Q(n13248) );
  AND2X1 U13818 ( .IN1(n9142), .IN2(g5813), .Q(n13242) );
  OR3X1 U13819 ( .IN1(n13148), .IN2(n13254), .IN3(n13255), .Q(g29291) );
  AND2X1 U13820 ( .IN1(n3765), .IN2(n13256), .Q(n13255) );
  OR2X1 U13821 ( .IN1(n10987), .IN2(n5737), .Q(n13256) );
  AND3X1 U13822 ( .IN1(n9449), .IN2(g5503), .IN3(n12338), .Q(n13254) );
  OR3X1 U13823 ( .IN1(n13257), .IN2(n13258), .IN3(n13259), .Q(g29290) );
  AND2X1 U13824 ( .IN1(n9142), .IN2(g5485), .Q(n13259) );
  AND2X1 U13825 ( .IN1(n5660), .IN2(n13260), .Q(n13258) );
  AND2X1 U13826 ( .IN1(n13261), .IN2(g5489), .Q(n13257) );
  OR3X1 U13827 ( .IN1(n13262), .IN2(n13263), .IN3(n13264), .Q(g29289) );
  AND2X1 U13828 ( .IN1(n13261), .IN2(g5485), .Q(n13264) );
  AND3X1 U13829 ( .IN1(n5425), .IN2(n13260), .IN3(n5805), .Q(n13263) );
  AND2X1 U13830 ( .IN1(n13265), .IN2(g5481), .Q(n13262) );
  OR2X1 U13831 ( .IN1(n9131), .IN2(n13266), .Q(n13265) );
  AND2X1 U13832 ( .IN1(n13267), .IN2(g5475), .Q(n13266) );
  OR2X1 U13833 ( .IN1(n13268), .IN2(n13269), .Q(g29288) );
  AND2X1 U13834 ( .IN1(n13270), .IN2(g5475), .Q(n13269) );
  AND2X1 U13835 ( .IN1(n13261), .IN2(g5481), .Q(n13268) );
  INVX0 U13836 ( .INP(n13270), .ZN(n13261) );
  OR2X1 U13837 ( .IN1(n9131), .IN2(n13267), .Q(n13270) );
  OR3X1 U13838 ( .IN1(n13271), .IN2(n13272), .IN3(n13273), .Q(g29287) );
  INVX0 U13839 ( .INP(n13274), .ZN(n13273) );
  OR2X1 U13840 ( .IN1(n12070), .IN2(n13267), .Q(n13274) );
  OR2X1 U13841 ( .IN1(n8780), .IN2(n9123), .Q(n12070) );
  AND3X1 U13842 ( .IN1(n13260), .IN2(g5467), .IN3(n5744), .Q(n13272) );
  AND2X1 U13843 ( .IN1(n9042), .IN2(n13267), .Q(n13260) );
  AND2X1 U13844 ( .IN1(n13275), .IN2(g5462), .Q(n13271) );
  OR2X1 U13845 ( .IN1(n9132), .IN2(n13276), .Q(n13275) );
  AND2X1 U13846 ( .IN1(n8725), .IN2(n13267), .Q(n13276) );
  OR3X1 U13847 ( .IN1(n13277), .IN2(n13278), .IN3(n13279), .Q(g29286) );
  AND2X1 U13848 ( .IN1(n11060), .IN2(g5462), .Q(n13279) );
  AND3X1 U13849 ( .IN1(n13280), .IN2(n13281), .IN3(n9079), .Q(n13278) );
  OR2X1 U13850 ( .IN1(n13282), .IN2(n13267), .Q(n13281) );
  AND2X1 U13851 ( .IN1(n11052), .IN2(n13283), .Q(n13267) );
  INVX0 U13852 ( .INP(n13284), .ZN(n13282) );
  OR2X1 U13853 ( .IN1(n11056), .IN2(n13285), .Q(n13284) );
  AND2X1 U13854 ( .IN1(g5462), .IN2(n13286), .Q(n13285) );
  OR2X1 U13855 ( .IN1(n13287), .IN2(n13286), .Q(n13280) );
  INVX0 U13856 ( .INP(n13288), .ZN(n13287) );
  OR2X1 U13857 ( .IN1(n13283), .IN2(n5744), .Q(n13288) );
  AND3X1 U13858 ( .IN1(g17604), .IN2(g5689), .IN3(n10237), .Q(n13283) );
  AND2X1 U13859 ( .IN1(n9141), .IN2(g5467), .Q(n13277) );
  OR3X1 U13860 ( .IN1(n13148), .IN2(n13289), .IN3(n13290), .Q(g29285) );
  AND2X1 U13861 ( .IN1(n3765), .IN2(n13291), .Q(n13290) );
  OR2X1 U13862 ( .IN1(g32975), .IN2(n5734), .Q(n13291) );
  AND3X1 U13863 ( .IN1(n9449), .IN2(g5156), .IN3(n9490), .Q(n13289) );
  OR3X1 U13864 ( .IN1(n13292), .IN2(n13293), .IN3(n13294), .Q(g29284) );
  AND2X1 U13865 ( .IN1(n9141), .IN2(g5138), .Q(n13294) );
  AND2X1 U13866 ( .IN1(n13295), .IN2(n5658), .Q(n13293) );
  AND2X1 U13867 ( .IN1(n13296), .IN2(g5142), .Q(n13292) );
  OR3X1 U13868 ( .IN1(n13297), .IN2(n13298), .IN3(n13299), .Q(g29283) );
  AND2X1 U13869 ( .IN1(n13296), .IN2(g5138), .Q(n13299) );
  AND3X1 U13870 ( .IN1(n13295), .IN2(n8848), .IN3(n5807), .Q(n13298) );
  AND2X1 U13871 ( .IN1(n13300), .IN2(g5134), .Q(n13297) );
  OR2X1 U13872 ( .IN1(n9132), .IN2(n13301), .Q(n13300) );
  AND2X1 U13873 ( .IN1(test_so96), .IN2(n13302), .Q(n13301) );
  OR2X1 U13874 ( .IN1(n13303), .IN2(n13304), .Q(g29282) );
  AND2X1 U13875 ( .IN1(test_so96), .IN2(n13305), .Q(n13304) );
  AND2X1 U13876 ( .IN1(n13296), .IN2(g5134), .Q(n13303) );
  INVX0 U13877 ( .INP(n13305), .ZN(n13296) );
  OR2X1 U13878 ( .IN1(n9132), .IN2(n13302), .Q(n13305) );
  OR3X1 U13879 ( .IN1(n13306), .IN2(n13307), .IN3(n13308), .Q(g29281) );
  INVX0 U13880 ( .INP(n13309), .ZN(n13308) );
  OR2X1 U13881 ( .IN1(n12067), .IN2(n13302), .Q(n13309) );
  OR2X1 U13882 ( .IN1(n8787), .IN2(n9123), .Q(n12067) );
  AND3X1 U13883 ( .IN1(n13295), .IN2(g5120), .IN3(n5743), .Q(n13307) );
  AND2X1 U13884 ( .IN1(n9042), .IN2(n13302), .Q(n13295) );
  AND2X1 U13885 ( .IN1(n13310), .IN2(g5115), .Q(n13306) );
  OR2X1 U13886 ( .IN1(n9132), .IN2(n13311), .Q(n13310) );
  AND2X1 U13887 ( .IN1(n8726), .IN2(n13302), .Q(n13311) );
  OR3X1 U13888 ( .IN1(n13312), .IN2(n13313), .IN3(n13314), .Q(g29280) );
  AND2X1 U13889 ( .IN1(n11072), .IN2(g5115), .Q(n13314) );
  AND3X1 U13890 ( .IN1(n13315), .IN2(n13316), .IN3(n9078), .Q(n13313) );
  OR2X1 U13891 ( .IN1(n13317), .IN2(n13302), .Q(n13316) );
  AND2X1 U13892 ( .IN1(g33959), .IN2(n13318), .Q(n13302) );
  INVX0 U13893 ( .INP(n13319), .ZN(n13317) );
  OR2X1 U13894 ( .IN1(n13320), .IN2(n8804), .Q(n13319) );
  AND2X1 U13895 ( .IN1(g5115), .IN2(n13321), .Q(n13320) );
  OR2X1 U13896 ( .IN1(n13322), .IN2(n13321), .Q(n13315) );
  INVX0 U13897 ( .INP(n13323), .ZN(n13322) );
  OR2X1 U13898 ( .IN1(n13318), .IN2(n5743), .Q(n13323) );
  AND3X1 U13899 ( .IN1(g17577), .IN2(g31860), .IN3(test_so10), .Q(n13318) );
  AND2X1 U13900 ( .IN1(n9141), .IN2(g5120), .Q(n13312) );
  OR2X1 U13901 ( .IN1(n13324), .IN2(g29279), .Q(g29278) );
  AND2X1 U13902 ( .IN1(n9141), .IN2(g4572), .Q(n13324) );
  OR2X1 U13903 ( .IN1(n13325), .IN2(g29277), .Q(g29276) );
  AND2X1 U13904 ( .IN1(test_so100), .IN2(n9138), .Q(n13325) );
  OR2X1 U13905 ( .IN1(n13326), .IN2(n13327), .Q(g29275) );
  AND2X1 U13906 ( .IN1(test_so11), .IN2(n9138), .Q(n13327) );
  AND3X1 U13907 ( .IN1(n3729), .IN2(g4169), .IN3(n13328), .Q(n13326) );
  OR2X1 U13908 ( .IN1(n13329), .IN2(n13330), .Q(n13328) );
  AND2X1 U13909 ( .IN1(n9043), .IN2(g4087), .Q(n13330) );
  AND2X1 U13910 ( .IN1(test_so11), .IN2(n12528), .Q(n13329) );
  INVX0 U13911 ( .INP(n12013), .ZN(n3729) );
  AND3X1 U13912 ( .IN1(g4087), .IN2(n12528), .IN3(test_so11), .Q(n12013) );
  OR3X1 U13913 ( .IN1(n13148), .IN2(n13331), .IN3(n13332), .Q(g29274) );
  AND2X1 U13914 ( .IN1(n3765), .IN2(n13333), .Q(n13332) );
  OR2X1 U13915 ( .IN1(n9376), .IN2(n5735), .Q(n13333) );
  AND3X1 U13916 ( .IN1(n9449), .IN2(g3849), .IN3(n9375), .Q(n13331) );
  OR3X1 U13917 ( .IN1(n13334), .IN2(n13335), .IN3(n13336), .Q(g29273) );
  AND2X1 U13918 ( .IN1(n9142), .IN2(g3831), .Q(n13336) );
  AND2X1 U13919 ( .IN1(n13337), .IN2(n5662), .Q(n13335) );
  AND2X1 U13920 ( .IN1(n13338), .IN2(g3835), .Q(n13334) );
  OR3X1 U13921 ( .IN1(n13339), .IN2(n13340), .IN3(n13341), .Q(g29272) );
  AND2X1 U13922 ( .IN1(n13338), .IN2(g3831), .Q(n13341) );
  AND3X1 U13923 ( .IN1(n5428), .IN2(n13337), .IN3(n5808), .Q(n13340) );
  AND2X1 U13924 ( .IN1(n13342), .IN2(g3827), .Q(n13339) );
  OR2X1 U13925 ( .IN1(n9132), .IN2(n13343), .Q(n13342) );
  AND2X1 U13926 ( .IN1(n13344), .IN2(g3821), .Q(n13343) );
  OR2X1 U13927 ( .IN1(n13345), .IN2(n13346), .Q(g29271) );
  AND2X1 U13928 ( .IN1(n13347), .IN2(g3821), .Q(n13346) );
  AND2X1 U13929 ( .IN1(n13338), .IN2(g3827), .Q(n13345) );
  INVX0 U13930 ( .INP(n13347), .ZN(n13338) );
  OR2X1 U13931 ( .IN1(n9132), .IN2(n13344), .Q(n13347) );
  OR3X1 U13932 ( .IN1(n13348), .IN2(n13349), .IN3(n13350), .Q(g29270) );
  INVX0 U13933 ( .INP(n13351), .ZN(n13350) );
  OR2X1 U13934 ( .IN1(n9888), .IN2(n13344), .Q(n13351) );
  OR2X1 U13935 ( .IN1(n8759), .IN2(n9123), .Q(n9888) );
  AND3X1 U13936 ( .IN1(n13337), .IN2(g3813), .IN3(n5745), .Q(n13349) );
  AND2X1 U13937 ( .IN1(n9043), .IN2(n13344), .Q(n13337) );
  AND2X1 U13938 ( .IN1(n13352), .IN2(g3808), .Q(n13348) );
  OR2X1 U13939 ( .IN1(n9132), .IN2(n13353), .Q(n13352) );
  AND2X1 U13940 ( .IN1(n8724), .IN2(n13344), .Q(n13353) );
  OR3X1 U13941 ( .IN1(n13354), .IN2(n13355), .IN3(n13356), .Q(g29269) );
  AND2X1 U13942 ( .IN1(n11099), .IN2(g3808), .Q(n13356) );
  AND3X1 U13943 ( .IN1(n13357), .IN2(n13358), .IN3(n9078), .Q(n13355) );
  OR2X1 U13944 ( .IN1(n13359), .IN2(n13344), .Q(n13358) );
  AND2X1 U13945 ( .IN1(n11091), .IN2(n13360), .Q(n13344) );
  INVX0 U13946 ( .INP(n13361), .ZN(n13359) );
  OR2X1 U13947 ( .IN1(n11095), .IN2(n13362), .Q(n13361) );
  AND2X1 U13948 ( .IN1(g3808), .IN2(n13363), .Q(n13362) );
  OR2X1 U13949 ( .IN1(n13364), .IN2(n13363), .Q(n13357) );
  INVX0 U13950 ( .INP(n13365), .ZN(n13364) );
  OR2X1 U13951 ( .IN1(n13360), .IN2(n5745), .Q(n13365) );
  AND3X1 U13952 ( .IN1(g16693), .IN2(g4040), .IN3(n10231), .Q(n13360) );
  AND2X1 U13953 ( .IN1(n9140), .IN2(g3813), .Q(n13354) );
  OR3X1 U13954 ( .IN1(n13148), .IN2(n13366), .IN3(n13367), .Q(g29268) );
  AND2X1 U13955 ( .IN1(n3765), .IN2(n13368), .Q(n13367) );
  OR2X1 U13956 ( .IN1(n10982), .IN2(n5740), .Q(n13368) );
  AND3X1 U13957 ( .IN1(n9449), .IN2(g3498), .IN3(n12616), .Q(n13366) );
  OR3X1 U13958 ( .IN1(n13369), .IN2(n13370), .IN3(n13371), .Q(g29267) );
  AND2X1 U13959 ( .IN1(n9141), .IN2(g3480), .Q(n13371) );
  AND2X1 U13960 ( .IN1(n5668), .IN2(n9502), .Q(n13370) );
  AND2X1 U13961 ( .IN1(n13372), .IN2(g3484), .Q(n13369) );
  OR3X1 U13962 ( .IN1(n13373), .IN2(n13374), .IN3(n13375), .Q(g29266) );
  AND2X1 U13963 ( .IN1(n13372), .IN2(g3480), .Q(n13375) );
  AND3X1 U13964 ( .IN1(n5424), .IN2(n9502), .IN3(n5786), .Q(n13374) );
  AND2X1 U13965 ( .IN1(n9043), .IN2(n9501), .Q(n9502) );
  AND2X1 U13966 ( .IN1(n13376), .IN2(g3476), .Q(n13373) );
  OR2X1 U13967 ( .IN1(n9132), .IN2(n13377), .Q(n13376) );
  AND2X1 U13968 ( .IN1(n9501), .IN2(g3470), .Q(n13377) );
  OR2X1 U13969 ( .IN1(n13378), .IN2(n13379), .Q(g29265) );
  AND2X1 U13970 ( .IN1(n13380), .IN2(g3470), .Q(n13379) );
  AND2X1 U13971 ( .IN1(n13372), .IN2(g3476), .Q(n13378) );
  INVX0 U13972 ( .INP(n13380), .ZN(n13372) );
  OR2X1 U13973 ( .IN1(n9132), .IN2(n9501), .Q(n13380) );
  OR3X1 U13974 ( .IN1(n13381), .IN2(n13382), .IN3(n13383), .Q(g29263) );
  AND2X1 U13975 ( .IN1(n11115), .IN2(test_so4), .Q(n13383) );
  AND3X1 U13976 ( .IN1(n13384), .IN2(n13385), .IN3(n9078), .Q(n13382) );
  INVX0 U13977 ( .INP(n13386), .ZN(n13385) );
  AND2X1 U13978 ( .IN1(n13387), .IN2(n13388), .Q(n13386) );
  OR2X1 U13979 ( .IN1(n8821), .IN2(n13389), .Q(n13387) );
  OR2X1 U13980 ( .IN1(n13390), .IN2(n9501), .Q(n13384) );
  AND2X1 U13981 ( .IN1(n13389), .IN2(n11107), .Q(n9501) );
  AND3X1 U13982 ( .IN1(g16656), .IN2(g3689), .IN3(n10244), .Q(n13389) );
  AND2X1 U13983 ( .IN1(n11107), .IN2(n13391), .Q(n13390) );
  OR2X1 U13984 ( .IN1(n13388), .IN2(n8821), .Q(n13391) );
  INVX0 U13985 ( .INP(n13392), .ZN(n13388) );
  AND2X1 U13986 ( .IN1(n9140), .IN2(g3462), .Q(n13381) );
  OR3X1 U13987 ( .IN1(n13148), .IN2(n13393), .IN3(n13394), .Q(g29262) );
  AND2X1 U13988 ( .IN1(n3765), .IN2(n13395), .Q(n13394) );
  OR2X1 U13989 ( .IN1(n10977), .IN2(n5738), .Q(n13395) );
  AND3X1 U13990 ( .IN1(n9449), .IN2(g3147), .IN3(n12701), .Q(n13393) );
  AND2X1 U13991 ( .IN1(n9449), .IN2(n3765), .Q(n13148) );
  AND2X1 U13992 ( .IN1(g4180), .IN2(n8361), .Q(n9449) );
  OR3X1 U13993 ( .IN1(n13396), .IN2(n13397), .IN3(n13398), .Q(g29261) );
  AND2X1 U13994 ( .IN1(n9141), .IN2(g3129), .Q(n13398) );
  AND2X1 U13995 ( .IN1(n5661), .IN2(n13399), .Q(n13397) );
  AND2X1 U13996 ( .IN1(n13400), .IN2(g3133), .Q(n13396) );
  OR3X1 U13997 ( .IN1(n13401), .IN2(n13402), .IN3(n13403), .Q(g29260) );
  AND2X1 U13998 ( .IN1(n13400), .IN2(g3129), .Q(n13403) );
  AND3X1 U13999 ( .IN1(n5423), .IN2(n13399), .IN3(n5781), .Q(n13402) );
  AND2X1 U14000 ( .IN1(n13404), .IN2(g3125), .Q(n13401) );
  OR2X1 U14001 ( .IN1(n9133), .IN2(n13405), .Q(n13404) );
  AND2X1 U14002 ( .IN1(n13406), .IN2(g3119), .Q(n13405) );
  OR2X1 U14003 ( .IN1(n13407), .IN2(n13408), .Q(g29259) );
  AND2X1 U14004 ( .IN1(n13409), .IN2(g3119), .Q(n13408) );
  AND2X1 U14005 ( .IN1(n13400), .IN2(g3125), .Q(n13407) );
  INVX0 U14006 ( .INP(n13409), .ZN(n13400) );
  OR2X1 U14007 ( .IN1(n9133), .IN2(n13406), .Q(n13409) );
  OR3X1 U14008 ( .IN1(n13410), .IN2(n13411), .IN3(n13412), .Q(g29258) );
  INVX0 U14009 ( .INP(n13413), .ZN(n13412) );
  OR2X1 U14010 ( .IN1(n12075), .IN2(n13406), .Q(n13413) );
  OR2X1 U14011 ( .IN1(n8738), .IN2(n9123), .Q(n12075) );
  AND3X1 U14012 ( .IN1(n13399), .IN2(g3111), .IN3(n5742), .Q(n13411) );
  AND2X1 U14013 ( .IN1(n9043), .IN2(n13406), .Q(n13399) );
  AND2X1 U14014 ( .IN1(n13414), .IN2(g3106), .Q(n13410) );
  OR2X1 U14015 ( .IN1(n9133), .IN2(n13415), .Q(n13414) );
  AND2X1 U14016 ( .IN1(n8727), .IN2(n13406), .Q(n13415) );
  OR3X1 U14017 ( .IN1(n13416), .IN2(n13417), .IN3(n13418), .Q(g29257) );
  AND2X1 U14018 ( .IN1(n11129), .IN2(g3106), .Q(n13418) );
  AND3X1 U14019 ( .IN1(n13419), .IN2(n13420), .IN3(n9077), .Q(n13417) );
  OR2X1 U14020 ( .IN1(n13421), .IN2(n13406), .Q(n13420) );
  AND2X1 U14021 ( .IN1(n11125), .IN2(n13422), .Q(n13406) );
  INVX0 U14022 ( .INP(n13423), .ZN(n13421) );
  OR2X1 U14023 ( .IN1(n11123), .IN2(n13424), .Q(n13423) );
  AND2X1 U14024 ( .IN1(g3106), .IN2(n13425), .Q(n13424) );
  OR2X1 U14025 ( .IN1(n13426), .IN2(n13425), .Q(n13419) );
  INVX0 U14026 ( .INP(n13427), .ZN(n13426) );
  OR2X1 U14027 ( .IN1(n13422), .IN2(n5742), .Q(n13427) );
  AND3X1 U14028 ( .IN1(g16624), .IN2(g3338), .IN3(n10236), .Q(n13422) );
  AND2X1 U14029 ( .IN1(n9140), .IN2(g3111), .Q(n13416) );
  OR4X1 U14030 ( .IN1(n2787), .IN2(n13428), .IN3(n13429), .IN4(n13430), .Q(
        g29256) );
  AND2X1 U14031 ( .IN1(n9141), .IN2(g2729), .Q(n13430) );
  AND3X1 U14032 ( .IN1(n13431), .IN2(g2735), .IN3(n9077), .Q(n13429) );
  AND2X1 U14033 ( .IN1(n5600), .IN2(n12824), .Q(n13428) );
  INVX0 U14034 ( .INP(n13431), .ZN(n12824) );
  OR2X1 U14035 ( .IN1(n13432), .IN2(n13433), .Q(g29255) );
  AND2X1 U14036 ( .IN1(n13434), .IN2(g2652), .Q(n13433) );
  OR2X1 U14037 ( .IN1(n13435), .IN2(n11747), .Q(n13434) );
  AND2X1 U14038 ( .IN1(n4379), .IN2(n9022), .Q(n13435) );
  AND2X1 U14039 ( .IN1(n13436), .IN2(g2638), .Q(n13432) );
  OR2X1 U14040 ( .IN1(n9133), .IN2(n13437), .Q(n13436) );
  AND2X1 U14041 ( .IN1(n11744), .IN2(n9388), .Q(n13437) );
  OR2X1 U14042 ( .IN1(n8808), .IN2(n8622), .Q(n9388) );
  OR4X1 U14043 ( .IN1(n13438), .IN2(n13439), .IN3(n13440), .IN4(n13441), .Q(
        g29254) );
  AND2X1 U14044 ( .IN1(n3517), .IN2(n13442), .Q(n13441) );
  OR4X1 U14045 ( .IN1(n13443), .IN2(n13444), .IN3(n13445), .IN4(n13446), .Q(
        n13442) );
  AND2X1 U14046 ( .IN1(n8772), .IN2(n13447), .Q(n13446) );
  OR2X1 U14047 ( .IN1(n13448), .IN2(n13449), .Q(n13447) );
  AND2X1 U14048 ( .IN1(g2619), .IN2(g2571), .Q(n13449) );
  AND2X1 U14049 ( .IN1(test_so61), .IN2(g2587), .Q(n13448) );
  AND3X1 U14050 ( .IN1(n5508), .IN2(n5372), .IN3(test_so66), .Q(n13445) );
  AND2X1 U14051 ( .IN1(n8808), .IN2(g2563), .Q(n13444) );
  INVX0 U14052 ( .INP(n11758), .ZN(n8808) );
  OR2X1 U14053 ( .IN1(n8772), .IN2(g2587), .Q(n11758) );
  AND2X1 U14054 ( .IN1(n10391), .IN2(g2583), .Q(n13443) );
  AND2X1 U14055 ( .IN1(g2610), .IN2(n5508), .Q(n10391) );
  AND2X1 U14056 ( .IN1(n9043), .IN2(n11744), .Q(n3517) );
  AND2X1 U14057 ( .IN1(n12829), .IN2(g2567), .Q(n13440) );
  AND2X1 U14058 ( .IN1(n9043), .IN2(n12832), .Q(n12829) );
  AND3X1 U14059 ( .IN1(g2619), .IN2(g2587), .IN3(n11744), .Q(n12832) );
  INVX0 U14060 ( .INP(n13450), .ZN(n11744) );
  AND2X1 U14061 ( .IN1(n9140), .IN2(g2619), .Q(n13439) );
  AND2X1 U14062 ( .IN1(n11747), .IN2(g2638), .Q(n13438) );
  AND2X1 U14063 ( .IN1(n9044), .IN2(n13450), .Q(n11747) );
  OR3X1 U14064 ( .IN1(n13451), .IN2(n13452), .IN3(n12798), .Q(n13450) );
  AND2X1 U14065 ( .IN1(n10197), .IN2(g2819), .Q(n13452) );
  OR2X1 U14066 ( .IN1(n13453), .IN2(n13454), .Q(g29253) );
  AND2X1 U14067 ( .IN1(n13455), .IN2(g2518), .Q(n13454) );
  OR2X1 U14068 ( .IN1(n13456), .IN2(n11766), .Q(n13455) );
  AND2X1 U14069 ( .IN1(n4391), .IN2(n9021), .Q(n13456) );
  AND2X1 U14070 ( .IN1(n13457), .IN2(g2504), .Q(n13453) );
  OR2X1 U14071 ( .IN1(n9133), .IN2(n13458), .Q(n13457) );
  AND2X1 U14072 ( .IN1(n11763), .IN2(n9387), .Q(n13458) );
  OR2X1 U14073 ( .IN1(n8815), .IN2(n8624), .Q(n9387) );
  OR4X1 U14074 ( .IN1(n13459), .IN2(n13460), .IN3(n13461), .IN4(n13462), .Q(
        g29252) );
  OR2X1 U14075 ( .IN1(n13463), .IN2(n13464), .Q(n13462) );
  AND2X1 U14076 ( .IN1(n3536), .IN2(n13465), .Q(n13464) );
  OR3X1 U14077 ( .IN1(n13466), .IN2(n13467), .IN3(n13468), .Q(n13465) );
  AND2X1 U14078 ( .IN1(n8815), .IN2(g2429), .Q(n13468) );
  INVX0 U14079 ( .INP(n11777), .ZN(n8815) );
  OR2X1 U14080 ( .IN1(n8773), .IN2(g2453), .Q(n11777) );
  AND2X1 U14081 ( .IN1(n8773), .IN2(n13469), .Q(n13467) );
  OR2X1 U14082 ( .IN1(n13470), .IN2(n13471), .Q(n13469) );
  AND2X1 U14083 ( .IN1(g2485), .IN2(g2437), .Q(n13471) );
  AND2X1 U14084 ( .IN1(g2453), .IN2(n9274), .Q(n13470) );
  AND3X1 U14085 ( .IN1(n5373), .IN2(g2441), .IN3(n5509), .Q(n13466) );
  AND2X1 U14086 ( .IN1(n9044), .IN2(n11763), .Q(n3536) );
  AND2X1 U14087 ( .IN1(n12857), .IN2(g2433), .Q(n13463) );
  AND2X1 U14088 ( .IN1(n9044), .IN2(n12860), .Q(n12857) );
  AND3X1 U14089 ( .IN1(g2485), .IN2(g2453), .IN3(n11763), .Q(n12860) );
  AND2X1 U14090 ( .IN1(n11766), .IN2(g2504), .Q(n13461) );
  AND2X1 U14091 ( .IN1(n9044), .IN2(n13472), .Q(n11766) );
  AND3X1 U14092 ( .IN1(n12880), .IN2(g2449), .IN3(n9077), .Q(n13460) );
  AND3X1 U14093 ( .IN1(g2476), .IN2(n11763), .IN3(n5509), .Q(n12880) );
  INVX0 U14094 ( .INP(n13472), .ZN(n11763) );
  OR3X1 U14095 ( .IN1(n13451), .IN2(n13473), .IN3(n12799), .Q(n13472) );
  AND2X1 U14096 ( .IN1(n10197), .IN2(g2815), .Q(n13473) );
  AND2X1 U14097 ( .IN1(n9140), .IN2(g2485), .Q(n13459) );
  OR2X1 U14098 ( .IN1(n13474), .IN2(n13475), .Q(g29251) );
  AND2X1 U14099 ( .IN1(n13476), .IN2(g2370), .Q(n13475) );
  OR2X1 U14100 ( .IN1(n9133), .IN2(n13477), .Q(n13476) );
  AND2X1 U14101 ( .IN1(n11782), .IN2(n9386), .Q(n13477) );
  OR2X1 U14102 ( .IN1(n8810), .IN2(n8629), .Q(n9386) );
  AND2X1 U14103 ( .IN1(n13478), .IN2(g2384), .Q(n13474) );
  OR2X1 U14104 ( .IN1(n13479), .IN2(n11785), .Q(n13478) );
  AND2X1 U14105 ( .IN1(n4402), .IN2(n9021), .Q(n13479) );
  OR4X1 U14106 ( .IN1(n13480), .IN2(n13481), .IN3(n13482), .IN4(n13483), .Q(
        g29250) );
  OR2X1 U14107 ( .IN1(n13484), .IN2(n13485), .Q(n13483) );
  AND2X1 U14108 ( .IN1(n3555), .IN2(n13486), .Q(n13485) );
  OR3X1 U14109 ( .IN1(n13487), .IN2(n13488), .IN3(n13489), .Q(n13486) );
  AND2X1 U14110 ( .IN1(n8810), .IN2(g2295), .Q(n13489) );
  INVX0 U14111 ( .INP(n11796), .ZN(n8810) );
  OR2X1 U14112 ( .IN1(g2319), .IN2(n8830), .Q(n11796) );
  AND2X1 U14113 ( .IN1(n13490), .IN2(n8830), .Q(n13488) );
  OR2X1 U14114 ( .IN1(n13491), .IN2(n13492), .Q(n13490) );
  AND2X1 U14115 ( .IN1(g2351), .IN2(g2303), .Q(n13492) );
  AND2X1 U14116 ( .IN1(g2319), .IN2(n9314), .Q(n13491) );
  AND3X1 U14117 ( .IN1(n5375), .IN2(g2307), .IN3(n5511), .Q(n13487) );
  AND2X1 U14118 ( .IN1(n9044), .IN2(n11782), .Q(n3555) );
  AND2X1 U14119 ( .IN1(n12887), .IN2(g2299), .Q(n13484) );
  AND2X1 U14120 ( .IN1(n9044), .IN2(n12890), .Q(n12887) );
  AND3X1 U14121 ( .IN1(g2351), .IN2(g2319), .IN3(n11782), .Q(n12890) );
  AND2X1 U14122 ( .IN1(n11785), .IN2(g2370), .Q(n13482) );
  AND2X1 U14123 ( .IN1(n9044), .IN2(n13493), .Q(n11785) );
  AND3X1 U14124 ( .IN1(n12910), .IN2(g2315), .IN3(n9077), .Q(n13481) );
  AND3X1 U14125 ( .IN1(test_so21), .IN2(n11782), .IN3(n5511), .Q(n12910) );
  INVX0 U14126 ( .INP(n13493), .ZN(n11782) );
  OR3X1 U14127 ( .IN1(n1256), .IN2(n13451), .IN3(n13494), .Q(n13493) );
  AND2X1 U14128 ( .IN1(n10197), .IN2(g2807), .Q(n13494) );
  AND2X1 U14129 ( .IN1(n9140), .IN2(g2351), .Q(n13480) );
  OR2X1 U14130 ( .IN1(n13495), .IN2(n13496), .Q(g29249) );
  AND2X1 U14131 ( .IN1(n13497), .IN2(g2236), .Q(n13496) );
  OR2X1 U14132 ( .IN1(n9133), .IN2(n13498), .Q(n13497) );
  AND2X1 U14133 ( .IN1(n11801), .IN2(n9385), .Q(n13498) );
  OR2X1 U14134 ( .IN1(n8816), .IN2(n8633), .Q(n9385) );
  AND2X1 U14135 ( .IN1(n13499), .IN2(g2250), .Q(n13495) );
  OR2X1 U14136 ( .IN1(n13500), .IN2(n11804), .Q(n13499) );
  AND2X1 U14137 ( .IN1(n4414), .IN2(n9021), .Q(n13500) );
  OR4X1 U14138 ( .IN1(n13501), .IN2(n13502), .IN3(n13503), .IN4(n13504), .Q(
        g29248) );
  OR2X1 U14139 ( .IN1(n13505), .IN2(n13506), .Q(n13504) );
  AND2X1 U14140 ( .IN1(n3574), .IN2(n13507), .Q(n13506) );
  OR3X1 U14141 ( .IN1(n13508), .IN2(n13509), .IN3(n13510), .Q(n13507) );
  AND2X1 U14142 ( .IN1(n8816), .IN2(g2161), .Q(n13510) );
  INVX0 U14143 ( .INP(n11815), .ZN(n8816) );
  OR2X1 U14144 ( .IN1(n8721), .IN2(g2185), .Q(n11815) );
  AND2X1 U14145 ( .IN1(n8721), .IN2(n13511), .Q(n13509) );
  OR2X1 U14146 ( .IN1(n13512), .IN2(n13513), .Q(n13511) );
  AND2X1 U14147 ( .IN1(g2217), .IN2(g2169), .Q(n13513) );
  AND2X1 U14148 ( .IN1(g2185), .IN2(n9352), .Q(n13512) );
  AND3X1 U14149 ( .IN1(n5376), .IN2(g2173), .IN3(n5512), .Q(n13508) );
  AND2X1 U14150 ( .IN1(n9044), .IN2(n11801), .Q(n3574) );
  AND2X1 U14151 ( .IN1(n12917), .IN2(g2165), .Q(n13505) );
  AND2X1 U14152 ( .IN1(n9044), .IN2(n12920), .Q(n12917) );
  AND3X1 U14153 ( .IN1(g2217), .IN2(g2185), .IN3(n11801), .Q(n12920) );
  AND2X1 U14154 ( .IN1(n11804), .IN2(g2236), .Q(n13503) );
  AND2X1 U14155 ( .IN1(n9044), .IN2(n13514), .Q(n11804) );
  AND3X1 U14156 ( .IN1(n12940), .IN2(g2181), .IN3(n9077), .Q(n13502) );
  AND3X1 U14157 ( .IN1(g2208), .IN2(n11801), .IN3(n5512), .Q(n12940) );
  INVX0 U14158 ( .INP(n13514), .ZN(n11801) );
  OR2X1 U14159 ( .IN1(n13515), .IN2(n13516), .Q(n13514) );
  AND2X1 U14160 ( .IN1(n10197), .IN2(g2803), .Q(n13515) );
  AND2X1 U14161 ( .IN1(n9141), .IN2(g2217), .Q(n13501) );
  OR2X1 U14162 ( .IN1(n13517), .IN2(n13518), .Q(g29247) );
  AND2X1 U14163 ( .IN1(test_so78), .IN2(n13519), .Q(n13518) );
  OR2X1 U14164 ( .IN1(n13520), .IN2(n11823), .Q(n13519) );
  AND2X1 U14165 ( .IN1(n4425), .IN2(n9020), .Q(n13520) );
  AND2X1 U14166 ( .IN1(n13521), .IN2(g2079), .Q(n13517) );
  OR2X1 U14167 ( .IN1(n9133), .IN2(n13522), .Q(n13521) );
  AND2X1 U14168 ( .IN1(n11820), .IN2(n9384), .Q(n13522) );
  OR2X1 U14169 ( .IN1(n8818), .IN2(n8833), .Q(n9384) );
  OR4X1 U14170 ( .IN1(n13523), .IN2(n13524), .IN3(n13525), .IN4(n13526), .Q(
        g29246) );
  AND2X1 U14171 ( .IN1(n3593), .IN2(n13527), .Q(n13526) );
  OR4X1 U14172 ( .IN1(n13528), .IN2(n13529), .IN3(n13530), .IN4(n13531), .Q(
        n13527) );
  AND2X1 U14173 ( .IN1(n8778), .IN2(n13532), .Q(n13531) );
  OR2X1 U14174 ( .IN1(n13533), .IN2(n13534), .Q(n13532) );
  AND2X1 U14175 ( .IN1(g2060), .IN2(g2012), .Q(n13534) );
  AND2X1 U14176 ( .IN1(g2028), .IN2(n9312), .Q(n13533) );
  AND3X1 U14177 ( .IN1(n5371), .IN2(g2016), .IN3(n5507), .Q(n13530) );
  AND2X1 U14178 ( .IN1(n8818), .IN2(g2004), .Q(n13529) );
  INVX0 U14179 ( .INP(n11834), .ZN(n8818) );
  OR2X1 U14180 ( .IN1(n8778), .IN2(g2028), .Q(n11834) );
  AND2X1 U14181 ( .IN1(n10394), .IN2(g2024), .Q(n13528) );
  AND2X1 U14182 ( .IN1(g2051), .IN2(n5507), .Q(n10394) );
  AND2X1 U14183 ( .IN1(n9045), .IN2(n11820), .Q(n3593) );
  AND2X1 U14184 ( .IN1(n12947), .IN2(g2008), .Q(n13525) );
  AND2X1 U14185 ( .IN1(n9045), .IN2(n12950), .Q(n12947) );
  AND3X1 U14186 ( .IN1(g2060), .IN2(g2028), .IN3(n11820), .Q(n12950) );
  INVX0 U14187 ( .INP(n13535), .ZN(n11820) );
  AND2X1 U14188 ( .IN1(n9141), .IN2(g2060), .Q(n13524) );
  AND2X1 U14189 ( .IN1(n11823), .IN2(g2079), .Q(n13523) );
  AND2X1 U14190 ( .IN1(n9045), .IN2(n13535), .Q(n11823) );
  OR3X1 U14191 ( .IN1(n13451), .IN2(n13536), .IN3(n12798), .Q(n13535) );
  AND2X1 U14192 ( .IN1(n10197), .IN2(g2787), .Q(n13536) );
  OR2X1 U14193 ( .IN1(n13537), .IN2(n13538), .Q(g29245) );
  AND2X1 U14194 ( .IN1(test_so53), .IN2(n13539), .Q(n13538) );
  OR2X1 U14195 ( .IN1(n9133), .IN2(n13540), .Q(n13539) );
  AND2X1 U14196 ( .IN1(n11839), .IN2(n9383), .Q(n13540) );
  OR2X1 U14197 ( .IN1(n8807), .IN2(n8625), .Q(n9383) );
  AND2X1 U14198 ( .IN1(n13541), .IN2(g1959), .Q(n13537) );
  OR2X1 U14199 ( .IN1(n13542), .IN2(n11842), .Q(n13541) );
  AND2X1 U14200 ( .IN1(n4436), .IN2(n9020), .Q(n13542) );
  OR4X1 U14201 ( .IN1(n13543), .IN2(n13544), .IN3(n13545), .IN4(n13546), .Q(
        g29244) );
  OR2X1 U14202 ( .IN1(n13547), .IN2(n13548), .Q(n13546) );
  AND2X1 U14203 ( .IN1(n3611), .IN2(n13549), .Q(n13548) );
  OR3X1 U14204 ( .IN1(n13550), .IN2(n13551), .IN3(n13552), .Q(n13549) );
  AND2X1 U14205 ( .IN1(n8807), .IN2(g1870), .Q(n13552) );
  INVX0 U14206 ( .INP(n11854), .ZN(n8807) );
  OR2X1 U14207 ( .IN1(n8779), .IN2(g1894), .Q(n11854) );
  AND2X1 U14208 ( .IN1(n8779), .IN2(n13553), .Q(n13551) );
  OR2X1 U14209 ( .IN1(n13554), .IN2(n13555), .Q(n13553) );
  AND2X1 U14210 ( .IN1(g1926), .IN2(g1878), .Q(n13555) );
  AND2X1 U14211 ( .IN1(g1894), .IN2(n9280), .Q(n13554) );
  AND3X1 U14212 ( .IN1(n5374), .IN2(g1882), .IN3(n5510), .Q(n13550) );
  AND2X1 U14213 ( .IN1(n9045), .IN2(n11839), .Q(n3611) );
  AND2X1 U14214 ( .IN1(n12974), .IN2(g1874), .Q(n13547) );
  AND2X1 U14215 ( .IN1(n9046), .IN2(n12977), .Q(n12974) );
  AND3X1 U14216 ( .IN1(g1926), .IN2(g1894), .IN3(n11839), .Q(n12977) );
  AND2X1 U14217 ( .IN1(n11842), .IN2(test_so53), .Q(n13545) );
  AND2X1 U14218 ( .IN1(n9046), .IN2(n13556), .Q(n11842) );
  AND3X1 U14219 ( .IN1(n12997), .IN2(g1890), .IN3(n9076), .Q(n13544) );
  AND3X1 U14220 ( .IN1(g1917), .IN2(n11839), .IN3(n5510), .Q(n12997) );
  INVX0 U14221 ( .INP(n13556), .ZN(n11839) );
  OR3X1 U14222 ( .IN1(n13451), .IN2(n13557), .IN3(n12799), .Q(n13556) );
  INVX0 U14223 ( .INP(n13558), .ZN(n12799) );
  AND2X1 U14224 ( .IN1(n10197), .IN2(g2783), .Q(n13557) );
  AND2X1 U14225 ( .IN1(n9141), .IN2(g1926), .Q(n13543) );
  OR2X1 U14226 ( .IN1(n13559), .IN2(n13560), .Q(g29243) );
  AND2X1 U14227 ( .IN1(n13561), .IN2(g1811), .Q(n13560) );
  OR2X1 U14228 ( .IN1(n9133), .IN2(n13562), .Q(n13561) );
  AND2X1 U14229 ( .IN1(n11859), .IN2(n9382), .Q(n13562) );
  OR2X1 U14230 ( .IN1(n8813), .IN2(n8631), .Q(n9382) );
  AND2X1 U14231 ( .IN1(n13563), .IN2(g1825), .Q(n13559) );
  OR2X1 U14232 ( .IN1(n13564), .IN2(n11862), .Q(n13563) );
  AND2X1 U14233 ( .IN1(n4447), .IN2(n9020), .Q(n13564) );
  OR4X1 U14234 ( .IN1(n13565), .IN2(n13566), .IN3(n13567), .IN4(n13568), .Q(
        g29242) );
  OR2X1 U14235 ( .IN1(n13569), .IN2(n13570), .Q(n13568) );
  AND2X1 U14236 ( .IN1(n3628), .IN2(n13571), .Q(n13570) );
  OR3X1 U14237 ( .IN1(n13572), .IN2(n13573), .IN3(n13574), .Q(n13571) );
  AND2X1 U14238 ( .IN1(n8813), .IN2(g1736), .Q(n13574) );
  INVX0 U14239 ( .INP(n11873), .ZN(n8813) );
  OR2X1 U14240 ( .IN1(n5596), .IN2(g1760), .Q(n11873) );
  AND2X1 U14241 ( .IN1(n5596), .IN2(n13575), .Q(n13573) );
  OR2X1 U14242 ( .IN1(n13576), .IN2(n13577), .Q(n13575) );
  AND2X1 U14243 ( .IN1(g1760), .IN2(g1752), .Q(n13577) );
  AND2X1 U14244 ( .IN1(g1792), .IN2(g1744), .Q(n13576) );
  AND3X1 U14245 ( .IN1(n5602), .IN2(g1748), .IN3(n5359), .Q(n13572) );
  AND2X1 U14246 ( .IN1(n9046), .IN2(n11859), .Q(n3628) );
  AND2X1 U14247 ( .IN1(n13004), .IN2(g1740), .Q(n13569) );
  AND2X1 U14248 ( .IN1(n9045), .IN2(n13007), .Q(n13004) );
  AND3X1 U14249 ( .IN1(g1760), .IN2(g1792), .IN3(n11859), .Q(n13007) );
  AND2X1 U14250 ( .IN1(n11862), .IN2(g1811), .Q(n13567) );
  AND2X1 U14251 ( .IN1(n9046), .IN2(n13578), .Q(n11862) );
  AND3X1 U14252 ( .IN1(n13027), .IN2(g1756), .IN3(n9076), .Q(n13566) );
  AND3X1 U14253 ( .IN1(g1783), .IN2(n11859), .IN3(n5359), .Q(n13027) );
  INVX0 U14254 ( .INP(n13578), .ZN(n11859) );
  OR3X1 U14255 ( .IN1(n1256), .IN2(n13451), .IN3(n13579), .Q(n13578) );
  AND2X1 U14256 ( .IN1(n10197), .IN2(g2775), .Q(n13579) );
  OR2X1 U14257 ( .IN1(n5299), .IN2(g2719), .Q(n1256) );
  AND2X1 U14258 ( .IN1(n9141), .IN2(g1792), .Q(n13565) );
  OR2X1 U14259 ( .IN1(n13580), .IN2(n13581), .Q(g29241) );
  AND2X1 U14260 ( .IN1(n13582), .IN2(g1677), .Q(n13581) );
  OR2X1 U14261 ( .IN1(n9134), .IN2(n13583), .Q(n13582) );
  AND2X1 U14262 ( .IN1(n11878), .IN2(n9381), .Q(n13583) );
  OR2X1 U14263 ( .IN1(n8817), .IN2(n8627), .Q(n9381) );
  AND2X1 U14264 ( .IN1(n13584), .IN2(g1691), .Q(n13580) );
  OR2X1 U14265 ( .IN1(n13585), .IN2(n11881), .Q(n13584) );
  AND2X1 U14266 ( .IN1(n4458), .IN2(n9020), .Q(n13585) );
  OR4X1 U14267 ( .IN1(n13586), .IN2(n13587), .IN3(n13588), .IN4(n13589), .Q(
        g29240) );
  AND2X1 U14268 ( .IN1(n11881), .IN2(g1677), .Q(n13589) );
  AND2X1 U14269 ( .IN1(n9047), .IN2(n13590), .Q(n11881) );
  AND2X1 U14270 ( .IN1(n3646), .IN2(n13591), .Q(n13588) );
  OR4X1 U14271 ( .IN1(n13592), .IN2(n13593), .IN3(n13594), .IN4(n13595), .Q(
        n13591) );
  AND2X1 U14272 ( .IN1(n13596), .IN2(n8831), .Q(n13595) );
  OR2X1 U14273 ( .IN1(n13597), .IN2(n13598), .Q(n13596) );
  AND2X1 U14274 ( .IN1(g1657), .IN2(g1608), .Q(n13598) );
  AND2X1 U14275 ( .IN1(g1624), .IN2(n9303), .Q(n13597) );
  AND3X1 U14276 ( .IN1(n5370), .IN2(g1612), .IN3(n5525), .Q(n13594) );
  AND2X1 U14277 ( .IN1(n8817), .IN2(g1600), .Q(n13593) );
  INVX0 U14278 ( .INP(n11898), .ZN(n8817) );
  OR2X1 U14279 ( .IN1(g1624), .IN2(n8831), .Q(n11898) );
  AND2X1 U14280 ( .IN1(g25167), .IN2(g1620), .Q(n13592) );
  AND2X1 U14281 ( .IN1(n9047), .IN2(n11878), .Q(n3646) );
  AND2X1 U14282 ( .IN1(n9141), .IN2(g1657), .Q(n13587) );
  AND2X1 U14283 ( .IN1(n13034), .IN2(g1604), .Q(n13586) );
  AND3X1 U14284 ( .IN1(g1657), .IN2(g1624), .IN3(n11878), .Q(n13034) );
  INVX0 U14285 ( .INP(n13590), .ZN(n11878) );
  OR2X1 U14286 ( .IN1(n13599), .IN2(n13516), .Q(n13590) );
  OR2X1 U14287 ( .IN1(n13451), .IN2(n12797), .Q(n13516) );
  OR2X1 U14288 ( .IN1(g2715), .IN2(g2719), .Q(n12797) );
  AND2X1 U14289 ( .IN1(n13600), .IN2(n10197), .Q(n13451) );
  INVX0 U14290 ( .INP(n4388), .ZN(n13600) );
  AND2X1 U14291 ( .IN1(n10197), .IN2(g2771), .Q(n13599) );
  AND2X1 U14292 ( .IN1(n5301), .IN2(n8676), .Q(n10197) );
  OR3X1 U14293 ( .IN1(n13601), .IN2(n13602), .IN3(n13603), .Q(g29239) );
  AND3X1 U14294 ( .IN1(n13604), .IN2(n11258), .IN3(n13605), .Q(n13603) );
  INVX0 U14295 ( .INP(n13606), .ZN(n11258) );
  AND3X1 U14296 ( .IN1(n13607), .IN2(g1454), .IN3(n9076), .Q(n13602) );
  OR3X1 U14297 ( .IN1(n8741), .IN2(n13604), .IN3(n13606), .Q(n13607) );
  INVX0 U14298 ( .INP(n13608), .ZN(n13604) );
  OR2X1 U14299 ( .IN1(n13609), .IN2(n13610), .Q(n13608) );
  AND2X1 U14300 ( .IN1(n13611), .IN2(g1448), .Q(n13610) );
  AND2X1 U14301 ( .IN1(n5343), .IN2(n13612), .Q(n13609) );
  AND2X1 U14302 ( .IN1(n9141), .IN2(g1478), .Q(n13601) );
  OR3X1 U14303 ( .IN1(n13613), .IN2(n13614), .IN3(n13615), .Q(g29238) );
  AND2X1 U14304 ( .IN1(n13616), .IN2(g1484), .Q(n13615) );
  AND4X1 U14305 ( .IN1(n13617), .IN2(n13618), .IN3(n13619), .IN4(n9049), .Q(
        n13614) );
  OR2X1 U14306 ( .IN1(n13620), .IN2(g1484), .Q(n13619) );
  AND3X1 U14307 ( .IN1(n8551), .IN2(n5850), .IN3(n13621), .Q(n13620) );
  OR2X1 U14308 ( .IN1(n13611), .IN2(g1300), .Q(n13618) );
  OR2X1 U14309 ( .IN1(n5483), .IN2(n13612), .Q(n13617) );
  AND2X1 U14310 ( .IN1(n9141), .IN2(g1472), .Q(n13613) );
  OR3X1 U14311 ( .IN1(n13622), .IN2(n13623), .IN3(n13624), .Q(g29237) );
  AND3X1 U14312 ( .IN1(n13605), .IN2(n11216), .IN3(n13625), .Q(n13624) );
  AND3X1 U14313 ( .IN1(n13626), .IN2(g1467), .IN3(n9076), .Q(n13623) );
  OR3X1 U14314 ( .IN1(n8741), .IN2(n13625), .IN3(n13627), .Q(n13626) );
  INVX0 U14315 ( .INP(n13628), .ZN(n13625) );
  OR2X1 U14316 ( .IN1(n13629), .IN2(n13630), .Q(n13628) );
  AND2X1 U14317 ( .IN1(n13611), .IN2(g1472), .Q(n13630) );
  AND2X1 U14318 ( .IN1(n5290), .IN2(n13612), .Q(n13629) );
  AND2X1 U14319 ( .IN1(n9151), .IN2(g1448), .Q(n13622) );
  OR3X1 U14320 ( .IN1(n13631), .IN2(n13632), .IN3(n13633), .Q(g29236) );
  AND3X1 U14321 ( .IN1(n13605), .IN2(n11300), .IN3(n13634), .Q(n13633) );
  INVX0 U14322 ( .INP(n13635), .ZN(n11300) );
  AND4X1 U14323 ( .IN1(n5850), .IN2(n8551), .IN3(g13272), .IN4(n9050), .Q(
        n13605) );
  AND3X1 U14324 ( .IN1(n13636), .IN2(g1437), .IN3(n9076), .Q(n13632) );
  OR3X1 U14325 ( .IN1(n8741), .IN2(n13634), .IN3(n13635), .Q(n13636) );
  INVX0 U14326 ( .INP(n13637), .ZN(n13634) );
  OR2X1 U14327 ( .IN1(n13638), .IN2(n13639), .Q(n13637) );
  AND2X1 U14328 ( .IN1(n13611), .IN2(g1478), .Q(n13639) );
  INVX0 U14329 ( .INP(n13612), .ZN(n13611) );
  AND2X1 U14330 ( .IN1(n5289), .IN2(n13612), .Q(n13638) );
  OR2X1 U14331 ( .IN1(n9854), .IN2(n9267), .Q(n13612) );
  AND2X1 U14332 ( .IN1(n9151), .IN2(g1442), .Q(n13631) );
  OR3X1 U14333 ( .IN1(n13640), .IN2(n13641), .IN3(n13642), .Q(g29235) );
  AND2X1 U14334 ( .IN1(n9151), .IN2(g1252), .Q(n13642) );
  AND2X1 U14335 ( .IN1(n4178), .IN2(n5558), .Q(n13641) );
  AND3X1 U14336 ( .IN1(n11485), .IN2(n13643), .IN3(g1256), .Q(n13640) );
  INVX0 U14337 ( .INP(n4178), .ZN(n13643) );
  OR3X1 U14338 ( .IN1(n13644), .IN2(n13645), .IN3(n13646), .Q(g29234) );
  AND3X1 U14339 ( .IN1(n13647), .IN2(n11430), .IN3(n13648), .Q(n13646) );
  AND3X1 U14340 ( .IN1(test_so90), .IN2(n13649), .IN3(n9076), .Q(n13645) );
  OR3X1 U14341 ( .IN1(n8748), .IN2(n13647), .IN3(n13650), .Q(n13649) );
  INVX0 U14342 ( .INP(n13651), .ZN(n13647) );
  OR2X1 U14343 ( .IN1(n13652), .IN2(n13653), .Q(n13651) );
  AND2X1 U14344 ( .IN1(n13654), .IN2(g1105), .Q(n13653) );
  AND2X1 U14345 ( .IN1(n5478), .IN2(n13655), .Q(n13652) );
  AND2X1 U14346 ( .IN1(n9151), .IN2(g1135), .Q(n13644) );
  OR3X1 U14347 ( .IN1(n13656), .IN2(n13657), .IN3(n13658), .Q(g29233) );
  AND2X1 U14348 ( .IN1(n13659), .IN2(g1141), .Q(n13658) );
  AND4X1 U14349 ( .IN1(n13660), .IN2(n13661), .IN3(n13662), .IN4(n9050), .Q(
        n13657) );
  OR2X1 U14350 ( .IN1(n13663), .IN2(g1141), .Q(n13662) );
  AND3X1 U14351 ( .IN1(n5851), .IN2(n8820), .IN3(n13664), .Q(n13663) );
  OR2X1 U14352 ( .IN1(n13654), .IN2(g956), .Q(n13661) );
  OR2X1 U14353 ( .IN1(n5341), .IN2(n13655), .Q(n13660) );
  AND2X1 U14354 ( .IN1(n9151), .IN2(g1129), .Q(n13656) );
  OR3X1 U14355 ( .IN1(n13665), .IN2(n13666), .IN3(n13667), .Q(g29232) );
  AND3X1 U14356 ( .IN1(n13648), .IN2(n11387), .IN3(n13668), .Q(n13667) );
  INVX0 U14357 ( .INP(n13669), .ZN(n13668) );
  AND3X1 U14358 ( .IN1(n13670), .IN2(g1124), .IN3(n9075), .Q(n13666) );
  INVX0 U14359 ( .INP(n13671), .ZN(n13670) );
  AND3X1 U14360 ( .IN1(g13259), .IN2(n13669), .IN3(n11387), .Q(n13671) );
  OR2X1 U14361 ( .IN1(n13672), .IN2(n13673), .Q(n13669) );
  AND2X1 U14362 ( .IN1(n13654), .IN2(g1129), .Q(n13673) );
  AND2X1 U14363 ( .IN1(n5329), .IN2(n13655), .Q(n13672) );
  AND2X1 U14364 ( .IN1(n9151), .IN2(g1105), .Q(n13665) );
  OR3X1 U14365 ( .IN1(n13674), .IN2(n13675), .IN3(n13676), .Q(g29231) );
  AND4X1 U14366 ( .IN1(n13677), .IN2(n13648), .IN3(n5599), .IN4(g1171), .Q(
        n13676) );
  AND4X1 U14367 ( .IN1(n9048), .IN2(n5851), .IN3(n8820), .IN4(g13259), .Q(
        n13648) );
  AND3X1 U14368 ( .IN1(n13678), .IN2(g1094), .IN3(n9074), .Q(n13675) );
  OR4X1 U14369 ( .IN1(n13677), .IN2(g1183), .IN3(n8748), .IN4(n5363), .Q(
        n13678) );
  INVX0 U14370 ( .INP(n13679), .ZN(n13677) );
  OR2X1 U14371 ( .IN1(n13680), .IN2(n13681), .Q(n13679) );
  AND2X1 U14372 ( .IN1(n13654), .IN2(g1135), .Q(n13681) );
  INVX0 U14373 ( .INP(n13655), .ZN(n13654) );
  AND2X1 U14374 ( .IN1(n5328), .IN2(n13655), .Q(n13680) );
  OR2X1 U14375 ( .IN1(n9855), .IN2(n9367), .Q(n13655) );
  INVX0 U14376 ( .INP(n11471), .ZN(n9855) );
  AND2X1 U14377 ( .IN1(test_so7), .IN2(n9140), .Q(n13674) );
  OR3X1 U14378 ( .IN1(n13682), .IN2(n13683), .IN3(n13684), .Q(g29230) );
  AND2X1 U14379 ( .IN1(n9151), .IN2(g907), .Q(n13684) );
  AND2X1 U14380 ( .IN1(n4196), .IN2(n5559), .Q(n13683) );
  AND3X1 U14381 ( .IN1(n11500), .IN2(n13685), .IN3(g911), .Q(n13682) );
  INVX0 U14382 ( .INP(n4196), .ZN(n13685) );
  OR3X1 U14383 ( .IN1(n13686), .IN2(n13687), .IN3(n13688), .Q(g29229) );
  AND2X1 U14384 ( .IN1(n9151), .IN2(g827), .Q(n13688) );
  AND3X1 U14385 ( .IN1(n4516), .IN2(n13689), .IN3(n5826), .Q(n13687) );
  AND2X1 U14386 ( .IN1(n4517), .IN2(g723), .Q(n13686) );
  OR2X1 U14387 ( .IN1(n13690), .IN2(n13691), .Q(g29228) );
  AND2X1 U14388 ( .IN1(n9151), .IN2(g736), .Q(n13691) );
  AND2X1 U14389 ( .IN1(n2404), .IN2(n13692), .Q(n13690) );
  OR2X1 U14390 ( .IN1(n13693), .IN2(n13694), .Q(n13692) );
  AND2X1 U14391 ( .IN1(n13133), .IN2(n8853), .Q(n13694) );
  INVX0 U14392 ( .INP(n13695), .ZN(n13133) );
  AND2X1 U14393 ( .IN1(test_so60), .IN2(n13695), .Q(n13693) );
  OR2X1 U14394 ( .IN1(n13696), .IN2(n13145), .Q(n13695) );
  AND2X1 U14395 ( .IN1(n5482), .IN2(g12184), .Q(n13696) );
  OR3X1 U14396 ( .IN1(n13697), .IN2(n13698), .IN3(n13699), .Q(g29227) );
  AND2X1 U14397 ( .IN1(n9151), .IN2(g676), .Q(n13699) );
  AND2X1 U14398 ( .IN1(n4524), .IN2(test_so70), .Q(n13698) );
  AND3X1 U14399 ( .IN1(n4523), .IN2(n13700), .IN3(n8852), .Q(n13697) );
  OR3X1 U14400 ( .IN1(n13701), .IN2(n13702), .IN3(n13703), .Q(g29226) );
  AND2X1 U14401 ( .IN1(n9151), .IN2(g671), .Q(n13703) );
  AND3X1 U14402 ( .IN1(n4526), .IN2(n13700), .IN3(n5751), .Q(n13702) );
  AND3X1 U14403 ( .IN1(n4525), .IN2(n13704), .IN3(g676), .Q(n13701) );
  INVX0 U14404 ( .INP(n4526), .ZN(n13704) );
  OR2X1 U14405 ( .IN1(n13705), .IN2(n13706), .Q(g29225) );
  AND2X1 U14406 ( .IN1(n9151), .IN2(g667), .Q(n13706) );
  AND3X1 U14407 ( .IN1(n13707), .IN2(n13708), .IN3(n4525), .Q(n13705) );
  AND2X1 U14408 ( .IN1(n9047), .IN2(n13700), .Q(n4525) );
  AND2X1 U14409 ( .IN1(g703), .IN2(n13709), .Q(n13700) );
  OR4X1 U14410 ( .IN1(n4535), .IN2(n13710), .IN3(n158), .IN4(n8678), .Q(n13709) );
  OR2X1 U14411 ( .IN1(n13711), .IN2(n13712), .Q(n4535) );
  AND2X1 U14412 ( .IN1(n8784), .IN2(g718), .Q(n13712) );
  AND2X1 U14413 ( .IN1(n8785), .IN2(g655), .Q(n13711) );
  OR2X1 U14414 ( .IN1(n13713), .IN2(g671), .Q(n13708) );
  OR2X1 U14415 ( .IN1(n8307), .IN2(n158), .Q(n13707) );
  INVX0 U14416 ( .INP(n13713), .ZN(n158) );
  OR3X1 U14417 ( .IN1(n13714), .IN2(n13715), .IN3(n13716), .Q(g29224) );
  AND2X1 U14418 ( .IN1(n9151), .IN2(g572), .Q(n13716) );
  AND2X1 U14419 ( .IN1(n4201), .IN2(n5336), .Q(n13715) );
  AND3X1 U14420 ( .IN1(n2421), .IN2(n13717), .IN3(g586), .Q(n13714) );
  INVX0 U14421 ( .INP(n4201), .ZN(n13717) );
  OR4X1 U14422 ( .IN1(n13718), .IN2(n13719), .IN3(n13720), .IN4(n13721), .Q(
        g29223) );
  AND2X1 U14423 ( .IN1(n9151), .IN2(g482), .Q(n13721) );
  AND3X1 U14424 ( .IN1(n13722), .IN2(g490), .IN3(n9074), .Q(n13720) );
  AND2X1 U14425 ( .IN1(n13723), .IN2(n5708), .Q(n13719) );
  INVX0 U14426 ( .INP(n13722), .ZN(n13723) );
  OR3X1 U14427 ( .IN1(n13724), .IN2(n13725), .IN3(n13726), .Q(g29222) );
  AND2X1 U14428 ( .IN1(n13727), .IN2(g411), .Q(n13726) );
  AND3X1 U14429 ( .IN1(n13728), .IN2(n517), .IN3(n5358), .Q(n13725) );
  INVX0 U14430 ( .INP(n13729), .ZN(n517) );
  AND2X1 U14431 ( .IN1(n13730), .IN2(g417), .Q(n13724) );
  OR2X1 U14432 ( .IN1(n9134), .IN2(n13731), .Q(n13730) );
  AND2X1 U14433 ( .IN1(n4948), .IN2(n13729), .Q(n13731) );
  AND2X1 U14434 ( .IN1(n13732), .IN2(n13733), .Q(n13729) );
  OR2X1 U14435 ( .IN1(n13734), .IN2(n5358), .Q(n13733) );
  INVX0 U14436 ( .INP(n13735), .ZN(n13734) );
  OR2X1 U14437 ( .IN1(n13735), .IN2(g417), .Q(n13732) );
  OR2X1 U14438 ( .IN1(n13736), .IN2(n13737), .Q(n13735) );
  AND2X1 U14439 ( .IN1(n13738), .IN2(n8674), .Q(n13737) );
  OR2X1 U14440 ( .IN1(n13739), .IN2(n13740), .Q(n13738) );
  AND2X1 U14441 ( .IN1(n8673), .IN2(g424), .Q(n13740) );
  AND2X1 U14442 ( .IN1(g437), .IN2(g392), .Q(n13739) );
  AND2X1 U14443 ( .IN1(n13741), .IN2(g405), .Q(n13736) );
  OR2X1 U14444 ( .IN1(n13742), .IN2(n13743), .Q(n13741) );
  AND2X1 U14445 ( .IN1(g401), .IN2(g392), .Q(n13743) );
  AND2X1 U14446 ( .IN1(n8673), .IN2(g437), .Q(n13742) );
  OR3X1 U14447 ( .IN1(n13744), .IN2(n13745), .IN3(n13746), .Q(g28105) );
  AND2X1 U14448 ( .IN1(n11010), .IN2(g5011), .Q(n13746) );
  AND3X1 U14449 ( .IN1(n13181), .IN2(n11004), .IN3(n9074), .Q(n13745) );
  INVX0 U14450 ( .INP(n8809), .ZN(n11004) );
  OR2X1 U14451 ( .IN1(n13747), .IN2(n13748), .Q(n13181) );
  AND2X1 U14452 ( .IN1(n13749), .IN2(g6727), .Q(n13748) );
  OR4X1 U14453 ( .IN1(n13750), .IN2(n13751), .IN3(n13752), .IN4(n13753), .Q(
        n13749) );
  OR3X1 U14454 ( .IN1(n13754), .IN2(n13755), .IN3(n13756), .Q(n13753) );
  AND2X1 U14455 ( .IN1(n9366), .IN2(n13757), .Q(n13756) );
  OR2X1 U14456 ( .IN1(n13758), .IN2(n13759), .Q(n13757) );
  AND2X1 U14457 ( .IN1(g6641), .IN2(g17764), .Q(n13759) );
  AND2X1 U14458 ( .IN1(g6657), .IN2(g17722), .Q(n13758) );
  AND3X1 U14459 ( .IN1(g6609), .IN2(g17871), .IN3(n9365), .Q(n13755) );
  AND3X1 U14460 ( .IN1(g14749), .IN2(g6625), .IN3(n9369), .Q(n13754) );
  AND2X1 U14461 ( .IN1(n9368), .IN2(n13760), .Q(n13752) );
  OR2X1 U14462 ( .IN1(n13761), .IN2(n13762), .Q(n13760) );
  AND2X1 U14463 ( .IN1(g6581), .IN2(g13099), .Q(n13762) );
  AND2X1 U14464 ( .IN1(g6589), .IN2(g6723), .Q(n13761) );
  AND2X1 U14465 ( .IN1(test_so80), .IN2(n13763), .Q(n13751) );
  OR2X1 U14466 ( .IN1(n13764), .IN2(n13765), .Q(n13763) );
  AND2X1 U14467 ( .IN1(test_so71), .IN2(n9365), .Q(n13764) );
  AND2X1 U14468 ( .IN1(n13766), .IN2(n8840), .Q(n13750) );
  AND2X1 U14469 ( .IN1(n5531), .IN2(n13767), .Q(n13747) );
  OR4X1 U14470 ( .IN1(n13768), .IN2(n13769), .IN3(n13770), .IN4(n13771), .Q(
        n13767) );
  OR3X1 U14471 ( .IN1(n13772), .IN2(n13773), .IN3(n13774), .Q(n13771) );
  AND2X1 U14472 ( .IN1(n9369), .IN2(n13775), .Q(n13774) );
  OR2X1 U14473 ( .IN1(n13776), .IN2(n13777), .Q(n13775) );
  AND2X1 U14474 ( .IN1(g6593), .IN2(g13099), .Q(n13777) );
  AND2X1 U14475 ( .IN1(g6723), .IN2(g6605), .Q(n13776) );
  AND3X1 U14476 ( .IN1(g14749), .IN2(g6633), .IN3(n9368), .Q(n13773) );
  AND3X1 U14477 ( .IN1(g17871), .IN2(g6617), .IN3(n9366), .Q(n13772) );
  AND2X1 U14478 ( .IN1(n9365), .IN2(n13778), .Q(n13770) );
  OR2X1 U14479 ( .IN1(n13779), .IN2(n13780), .Q(n13778) );
  AND2X1 U14480 ( .IN1(g6597), .IN2(g17722), .Q(n13780) );
  AND2X1 U14481 ( .IN1(g17764), .IN2(g6649), .Q(n13779) );
  AND2X1 U14482 ( .IN1(test_so80), .IN2(n13781), .Q(n13769) );
  OR2X1 U14483 ( .IN1(n13782), .IN2(n13766), .Q(n13781) );
  OR3X1 U14484 ( .IN1(n13783), .IN2(n13784), .IN3(n13785), .Q(n13766) );
  AND3X1 U14485 ( .IN1(g14828), .IN2(g6621), .IN3(n9368), .Q(n13785) );
  AND3X1 U14486 ( .IN1(g6637), .IN2(g17778), .IN3(n9365), .Q(n13784) );
  AND2X1 U14487 ( .IN1(g6741), .IN2(n5590), .Q(n9365) );
  AND3X1 U14488 ( .IN1(g6653), .IN2(g17688), .IN3(n9369), .Q(n13783) );
  AND2X1 U14489 ( .IN1(n9366), .IN2(g6601), .Q(n13782) );
  AND2X1 U14490 ( .IN1(n13765), .IN2(n8840), .Q(n13768) );
  OR3X1 U14491 ( .IN1(n13786), .IN2(n13787), .IN3(n13788), .Q(n13765) );
  AND3X1 U14492 ( .IN1(g6645), .IN2(g17688), .IN3(n9368), .Q(n13788) );
  AND2X1 U14493 ( .IN1(n5590), .IN2(n5398), .Q(n9368) );
  AND3X1 U14494 ( .IN1(g14828), .IN2(g6613), .IN3(n9369), .Q(n13787) );
  AND2X1 U14495 ( .IN1(g6682), .IN2(n5398), .Q(n9369) );
  AND3X1 U14496 ( .IN1(g6629), .IN2(g17778), .IN3(n9366), .Q(n13786) );
  AND2X1 U14497 ( .IN1(g6682), .IN2(g6741), .Q(n9366) );
  AND2X1 U14498 ( .IN1(n9151), .IN2(g6657), .Q(n13744) );
  OR3X1 U14499 ( .IN1(n13789), .IN2(n13790), .IN3(n13791), .Q(g28102) );
  AND2X1 U14500 ( .IN1(n11027), .IN2(g4826), .Q(n13791) );
  AND3X1 U14501 ( .IN1(n11019), .IN2(n13216), .IN3(n9077), .Q(n13790) );
  OR2X1 U14502 ( .IN1(n13792), .IN2(n13793), .Q(n13216) );
  AND2X1 U14503 ( .IN1(n13794), .IN2(n8829), .Q(n13793) );
  OR4X1 U14504 ( .IN1(n13795), .IN2(n13796), .IN3(n13797), .IN4(n13798), .Q(
        n13794) );
  OR3X1 U14505 ( .IN1(n13799), .IN2(n13800), .IN3(n13801), .Q(n13798) );
  AND2X1 U14506 ( .IN1(n11018), .IN2(n13802), .Q(n13801) );
  OR2X1 U14507 ( .IN1(n13803), .IN2(n13804), .Q(n13802) );
  AND2X1 U14508 ( .IN1(g6251), .IN2(g17685), .Q(n13804) );
  AND2X1 U14509 ( .IN1(g17743), .IN2(g6303), .Q(n13803) );
  AND3X1 U14510 ( .IN1(g17845), .IN2(g6271), .IN3(n10232), .Q(n13800) );
  AND3X1 U14511 ( .IN1(g14705), .IN2(g6287), .IN3(n13805), .Q(n13799) );
  AND2X1 U14512 ( .IN1(n11022), .IN2(n13806), .Q(n13797) );
  OR2X1 U14513 ( .IN1(n13807), .IN2(n13808), .Q(n13806) );
  AND2X1 U14514 ( .IN1(g6247), .IN2(g13085), .Q(n13808) );
  AND2X1 U14515 ( .IN1(g6377), .IN2(g6259), .Q(n13807) );
  AND2X1 U14516 ( .IN1(n13809), .IN2(g12422), .Q(n13796) );
  OR2X1 U14517 ( .IN1(n13810), .IN2(n13811), .Q(n13809) );
  AND2X1 U14518 ( .IN1(n10232), .IN2(g6255), .Q(n13810) );
  AND2X1 U14519 ( .IN1(n5437), .IN2(n13812), .Q(n13795) );
  AND2X1 U14520 ( .IN1(test_so69), .IN2(n13813), .Q(n13792) );
  OR4X1 U14521 ( .IN1(n13814), .IN2(n13815), .IN3(n13816), .IN4(n13817), .Q(
        n13813) );
  OR3X1 U14522 ( .IN1(n13818), .IN2(n13819), .IN3(n13820), .Q(n13817) );
  AND2X1 U14523 ( .IN1(n13805), .IN2(n13821), .Q(n13820) );
  OR2X1 U14524 ( .IN1(n13822), .IN2(n13823), .Q(n13821) );
  AND2X1 U14525 ( .IN1(g6235), .IN2(g13085), .Q(n13823) );
  AND2X1 U14526 ( .IN1(g6243), .IN2(g6377), .Q(n13822) );
  AND3X1 U14527 ( .IN1(g14705), .IN2(g6279), .IN3(n11022), .Q(n13819) );
  AND3X1 U14528 ( .IN1(g6263), .IN2(g17845), .IN3(n11018), .Q(n13818) );
  AND2X1 U14529 ( .IN1(n10232), .IN2(n13824), .Q(n13816) );
  OR2X1 U14530 ( .IN1(n13825), .IN2(n13826), .Q(n13824) );
  AND2X1 U14531 ( .IN1(g6295), .IN2(g17743), .Q(n13826) );
  AND2X1 U14532 ( .IN1(g6311), .IN2(g17685), .Q(n13825) );
  AND2X1 U14533 ( .IN1(n13827), .IN2(g12422), .Q(n13815) );
  OR2X1 U14534 ( .IN1(n13828), .IN2(n13812), .Q(n13827) );
  OR3X1 U14535 ( .IN1(n13829), .IN2(n13830), .IN3(n13831), .Q(n13812) );
  AND3X1 U14536 ( .IN1(g14779), .IN2(g6267), .IN3(n11022), .Q(n13831) );
  AND3X1 U14537 ( .IN1(g6283), .IN2(g17760), .IN3(n10232), .Q(n13830) );
  AND3X1 U14538 ( .IN1(g6299), .IN2(g17649), .IN3(n13805), .Q(n13829) );
  AND2X1 U14539 ( .IN1(n11018), .IN2(g6239), .Q(n13828) );
  AND2X1 U14540 ( .IN1(n5437), .IN2(n13811), .Q(n13814) );
  OR3X1 U14541 ( .IN1(n13832), .IN2(n13833), .IN3(n13834), .Q(n13811) );
  AND3X1 U14542 ( .IN1(g6307), .IN2(g17649), .IN3(n11022), .Q(n13834) );
  AND3X1 U14543 ( .IN1(g6291), .IN2(g17760), .IN3(n11018), .Q(n13833) );
  AND3X1 U14544 ( .IN1(g14779), .IN2(g6275), .IN3(n13805), .Q(n13832) );
  AND2X1 U14545 ( .IN1(n9150), .IN2(g6311), .Q(n13789) );
  OR3X1 U14546 ( .IN1(n13835), .IN2(n13836), .IN3(n13837), .Q(g28099) );
  AND2X1 U14547 ( .IN1(n11044), .IN2(g4831), .Q(n13837) );
  AND3X1 U14548 ( .IN1(n11036), .IN2(n13251), .IN3(n9057), .Q(n13836) );
  OR2X1 U14549 ( .IN1(n13838), .IN2(n13839), .Q(n13251) );
  AND2X1 U14550 ( .IN1(n13840), .IN2(g6035), .Q(n13839) );
  OR4X1 U14551 ( .IN1(n13841), .IN2(n13842), .IN3(n13843), .IN4(n13844), .Q(
        n13840) );
  OR3X1 U14552 ( .IN1(n13845), .IN2(n13846), .IN3(n13847), .Q(n13844) );
  AND2X1 U14553 ( .IN1(n13848), .IN2(n13849), .Q(n13847) );
  OR2X1 U14554 ( .IN1(n13850), .IN2(n13851), .Q(n13849) );
  AND2X1 U14555 ( .IN1(g5889), .IN2(g13068), .Q(n13851) );
  AND2X1 U14556 ( .IN1(g5897), .IN2(g6031), .Q(n13850) );
  AND3X1 U14557 ( .IN1(g14673), .IN2(g5933), .IN3(n11039), .Q(n13846) );
  AND3X1 U14558 ( .IN1(n11035), .IN2(g17819), .IN3(test_so28), .Q(n13845) );
  AND2X1 U14559 ( .IN1(n10245), .IN2(n13852), .Q(n13843) );
  OR2X1 U14560 ( .IN1(n13853), .IN2(n13854), .Q(n13852) );
  AND2X1 U14561 ( .IN1(test_so13), .IN2(g17646), .Q(n13854) );
  AND2X1 U14562 ( .IN1(g5949), .IN2(g17715), .Q(n13853) );
  AND2X1 U14563 ( .IN1(n13855), .IN2(g12350), .Q(n13842) );
  OR2X1 U14564 ( .IN1(n13856), .IN2(n13857), .Q(n13855) );
  AND2X1 U14565 ( .IN1(n11035), .IN2(g5893), .Q(n13856) );
  AND2X1 U14566 ( .IN1(n5432), .IN2(n13858), .Q(n13841) );
  AND2X1 U14567 ( .IN1(n5528), .IN2(n13859), .Q(n13838) );
  OR4X1 U14568 ( .IN1(n13860), .IN2(n13861), .IN3(n13862), .IN4(n13863), .Q(
        n13859) );
  OR3X1 U14569 ( .IN1(n13864), .IN2(n13865), .IN3(n13866), .Q(n13863) );
  AND2X1 U14570 ( .IN1(n11035), .IN2(n13867), .Q(n13866) );
  OR2X1 U14571 ( .IN1(n13868), .IN2(n13869), .Q(n13867) );
  AND2X1 U14572 ( .IN1(g5905), .IN2(g17646), .Q(n13869) );
  AND2X1 U14573 ( .IN1(g17715), .IN2(g5957), .Q(n13868) );
  AND3X1 U14574 ( .IN1(g17819), .IN2(g5925), .IN3(n10245), .Q(n13865) );
  AND3X1 U14575 ( .IN1(g14673), .IN2(g5941), .IN3(n13848), .Q(n13864) );
  AND2X1 U14576 ( .IN1(n11039), .IN2(n13870), .Q(n13862) );
  OR2X1 U14577 ( .IN1(n13871), .IN2(n13872), .Q(n13870) );
  AND2X1 U14578 ( .IN1(g5901), .IN2(g13068), .Q(n13872) );
  AND2X1 U14579 ( .IN1(g6031), .IN2(g5913), .Q(n13871) );
  AND2X1 U14580 ( .IN1(n13873), .IN2(g12350), .Q(n13861) );
  OR2X1 U14581 ( .IN1(n13874), .IN2(n13858), .Q(n13873) );
  OR3X1 U14582 ( .IN1(n13875), .IN2(n13876), .IN3(n13877), .Q(n13858) );
  AND3X1 U14583 ( .IN1(g5961), .IN2(g17607), .IN3(n11039), .Q(n13877) );
  AND3X1 U14584 ( .IN1(g5945), .IN2(g17739), .IN3(n11035), .Q(n13876) );
  AND3X1 U14585 ( .IN1(g14738), .IN2(g5929), .IN3(n13848), .Q(n13875) );
  AND2X1 U14586 ( .IN1(n10245), .IN2(g5909), .Q(n13874) );
  AND2X1 U14587 ( .IN1(n5432), .IN2(n13857), .Q(n13860) );
  OR3X1 U14588 ( .IN1(n13878), .IN2(n13879), .IN3(n13880), .Q(n13857) );
  AND3X1 U14589 ( .IN1(g14738), .IN2(g5921), .IN3(n11039), .Q(n13880) );
  AND3X1 U14590 ( .IN1(g5937), .IN2(g17739), .IN3(n10245), .Q(n13879) );
  AND3X1 U14591 ( .IN1(g5953), .IN2(g17607), .IN3(n13848), .Q(n13878) );
  AND2X1 U14592 ( .IN1(test_so13), .IN2(n9138), .Q(n13835) );
  OR3X1 U14593 ( .IN1(n13881), .IN2(n13882), .IN3(n13883), .Q(g28096) );
  AND2X1 U14594 ( .IN1(n11060), .IN2(g4821), .Q(n13883) );
  AND3X1 U14595 ( .IN1(n11052), .IN2(n13286), .IN3(n9058), .Q(n13882) );
  OR2X1 U14596 ( .IN1(n13884), .IN2(n13885), .Q(n13286) );
  AND2X1 U14597 ( .IN1(n13886), .IN2(g5689), .Q(n13885) );
  OR4X1 U14598 ( .IN1(n13887), .IN2(n13888), .IN3(n13889), .IN4(n13890), .Q(
        n13886) );
  OR3X1 U14599 ( .IN1(n13891), .IN2(n13892), .IN3(n13893), .Q(n13890) );
  AND2X1 U14600 ( .IN1(n13894), .IN2(n13895), .Q(n13893) );
  OR2X1 U14601 ( .IN1(n13896), .IN2(n13897), .Q(n13895) );
  AND2X1 U14602 ( .IN1(g5543), .IN2(g13049), .Q(n13897) );
  AND2X1 U14603 ( .IN1(g5551), .IN2(g5685), .Q(n13896) );
  AND3X1 U14604 ( .IN1(g14635), .IN2(g5587), .IN3(n11055), .Q(n13892) );
  AND3X1 U14605 ( .IN1(g5571), .IN2(g17813), .IN3(n11051), .Q(n13891) );
  AND2X1 U14606 ( .IN1(n10237), .IN2(n13898), .Q(n13889) );
  OR2X1 U14607 ( .IN1(n13899), .IN2(n13900), .Q(n13898) );
  AND2X1 U14608 ( .IN1(g5603), .IN2(g17678), .Q(n13900) );
  AND2X1 U14609 ( .IN1(g5619), .IN2(g17604), .Q(n13899) );
  AND2X1 U14610 ( .IN1(n13901), .IN2(g12300), .Q(n13888) );
  OR2X1 U14611 ( .IN1(n13902), .IN2(n13903), .Q(n13901) );
  AND2X1 U14612 ( .IN1(n11051), .IN2(g5547), .Q(n13902) );
  AND2X1 U14613 ( .IN1(n5439), .IN2(n13904), .Q(n13887) );
  AND2X1 U14614 ( .IN1(n5529), .IN2(n13905), .Q(n13884) );
  OR4X1 U14615 ( .IN1(n13906), .IN2(n13907), .IN3(n13908), .IN4(n13909), .Q(
        n13905) );
  OR3X1 U14616 ( .IN1(n13910), .IN2(n13911), .IN3(n13912), .Q(n13909) );
  AND2X1 U14617 ( .IN1(n11051), .IN2(n13913), .Q(n13912) );
  OR2X1 U14618 ( .IN1(n13914), .IN2(n13915), .Q(n13913) );
  AND2X1 U14619 ( .IN1(test_so6), .IN2(g17604), .Q(n13915) );
  AND2X1 U14620 ( .IN1(g17678), .IN2(g5611), .Q(n13914) );
  AND3X1 U14621 ( .IN1(g17813), .IN2(g5579), .IN3(n10237), .Q(n13911) );
  AND3X1 U14622 ( .IN1(g14635), .IN2(g5595), .IN3(n13894), .Q(n13910) );
  AND2X1 U14623 ( .IN1(n11055), .IN2(n13916), .Q(n13908) );
  OR2X1 U14624 ( .IN1(n13917), .IN2(n13918), .Q(n13916) );
  AND2X1 U14625 ( .IN1(g5555), .IN2(g13049), .Q(n13918) );
  AND2X1 U14626 ( .IN1(g5685), .IN2(g5567), .Q(n13917) );
  AND2X1 U14627 ( .IN1(n13919), .IN2(g12300), .Q(n13907) );
  OR2X1 U14628 ( .IN1(n13920), .IN2(n13904), .Q(n13919) );
  OR3X1 U14629 ( .IN1(n13921), .IN2(n13922), .IN3(n13923), .Q(n13904) );
  AND3X1 U14630 ( .IN1(g5615), .IN2(g17580), .IN3(n11055), .Q(n13923) );
  AND3X1 U14631 ( .IN1(g5599), .IN2(g17711), .IN3(n11051), .Q(n13922) );
  AND3X1 U14632 ( .IN1(g14694), .IN2(g5583), .IN3(n13894), .Q(n13921) );
  AND2X1 U14633 ( .IN1(n10237), .IN2(g5563), .Q(n13920) );
  AND2X1 U14634 ( .IN1(n5439), .IN2(n13903), .Q(n13906) );
  OR3X1 U14635 ( .IN1(n13924), .IN2(n13925), .IN3(n13926), .Q(n13903) );
  AND3X1 U14636 ( .IN1(g14694), .IN2(g5575), .IN3(n11055), .Q(n13926) );
  AND3X1 U14637 ( .IN1(n10237), .IN2(g17711), .IN3(test_so5), .Q(n13925) );
  AND3X1 U14638 ( .IN1(g5607), .IN2(g17580), .IN3(n13894), .Q(n13924) );
  AND2X1 U14639 ( .IN1(n9150), .IN2(g5619), .Q(n13881) );
  OR3X1 U14640 ( .IN1(n13927), .IN2(n13928), .IN3(n13929), .Q(g28093) );
  AND2X1 U14641 ( .IN1(n11072), .IN2(g29220), .Q(n13929) );
  AND3X1 U14642 ( .IN1(n13321), .IN2(g33959), .IN3(n9058), .Q(n13928) );
  INVX0 U14643 ( .INP(n8804), .ZN(g33959) );
  OR2X1 U14644 ( .IN1(n13930), .IN2(n13931), .Q(n13321) );
  AND2X1 U14645 ( .IN1(n13932), .IN2(n8828), .Q(n13931) );
  OR4X1 U14646 ( .IN1(n13933), .IN2(n13934), .IN3(n13935), .IN4(n13936), .Q(
        n13932) );
  OR3X1 U14647 ( .IN1(n13937), .IN2(n13938), .IN3(n13939), .Q(n13936) );
  AND2X1 U14648 ( .IN1(n9359), .IN2(n13940), .Q(n13939) );
  OR2X1 U14649 ( .IN1(n13941), .IN2(n13942), .Q(n13940) );
  AND2X1 U14650 ( .IN1(g5208), .IN2(g13039), .Q(n13942) );
  AND2X1 U14651 ( .IN1(g5220), .IN2(g5339), .Q(n13941) );
  AND3X1 U14652 ( .IN1(g17787), .IN2(g5232), .IN3(g31860), .Q(n13938) );
  AND3X1 U14653 ( .IN1(g14597), .IN2(g5248), .IN3(n9358), .Q(n13937) );
  AND2X1 U14654 ( .IN1(n9360), .IN2(n13943), .Q(n13935) );
  OR2X1 U14655 ( .IN1(n13944), .IN2(n13945), .Q(n13943) );
  AND2X1 U14656 ( .IN1(g5212), .IN2(g17577), .Q(n13945) );
  AND2X1 U14657 ( .IN1(g17639), .IN2(g5264), .Q(n13944) );
  AND2X1 U14658 ( .IN1(n13946), .IN2(g12238), .Q(n13934) );
  OR2X1 U14659 ( .IN1(n13947), .IN2(n13948), .Q(n13946) );
  AND2X1 U14660 ( .IN1(g31860), .IN2(g5216), .Q(n13947) );
  AND2X1 U14661 ( .IN1(n5438), .IN2(n13949), .Q(n13933) );
  AND2X1 U14662 ( .IN1(test_so10), .IN2(n13950), .Q(n13930) );
  OR4X1 U14663 ( .IN1(n13951), .IN2(n13952), .IN3(n13953), .IN4(n13954), .Q(
        n13950) );
  OR3X1 U14664 ( .IN1(n13955), .IN2(n13956), .IN3(n13957), .Q(n13954) );
  AND2X1 U14665 ( .IN1(n9358), .IN2(n13958), .Q(n13957) );
  OR2X1 U14666 ( .IN1(n13959), .IN2(n13960), .Q(n13958) );
  AND2X1 U14667 ( .IN1(g5196), .IN2(g13039), .Q(n13960) );
  AND2X1 U14668 ( .IN1(g5339), .IN2(g5204), .Q(n13959) );
  AND3X1 U14669 ( .IN1(g5224), .IN2(g17787), .IN3(n9360), .Q(n13956) );
  AND3X1 U14670 ( .IN1(g14597), .IN2(g5240), .IN3(n9359), .Q(n13955) );
  AND2X1 U14671 ( .IN1(g31860), .IN2(n13961), .Q(n13953) );
  OR2X1 U14672 ( .IN1(n13962), .IN2(n13963), .Q(n13961) );
  AND2X1 U14673 ( .IN1(g5256), .IN2(g17639), .Q(n13963) );
  AND2X1 U14674 ( .IN1(g5272), .IN2(g17577), .Q(n13962) );
  AND2X1 U14675 ( .IN1(n13964), .IN2(g12238), .Q(n13952) );
  OR2X1 U14676 ( .IN1(n13965), .IN2(n13949), .Q(n13964) );
  OR3X1 U14677 ( .IN1(n13966), .IN2(n13967), .IN3(n13968), .Q(n13949) );
  AND3X1 U14678 ( .IN1(g5244), .IN2(g17674), .IN3(g31860), .Q(n13968) );
  AND2X1 U14679 ( .IN1(g5297), .IN2(g5357), .Q(g31860) );
  AND3X1 U14680 ( .IN1(g5260), .IN2(g17519), .IN3(n9358), .Q(n13967) );
  AND3X1 U14681 ( .IN1(n9359), .IN2(g14662), .IN3(test_so82), .Q(n13966) );
  AND2X1 U14682 ( .IN1(n9360), .IN2(g5200), .Q(n13965) );
  AND2X1 U14683 ( .IN1(n5438), .IN2(n13948), .Q(n13951) );
  OR3X1 U14684 ( .IN1(n13969), .IN2(n13970), .IN3(n13971), .Q(n13948) );
  AND3X1 U14685 ( .IN1(g5252), .IN2(g17674), .IN3(n9360), .Q(n13971) );
  AND2X1 U14686 ( .IN1(g5357), .IN2(n5588), .Q(n9360) );
  AND3X1 U14687 ( .IN1(g14662), .IN2(g5236), .IN3(n9358), .Q(n13970) );
  AND2X1 U14688 ( .IN1(n5393), .IN2(n5588), .Q(n9358) );
  AND3X1 U14689 ( .IN1(g5268), .IN2(g17519), .IN3(n9359), .Q(n13969) );
  AND2X1 U14690 ( .IN1(g5297), .IN2(n5393), .Q(n9359) );
  AND2X1 U14691 ( .IN1(n9150), .IN2(g5272), .Q(n13927) );
  OR2X1 U14692 ( .IN1(n13972), .IN2(n13973), .Q(g28092) );
  AND3X1 U14693 ( .IN1(n11996), .IN2(n11995), .IN3(n9058), .Q(n13973) );
  OR3X1 U14694 ( .IN1(g84), .IN2(n13974), .IN3(g5052), .Q(n11995) );
  OR3X1 U14695 ( .IN1(n13975), .IN2(n13974), .IN3(g5041), .Q(n11996) );
  OR3X1 U14696 ( .IN1(n8767), .IN2(n5615), .IN3(g5046), .Q(n13974) );
  AND2X1 U14697 ( .IN1(n9150), .IN2(g5057), .Q(n13972) );
  OR2X1 U14698 ( .IN1(n13976), .IN2(n13977), .Q(g28091) );
  AND3X1 U14699 ( .IN1(n11997), .IN2(n11999), .IN3(n9059), .Q(n13977) );
  OR3X1 U14700 ( .IN1(n5607), .IN2(g84), .IN3(n13978), .Q(n11999) );
  OR3X1 U14701 ( .IN1(n5605), .IN2(n13978), .IN3(n13975), .Q(n11997) );
  INVX0 U14702 ( .INP(g84), .ZN(n13975) );
  OR3X1 U14703 ( .IN1(n8768), .IN2(n5578), .IN3(g5057), .Q(n13978) );
  AND2X1 U14704 ( .IN1(n9150), .IN2(g5069), .Q(n13976) );
  OR2X1 U14705 ( .IN1(n13979), .IN2(n13980), .Q(g28090) );
  AND2X1 U14706 ( .IN1(n11099), .IN2(g4961), .Q(n13980) );
  AND3X1 U14707 ( .IN1(n13981), .IN2(n9050), .IN3(n10280), .Q(n13979) );
  AND2X1 U14708 ( .IN1(n9435), .IN2(n9427), .Q(n10280) );
  OR2X1 U14709 ( .IN1(n13982), .IN2(g4961), .Q(n13981) );
  AND2X1 U14710 ( .IN1(n11091), .IN2(n13983), .Q(n13982) );
  OR4X1 U14711 ( .IN1(n13984), .IN2(n13985), .IN3(n13986), .IN4(n13987), .Q(
        n13983) );
  AND2X1 U14712 ( .IN1(n8746), .IN2(n11090), .Q(n13987) );
  AND2X1 U14713 ( .IN1(n10231), .IN2(g4049), .Q(n13986) );
  AND2X1 U14714 ( .IN1(n8416), .IN2(n13988), .Q(n13985) );
  AND2X1 U14715 ( .IN1(n11094), .IN2(g4045), .Q(n13984) );
  OR2X1 U14716 ( .IN1(n13989), .IN2(n13990), .Q(g28089) );
  AND2X1 U14717 ( .IN1(n11115), .IN2(g4950), .Q(n13990) );
  AND3X1 U14718 ( .IN1(n13991), .IN2(n9050), .IN3(n10288), .Q(n13989) );
  AND2X1 U14719 ( .IN1(n9434), .IN2(n9427), .Q(n10288) );
  OR2X1 U14720 ( .IN1(n13992), .IN2(g4950), .Q(n13991) );
  AND2X1 U14721 ( .IN1(n11107), .IN2(n13993), .Q(n13992) );
  OR4X1 U14722 ( .IN1(n13994), .IN2(n13995), .IN3(n13996), .IN4(n13997), .Q(
        n13993) );
  AND2X1 U14723 ( .IN1(n8755), .IN2(n11106), .Q(n13997) );
  AND2X1 U14724 ( .IN1(n10244), .IN2(g3698), .Q(n13996) );
  AND2X1 U14725 ( .IN1(n8414), .IN2(n13998), .Q(n13995) );
  AND2X1 U14726 ( .IN1(n11110), .IN2(g3694), .Q(n13994) );
  OR2X1 U14727 ( .IN1(n13999), .IN2(n14000), .Q(g28088) );
  AND2X1 U14728 ( .IN1(n11129), .IN2(g4939), .Q(n14000) );
  AND3X1 U14729 ( .IN1(n14001), .IN2(n9051), .IN3(n10295), .Q(n13999) );
  AND3X1 U14730 ( .IN1(n5360), .IN2(n5517), .IN3(n9427), .Q(n10295) );
  OR2X1 U14731 ( .IN1(n14002), .IN2(g4939), .Q(n14001) );
  AND2X1 U14732 ( .IN1(n11125), .IN2(n14003), .Q(n14002) );
  OR4X1 U14733 ( .IN1(n14004), .IN2(n14005), .IN3(n14006), .IN4(n14007), .Q(
        n14003) );
  AND2X1 U14734 ( .IN1(n8743), .IN2(n11124), .Q(n14007) );
  AND2X1 U14735 ( .IN1(n10236), .IN2(g3347), .Q(n14006) );
  AND2X1 U14736 ( .IN1(n8411), .IN2(n14008), .Q(n14005) );
  AND2X1 U14737 ( .IN1(n11122), .IN2(g3343), .Q(n14004) );
  OR2X1 U14738 ( .IN1(n14009), .IN2(n14010), .Q(g28087) );
  AND2X1 U14739 ( .IN1(n11010), .IN2(g4894), .Q(n14010) );
  AND2X1 U14740 ( .IN1(n9047), .IN2(n8809), .Q(n11010) );
  OR2X1 U14741 ( .IN1(n14011), .IN2(n5713), .Q(n8809) );
  AND2X1 U14742 ( .IN1(n14012), .IN2(n10963), .Q(n14011) );
  AND3X1 U14743 ( .IN1(g4888), .IN2(n5360), .IN3(n5517), .Q(n10963) );
  AND3X1 U14744 ( .IN1(n14013), .IN2(n9051), .IN3(n9914), .Q(n14009) );
  AND2X1 U14745 ( .IN1(n9437), .IN2(n9427), .Q(n9914) );
  AND2X1 U14746 ( .IN1(g4983), .IN2(n9438), .Q(n9427) );
  OR2X1 U14747 ( .IN1(n4689), .IN2(g4894), .Q(n14013) );
  OR2X1 U14748 ( .IN1(n14014), .IN2(n14015), .Q(g28086) );
  AND2X1 U14749 ( .IN1(n11027), .IN2(g4771), .Q(n14015) );
  AND2X1 U14750 ( .IN1(n9046), .IN2(n11023), .Q(n11027) );
  AND3X1 U14751 ( .IN1(n14016), .IN2(n9051), .IN3(n10316), .Q(n14014) );
  AND2X1 U14752 ( .IN1(n9405), .IN2(n9397), .Q(n10316) );
  OR2X1 U14753 ( .IN1(n14017), .IN2(g4771), .Q(n14016) );
  AND2X1 U14754 ( .IN1(n11019), .IN2(n14018), .Q(n14017) );
  OR4X1 U14755 ( .IN1(n14019), .IN2(n14020), .IN3(n14021), .IN4(n14022), .Q(
        n14018) );
  AND2X1 U14756 ( .IN1(n8412), .IN2(n13805), .Q(n14022) );
  AND2X1 U14757 ( .IN1(n5396), .IN2(n5592), .Q(n13805) );
  AND2X1 U14758 ( .IN1(n11022), .IN2(g6386), .Q(n14021) );
  AND2X1 U14759 ( .IN1(g6336), .IN2(n5396), .Q(n11022) );
  AND2X1 U14760 ( .IN1(n8744), .IN2(n11018), .Q(n14020) );
  AND2X1 U14761 ( .IN1(g6395), .IN2(n5592), .Q(n11018) );
  AND2X1 U14762 ( .IN1(n10232), .IN2(g6390), .Q(n14019) );
  AND2X1 U14763 ( .IN1(g6336), .IN2(g6395), .Q(n10232) );
  INVX0 U14764 ( .INP(n11023), .ZN(n11019) );
  OR2X1 U14765 ( .IN1(n14023), .IN2(n5656), .Q(n11023) );
  AND3X1 U14766 ( .IN1(n14024), .IN2(g4765), .IN3(n9407), .Q(n14023) );
  OR2X1 U14767 ( .IN1(n14025), .IN2(n14026), .Q(g28085) );
  AND2X1 U14768 ( .IN1(n11044), .IN2(g4760), .Q(n14026) );
  AND2X1 U14769 ( .IN1(n9046), .IN2(n11040), .Q(n11044) );
  AND3X1 U14770 ( .IN1(n14027), .IN2(n9052), .IN3(n10324), .Q(n14025) );
  AND2X1 U14771 ( .IN1(n9404), .IN2(n9397), .Q(n10324) );
  OR2X1 U14772 ( .IN1(n14028), .IN2(g4760), .Q(n14027) );
  AND2X1 U14773 ( .IN1(n11036), .IN2(n14029), .Q(n14028) );
  OR4X1 U14774 ( .IN1(n14030), .IN2(n14031), .IN3(n14032), .IN4(n14033), .Q(
        n14029) );
  AND2X1 U14775 ( .IN1(n8413), .IN2(n13848), .Q(n14033) );
  AND2X1 U14776 ( .IN1(n8835), .IN2(n5589), .Q(n13848) );
  AND2X1 U14777 ( .IN1(n11039), .IN2(g6040), .Q(n14032) );
  AND2X1 U14778 ( .IN1(n8835), .IN2(g5990), .Q(n11039) );
  AND2X1 U14779 ( .IN1(test_so50), .IN2(n10245), .Q(n14031) );
  AND2X1 U14780 ( .IN1(g5990), .IN2(test_so57), .Q(n10245) );
  AND2X1 U14781 ( .IN1(n11035), .IN2(n8844), .Q(n14030) );
  AND2X1 U14782 ( .IN1(test_so57), .IN2(n5589), .Q(n11035) );
  INVX0 U14783 ( .INP(n11040), .ZN(n11036) );
  OR2X1 U14784 ( .IN1(n14034), .IN2(n8553), .Q(n11040) );
  AND3X1 U14785 ( .IN1(n14024), .IN2(g4754), .IN3(n9405), .Q(n14034) );
  AND2X1 U14786 ( .IN1(g4709), .IN2(n5361), .Q(n9405) );
  OR2X1 U14787 ( .IN1(n14035), .IN2(n14036), .Q(g28084) );
  AND2X1 U14788 ( .IN1(n11060), .IN2(test_so18), .Q(n14036) );
  AND2X1 U14789 ( .IN1(n9046), .IN2(n11056), .Q(n11060) );
  AND3X1 U14790 ( .IN1(n14037), .IN2(n9052), .IN3(n10331), .Q(n14035) );
  AND3X1 U14791 ( .IN1(n5361), .IN2(n5518), .IN3(n9397), .Q(n10331) );
  OR2X1 U14792 ( .IN1(n14038), .IN2(test_so18), .Q(n14037) );
  AND2X1 U14793 ( .IN1(n11052), .IN2(n14039), .Q(n14038) );
  OR4X1 U14794 ( .IN1(n14040), .IN2(n14041), .IN3(n14042), .IN4(n14043), .Q(
        n14039) );
  AND2X1 U14795 ( .IN1(n8415), .IN2(n13894), .Q(n14043) );
  AND2X1 U14796 ( .IN1(n5397), .IN2(n5593), .Q(n13894) );
  AND2X1 U14797 ( .IN1(n11055), .IN2(g5694), .Q(n14042) );
  AND2X1 U14798 ( .IN1(g5644), .IN2(n5397), .Q(n11055) );
  AND2X1 U14799 ( .IN1(n8754), .IN2(n11051), .Q(n14041) );
  AND2X1 U14800 ( .IN1(g5703), .IN2(n5593), .Q(n11051) );
  AND2X1 U14801 ( .IN1(n10237), .IN2(g5698), .Q(n14040) );
  AND2X1 U14802 ( .IN1(g5644), .IN2(g5703), .Q(n10237) );
  INVX0 U14803 ( .INP(n11056), .ZN(n11052) );
  OR2X1 U14804 ( .IN1(n14044), .IN2(n5440), .Q(n11056) );
  AND3X1 U14805 ( .IN1(n14024), .IN2(g4743), .IN3(n9404), .Q(n14044) );
  AND2X1 U14806 ( .IN1(g4785), .IN2(n5518), .Q(n9404) );
  OR2X1 U14807 ( .IN1(n14045), .IN2(n14046), .Q(g28083) );
  AND2X1 U14808 ( .IN1(n11072), .IN2(g4704), .Q(n14046) );
  AND2X1 U14809 ( .IN1(n9045), .IN2(n8804), .Q(n11072) );
  OR2X1 U14810 ( .IN1(n14047), .IN2(n5712), .Q(n8804) );
  AND2X1 U14811 ( .IN1(n14024), .IN2(n10996), .Q(n14047) );
  AND3X1 U14812 ( .IN1(g4698), .IN2(n5361), .IN3(n5518), .Q(n10996) );
  AND3X1 U14813 ( .IN1(n10452), .IN2(n9408), .IN3(n5368), .Q(n14024) );
  AND3X1 U14814 ( .IN1(g4659), .IN2(g4669), .IN3(test_so19), .Q(n10452) );
  AND3X1 U14815 ( .IN1(n14048), .IN2(n9052), .IN3(n9917), .Q(n14045) );
  AND2X1 U14816 ( .IN1(n9407), .IN2(n9397), .Q(n9917) );
  AND2X1 U14817 ( .IN1(g4793), .IN2(n9408), .Q(n9397) );
  AND2X1 U14818 ( .IN1(n8836), .IN2(g4776), .Q(n9408) );
  AND2X1 U14819 ( .IN1(g4709), .IN2(g4785), .Q(n9407) );
  OR2X1 U14820 ( .IN1(n4708), .IN2(g4704), .Q(n14048) );
  OR2X1 U14821 ( .IN1(n14049), .IN2(n14050), .Q(g28082) );
  AND3X1 U14822 ( .IN1(n9795), .IN2(n9052), .IN3(n5752), .Q(n14050) );
  AND2X1 U14823 ( .IN1(n14051), .IN2(g4521), .Q(n14049) );
  OR2X1 U14824 ( .IN1(n9134), .IN2(n14052), .Q(n14051) );
  AND2X1 U14825 ( .IN1(n14053), .IN2(n14054), .Q(n14052) );
  OR2X1 U14826 ( .IN1(n10459), .IN2(g4527), .Q(n14054) );
  OR2X1 U14827 ( .IN1(n8514), .IN2(n14055), .Q(n14053) );
  OR3X1 U14828 ( .IN1(n14056), .IN2(n14057), .IN3(n14058), .Q(g28074) );
  AND2X1 U14829 ( .IN1(n9150), .IN2(g4119), .Q(n14058) );
  AND2X1 U14830 ( .IN1(n4714), .IN2(n4721), .Q(n14057) );
  AND3X1 U14831 ( .IN1(n9054), .IN2(g4122), .IN3(n14059), .Q(n14056) );
  INVX0 U14832 ( .INP(n4714), .ZN(n14059) );
  OR3X1 U14833 ( .IN1(n14060), .IN2(n14061), .IN3(n14062), .Q(g28073) );
  AND2X1 U14834 ( .IN1(n14063), .IN2(n4721), .Q(n14062) );
  AND2X1 U14835 ( .IN1(n9150), .IN2(g4116), .Q(n14061) );
  AND3X1 U14836 ( .IN1(n14064), .IN2(g4119), .IN3(n9064), .Q(n14060) );
  INVX0 U14837 ( .INP(n14063), .ZN(n14064) );
  AND2X1 U14838 ( .IN1(g4057), .IN2(n14065), .Q(n14063) );
  OR3X1 U14839 ( .IN1(n14066), .IN2(n14067), .IN3(n14068), .Q(g28072) );
  AND2X1 U14840 ( .IN1(n14069), .IN2(n4721), .Q(n14068) );
  AND2X1 U14841 ( .IN1(n9150), .IN2(g4112), .Q(n14067) );
  AND3X1 U14842 ( .IN1(n14070), .IN2(g4116), .IN3(n9064), .Q(n14066) );
  INVX0 U14843 ( .INP(n14069), .ZN(n14070) );
  AND3X1 U14844 ( .IN1(g4064), .IN2(n5711), .IN3(n4722), .Q(n14069) );
  OR2X1 U14845 ( .IN1(n14071), .IN2(n14072), .Q(g28071) );
  INVX0 U14846 ( .INP(n14073), .ZN(n14072) );
  OR2X1 U14847 ( .IN1(n14074), .IN2(n8515), .Q(n14073) );
  AND2X1 U14848 ( .IN1(n14074), .IN2(g4112), .Q(n14071) );
  AND2X1 U14849 ( .IN1(n9043), .IN2(n14075), .Q(n14074) );
  INVX0 U14850 ( .INP(n14076), .ZN(n14075) );
  AND2X1 U14851 ( .IN1(n14065), .IN2(n5711), .Q(n14076) );
  AND2X1 U14852 ( .IN1(n5416), .IN2(n4722), .Q(n14065) );
  AND4X1 U14853 ( .IN1(n8825), .IN2(n10218), .IN3(n5350), .IN4(n14077), .Q(
        n4722) );
  AND2X1 U14854 ( .IN1(n5612), .IN2(n8677), .Q(n14077) );
  INVX0 U14855 ( .INP(n12162), .ZN(n10218) );
  OR2X1 U14856 ( .IN1(g4087), .IN2(g4093), .Q(n12162) );
  OR4X1 U14857 ( .IN1(n8811), .IN2(n14078), .IN3(n14079), .IN4(n14080), .Q(
        g28070) );
  AND2X1 U14858 ( .IN1(n9150), .IN2(g4082), .Q(n14080) );
  AND3X1 U14859 ( .IN1(test_so11), .IN2(n14081), .IN3(n9065), .Q(n14079) );
  AND2X1 U14860 ( .IN1(n12528), .IN2(n8825), .Q(n14078) );
  OR3X1 U14861 ( .IN1(n14082), .IN2(n14083), .IN3(n14084), .Q(g28069) );
  AND2X1 U14862 ( .IN1(n11099), .IN2(g4035), .Q(n14084) );
  AND2X1 U14863 ( .IN1(n9042), .IN2(n11095), .Q(n11099) );
  AND3X1 U14864 ( .IN1(n11091), .IN2(n13363), .IN3(n9065), .Q(n14083) );
  OR2X1 U14865 ( .IN1(n14085), .IN2(n14086), .Q(n13363) );
  AND2X1 U14866 ( .IN1(n14087), .IN2(g4040), .Q(n14086) );
  OR4X1 U14867 ( .IN1(n14088), .IN2(n14089), .IN3(n14090), .IN4(n14091), .Q(
        n14087) );
  OR3X1 U14868 ( .IN1(n14092), .IN2(n14093), .IN3(n14094), .Q(n14091) );
  AND2X1 U14869 ( .IN1(n10231), .IN2(n14095), .Q(n14094) );
  OR2X1 U14870 ( .IN1(n14096), .IN2(n14097), .Q(n14095) );
  AND2X1 U14871 ( .IN1(test_so65), .IN2(g16748), .Q(n14097) );
  AND2X1 U14872 ( .IN1(g3965), .IN2(g16693), .Q(n14096) );
  AND3X1 U14873 ( .IN1(g3917), .IN2(g16955), .IN3(n11090), .Q(n14093) );
  AND3X1 U14874 ( .IN1(g13906), .IN2(g3933), .IN3(n11094), .Q(n14092) );
  AND2X1 U14875 ( .IN1(n13988), .IN2(n14098), .Q(n14090) );
  OR2X1 U14876 ( .IN1(n14099), .IN2(n14100), .Q(n14098) );
  AND2X1 U14877 ( .IN1(test_so24), .IN2(g14518), .Q(n14100) );
  AND2X1 U14878 ( .IN1(g3897), .IN2(g4031), .Q(n14099) );
  AND2X1 U14879 ( .IN1(n14101), .IN2(g11418), .Q(n14089) );
  OR2X1 U14880 ( .IN1(n14102), .IN2(n14103), .Q(n14101) );
  AND2X1 U14881 ( .IN1(n11090), .IN2(g3893), .Q(n14102) );
  AND2X1 U14882 ( .IN1(n5435), .IN2(n14104), .Q(n14088) );
  AND2X1 U14883 ( .IN1(n5530), .IN2(n14105), .Q(n14085) );
  OR4X1 U14884 ( .IN1(n14106), .IN2(n14107), .IN3(n14108), .IN4(n14109), .Q(
        n14105) );
  OR3X1 U14885 ( .IN1(n14110), .IN2(n14111), .IN3(n14112), .Q(n14109) );
  AND2X1 U14886 ( .IN1(n11094), .IN2(n14113), .Q(n14112) );
  OR2X1 U14887 ( .IN1(n14114), .IN2(n14115), .Q(n14113) );
  AND2X1 U14888 ( .IN1(g3901), .IN2(g14518), .Q(n14115) );
  AND2X1 U14889 ( .IN1(g4031), .IN2(g3913), .Q(n14114) );
  AND3X1 U14890 ( .IN1(g13906), .IN2(g3941), .IN3(n13988), .Q(n14111) );
  AND3X1 U14891 ( .IN1(g16955), .IN2(g3925), .IN3(n10231), .Q(n14110) );
  AND2X1 U14892 ( .IN1(n11090), .IN2(n14116), .Q(n14108) );
  OR2X1 U14893 ( .IN1(n14117), .IN2(n14118), .Q(n14116) );
  AND2X1 U14894 ( .IN1(g3905), .IN2(g16693), .Q(n14118) );
  AND2X1 U14895 ( .IN1(g16748), .IN2(g3957), .Q(n14117) );
  AND2X1 U14896 ( .IN1(n14119), .IN2(g11418), .Q(n14107) );
  OR2X1 U14897 ( .IN1(n14120), .IN2(n14104), .Q(n14119) );
  OR3X1 U14898 ( .IN1(n14121), .IN2(n14122), .IN3(n14123), .Q(n14104) );
  AND3X1 U14899 ( .IN1(g13966), .IN2(g3929), .IN3(n13988), .Q(n14123) );
  AND3X1 U14900 ( .IN1(g3945), .IN2(g16775), .IN3(n11090), .Q(n14122) );
  AND2X1 U14901 ( .IN1(g4054), .IN2(n5594), .Q(n11090) );
  AND3X1 U14902 ( .IN1(g3961), .IN2(g16659), .IN3(n11094), .Q(n14121) );
  AND2X1 U14903 ( .IN1(n10231), .IN2(g3909), .Q(n14120) );
  AND2X1 U14904 ( .IN1(n5435), .IN2(n14103), .Q(n14106) );
  OR3X1 U14905 ( .IN1(n14124), .IN2(n14125), .IN3(n14126), .Q(n14103) );
  AND3X1 U14906 ( .IN1(g3953), .IN2(g16659), .IN3(n13988), .Q(n14126) );
  AND2X1 U14907 ( .IN1(n5395), .IN2(n5594), .Q(n13988) );
  AND3X1 U14908 ( .IN1(g13966), .IN2(g3921), .IN3(n11094), .Q(n14125) );
  AND2X1 U14909 ( .IN1(g3990), .IN2(n5395), .Q(n11094) );
  AND3X1 U14910 ( .IN1(g3937), .IN2(g16775), .IN3(n10231), .Q(n14124) );
  AND2X1 U14911 ( .IN1(g3990), .IN2(g4054), .Q(n10231) );
  INVX0 U14912 ( .INP(n11095), .ZN(n11091) );
  OR2X1 U14913 ( .IN1(n14127), .IN2(n5283), .Q(n11095) );
  AND3X1 U14914 ( .IN1(n14012), .IN2(g4955), .IN3(n9437), .Q(n14127) );
  AND2X1 U14915 ( .IN1(g4899), .IN2(g4975), .Q(n9437) );
  AND2X1 U14916 ( .IN1(n9150), .IN2(g3965), .Q(n14082) );
  OR3X1 U14917 ( .IN1(n14128), .IN2(n14129), .IN3(n14130), .Q(g28066) );
  AND2X1 U14918 ( .IN1(n11115), .IN2(g3684), .Q(n14130) );
  AND2X1 U14919 ( .IN1(n9042), .IN2(n11111), .Q(n11115) );
  AND3X1 U14920 ( .IN1(n11107), .IN2(n13392), .IN3(n9066), .Q(n14129) );
  OR2X1 U14921 ( .IN1(n14131), .IN2(n14132), .Q(n13392) );
  AND2X1 U14922 ( .IN1(n14133), .IN2(g3689), .Q(n14132) );
  OR4X1 U14923 ( .IN1(n14134), .IN2(n14135), .IN3(n14136), .IN4(n14137), .Q(
        n14133) );
  OR3X1 U14924 ( .IN1(n14138), .IN2(n14139), .IN3(n14140), .Q(n14137) );
  AND2X1 U14925 ( .IN1(n10244), .IN2(n14141), .Q(n14140) );
  OR2X1 U14926 ( .IN1(n14142), .IN2(n14143), .Q(n14141) );
  AND2X1 U14927 ( .IN1(g3598), .IN2(g16722), .Q(n14143) );
  AND2X1 U14928 ( .IN1(g3614), .IN2(g16656), .Q(n14142) );
  AND3X1 U14929 ( .IN1(g3566), .IN2(g16924), .IN3(n11106), .Q(n14139) );
  AND3X1 U14930 ( .IN1(n11110), .IN2(g3582), .IN3(test_so26), .Q(n14138) );
  AND2X1 U14931 ( .IN1(n13998), .IN2(n14144), .Q(n14136) );
  OR2X1 U14932 ( .IN1(n14145), .IN2(n14146), .Q(n14144) );
  AND2X1 U14933 ( .IN1(g3538), .IN2(g14451), .Q(n14146) );
  AND2X1 U14934 ( .IN1(g3546), .IN2(g3680), .Q(n14145) );
  AND2X1 U14935 ( .IN1(n14147), .IN2(g11388), .Q(n14135) );
  OR2X1 U14936 ( .IN1(n14148), .IN2(n14149), .Q(n14147) );
  AND2X1 U14937 ( .IN1(n11106), .IN2(g3542), .Q(n14148) );
  AND2X1 U14938 ( .IN1(n5433), .IN2(n14150), .Q(n14134) );
  AND2X1 U14939 ( .IN1(n5532), .IN2(n14151), .Q(n14131) );
  OR4X1 U14940 ( .IN1(n14152), .IN2(n14153), .IN3(n14154), .IN4(n14155), .Q(
        n14151) );
  OR3X1 U14941 ( .IN1(n14156), .IN2(n14157), .IN3(n14158), .Q(n14155) );
  AND2X1 U14942 ( .IN1(n11110), .IN2(n14159), .Q(n14158) );
  OR2X1 U14943 ( .IN1(n14160), .IN2(n14161), .Q(n14159) );
  AND2X1 U14944 ( .IN1(g3550), .IN2(g14451), .Q(n14161) );
  AND2X1 U14945 ( .IN1(g3680), .IN2(g3562), .Q(n14160) );
  AND3X1 U14946 ( .IN1(test_so26), .IN2(g3590), .IN3(n13998), .Q(n14157) );
  AND3X1 U14947 ( .IN1(g16924), .IN2(g3574), .IN3(n10244), .Q(n14156) );
  AND2X1 U14948 ( .IN1(n11106), .IN2(n14162), .Q(n14154) );
  OR2X1 U14949 ( .IN1(n14163), .IN2(n14164), .Q(n14162) );
  AND2X1 U14950 ( .IN1(g3554), .IN2(g16656), .Q(n14164) );
  AND2X1 U14951 ( .IN1(g16722), .IN2(g3606), .Q(n14163) );
  AND2X1 U14952 ( .IN1(n14165), .IN2(g11388), .Q(n14153) );
  OR2X1 U14953 ( .IN1(n14166), .IN2(n14150), .Q(n14165) );
  OR3X1 U14954 ( .IN1(n14167), .IN2(n14168), .IN3(n14169), .Q(n14150) );
  AND3X1 U14955 ( .IN1(g13926), .IN2(g3578), .IN3(n13998), .Q(n14169) );
  AND3X1 U14956 ( .IN1(g3594), .IN2(g16744), .IN3(n11106), .Q(n14168) );
  AND2X1 U14957 ( .IN1(g3703), .IN2(n5591), .Q(n11106) );
  AND3X1 U14958 ( .IN1(g3610), .IN2(g16627), .IN3(n11110), .Q(n14167) );
  AND2X1 U14959 ( .IN1(n10244), .IN2(g3558), .Q(n14166) );
  AND2X1 U14960 ( .IN1(n5433), .IN2(n14149), .Q(n14152) );
  OR3X1 U14961 ( .IN1(n14170), .IN2(n14171), .IN3(n14172), .Q(n14149) );
  AND3X1 U14962 ( .IN1(test_so43), .IN2(g16627), .IN3(n13998), .Q(n14172) );
  AND2X1 U14963 ( .IN1(n5399), .IN2(n5591), .Q(n13998) );
  AND3X1 U14964 ( .IN1(g13926), .IN2(g3570), .IN3(n11110), .Q(n14171) );
  AND2X1 U14965 ( .IN1(g3639), .IN2(n5399), .Q(n11110) );
  AND3X1 U14966 ( .IN1(g3586), .IN2(g16744), .IN3(n10244), .Q(n14170) );
  AND2X1 U14967 ( .IN1(g3639), .IN2(g3703), .Q(n10244) );
  INVX0 U14968 ( .INP(n11111), .ZN(n11107) );
  OR2X1 U14969 ( .IN1(n14173), .IN2(n5443), .Q(n11111) );
  AND3X1 U14970 ( .IN1(n14012), .IN2(g4944), .IN3(n9435), .Q(n14173) );
  AND2X1 U14971 ( .IN1(g4899), .IN2(n5360), .Q(n9435) );
  AND2X1 U14972 ( .IN1(n9150), .IN2(g3614), .Q(n14128) );
  OR3X1 U14973 ( .IN1(n14174), .IN2(n14175), .IN3(n14176), .Q(g28063) );
  AND2X1 U14974 ( .IN1(n11129), .IN2(g3333), .Q(n14176) );
  AND2X1 U14975 ( .IN1(n9042), .IN2(n11123), .Q(n11129) );
  AND3X1 U14976 ( .IN1(n11125), .IN2(n13425), .IN3(n9066), .Q(n14175) );
  OR2X1 U14977 ( .IN1(n14177), .IN2(n14178), .Q(n13425) );
  AND2X1 U14978 ( .IN1(n14179), .IN2(g3338), .Q(n14178) );
  OR4X1 U14979 ( .IN1(n14180), .IN2(n14181), .IN3(n14182), .IN4(n14183), .Q(
        n14179) );
  OR3X1 U14980 ( .IN1(n14184), .IN2(n14185), .IN3(n14186), .Q(n14183) );
  AND2X1 U14981 ( .IN1(n10236), .IN2(n14187), .Q(n14186) );
  OR2X1 U14982 ( .IN1(n14188), .IN2(n14189), .Q(n14187) );
  AND2X1 U14983 ( .IN1(g3247), .IN2(g16686), .Q(n14189) );
  AND2X1 U14984 ( .IN1(g3263), .IN2(g16624), .Q(n14188) );
  AND3X1 U14985 ( .IN1(g3215), .IN2(g16874), .IN3(n11124), .Q(n14185) );
  AND3X1 U14986 ( .IN1(g13865), .IN2(g3231), .IN3(n11122), .Q(n14184) );
  AND2X1 U14987 ( .IN1(n14008), .IN2(n14190), .Q(n14182) );
  OR2X1 U14988 ( .IN1(n14191), .IN2(n14192), .Q(n14190) );
  AND2X1 U14989 ( .IN1(test_so91), .IN2(test_so88), .Q(n14192) );
  AND2X1 U14990 ( .IN1(g3187), .IN2(g14421), .Q(n14191) );
  AND2X1 U14991 ( .IN1(n14193), .IN2(g11349), .Q(n14181) );
  OR2X1 U14992 ( .IN1(n14194), .IN2(n14195), .Q(n14193) );
  AND2X1 U14993 ( .IN1(n11124), .IN2(g3191), .Q(n14194) );
  AND2X1 U14994 ( .IN1(n5436), .IN2(n14196), .Q(n14180) );
  AND2X1 U14995 ( .IN1(n5527), .IN2(n14197), .Q(n14177) );
  OR4X1 U14996 ( .IN1(n14198), .IN2(n14199), .IN3(n14200), .IN4(n14201), .Q(
        n14197) );
  OR3X1 U14997 ( .IN1(n14202), .IN2(n14203), .IN3(n14204), .Q(n14201) );
  AND2X1 U14998 ( .IN1(n11122), .IN2(n14205), .Q(n14204) );
  OR2X1 U14999 ( .IN1(n14206), .IN2(n14207), .Q(n14205) );
  AND2X1 U15000 ( .IN1(g3199), .IN2(g14421), .Q(n14207) );
  AND2X1 U15001 ( .IN1(test_so91), .IN2(g3211), .Q(n14206) );
  AND3X1 U15002 ( .IN1(g13865), .IN2(g3239), .IN3(n14008), .Q(n14203) );
  AND3X1 U15003 ( .IN1(g16874), .IN2(g3223), .IN3(n10236), .Q(n14202) );
  AND2X1 U15004 ( .IN1(n11124), .IN2(n14208), .Q(n14200) );
  OR2X1 U15005 ( .IN1(n14209), .IN2(n14210), .Q(n14208) );
  AND2X1 U15006 ( .IN1(g3203), .IN2(g16624), .Q(n14210) );
  AND2X1 U15007 ( .IN1(g16686), .IN2(g3255), .Q(n14209) );
  AND2X1 U15008 ( .IN1(n14211), .IN2(g11349), .Q(n14199) );
  OR2X1 U15009 ( .IN1(n14212), .IN2(n14196), .Q(n14211) );
  OR3X1 U15010 ( .IN1(n14213), .IN2(n14214), .IN3(n14215), .Q(n14196) );
  AND3X1 U15011 ( .IN1(g13895), .IN2(g3227), .IN3(n14008), .Q(n14215) );
  AND3X1 U15012 ( .IN1(g3243), .IN2(g16718), .IN3(n11124), .Q(n14214) );
  AND2X1 U15013 ( .IN1(g3352), .IN2(n5400), .Q(n11124) );
  AND3X1 U15014 ( .IN1(test_so84), .IN2(g16603), .IN3(n11122), .Q(n14213) );
  AND2X1 U15015 ( .IN1(n10236), .IN2(g3207), .Q(n14212) );
  AND2X1 U15016 ( .IN1(n5436), .IN2(n14195), .Q(n14198) );
  OR3X1 U15017 ( .IN1(n14216), .IN2(n14217), .IN3(n14218), .Q(n14195) );
  AND3X1 U15018 ( .IN1(g3251), .IN2(g16603), .IN3(n14008), .Q(n14218) );
  AND2X1 U15019 ( .IN1(n5604), .IN2(n5400), .Q(n14008) );
  AND3X1 U15020 ( .IN1(g13895), .IN2(g3219), .IN3(n11122), .Q(n14217) );
  AND2X1 U15021 ( .IN1(g3288), .IN2(n5604), .Q(n11122) );
  AND3X1 U15022 ( .IN1(g3235), .IN2(g16718), .IN3(n10236), .Q(n14216) );
  AND2X1 U15023 ( .IN1(g3352), .IN2(g3288), .Q(n10236) );
  INVX0 U15024 ( .INP(n11123), .ZN(n11125) );
  OR2X1 U15025 ( .IN1(n14219), .IN2(n5318), .Q(n11123) );
  AND3X1 U15026 ( .IN1(n14012), .IN2(g4933), .IN3(n9434), .Q(n14219) );
  AND2X1 U15027 ( .IN1(g4975), .IN2(n5517), .Q(n9434) );
  AND3X1 U15028 ( .IN1(n10427), .IN2(n9438), .IN3(n5367), .Q(n14012) );
  AND2X1 U15029 ( .IN1(n8837), .IN2(g4966), .Q(n9438) );
  AND3X1 U15030 ( .IN1(g4849), .IN2(g4843), .IN3(g4859), .Q(n10427) );
  AND2X1 U15031 ( .IN1(n9150), .IN2(g3263), .Q(n14174) );
  OR3X1 U15032 ( .IN1(n2787), .IN2(n14220), .IN3(n14221), .Q(g28060) );
  AND2X1 U15033 ( .IN1(n14222), .IN2(g2724), .Q(n14221) );
  OR2X1 U15034 ( .IN1(n9134), .IN2(n14223), .Q(n14222) );
  AND2X1 U15035 ( .IN1(n14224), .IN2(n13431), .Q(n14223) );
  AND3X1 U15036 ( .IN1(n9055), .IN2(g2729), .IN3(n13431), .Q(n14220) );
  OR2X1 U15037 ( .IN1(n12798), .IN2(n10178), .Q(n13431) );
  OR2X1 U15038 ( .IN1(n5301), .IN2(n8676), .Q(n10178) );
  OR3X1 U15039 ( .IN1(n14225), .IN2(n14226), .IN3(n14227), .Q(g28059) );
  AND2X1 U15040 ( .IN1(n9150), .IN2(g1351), .Q(n14227) );
  AND2X1 U15041 ( .IN1(n4798), .IN2(n13089), .Q(n14226) );
  AND3X1 U15042 ( .IN1(n11902), .IN2(n8799), .IN3(n14228), .Q(n14225) );
  AND2X1 U15043 ( .IN1(n9042), .IN2(n11477), .Q(n11902) );
  AND4X1 U15044 ( .IN1(n14229), .IN2(n5466), .IN3(n14230), .IN4(n14231), .Q(
        n11477) );
  INVX0 U15045 ( .INP(n14232), .ZN(n14231) );
  AND3X1 U15046 ( .IN1(n14233), .IN2(g1351), .IN3(n14234), .Q(n14232) );
  OR2X1 U15047 ( .IN1(n14234), .IN2(g1351), .Q(n14230) );
  OR3X1 U15048 ( .IN1(n14235), .IN2(n14236), .IN3(n14237), .Q(g28058) );
  AND2X1 U15049 ( .IN1(test_so77), .IN2(n9138), .Q(n14237) );
  AND2X1 U15050 ( .IN1(n4490), .IN2(n5554), .Q(n14236) );
  AND3X1 U15051 ( .IN1(n11485), .IN2(n14238), .IN3(g1252), .Q(n14235) );
  INVX0 U15052 ( .INP(n4490), .ZN(n14238) );
  OR3X1 U15053 ( .IN1(n14239), .IN2(n14240), .IN3(n14241), .Q(g28057) );
  AND2X1 U15054 ( .IN1(n9150), .IN2(g1008), .Q(n14241) );
  AND2X1 U15055 ( .IN1(n4805), .IN2(n13124), .Q(n14240) );
  AND3X1 U15056 ( .IN1(n11913), .IN2(n8796), .IN3(n14242), .Q(n14239) );
  AND2X1 U15057 ( .IN1(n9042), .IN2(n11492), .Q(n11913) );
  INVX0 U15058 ( .INP(n14243), .ZN(n11492) );
  OR4X1 U15059 ( .IN1(test_so20), .IN2(n14244), .IN3(n14245), .IN4(n14246), 
        .Q(n14243) );
  AND2X1 U15060 ( .IN1(n14247), .IN2(n5321), .Q(n14246) );
  AND3X1 U15061 ( .IN1(n14248), .IN2(n14249), .IN3(g1008), .Q(n14245) );
  INVX0 U15062 ( .INP(n14250), .ZN(n14244) );
  OR3X1 U15063 ( .IN1(n14251), .IN2(n14252), .IN3(n14253), .Q(g28056) );
  AND2X1 U15064 ( .IN1(n9150), .IN2(g936), .Q(n14253) );
  AND2X1 U15065 ( .IN1(n4514), .IN2(n5555), .Q(n14252) );
  AND3X1 U15066 ( .IN1(n11500), .IN2(n14254), .IN3(g907), .Q(n14251) );
  INVX0 U15067 ( .INP(n4514), .ZN(n14254) );
  OR3X1 U15068 ( .IN1(n14255), .IN2(n14256), .IN3(n14257), .Q(g28055) );
  AND2X1 U15069 ( .IN1(n9150), .IN2(g822), .Q(n14257) );
  AND3X1 U15070 ( .IN1(n4519), .IN2(n13689), .IN3(n5728), .Q(n14256) );
  AND3X1 U15071 ( .IN1(n4518), .IN2(n14258), .IN3(g827), .Q(n14255) );
  INVX0 U15072 ( .INP(n4519), .ZN(n14258) );
  OR2X1 U15073 ( .IN1(n14259), .IN2(n14260), .Q(g28054) );
  AND2X1 U15074 ( .IN1(n14261), .IN2(g661), .Q(n14260) );
  AND2X1 U15075 ( .IN1(n14262), .IN2(g728), .Q(n14259) );
  OR3X1 U15076 ( .IN1(n14263), .IN2(n14264), .IN3(n14265), .Q(g28053) );
  AND2X1 U15077 ( .IN1(n9150), .IN2(g681), .Q(n14265) );
  AND2X1 U15078 ( .IN1(n13727), .IN2(test_so87), .Q(n14264) );
  OR2X1 U15079 ( .IN1(n14266), .IN2(n14267), .Q(g28052) );
  AND2X1 U15080 ( .IN1(n14261), .IN2(g718), .Q(n14267) );
  AND2X1 U15081 ( .IN1(n14262), .IN2(g661), .Q(n14266) );
  OR2X1 U15082 ( .IN1(n14268), .IN2(n14269), .Q(g28051) );
  AND2X1 U15083 ( .IN1(n14261), .IN2(g655), .Q(n14269) );
  AND2X1 U15084 ( .IN1(n14262), .IN2(g718), .Q(n14268) );
  OR2X1 U15085 ( .IN1(n14270), .IN2(n14271), .Q(g28050) );
  AND2X1 U15086 ( .IN1(n14261), .IN2(g650), .Q(n14271) );
  AND2X1 U15087 ( .IN1(n14262), .IN2(g655), .Q(n14270) );
  OR3X1 U15088 ( .IN1(n14272), .IN2(n14273), .IN3(n14274), .Q(g28049) );
  AND2X1 U15089 ( .IN1(test_so87), .IN2(n9138), .Q(n14274) );
  AND2X1 U15090 ( .IN1(n14262), .IN2(g650), .Q(n14273) );
  AND2X1 U15091 ( .IN1(n14263), .IN2(g681), .Q(n14272) );
  OR3X1 U15092 ( .IN1(n14275), .IN2(n14276), .IN3(n14277), .Q(g28048) );
  AND2X1 U15093 ( .IN1(n14278), .IN2(g691), .Q(n14277) );
  OR2X1 U15094 ( .IN1(n14279), .IN2(n14280), .Q(n14278) );
  AND3X1 U15095 ( .IN1(g703), .IN2(n8852), .IN3(n9066), .Q(n14279) );
  AND3X1 U15096 ( .IN1(n14281), .IN2(n14282), .IN3(n9066), .Q(n14276) );
  INVX0 U15097 ( .INP(n939), .ZN(n14282) );
  OR4X1 U15098 ( .IN1(n14283), .IN2(g691), .IN3(n5821), .IN4(n13710), .Q(n939)
         );
  OR4X1 U15099 ( .IN1(n14284), .IN2(n14285), .IN3(n8845), .IN4(n14286), .Q(
        n13710) );
  OR2X1 U15100 ( .IN1(g645), .IN2(g650), .Q(n14286) );
  AND2X1 U15101 ( .IN1(n8381), .IN2(g728), .Q(n14285) );
  AND2X1 U15102 ( .IN1(n8382), .IN2(g661), .Q(n14284) );
  INVX0 U15103 ( .INP(n5112), .ZN(n14283) );
  AND2X1 U15104 ( .IN1(n9150), .IN2(g29212), .Q(n14275) );
  OR2X1 U15105 ( .IN1(n14287), .IN2(n14288), .Q(g28047) );
  AND2X1 U15106 ( .IN1(n14261), .IN2(g645), .Q(n14288) );
  INVX0 U15107 ( .INP(n14262), .ZN(n14261) );
  AND2X1 U15108 ( .IN1(n14262), .IN2(g681), .Q(n14287) );
  OR2X1 U15109 ( .IN1(n14289), .IN2(n14290), .Q(g28046) );
  AND2X1 U15110 ( .IN1(n14262), .IN2(g645), .Q(n14290) );
  AND2X1 U15111 ( .IN1(n9042), .IN2(n14291), .Q(n14262) );
  AND2X1 U15112 ( .IN1(n14263), .IN2(g446), .Q(n14289) );
  AND2X1 U15113 ( .IN1(n9041), .IN2(n14292), .Q(n14263) );
  INVX0 U15114 ( .INP(n14291), .ZN(n14292) );
  OR3X1 U15115 ( .IN1(n14293), .IN2(n14294), .IN3(n14295), .Q(n14291) );
  AND2X1 U15116 ( .IN1(n5520), .IN2(n14296), .Q(n14294) );
  OR3X1 U15117 ( .IN1(n5358), .IN2(g411), .IN3(g424), .Q(n14296) );
  AND2X1 U15118 ( .IN1(n14297), .IN2(g691), .Q(n14293) );
  OR3X1 U15119 ( .IN1(n14298), .IN2(n14299), .IN3(n14300), .Q(g28045) );
  AND2X1 U15120 ( .IN1(n9149), .IN2(g568), .Q(n14300) );
  AND2X1 U15121 ( .IN1(n4537), .IN2(n5337), .Q(n14299) );
  AND3X1 U15122 ( .IN1(n2421), .IN2(n14301), .IN3(g572), .Q(n14298) );
  INVX0 U15123 ( .INP(n4537), .ZN(n14301) );
  OR3X1 U15124 ( .IN1(n14302), .IN2(n14303), .IN3(n13718), .Q(g28044) );
  AND3X1 U15125 ( .IN1(n14304), .IN2(n13722), .IN3(n9065), .Q(n14303) );
  OR3X1 U15126 ( .IN1(n5820), .IN2(n14305), .IN3(n14306), .Q(n13722) );
  AND2X1 U15127 ( .IN1(n5327), .IN2(n14307), .Q(n14305) );
  OR2X1 U15128 ( .IN1(n14308), .IN2(g482), .Q(n14304) );
  AND2X1 U15129 ( .IN1(n14309), .IN2(g528), .Q(n14308) );
  AND2X1 U15130 ( .IN1(n9149), .IN2(g528), .Q(n14302) );
  OR2X1 U15131 ( .IN1(n14310), .IN2(n14311), .Q(g28043) );
  AND2X1 U15132 ( .IN1(n9149), .IN2(g278), .Q(n14311) );
  AND2X1 U15133 ( .IN1(n8803), .IN2(n8847), .Q(n14310) );
  AND2X1 U15134 ( .IN1(n9041), .IN2(n11937), .Q(n8803) );
  AND4X1 U15135 ( .IN1(g691), .IN2(n13145), .IN3(n14312), .IN4(n14313), .Q(
        n11937) );
  OR2X1 U15136 ( .IN1(n14314), .IN2(n5627), .Q(n14312) );
  INVX0 U15137 ( .INP(n14315), .ZN(n14314) );
  OR4X1 U15138 ( .IN1(n14316), .IN2(n14317), .IN3(n14318), .IN4(n14319), .Q(
        n13145) );
  AND3X1 U15139 ( .IN1(n8784), .IN2(n8783), .IN3(n8785), .Q(n14319) );
  AND3X1 U15140 ( .IN1(g753), .IN2(g655), .IN3(g718), .Q(n14318) );
  AND2X1 U15141 ( .IN1(g807), .IN2(g554), .Q(n14316) );
  OR3X1 U15142 ( .IN1(n9121), .IN2(g1306), .IN3(g962), .Q(g28042) );
  OR3X1 U15143 ( .IN1(n9121), .IN2(n11471), .IN3(n11298), .Q(g28041) );
  INVX0 U15144 ( .INP(n9854), .ZN(n11298) );
  OR2X1 U15145 ( .IN1(n8279), .IN2(n14320), .Q(n9854) );
  AND2X1 U15146 ( .IN1(g1193), .IN2(n4837), .Q(n11471) );
  OR2X1 U15147 ( .IN1(n14321), .IN2(n14322), .Q(g28030) );
  AND3X1 U15148 ( .IN1(n9881), .IN2(n9880), .IN3(n9882), .Q(n14322) );
  AND3X1 U15149 ( .IN1(n5861), .IN2(n14323), .IN3(n5882), .Q(n14321) );
  OR2X1 U15150 ( .IN1(n14324), .IN2(n14325), .Q(n14323) );
  AND2X1 U15151 ( .IN1(n9882), .IN2(n9881), .Q(n14325) );
  AND2X1 U15152 ( .IN1(n14326), .IN2(n9880), .Q(n14324) );
  OR2X1 U15153 ( .IN1(n9135), .IN2(n14327), .Q(n9880) );
  AND2X1 U15154 ( .IN1(n5889), .IN2(n5868), .Q(n14327) );
  OR2X1 U15155 ( .IN1(n14328), .IN2(n14329), .Q(n14326) );
  AND2X1 U15156 ( .IN1(n9882), .IN2(n14330), .Q(n14329) );
  OR2X1 U15157 ( .IN1(n14331), .IN2(n14332), .Q(n14330) );
  AND4X1 U15158 ( .IN1(n5885), .IN2(n5869), .IN3(n14333), .IN4(n14334), .Q(
        n14331) );
  OR2X1 U15159 ( .IN1(n14335), .IN2(n14336), .Q(n14334) );
  OR2X1 U15160 ( .IN1(n14337), .IN2(n14338), .Q(n14333) );
  AND2X1 U15161 ( .IN1(n14339), .IN2(n14340), .Q(n9882) );
  AND2X1 U15162 ( .IN1(n9881), .IN2(n14341), .Q(n14328) );
  OR2X1 U15163 ( .IN1(n14340), .IN2(n14339), .Q(n14341) );
  OR2X1 U15164 ( .IN1(n9135), .IN2(n14342), .Q(n14339) );
  AND2X1 U15165 ( .IN1(n5883), .IN2(n5871), .Q(n14342) );
  OR2X1 U15166 ( .IN1(n9135), .IN2(n14343), .Q(n14340) );
  AND2X1 U15167 ( .IN1(n5886), .IN2(n5872), .Q(n14343) );
  AND2X1 U15168 ( .IN1(n14344), .IN2(n14332), .Q(n9881) );
  AND2X1 U15169 ( .IN1(n14336), .IN2(n14335), .Q(n14332) );
  AND2X1 U15170 ( .IN1(n14338), .IN2(n14337), .Q(n14335) );
  INVX0 U15171 ( .INP(n14345), .ZN(n14337) );
  AND2X1 U15172 ( .IN1(n9041), .IN2(n14346), .Q(n14345) );
  OR2X1 U15173 ( .IN1(g5831), .IN2(test_so83), .Q(n14346) );
  OR2X1 U15174 ( .IN1(n9136), .IN2(n14347), .Q(n14338) );
  AND2X1 U15175 ( .IN1(n5888), .IN2(n5874), .Q(n14347) );
  OR2X1 U15176 ( .IN1(n9126), .IN2(n14348), .Q(n14336) );
  AND2X1 U15177 ( .IN1(n5884), .IN2(n5870), .Q(n14348) );
  OR2X1 U15178 ( .IN1(n14349), .IN2(n9122), .Q(n14344) );
  AND2X1 U15179 ( .IN1(n5869), .IN2(n5885), .Q(n14349) );
  OR2X1 U15180 ( .IN1(n14350), .IN2(n14351), .Q(g26971) );
  AND2X1 U15181 ( .IN1(n14352), .IN2(n9016), .Q(n14351) );
  OR2X1 U15182 ( .IN1(n5670), .IN2(n8742), .Q(n14352) );
  AND2X1 U15183 ( .IN1(n9149), .IN2(g4512), .Q(n14350) );
  OR2X1 U15184 ( .IN1(n14353), .IN2(n14354), .Q(g26970) );
  AND2X1 U15185 ( .IN1(n9149), .IN2(g4459), .Q(n14354) );
  AND2X1 U15186 ( .IN1(n9041), .IN2(g4473), .Q(n14353) );
  OR2X1 U15187 ( .IN1(n14355), .IN2(n14356), .Q(g26969) );
  AND3X1 U15188 ( .IN1(n8752), .IN2(n8838), .IN3(n9065), .Q(n14356) );
  AND2X1 U15189 ( .IN1(n9149), .IN2(g4462), .Q(n14355) );
  OR2X1 U15190 ( .IN1(n14357), .IN2(n14358), .Q(g26968) );
  AND2X1 U15191 ( .IN1(n9149), .IN2(g4558), .Q(n14358) );
  OR2X1 U15192 ( .IN1(n14359), .IN2(n14360), .Q(g26967) );
  AND2X1 U15193 ( .IN1(n9149), .IN2(g4561), .Q(n14360) );
  OR2X1 U15194 ( .IN1(n14361), .IN2(n14362), .Q(g26966) );
  AND2X1 U15195 ( .IN1(n9148), .IN2(g4555), .Q(n14362) );
  AND2X1 U15196 ( .IN1(n14363), .IN2(n14364), .Q(g26965) );
  INVX0 U15197 ( .INP(n14365), .ZN(n14364) );
  AND2X1 U15198 ( .IN1(n14366), .IN2(n15422), .Q(n14365) );
  OR2X1 U15199 ( .IN1(n15422), .IN2(n14366), .Q(n14363) );
  OR2X1 U15200 ( .IN1(n8691), .IN2(n9122), .Q(n14366) );
  OR2X1 U15201 ( .IN1(n14367), .IN2(n14368), .Q(g26964) );
  AND2X1 U15202 ( .IN1(n14369), .IN2(g4527), .Q(n14368) );
  OR2X1 U15203 ( .IN1(n9124), .IN2(n14370), .Q(n14369) );
  AND2X1 U15204 ( .IN1(n5752), .IN2(n14055), .Q(n14370) );
  INVX0 U15205 ( .INP(n10459), .ZN(n14055) );
  AND3X1 U15206 ( .IN1(n14371), .IN2(n14372), .IN3(n9064), .Q(n14367) );
  OR2X1 U15207 ( .IN1(n5752), .IN2(g4515), .Q(n14372) );
  OR2X1 U15208 ( .IN1(n14373), .IN2(g4521), .Q(n14371) );
  AND2X1 U15209 ( .IN1(n10459), .IN2(n8514), .Q(n14373) );
  AND4X1 U15210 ( .IN1(g4483), .IN2(test_so27), .IN3(g4492), .IN4(g4489), .Q(
        n10459) );
  OR2X1 U15211 ( .IN1(n14359), .IN2(n14374), .Q(g26963) );
  AND2X1 U15212 ( .IN1(n9148), .IN2(g4489), .Q(n14374) );
  AND2X1 U15213 ( .IN1(g6750), .IN2(n9017), .Q(n14359) );
  OR2X1 U15214 ( .IN1(n14375), .IN2(n14357), .Q(g26962) );
  AND2X1 U15215 ( .IN1(g6749), .IN2(n9016), .Q(n14357) );
  AND2X1 U15216 ( .IN1(test_so27), .IN2(n9137), .Q(n14375) );
  OR2X1 U15217 ( .IN1(n14361), .IN2(n14376), .Q(g26961) );
  AND2X1 U15218 ( .IN1(n9148), .IN2(g4483), .Q(n14376) );
  AND2X1 U15219 ( .IN1(g6748), .IN2(n9016), .Q(n14361) );
  OR2X1 U15220 ( .IN1(n14377), .IN2(n14378), .Q(g26958) );
  AND2X1 U15221 ( .IN1(n9148), .IN2(g4455), .Q(n14377) );
  OR2X1 U15222 ( .IN1(n14379), .IN2(n14380), .Q(g26957) );
  AND2X1 U15223 ( .IN1(test_so47), .IN2(n9016), .Q(n14380) );
  AND2X1 U15224 ( .IN1(n14381), .IN2(g4434), .Q(n14379) );
  OR2X1 U15225 ( .IN1(n9125), .IN2(n14382), .Q(n14381) );
  AND2X1 U15226 ( .IN1(n14383), .IN2(g4392), .Q(n14382) );
  OR2X1 U15227 ( .IN1(n14384), .IN2(n9336), .Q(g26956) );
  AND3X1 U15228 ( .IN1(n14383), .IN2(g4430), .IN3(n14385), .Q(n14384) );
  OR2X1 U15229 ( .IN1(n14386), .IN2(n14387), .Q(g26955) );
  AND2X1 U15230 ( .IN1(n14388), .IN2(g4438), .Q(n14387) );
  AND2X1 U15231 ( .IN1(n14383), .IN2(n14389), .Q(n14386) );
  OR3X1 U15232 ( .IN1(n14390), .IN2(n14391), .IN3(n14392), .Q(g26954) );
  AND2X1 U15233 ( .IN1(test_so47), .IN2(n9138), .Q(n14392) );
  AND2X1 U15234 ( .IN1(n14393), .IN2(g4438), .Q(n14391) );
  AND2X1 U15235 ( .IN1(n14385), .IN2(n14383), .Q(n14390) );
  INVX0 U15236 ( .INP(n14394), .ZN(n14383) );
  OR4X1 U15237 ( .IN1(test_so47), .IN2(g4438), .IN3(n9336), .IN4(n14395), .Q(
        n14394) );
  OR2X1 U15238 ( .IN1(g7245), .IN2(g7260), .Q(n14395) );
  OR2X1 U15239 ( .IN1(n14396), .IN2(n14397), .Q(g26952) );
  AND2X1 U15240 ( .IN1(n14398), .IN2(g4430), .Q(n14397) );
  AND2X1 U15241 ( .IN1(n14399), .IN2(n9015), .Q(n14396) );
  OR3X1 U15242 ( .IN1(n14400), .IN2(n14401), .IN3(n14402), .Q(n14399) );
  AND2X1 U15243 ( .IN1(n14398), .IN2(g4388), .Q(n14402) );
  OR3X1 U15244 ( .IN1(n8731), .IN2(n8728), .IN3(n9121), .Q(n14398) );
  AND2X1 U15245 ( .IN1(n8342), .IN2(g4434), .Q(n14401) );
  AND2X1 U15246 ( .IN1(n8343), .IN2(g4401), .Q(n14400) );
  OR2X1 U15247 ( .IN1(n14403), .IN2(g26953), .Q(g26951) );
  AND2X1 U15248 ( .IN1(n9148), .IN2(g4427), .Q(n14403) );
  OR2X1 U15249 ( .IN1(n14404), .IN2(n14378), .Q(g26950) );
  OR2X1 U15250 ( .IN1(n14405), .IN2(n14406), .Q(n14378) );
  AND2X1 U15251 ( .IN1(n14407), .IN2(n9015), .Q(n14406) );
  AND2X1 U15252 ( .IN1(n14389), .IN2(n14408), .Q(n14405) );
  AND2X1 U15253 ( .IN1(n9145), .IN2(g4417), .Q(n14404) );
  OR2X1 U15254 ( .IN1(n14409), .IN2(n14410), .Q(g26949) );
  AND2X1 U15255 ( .IN1(n9041), .IN2(g4411), .Q(n14410) );
  AND2X1 U15256 ( .IN1(n14411), .IN2(g4401), .Q(n14409) );
  OR2X1 U15257 ( .IN1(n9126), .IN2(n14412), .Q(n14411) );
  AND2X1 U15258 ( .IN1(n14413), .IN2(g4392), .Q(n14412) );
  OR2X1 U15259 ( .IN1(n14414), .IN2(g4405), .Q(g26948) );
  AND3X1 U15260 ( .IN1(n14413), .IN2(g4388), .IN3(n14385), .Q(n14414) );
  OR3X1 U15261 ( .IN1(n14415), .IN2(n14416), .IN3(n14417), .Q(g26947) );
  AND2X1 U15262 ( .IN1(n14418), .IN2(n9015), .Q(n14416) );
  OR2X1 U15263 ( .IN1(n14419), .IN2(n14407), .Q(n14418) );
  AND3X1 U15264 ( .IN1(n14413), .IN2(n5710), .IN3(n8790), .Q(n14407) );
  AND3X1 U15265 ( .IN1(n14408), .IN2(g4382), .IN3(n8277), .Q(n14419) );
  AND2X1 U15266 ( .IN1(n9148), .IN2(g4388), .Q(n14415) );
  OR2X1 U15267 ( .IN1(n14420), .IN2(n14421), .Q(g26946) );
  AND2X1 U15268 ( .IN1(n14388), .IN2(g4375), .Q(n14421) );
  AND2X1 U15269 ( .IN1(n14413), .IN2(n14389), .Q(n14420) );
  AND2X1 U15270 ( .IN1(g4392), .IN2(n9015), .Q(n14389) );
  OR3X1 U15271 ( .IN1(n14422), .IN2(n14417), .IN3(n14423), .Q(g26945) );
  AND2X1 U15272 ( .IN1(n9148), .IN2(g4411), .Q(n14423) );
  AND2X1 U15273 ( .IN1(n14393), .IN2(g4375), .Q(n14417) );
  INVX0 U15274 ( .INP(n14388), .ZN(n14393) );
  OR2X1 U15275 ( .IN1(n9126), .IN2(g4382), .Q(n14388) );
  AND2X1 U15276 ( .IN1(n14385), .IN2(n14413), .Q(n14422) );
  INVX0 U15277 ( .INP(n14408), .ZN(n14413) );
  OR4X1 U15278 ( .IN1(g4405), .IN2(g4375), .IN3(g4411), .IN4(n14424), .Q(
        n14408) );
  OR2X1 U15279 ( .IN1(g7257), .IN2(g7243), .Q(n14424) );
  AND2X1 U15280 ( .IN1(n9041), .IN2(n5710), .Q(n14385) );
  AND2X1 U15281 ( .IN1(n14425), .IN2(n9015), .Q(g26944) );
  INVX0 U15282 ( .INP(n14426), .ZN(n14425) );
  AND4X1 U15283 ( .IN1(n9795), .IN2(n14427), .IN3(g4358), .IN4(test_so81), .Q(
        n14426) );
  INVX0 U15284 ( .INP(n14428), .ZN(n9795) );
  OR2X1 U15285 ( .IN1(n14429), .IN2(g135), .Q(n14428) );
  AND3X1 U15286 ( .IN1(n14430), .IN2(n14431), .IN3(n14432), .Q(n14429) );
  OR4X1 U15287 ( .IN1(g4616), .IN2(n14433), .IN3(n14434), .IN4(n14435), .Q(
        n14432) );
  AND2X1 U15288 ( .IN1(n5274), .IN2(g4584), .Q(n14435) );
  AND2X1 U15289 ( .IN1(n5539), .IN2(g4608), .Q(n14434) );
  OR2X1 U15290 ( .IN1(n14436), .IN2(n14437), .Q(n14433) );
  AND2X1 U15291 ( .IN1(n5303), .IN2(g4601), .Q(n14437) );
  AND2X1 U15292 ( .IN1(n5365), .IN2(g4593), .Q(n14436) );
  OR4X1 U15293 ( .IN1(n5303), .IN2(g4601), .IN3(g4608), .IN4(n5539), .Q(n14431) );
  OR3X1 U15294 ( .IN1(n5274), .IN2(g4593), .IN3(g4584), .Q(n14430) );
  OR2X1 U15295 ( .IN1(n14438), .IN2(n14439), .Q(g26940) );
  AND2X1 U15296 ( .IN1(n12516), .IN2(n9015), .Q(n14439) );
  OR2X1 U15297 ( .IN1(n14440), .IN2(n14441), .Q(n12516) );
  AND2X1 U15298 ( .IN1(g114), .IN2(n5983), .Q(n14441) );
  AND2X1 U15299 ( .IN1(g116), .IN2(g4157), .Q(n14440) );
  AND2X1 U15300 ( .IN1(n9148), .IN2(g4153), .Q(n14438) );
  OR2X1 U15301 ( .IN1(n14442), .IN2(n14443), .Q(g26939) );
  AND2X1 U15302 ( .IN1(n12521), .IN2(n9016), .Q(n14443) );
  OR2X1 U15303 ( .IN1(n14444), .IN2(n14445), .Q(n12521) );
  AND2X1 U15304 ( .IN1(g120), .IN2(n5981), .Q(n14445) );
  AND2X1 U15305 ( .IN1(g124), .IN2(g4146), .Q(n14444) );
  AND2X1 U15306 ( .IN1(n9147), .IN2(g4104), .Q(n14442) );
  OR3X1 U15307 ( .IN1(n8811), .IN2(n14446), .IN3(n14447), .Q(g26938) );
  AND2X1 U15308 ( .IN1(n14448), .IN2(g4141), .Q(n14447) );
  OR2X1 U15309 ( .IN1(n9126), .IN2(n14449), .Q(n14448) );
  AND2X1 U15310 ( .IN1(n14081), .IN2(n14450), .Q(n14449) );
  AND3X1 U15311 ( .IN1(n9057), .IN2(g4082), .IN3(n14081), .Q(n14446) );
  INVX0 U15312 ( .INP(n12528), .ZN(n14081) );
  AND3X1 U15313 ( .IN1(g4082), .IN2(g4141), .IN3(n14450), .Q(n12528) );
  OR3X1 U15314 ( .IN1(n14451), .IN2(n14452), .IN3(n14453), .Q(g26934) );
  AND2X1 U15315 ( .IN1(n4888), .IN2(g2827), .Q(n14453) );
  AND2X1 U15316 ( .IN1(test_so37), .IN2(n9138), .Q(n14452) );
  AND2X1 U15317 ( .IN1(n14454), .IN2(n8856), .Q(n14451) );
  OR3X1 U15318 ( .IN1(n14455), .IN2(n14456), .IN3(n14457), .Q(g26933) );
  AND2X1 U15319 ( .IN1(test_so37), .IN2(n4888), .Q(n14457) );
  AND2X1 U15320 ( .IN1(n9147), .IN2(g2811), .Q(n14456) );
  AND2X1 U15321 ( .IN1(n5840), .IN2(n14454), .Q(n14455) );
  OR3X1 U15322 ( .IN1(n14458), .IN2(n14459), .IN3(n14460), .Q(g26932) );
  AND2X1 U15323 ( .IN1(n4888), .IN2(g2811), .Q(n14460) );
  AND2X1 U15324 ( .IN1(n9147), .IN2(g2799), .Q(n14459) );
  AND2X1 U15325 ( .IN1(n5841), .IN2(n14454), .Q(n14458) );
  OR3X1 U15326 ( .IN1(n14461), .IN2(n14462), .IN3(n14463), .Q(g26931) );
  AND2X1 U15327 ( .IN1(n4888), .IN2(g2799), .Q(n14463) );
  AND2X1 U15328 ( .IN1(n9147), .IN2(g29219), .Q(n14462) );
  AND2X1 U15329 ( .IN1(n5839), .IN2(n14454), .Q(n14461) );
  OR3X1 U15330 ( .IN1(n14464), .IN2(n14465), .IN3(n14466), .Q(g26930) );
  AND2X1 U15331 ( .IN1(n4888), .IN2(g2795), .Q(n14466) );
  AND2X1 U15332 ( .IN1(n9147), .IN2(g2791), .Q(n14465) );
  AND2X1 U15333 ( .IN1(n14454), .IN2(n8857), .Q(n14464) );
  OR3X1 U15334 ( .IN1(n14467), .IN2(n14468), .IN3(n14469), .Q(g26929) );
  AND2X1 U15335 ( .IN1(n4888), .IN2(g2791), .Q(n14469) );
  AND2X1 U15336 ( .IN1(n9147), .IN2(g2779), .Q(n14468) );
  AND2X1 U15337 ( .IN1(n5837), .IN2(n14454), .Q(n14467) );
  OR3X1 U15338 ( .IN1(n14470), .IN2(n14471), .IN3(n14472), .Q(g26928) );
  AND2X1 U15339 ( .IN1(n4888), .IN2(g2779), .Q(n14472) );
  AND2X1 U15340 ( .IN1(n9147), .IN2(g2767), .Q(n14471) );
  AND2X1 U15341 ( .IN1(n5834), .IN2(n14454), .Q(n14470) );
  OR3X1 U15342 ( .IN1(n14473), .IN2(n14474), .IN3(n14475), .Q(g26927) );
  AND2X1 U15343 ( .IN1(n4888), .IN2(g2767), .Q(n14475) );
  AND2X1 U15344 ( .IN1(n9147), .IN2(g2763), .Q(n14474) );
  AND2X1 U15345 ( .IN1(n5836), .IN2(n14454), .Q(n14473) );
  AND3X1 U15346 ( .IN1(n10179), .IN2(n9463), .IN3(n4888), .Q(n14454) );
  OR2X1 U15347 ( .IN1(test_so30), .IN2(g2748), .Q(n9463) );
  INVX0 U15348 ( .INP(n10185), .ZN(n10179) );
  AND3X1 U15349 ( .IN1(g2735), .IN2(n3505), .IN3(test_so30), .Q(n10185) );
  AND2X1 U15350 ( .IN1(g2748), .IN2(g2741), .Q(n3505) );
  OR2X1 U15351 ( .IN1(n14476), .IN2(n14477), .Q(g26926) );
  AND2X1 U15352 ( .IN1(n9147), .IN2(g2719), .Q(n14477) );
  AND3X1 U15353 ( .IN1(n14478), .IN2(n14479), .IN3(n3730), .Q(n14476) );
  OR2X1 U15354 ( .IN1(n14224), .IN2(g2724), .Q(n14479) );
  INVX0 U15355 ( .INP(n12798), .ZN(n14224) );
  OR2X1 U15356 ( .IN1(n5301), .IN2(n12798), .Q(n14478) );
  OR2X1 U15357 ( .IN1(n5465), .IN2(n5299), .Q(n12798) );
  OR2X1 U15358 ( .IN1(n14480), .IN2(n14481), .Q(g26925) );
  AND2X1 U15359 ( .IN1(n14482), .IN2(n9014), .Q(n14481) );
  OR2X1 U15360 ( .IN1(n14483), .IN2(n4173), .Q(n14482) );
  AND2X1 U15361 ( .IN1(n13062), .IN2(g1536), .Q(n14483) );
  OR2X1 U15362 ( .IN1(n8791), .IN2(n13065), .Q(n13062) );
  OR2X1 U15363 ( .IN1(n8378), .IN2(n13072), .Q(n13065) );
  OR3X1 U15364 ( .IN1(n5302), .IN2(n13084), .IN3(n13606), .Q(n13072) );
  AND3X1 U15365 ( .IN1(g1521), .IN2(g1339), .IN3(n8573), .Q(n13084) );
  AND2X1 U15366 ( .IN1(n9147), .IN2(g1532), .Q(n14480) );
  OR3X1 U15367 ( .IN1(n14484), .IN2(n14485), .IN3(n14486), .Q(g26924) );
  AND2X1 U15368 ( .IN1(n14487), .IN2(n5289), .Q(n14486) );
  INVX0 U15369 ( .INP(n14488), .ZN(n14487) );
  AND2X1 U15370 ( .IN1(n9147), .IN2(g1437), .Q(n14485) );
  AND3X1 U15371 ( .IN1(n14488), .IN2(g1478), .IN3(n9063), .Q(n14484) );
  OR3X1 U15372 ( .IN1(n5696), .IN2(n13635), .IN3(n14489), .Q(n14488) );
  OR2X1 U15373 ( .IN1(test_so49), .IN2(n5364), .Q(n13635) );
  OR3X1 U15374 ( .IN1(n14490), .IN2(n14491), .IN3(n14492), .Q(g26923) );
  AND2X1 U15375 ( .IN1(n14493), .IN2(n5290), .Q(n14492) );
  INVX0 U15376 ( .INP(n14494), .ZN(n14493) );
  AND2X1 U15377 ( .IN1(n9146), .IN2(g1467), .Q(n14491) );
  AND3X1 U15378 ( .IN1(n14494), .IN2(g1472), .IN3(n9063), .Q(n14490) );
  OR3X1 U15379 ( .IN1(n5693), .IN2(n13627), .IN3(n14489), .Q(n14494) );
  OR3X1 U15380 ( .IN1(n14495), .IN2(n14496), .IN3(n14497), .Q(g26922) );
  AND2X1 U15381 ( .IN1(n14498), .IN2(n5343), .Q(n14497) );
  INVX0 U15382 ( .INP(n14499), .ZN(n14498) );
  AND2X1 U15383 ( .IN1(n9146), .IN2(g1454), .Q(n14496) );
  AND3X1 U15384 ( .IN1(n14499), .IN2(g1448), .IN3(n9063), .Q(n14495) );
  OR3X1 U15385 ( .IN1(n5866), .IN2(n13606), .IN3(n14489), .Q(n14499) );
  OR2X1 U15386 ( .IN1(n8741), .IN2(n14500), .Q(n14489) );
  OR2X1 U15387 ( .IN1(n8819), .IN2(g1514), .Q(n13606) );
  OR2X1 U15388 ( .IN1(n14501), .IN2(n14502), .Q(g26921) );
  AND4X1 U15389 ( .IN1(n14503), .IN2(n14504), .IN3(n8824), .IN4(n9049), .Q(
        n14502) );
  OR2X1 U15390 ( .IN1(n14505), .IN2(g1404), .Q(n14504) );
  OR2X1 U15391 ( .IN1(n8757), .IN2(n14506), .Q(n14503) );
  AND2X1 U15392 ( .IN1(n9146), .IN2(g1395), .Q(n14501) );
  OR3X1 U15393 ( .IN1(n14507), .IN2(n14508), .IN3(n14509), .Q(g26920) );
  AND2X1 U15394 ( .IN1(n4913), .IN2(n14510), .Q(n14509) );
  AND3X1 U15395 ( .IN1(n9495), .IN2(g1389), .IN3(n9063), .Q(n14508) );
  OR2X1 U15396 ( .IN1(n14511), .IN2(n14512), .Q(n9495) );
  AND2X1 U15397 ( .IN1(n8764), .IN2(g1351), .Q(n14511) );
  AND2X1 U15398 ( .IN1(n9146), .IN2(g1384), .Q(n14507) );
  OR3X1 U15399 ( .IN1(n14513), .IN2(n14514), .IN3(n14515), .Q(g26919) );
  AND2X1 U15400 ( .IN1(n9146), .IN2(g1266), .Q(n14515) );
  AND2X1 U15401 ( .IN1(n4804), .IN2(n5556), .Q(n14514) );
  AND3X1 U15402 ( .IN1(test_so77), .IN2(n11485), .IN3(n14516), .Q(n14513) );
  INVX0 U15403 ( .INP(n4804), .ZN(n14516) );
  AND3X1 U15404 ( .IN1(g1249), .IN2(g1266), .IN3(g12923), .Q(n4804) );
  OR2X1 U15405 ( .IN1(n14517), .IN2(n14518), .Q(g26918) );
  AND2X1 U15406 ( .IN1(n14519), .IN2(n9014), .Q(n14518) );
  OR2X1 U15407 ( .IN1(n14520), .IN2(n4191), .Q(n14519) );
  AND2X1 U15408 ( .IN1(n13098), .IN2(g1193), .Q(n14520) );
  OR2X1 U15409 ( .IN1(n8792), .IN2(n13101), .Q(n13098) );
  OR2X1 U15410 ( .IN1(n8379), .IN2(n13108), .Q(n13101) );
  OR3X1 U15411 ( .IN1(n5304), .IN2(n13119), .IN3(n13650), .Q(n13108) );
  AND3X1 U15412 ( .IN1(g996), .IN2(g1178), .IN3(n5642), .Q(n13119) );
  AND2X1 U15413 ( .IN1(n9146), .IN2(g1189), .Q(n14517) );
  OR3X1 U15414 ( .IN1(n14521), .IN2(n14522), .IN3(n14523), .Q(g26917) );
  AND2X1 U15415 ( .IN1(n14524), .IN2(n5328), .Q(n14523) );
  INVX0 U15416 ( .INP(n14525), .ZN(n14524) );
  AND2X1 U15417 ( .IN1(n9146), .IN2(g1094), .Q(n14522) );
  AND3X1 U15418 ( .IN1(n14525), .IN2(g1135), .IN3(n9063), .Q(n14521) );
  OR3X1 U15419 ( .IN1(n5697), .IN2(g1183), .IN3(n14526), .Q(n14525) );
  OR3X1 U15420 ( .IN1(n14527), .IN2(n14528), .IN3(n14529), .Q(g26916) );
  AND2X1 U15421 ( .IN1(n14530), .IN2(n5329), .Q(n14529) );
  INVX0 U15422 ( .INP(n14531), .ZN(n14530) );
  AND2X1 U15423 ( .IN1(n9146), .IN2(g1124), .Q(n14528) );
  AND3X1 U15424 ( .IN1(n14531), .IN2(g1129), .IN3(n9063), .Q(n14527) );
  OR3X1 U15425 ( .IN1(n5692), .IN2(n5599), .IN3(n14526), .Q(n14531) );
  OR3X1 U15426 ( .IN1(n8748), .IN2(n5363), .IN3(n14532), .Q(n14526) );
  OR3X1 U15427 ( .IN1(n14533), .IN2(n14534), .IN3(n14535), .Q(g26915) );
  AND2X1 U15428 ( .IN1(n14536), .IN2(n5478), .Q(n14535) );
  AND2X1 U15429 ( .IN1(test_so90), .IN2(n9140), .Q(n14534) );
  AND3X1 U15430 ( .IN1(n14537), .IN2(g1105), .IN3(n9063), .Q(n14533) );
  INVX0 U15431 ( .INP(n14536), .ZN(n14537) );
  AND4X1 U15432 ( .IN1(test_so90), .IN2(n14538), .IN3(g13259), .IN4(n11430), 
        .Q(n14536) );
  INVX0 U15433 ( .INP(n13650), .ZN(n11430) );
  OR2X1 U15434 ( .IN1(n5599), .IN2(g1171), .Q(n13650) );
  OR2X1 U15435 ( .IN1(n14539), .IN2(n14540), .Q(g26914) );
  AND4X1 U15436 ( .IN1(n14541), .IN2(n14542), .IN3(n5320), .IN4(n9049), .Q(
        n14540) );
  OR2X1 U15437 ( .IN1(n14543), .IN2(g1061), .Q(n14542) );
  OR2X1 U15438 ( .IN1(n8756), .IN2(n14544), .Q(n14541) );
  AND2X1 U15439 ( .IN1(n9145), .IN2(g1052), .Q(n14539) );
  OR3X1 U15440 ( .IN1(n14545), .IN2(n14546), .IN3(n14547), .Q(g26913) );
  AND2X1 U15441 ( .IN1(n4938), .IN2(n14548), .Q(n14547) );
  AND3X1 U15442 ( .IN1(n9341), .IN2(g1046), .IN3(n9062), .Q(n14546) );
  OR2X1 U15443 ( .IN1(n14549), .IN2(n14550), .Q(n9341) );
  AND2X1 U15444 ( .IN1(n8765), .IN2(g1008), .Q(n14549) );
  AND2X1 U15445 ( .IN1(n9145), .IN2(g1041), .Q(n14545) );
  OR3X1 U15446 ( .IN1(n14551), .IN2(n14552), .IN3(n14553), .Q(g26912) );
  AND2X1 U15447 ( .IN1(n9145), .IN2(g921), .Q(n14553) );
  AND2X1 U15448 ( .IN1(n4811), .IN2(n5557), .Q(n14552) );
  AND3X1 U15449 ( .IN1(n11500), .IN2(n14554), .IN3(g936), .Q(n14551) );
  INVX0 U15450 ( .INP(n4811), .ZN(n14554) );
  AND3X1 U15451 ( .IN1(g904), .IN2(g921), .IN3(g12919), .Q(n4811) );
  OR2X1 U15452 ( .IN1(n14555), .IN2(n14556), .Q(g26910) );
  AND3X1 U15453 ( .IN1(n5305), .IN2(n9052), .IN3(n5682), .Q(n14556) );
  AND2X1 U15454 ( .IN1(n14557), .IN2(g862), .Q(n14555) );
  OR2X1 U15455 ( .IN1(n9129), .IN2(g890), .Q(n14557) );
  OR2X1 U15456 ( .IN1(n14558), .IN2(n14559), .Q(g26909) );
  AND2X1 U15457 ( .IN1(n14560), .IN2(n9014), .Q(n14559) );
  OR2X1 U15458 ( .IN1(n14561), .IN2(n14562), .Q(n14560) );
  AND2X1 U15459 ( .IN1(n5305), .IN2(g896), .Q(n14562) );
  AND2X1 U15460 ( .IN1(n5431), .IN2(g862), .Q(n14561) );
  AND2X1 U15461 ( .IN1(n9145), .IN2(g890), .Q(n14558) );
  OR3X1 U15462 ( .IN1(n14563), .IN2(n14564), .IN3(n14565), .Q(g26908) );
  AND2X1 U15463 ( .IN1(n4945), .IN2(g446), .Q(n14565) );
  AND2X1 U15464 ( .IN1(n9145), .IN2(g246), .Q(n14564) );
  AND2X1 U15465 ( .IN1(n14566), .IN2(g872), .Q(n14563) );
  OR3X1 U15466 ( .IN1(n14567), .IN2(n14568), .IN3(n14569), .Q(g26907) );
  AND2X1 U15467 ( .IN1(n4945), .IN2(g246), .Q(n14569) );
  AND2X1 U15468 ( .IN1(n9145), .IN2(g269), .Q(n14568) );
  AND2X1 U15469 ( .IN1(n14566), .IN2(g14167), .Q(n14567) );
  OR3X1 U15470 ( .IN1(n14570), .IN2(n14571), .IN3(n14572), .Q(g26906) );
  AND2X1 U15471 ( .IN1(n4945), .IN2(g269), .Q(n14572) );
  AND2X1 U15472 ( .IN1(n9145), .IN2(g239), .Q(n14571) );
  AND2X1 U15473 ( .IN1(n14566), .IN2(g14147), .Q(n14570) );
  OR3X1 U15474 ( .IN1(n14573), .IN2(n14574), .IN3(n14575), .Q(g26905) );
  AND2X1 U15475 ( .IN1(n4945), .IN2(g239), .Q(n14575) );
  AND2X1 U15476 ( .IN1(n9145), .IN2(g262), .Q(n14574) );
  AND2X1 U15477 ( .IN1(n14566), .IN2(g14125), .Q(n14573) );
  OR3X1 U15478 ( .IN1(n14576), .IN2(n14577), .IN3(n14578), .Q(g26904) );
  AND2X1 U15479 ( .IN1(n4945), .IN2(g262), .Q(n14578) );
  AND2X1 U15480 ( .IN1(n9145), .IN2(g232), .Q(n14577) );
  AND2X1 U15481 ( .IN1(n14566), .IN2(g14096), .Q(n14576) );
  OR3X1 U15482 ( .IN1(n14579), .IN2(n14580), .IN3(n14581), .Q(g26903) );
  AND2X1 U15483 ( .IN1(n4945), .IN2(g232), .Q(n14581) );
  AND2X1 U15484 ( .IN1(n9145), .IN2(g255), .Q(n14580) );
  AND2X1 U15485 ( .IN1(n14566), .IN2(g14217), .Q(n14579) );
  OR3X1 U15486 ( .IN1(n14582), .IN2(n14583), .IN3(n14584), .Q(g26902) );
  AND2X1 U15487 ( .IN1(n4945), .IN2(g255), .Q(n14584) );
  AND2X1 U15488 ( .IN1(n9145), .IN2(g225), .Q(n14583) );
  AND2X1 U15489 ( .IN1(n14566), .IN2(g14201), .Q(n14582) );
  OR3X1 U15490 ( .IN1(n14585), .IN2(n14586), .IN3(n14587), .Q(g26901) );
  AND2X1 U15491 ( .IN1(n4945), .IN2(g225), .Q(n14587) );
  AND2X1 U15492 ( .IN1(n9145), .IN2(g872), .Q(n14586) );
  AND2X1 U15493 ( .IN1(n14566), .IN2(g14189), .Q(n14585) );
  AND2X1 U15494 ( .IN1(n9041), .IN2(n9511), .Q(n14566) );
  AND3X1 U15495 ( .IN1(g890), .IN2(n5431), .IN3(n5682), .Q(n9511) );
  OR2X1 U15496 ( .IN1(n14588), .IN2(n14589), .Q(g26899) );
  AND2X1 U15497 ( .IN1(n9145), .IN2(g832), .Q(n14589) );
  AND2X1 U15498 ( .IN1(n14590), .IN2(n14591), .Q(n14588) );
  OR2X1 U15499 ( .IN1(n5422), .IN2(n14592), .Q(n14591) );
  INVX0 U15500 ( .INP(n4814), .ZN(n14592) );
  OR2X1 U15501 ( .IN1(n14593), .IN2(n14594), .Q(n14590) );
  AND2X1 U15502 ( .IN1(n4518), .IN2(g822), .Q(n14594) );
  AND2X1 U15503 ( .IN1(n4814), .IN2(n13689), .Q(n14593) );
  AND3X1 U15504 ( .IN1(g832), .IN2(g817), .IN3(n4948), .Q(n4814) );
  OR2X1 U15505 ( .IN1(n14595), .IN2(n14596), .Q(g26898) );
  AND2X1 U15506 ( .IN1(n14597), .IN2(g843), .Q(n14596) );
  OR2X1 U15507 ( .IN1(n9129), .IN2(n14598), .Q(n14597) );
  AND3X1 U15508 ( .IN1(n5733), .IN2(g837), .IN3(n14599), .Q(n14598) );
  AND3X1 U15509 ( .IN1(g837), .IN2(g812), .IN3(n14600), .Q(n14595) );
  OR2X1 U15510 ( .IN1(n14601), .IN2(n13727), .Q(n14600) );
  AND2X1 U15511 ( .IN1(n14602), .IN2(n9014), .Q(n14601) );
  OR2X1 U15512 ( .IN1(n5709), .IN2(n8356), .Q(n14602) );
  OR2X1 U15513 ( .IN1(n14603), .IN2(n14604), .Q(g26897) );
  AND2X1 U15514 ( .IN1(n14605), .IN2(g732), .Q(n14604) );
  INVX0 U15515 ( .INP(n14606), .ZN(n14605) );
  AND2X1 U15516 ( .IN1(n14606), .IN2(g753), .Q(n14603) );
  AND2X1 U15517 ( .IN1(n9040), .IN2(n14317), .Q(n14606) );
  OR3X1 U15518 ( .IN1(n14607), .IN2(n14608), .IN3(n14609), .Q(g26896) );
  AND2X1 U15519 ( .IN1(n4956), .IN2(n13713), .Q(n14609) );
  AND2X1 U15520 ( .IN1(n14610), .IN2(g728), .Q(n14608) );
  AND2X1 U15521 ( .IN1(n14611), .IN2(g29212), .Q(n14607) );
  INVX0 U15522 ( .INP(n14610), .ZN(n14611) );
  OR2X1 U15523 ( .IN1(n9129), .IN2(n13713), .Q(n14610) );
  AND4X1 U15524 ( .IN1(n14612), .IN2(test_so54), .IN3(n5519), .IN4(n4948), .Q(
        n13713) );
  OR3X1 U15525 ( .IN1(n14613), .IN2(n14614), .IN3(n14615), .Q(g26895) );
  AND2X1 U15526 ( .IN1(n9145), .IN2(g562), .Q(n14615) );
  AND2X1 U15527 ( .IN1(n4826), .IN2(n5335), .Q(n14614) );
  INVX0 U15528 ( .INP(n14616), .ZN(n4826) );
  AND3X1 U15529 ( .IN1(n2421), .IN2(n14616), .IN3(g568), .Q(n14613) );
  OR2X1 U15530 ( .IN1(n14617), .IN2(n14618), .Q(n14616) );
  INVX0 U15531 ( .INP(n4959), .ZN(n14618) );
  OR2X1 U15532 ( .IN1(n14619), .IN2(n14620), .Q(g26894) );
  AND4X1 U15533 ( .IN1(n14621), .IN2(n14622), .IN3(n14623), .IN4(n9049), .Q(
        n14620) );
  OR2X1 U15534 ( .IN1(n5327), .IN2(n14306), .Q(n14622) );
  INVX0 U15535 ( .INP(n14309), .ZN(n14306) );
  OR2X1 U15536 ( .IN1(n14624), .IN2(g528), .Q(n14621) );
  AND2X1 U15537 ( .IN1(n14309), .IN2(n14307), .Q(n14624) );
  INVX0 U15538 ( .INP(n14612), .ZN(n14307) );
  AND3X1 U15539 ( .IN1(g482), .IN2(g490), .IN3(n5327), .Q(n14612) );
  AND3X1 U15540 ( .IN1(g518), .IN2(n5548), .IN3(n14281), .Q(n14309) );
  AND2X1 U15541 ( .IN1(n9148), .IN2(g518), .Q(n14619) );
  OR2X1 U15542 ( .IN1(n14625), .IN2(n14626), .Q(g26893) );
  AND2X1 U15543 ( .IN1(n14627), .IN2(n9007), .Q(n14626) );
  OR2X1 U15544 ( .IN1(n14628), .IN2(n14629), .Q(n14627) );
  AND2X1 U15545 ( .IN1(test_so17), .IN2(n14630), .Q(n14629) );
  AND2X1 U15546 ( .IN1(g29211), .IN2(n8846), .Q(n14628) );
  AND2X1 U15547 ( .IN1(n9141), .IN2(g355), .Q(n14625) );
  OR2X1 U15548 ( .IN1(n14631), .IN2(n14632), .Q(g26892) );
  AND2X1 U15549 ( .IN1(test_so17), .IN2(n9137), .Q(n14632) );
  AND3X1 U15550 ( .IN1(n9056), .IN2(n14630), .IN3(n8846), .Q(n14631) );
  OR2X1 U15551 ( .IN1(g333), .IN2(g355), .Q(n14630) );
  OR2X1 U15552 ( .IN1(n14633), .IN2(n14634), .Q(g26891) );
  AND3X1 U15553 ( .IN1(n9057), .IN2(g7540), .IN3(n5860), .Q(n14634) );
  AND2X1 U15554 ( .IN1(n9145), .IN2(g347), .Q(n14633) );
  OR2X1 U15555 ( .IN1(n14635), .IN2(n14636), .Q(g26890) );
  AND2X1 U15556 ( .IN1(n9145), .IN2(g333), .Q(n14636) );
  AND2X1 U15557 ( .IN1(n5860), .IN2(n9014), .Q(n14635) );
  OR2X1 U15558 ( .IN1(n14637), .IN2(n14638), .Q(g26889) );
  AND4X1 U15559 ( .IN1(g329), .IN2(DFF_709_n1), .IN3(n14639), .IN4(n9049), .Q(
        n14638) );
  AND2X1 U15560 ( .IN1(n9145), .IN2(g29211), .Q(n14637) );
  OR2X1 U15561 ( .IN1(n14640), .IN2(n14641), .Q(g26888) );
  AND2X1 U15562 ( .IN1(n9145), .IN2(g29216), .Q(n14641) );
  AND2X1 U15563 ( .IN1(n9040), .IN2(g316), .Q(n14640) );
  OR3X1 U15564 ( .IN1(n14642), .IN2(n14643), .IN3(n14644), .Q(g26887) );
  AND3X1 U15565 ( .IN1(n5317), .IN2(g324), .IN3(n9061), .Q(n14643) );
  AND2X1 U15566 ( .IN1(n9145), .IN2(g336), .Q(n14642) );
  OR3X1 U15567 ( .IN1(n14645), .IN2(n14646), .IN3(n14647), .Q(g26886) );
  AND2X1 U15568 ( .IN1(n14644), .IN2(n14648), .Q(n14647) );
  AND2X1 U15569 ( .IN1(n9145), .IN2(g311), .Q(n14646) );
  AND3X1 U15570 ( .IN1(n14639), .IN2(g336), .IN3(n9061), .Q(n14645) );
  OR2X1 U15571 ( .IN1(n14649), .IN2(n14650), .Q(g26884) );
  AND2X1 U15572 ( .IN1(n14651), .IN2(n9030), .Q(n14650) );
  OR2X1 U15573 ( .IN1(n14652), .IN2(n14653), .Q(n14651) );
  AND2X1 U15574 ( .IN1(n14648), .IN2(n14654), .Q(n14653) );
  OR3X1 U15575 ( .IN1(n14655), .IN2(n14656), .IN3(g26885), .Q(n14654) );
  AND2X1 U15576 ( .IN1(g305), .IN2(g336), .Q(n14656) );
  AND2X1 U15577 ( .IN1(n5824), .IN2(g311), .Q(n14655) );
  AND4X1 U15578 ( .IN1(n5766), .IN2(n5456), .IN3(n5282), .IN4(n5317), .Q(
        n14652) );
  AND2X1 U15579 ( .IN1(n9146), .IN2(g329), .Q(n14649) );
  OR2X1 U15580 ( .IN1(n14657), .IN2(n14658), .Q(g26883) );
  AND2X1 U15581 ( .IN1(n14648), .IN2(n9030), .Q(n14658) );
  INVX0 U15582 ( .INP(n14639), .ZN(n14648) );
  OR2X1 U15583 ( .IN1(n14659), .IN2(n14660), .Q(n14639) );
  AND2X1 U15584 ( .IN1(n5827), .IN2(n5317), .Q(n14660) );
  AND2X1 U15585 ( .IN1(n5282), .IN2(g324), .Q(n14659) );
  AND2X1 U15586 ( .IN1(n9146), .IN2(g324), .Q(n14657) );
  OR3X1 U15587 ( .IN1(n14661), .IN2(n14662), .IN3(n14644), .Q(g26882) );
  AND2X1 U15588 ( .IN1(g305), .IN2(n9030), .Q(n14644) );
  AND2X1 U15589 ( .IN1(n9146), .IN2(g316), .Q(n14662) );
  AND2X1 U15590 ( .IN1(n9040), .IN2(g311), .Q(n14661) );
  OR2X1 U15591 ( .IN1(n14663), .IN2(n14664), .Q(g26881) );
  AND2X1 U15592 ( .IN1(n9146), .IN2(g305), .Q(n14664) );
  AND2X1 U15593 ( .IN1(g6744), .IN2(n9031), .Q(n14663) );
  INVX0 U15594 ( .INP(n14665), .ZN(g26877) );
  AND3X1 U15595 ( .IN1(n9057), .IN2(n9875), .IN3(n9874), .Q(n14665) );
  OR2X1 U15596 ( .IN1(n14666), .IN2(n14667), .Q(n9874) );
  OR4X1 U15597 ( .IN1(g2472), .IN2(g2204), .IN3(g2491), .IN4(g2223), .Q(n14667) );
  OR4X1 U15598 ( .IN1(g2338), .IN2(g2606), .IN3(test_so40), .IN4(g2357), .Q(
        n14666) );
  OR2X1 U15599 ( .IN1(n14668), .IN2(n14669), .Q(n9875) );
  OR4X1 U15600 ( .IN1(g2066), .IN2(g1798), .IN3(g1779), .IN4(g2047), .Q(n14669) );
  OR4X1 U15601 ( .IN1(g1913), .IN2(g1932), .IN3(test_so75), .IN4(g1664), .Q(
        n14668) );
  INVX0 U15602 ( .INP(n14670), .ZN(g26876) );
  AND3X1 U15603 ( .IN1(n9057), .IN2(n9895), .IN3(n9894), .Q(n14670) );
  OR2X1 U15604 ( .IN1(n14671), .IN2(n14672), .Q(n9894) );
  OR4X1 U15605 ( .IN1(n9324), .IN2(n9262), .IN3(n9295), .IN4(n9273), .Q(n14672) );
  OR4X1 U15606 ( .IN1(g2269), .IN2(g2537), .IN3(test_so31), .IN4(g2671), .Q(
        n14671) );
  OR2X1 U15607 ( .IN1(n14673), .IN2(n14674), .Q(n9895) );
  OR4X1 U15608 ( .IN1(g1858), .IN2(n9236), .IN3(g1992), .IN4(g2126), .Q(n14674) );
  OR4X1 U15609 ( .IN1(g1844), .IN2(g2112), .IN3(g1710), .IN4(g1978), .Q(n14673) );
  OR3X1 U15610 ( .IN1(n9121), .IN2(n9901), .IN3(n9900), .Q(g26875) );
  AND4X1 U15611 ( .IN1(n5414), .IN2(n5631), .IN3(n5281), .IN4(n5316), .Q(n9900) );
  AND4X1 U15612 ( .IN1(n5413), .IN2(n5628), .IN3(n5280), .IN4(n5315), .Q(n9901) );
  OR2X1 U15613 ( .IN1(n14675), .IN2(n14676), .Q(g25764) );
  AND2X1 U15614 ( .IN1(n14677), .IN2(g6541), .Q(n14676) );
  AND2X1 U15615 ( .IN1(n12080), .IN2(g6505), .Q(n14675) );
  OR3X1 U15616 ( .IN1(n14678), .IN2(n14679), .IN3(n14680), .Q(g25763) );
  AND2X1 U15617 ( .IN1(n12080), .IN2(g6537), .Q(n14680) );
  AND4X1 U15618 ( .IN1(n10979), .IN2(n9082), .IN3(n5659), .IN4(n5445), .Q(
        n14679) );
  AND2X1 U15619 ( .IN1(n14681), .IN2(g6533), .Q(n14678) );
  OR2X1 U15620 ( .IN1(n9129), .IN2(n14682), .Q(n14681) );
  AND2X1 U15621 ( .IN1(n10979), .IN2(g6527), .Q(n14682) );
  OR2X1 U15622 ( .IN1(n14683), .IN2(n14684), .Q(g25762) );
  AND2X1 U15623 ( .IN1(n14677), .IN2(g6527), .Q(n14684) );
  AND2X1 U15624 ( .IN1(n12080), .IN2(g6533), .Q(n14683) );
  OR3X1 U15625 ( .IN1(n14685), .IN2(n14686), .IN3(n14687), .Q(g25761) );
  AND2X1 U15626 ( .IN1(n12080), .IN2(g6513), .Q(n14687) );
  INVX0 U15627 ( .INP(n14677), .ZN(n12080) );
  OR2X1 U15628 ( .IN1(n9129), .IN2(n10979), .Q(n14677) );
  AND2X1 U15629 ( .IN1(n9146), .IN2(g6509), .Q(n14686) );
  AND3X1 U15630 ( .IN1(n5426), .IN2(n10979), .IN3(n9060), .Q(n14685) );
  AND2X1 U15631 ( .IN1(g6561), .IN2(n12098), .Q(n10979) );
  INVX0 U15632 ( .INP(n1422), .ZN(n12098) );
  OR2X1 U15633 ( .IN1(n5563), .IN2(n5386), .Q(n1422) );
  OR2X1 U15634 ( .IN1(n14688), .IN2(n14689), .Q(g25758) );
  AND3X1 U15635 ( .IN1(n8313), .IN2(n14690), .IN3(n9060), .Q(n14689) );
  OR2X1 U15636 ( .IN1(n14691), .IN2(g6444), .Q(n14690) );
  AND2X1 U15637 ( .IN1(n8314), .IN2(g9743), .Q(n14691) );
  AND2X1 U15638 ( .IN1(n9146), .IN2(g6494), .Q(n14688) );
  OR2X1 U15639 ( .IN1(n14692), .IN2(n14693), .Q(g25757) );
  AND2X1 U15640 ( .IN1(n9146), .IN2(g6444), .Q(n14693) );
  AND2X1 U15641 ( .IN1(n9040), .IN2(g6727), .Q(n14692) );
  AND2X1 U15642 ( .IN1(g6573), .IN2(n9031), .Q(g25756) );
  OR2X1 U15643 ( .IN1(n14694), .IN2(n14695), .Q(g25750) );
  AND2X1 U15644 ( .IN1(n14696), .IN2(g6195), .Q(n14695) );
  AND2X1 U15645 ( .IN1(n12167), .IN2(g6159), .Q(n14694) );
  OR3X1 U15646 ( .IN1(n14697), .IN2(n14698), .IN3(n14699), .Q(g25749) );
  AND2X1 U15647 ( .IN1(n12167), .IN2(g6191), .Q(n14699) );
  AND4X1 U15648 ( .IN1(n10991), .IN2(n9081), .IN3(n5667), .IN4(n5453), .Q(
        n14698) );
  AND2X1 U15649 ( .IN1(n14700), .IN2(g6187), .Q(n14697) );
  OR2X1 U15650 ( .IN1(n9128), .IN2(n14701), .Q(n14700) );
  AND2X1 U15651 ( .IN1(n10991), .IN2(g6181), .Q(n14701) );
  OR2X1 U15652 ( .IN1(n14702), .IN2(n14703), .Q(g25748) );
  AND2X1 U15653 ( .IN1(n14696), .IN2(g6181), .Q(n14703) );
  AND2X1 U15654 ( .IN1(n12167), .IN2(g6187), .Q(n14702) );
  OR3X1 U15655 ( .IN1(n14704), .IN2(n14705), .IN3(n14706), .Q(g25747) );
  AND2X1 U15656 ( .IN1(n12167), .IN2(g6167), .Q(n14706) );
  INVX0 U15657 ( .INP(n14696), .ZN(n12167) );
  OR2X1 U15658 ( .IN1(n9128), .IN2(n10991), .Q(n14696) );
  AND2X1 U15659 ( .IN1(n9146), .IN2(g6163), .Q(n14705) );
  AND3X1 U15660 ( .IN1(n5430), .IN2(n10991), .IN3(n9059), .Q(n14704) );
  AND2X1 U15661 ( .IN1(g6215), .IN2(n12185), .Q(n10991) );
  INVX0 U15662 ( .INP(n92), .ZN(n12185) );
  OR2X1 U15663 ( .IN1(n5568), .IN2(n5385), .Q(n92) );
  OR2X1 U15664 ( .IN1(n14707), .IN2(n14708), .Q(g25744) );
  AND3X1 U15665 ( .IN1(n8310), .IN2(n14709), .IN3(n9060), .Q(n14708) );
  OR2X1 U15666 ( .IN1(n14710), .IN2(g6098), .Q(n14709) );
  AND2X1 U15667 ( .IN1(test_so92), .IN2(n8311), .Q(n14710) );
  AND2X1 U15668 ( .IN1(n9146), .IN2(g6148), .Q(n14707) );
  OR2X1 U15669 ( .IN1(n14711), .IN2(n14712), .Q(g25743) );
  AND2X1 U15670 ( .IN1(n9146), .IN2(g6098), .Q(n14712) );
  AND2X1 U15671 ( .IN1(test_so69), .IN2(n9032), .Q(n14711) );
  AND2X1 U15672 ( .IN1(g6227), .IN2(n9031), .Q(g25742) );
  OR2X1 U15673 ( .IN1(n14713), .IN2(n14714), .Q(g25736) );
  AND2X1 U15674 ( .IN1(n14715), .IN2(g5849), .Q(n14714) );
  AND2X1 U15675 ( .IN1(n12253), .IN2(g5813), .Q(n14713) );
  OR3X1 U15676 ( .IN1(n14716), .IN2(n14717), .IN3(n14718), .Q(g25735) );
  AND2X1 U15677 ( .IN1(test_so83), .IN2(n12253), .Q(n14718) );
  AND4X1 U15678 ( .IN1(n10990), .IN2(n9081), .IN3(n5663), .IN4(n5449), .Q(
        n14717) );
  AND2X1 U15679 ( .IN1(n14719), .IN2(g5841), .Q(n14716) );
  OR2X1 U15680 ( .IN1(n9128), .IN2(n14720), .Q(n14719) );
  AND2X1 U15681 ( .IN1(n10990), .IN2(g5835), .Q(n14720) );
  OR2X1 U15682 ( .IN1(n14721), .IN2(n14722), .Q(g25734) );
  AND2X1 U15683 ( .IN1(n14715), .IN2(g5835), .Q(n14722) );
  AND2X1 U15684 ( .IN1(n12253), .IN2(g5841), .Q(n14721) );
  OR3X1 U15685 ( .IN1(n14723), .IN2(n14724), .IN3(n14725), .Q(g25733) );
  AND2X1 U15686 ( .IN1(n12253), .IN2(g5821), .Q(n14725) );
  INVX0 U15687 ( .INP(n14715), .ZN(n12253) );
  OR2X1 U15688 ( .IN1(n9128), .IN2(n10990), .Q(n14715) );
  AND2X1 U15689 ( .IN1(n9146), .IN2(g5817), .Q(n14724) );
  AND3X1 U15690 ( .IN1(n5429), .IN2(n10990), .IN3(n9060), .Q(n14723) );
  AND2X1 U15691 ( .IN1(g5869), .IN2(n12271), .Q(n10990) );
  INVX0 U15692 ( .INP(n735), .ZN(n12271) );
  OR2X1 U15693 ( .IN1(n5388), .IN2(n8832), .Q(n735) );
  OR2X1 U15694 ( .IN1(n14726), .IN2(n14727), .Q(g25730) );
  AND3X1 U15695 ( .IN1(n8321), .IN2(n14728), .IN3(n9059), .Q(n14727) );
  OR2X1 U15696 ( .IN1(n14729), .IN2(g5752), .Q(n14728) );
  AND2X1 U15697 ( .IN1(n8322), .IN2(g9617), .Q(n14729) );
  AND2X1 U15698 ( .IN1(n9146), .IN2(g5802), .Q(n14726) );
  OR2X1 U15699 ( .IN1(n14730), .IN2(n14731), .Q(g25729) );
  AND2X1 U15700 ( .IN1(n9146), .IN2(g5752), .Q(n14731) );
  AND2X1 U15701 ( .IN1(n9040), .IN2(g6035), .Q(n14730) );
  AND2X1 U15702 ( .IN1(n9040), .IN2(test_so36), .Q(g25728) );
  OR2X1 U15703 ( .IN1(n14732), .IN2(n14733), .Q(g25722) );
  AND2X1 U15704 ( .IN1(n14734), .IN2(g5503), .Q(n14733) );
  AND2X1 U15705 ( .IN1(n12338), .IN2(g5467), .Q(n14732) );
  OR3X1 U15706 ( .IN1(n14735), .IN2(n14736), .IN3(n14737), .Q(g25721) );
  AND2X1 U15707 ( .IN1(n12338), .IN2(g5499), .Q(n14737) );
  AND4X1 U15708 ( .IN1(n10987), .IN2(n9081), .IN3(n5660), .IN4(n5446), .Q(
        n14736) );
  AND2X1 U15709 ( .IN1(n14738), .IN2(g5495), .Q(n14735) );
  OR2X1 U15710 ( .IN1(n9128), .IN2(n14739), .Q(n14738) );
  AND2X1 U15711 ( .IN1(n10987), .IN2(g5489), .Q(n14739) );
  OR2X1 U15712 ( .IN1(n14740), .IN2(n14741), .Q(g25720) );
  AND2X1 U15713 ( .IN1(n14734), .IN2(g5489), .Q(n14741) );
  AND2X1 U15714 ( .IN1(n12338), .IN2(g5495), .Q(n14740) );
  OR3X1 U15715 ( .IN1(n14742), .IN2(n14743), .IN3(n14744), .Q(g25719) );
  AND2X1 U15716 ( .IN1(n12338), .IN2(g5475), .Q(n14744) );
  INVX0 U15717 ( .INP(n14734), .ZN(n12338) );
  OR2X1 U15718 ( .IN1(n9127), .IN2(n10987), .Q(n14734) );
  AND2X1 U15719 ( .IN1(n9146), .IN2(g5471), .Q(n14743) );
  AND3X1 U15720 ( .IN1(n5425), .IN2(n10987), .IN3(n9061), .Q(n14742) );
  AND2X1 U15721 ( .IN1(g5523), .IN2(n12356), .Q(n10987) );
  INVX0 U15722 ( .INP(n945), .ZN(n12356) );
  OR2X1 U15723 ( .IN1(n5566), .IN2(n5389), .Q(n945) );
  OR2X1 U15724 ( .IN1(n14745), .IN2(n14746), .Q(g25716) );
  AND3X1 U15725 ( .IN1(n14747), .IN2(n8315), .IN3(n9059), .Q(n14746) );
  OR2X1 U15726 ( .IN1(n14748), .IN2(g5406), .Q(n14747) );
  AND2X1 U15727 ( .IN1(n8316), .IN2(g9555), .Q(n14748) );
  AND2X1 U15728 ( .IN1(n9147), .IN2(g5456), .Q(n14745) );
  OR2X1 U15729 ( .IN1(n14749), .IN2(n14750), .Q(g25715) );
  AND2X1 U15730 ( .IN1(n9147), .IN2(g5406), .Q(n14750) );
  AND2X1 U15731 ( .IN1(n9045), .IN2(g5689), .Q(n14749) );
  AND2X1 U15732 ( .IN1(g5535), .IN2(n9031), .Q(g25714) );
  OR2X1 U15733 ( .IN1(n14751), .IN2(n14752), .Q(g25708) );
  AND2X1 U15734 ( .IN1(n14753), .IN2(g5156), .Q(n14752) );
  AND2X1 U15735 ( .IN1(n9490), .IN2(g5120), .Q(n14751) );
  OR2X1 U15736 ( .IN1(n14754), .IN2(n14755), .Q(g25706) );
  AND2X1 U15737 ( .IN1(n14753), .IN2(g5142), .Q(n14755) );
  AND2X1 U15738 ( .IN1(test_so98), .IN2(n9490), .Q(n14754) );
  OR3X1 U15739 ( .IN1(n14756), .IN2(n14757), .IN3(n14758), .Q(g25705) );
  AND2X1 U15740 ( .IN1(test_so96), .IN2(n9490), .Q(n14758) );
  INVX0 U15741 ( .INP(n14753), .ZN(n9490) );
  OR2X1 U15742 ( .IN1(n9127), .IN2(g32975), .Q(n14753) );
  AND2X1 U15743 ( .IN1(n9147), .IN2(g5124), .Q(n14757) );
  AND3X1 U15744 ( .IN1(g32975), .IN2(n8848), .IN3(n9058), .Q(n14756) );
  AND2X1 U15745 ( .IN1(g5176), .IN2(n12441), .Q(g32975) );
  INVX0 U15746 ( .INP(n231), .ZN(n12441) );
  OR2X1 U15747 ( .IN1(n5567), .IN2(n5384), .Q(n231) );
  AND2X1 U15748 ( .IN1(n14759), .IN2(g5073), .Q(g25704) );
  OR2X1 U15749 ( .IN1(n9127), .IN2(g5069), .Q(n14759) );
  OR2X1 U15750 ( .IN1(n14760), .IN2(n14761), .Q(g25703) );
  AND3X1 U15751 ( .IN1(n5689), .IN2(n14762), .IN3(n9059), .Q(n14761) );
  INVX0 U15752 ( .INP(n14763), .ZN(n14762) );
  AND2X1 U15753 ( .IN1(n14764), .IN2(n8767), .Q(n14763) );
  OR2X1 U15754 ( .IN1(g5112), .IN2(n5690), .Q(n14764) );
  AND2X1 U15755 ( .IN1(n9147), .IN2(g5112), .Q(n14760) );
  OR2X1 U15756 ( .IN1(n14765), .IN2(n14766), .Q(g25702) );
  AND3X1 U15757 ( .IN1(n5690), .IN2(n14767), .IN3(n9061), .Q(n14766) );
  OR2X1 U15758 ( .IN1(n14768), .IN2(g5062), .Q(n14767) );
  INVX0 U15759 ( .INP(n14769), .ZN(n14768) );
  OR2X1 U15760 ( .IN1(n5689), .IN2(test_so32), .Q(n14769) );
  AND2X1 U15761 ( .IN1(test_so32), .IN2(n9139), .Q(n14765) );
  OR2X1 U15762 ( .IN1(n14770), .IN2(n14771), .Q(g25701) );
  AND2X1 U15763 ( .IN1(n9147), .IN2(g5062), .Q(n14771) );
  AND2X1 U15764 ( .IN1(test_so10), .IN2(n9030), .Q(n14770) );
  AND2X1 U15765 ( .IN1(g5188), .IN2(n9030), .Q(g25700) );
  OR3X1 U15766 ( .IN1(n14772), .IN2(n14773), .IN3(n14774), .Q(g25699) );
  AND2X1 U15767 ( .IN1(n9147), .IN2(g5097), .Q(n14774) );
  AND2X1 U15768 ( .IN1(n5014), .IN2(n5669), .Q(n14773) );
  INVX0 U15769 ( .INP(n14775), .ZN(n14772) );
  OR3X1 U15770 ( .IN1(n9121), .IN2(n5014), .IN3(n5669), .Q(n14775) );
  OR3X1 U15771 ( .IN1(n14776), .IN2(n14777), .IN3(n14778), .Q(g25698) );
  AND2X1 U15772 ( .IN1(n9147), .IN2(g5092), .Q(n14778) );
  AND2X1 U15773 ( .IN1(n5016), .IN2(n5753), .Q(n14777) );
  AND3X1 U15774 ( .IN1(n9056), .IN2(n14779), .IN3(g5097), .Q(n14776) );
  INVX0 U15775 ( .INP(n5016), .ZN(n14779) );
  AND2X1 U15776 ( .IN1(n14780), .IN2(n14781), .Q(g25697) );
  INVX0 U15777 ( .INP(n14782), .ZN(n14781) );
  AND2X1 U15778 ( .IN1(n14783), .IN2(n5681), .Q(n14782) );
  OR2X1 U15779 ( .IN1(n5681), .IN2(n14783), .Q(n14780) );
  OR2X1 U15780 ( .IN1(n8697), .IN2(n9123), .Q(n14783) );
  OR3X1 U15781 ( .IN1(n14784), .IN2(n14785), .IN3(n14786), .Q(g25696) );
  AND3X1 U15782 ( .IN1(n9056), .IN2(g5077), .IN3(n8722), .Q(n14786) );
  AND3X1 U15783 ( .IN1(n14787), .IN2(n14788), .IN3(n5893), .Q(n14785) );
  OR2X1 U15784 ( .IN1(n5455), .IN2(g5069), .Q(n14788) );
  INVX0 U15785 ( .INP(n14789), .ZN(n14784) );
  OR2X1 U15786 ( .IN1(n14787), .IN2(n5893), .Q(n14789) );
  AND2X1 U15787 ( .IN1(n9040), .IN2(n5681), .Q(n14787) );
  AND2X1 U15788 ( .IN1(n14790), .IN2(g5077), .Q(g25695) );
  OR3X1 U15789 ( .IN1(n14791), .IN2(n14792), .IN3(n9122), .Q(n14790) );
  AND2X1 U15790 ( .IN1(n8722), .IN2(n5681), .Q(n14792) );
  AND2X1 U15791 ( .IN1(n8344), .IN2(g5084), .Q(n14791) );
  OR2X1 U15792 ( .IN1(n14793), .IN2(n14794), .Q(g25691) );
  AND2X1 U15793 ( .IN1(n9147), .IN2(g4125), .Q(n14794) );
  AND2X1 U15794 ( .IN1(n8811), .IN2(n14795), .Q(n14793) );
  OR4X1 U15795 ( .IN1(n8825), .IN2(g4064), .IN3(g4057), .IN4(n14796), .Q(
        n14795) );
  OR4X1 U15796 ( .IN1(g4141), .IN2(g4082), .IN3(n5350), .IN4(n12420), .Q(
        n14796) );
  INVX0 U15797 ( .INP(n10978), .ZN(n12420) );
  AND2X1 U15798 ( .IN1(g4087), .IN2(n5340), .Q(n10978) );
  OR2X1 U15799 ( .IN1(n14797), .IN2(n14798), .Q(g25690) );
  AND3X1 U15800 ( .IN1(n8555), .IN2(g25689), .IN3(n9061), .Q(n14798) );
  AND2X1 U15801 ( .IN1(n9147), .IN2(g4169), .Q(n14797) );
  OR3X1 U15802 ( .IN1(n14799), .IN2(n14800), .IN3(n14801), .Q(g25687) );
  AND2X1 U15803 ( .IN1(n9147), .IN2(g4057), .Q(n14801) );
  AND2X1 U15804 ( .IN1(n5026), .IN2(n12527), .Q(n14800) );
  AND3X1 U15805 ( .IN1(n14450), .IN2(g4169), .IN3(n5612), .Q(n14799) );
  INVX0 U15806 ( .INP(n1253), .ZN(n14450) );
  OR2X1 U15807 ( .IN1(n5416), .IN2(n5711), .Q(n1253) );
  OR2X1 U15808 ( .IN1(n14802), .IN2(n14803), .Q(g25686) );
  AND3X1 U15809 ( .IN1(n12527), .IN2(g4057), .IN3(n5416), .Q(n14803) );
  AND2X1 U15810 ( .IN1(g4169), .IN2(n9029), .Q(n12527) );
  AND2X1 U15811 ( .IN1(n14804), .IN2(g4064), .Q(n14802) );
  OR2X1 U15812 ( .IN1(n9126), .IN2(n14805), .Q(n14804) );
  AND2X1 U15813 ( .IN1(n5711), .IN2(g4169), .Q(n14805) );
  OR3X1 U15814 ( .IN1(n14806), .IN2(n14807), .IN3(n8811), .Q(g25685) );
  AND2X1 U15815 ( .IN1(n9040), .IN2(n5729), .Q(n8811) );
  AND2X1 U15816 ( .IN1(n9147), .IN2(g4072), .Q(n14807) );
  AND2X1 U15817 ( .IN1(n5416), .IN2(n9029), .Q(n14806) );
  OR2X1 U15818 ( .IN1(n14808), .IN2(n14809), .Q(g25684) );
  AND2X1 U15819 ( .IN1(n14810), .IN2(g3849), .Q(n14809) );
  AND2X1 U15820 ( .IN1(n9375), .IN2(g3813), .Q(n14808) );
  OR2X1 U15821 ( .IN1(n14811), .IN2(n14812), .Q(g25682) );
  AND2X1 U15822 ( .IN1(n14810), .IN2(g3835), .Q(n14812) );
  AND2X1 U15823 ( .IN1(test_so97), .IN2(n9375), .Q(n14811) );
  OR3X1 U15824 ( .IN1(n14813), .IN2(n14814), .IN3(n14815), .Q(g25681) );
  AND2X1 U15825 ( .IN1(n9375), .IN2(g3821), .Q(n14815) );
  INVX0 U15826 ( .INP(n14810), .ZN(n9375) );
  OR2X1 U15827 ( .IN1(n9126), .IN2(n9376), .Q(n14810) );
  AND2X1 U15828 ( .IN1(n9148), .IN2(g3817), .Q(n14814) );
  AND3X1 U15829 ( .IN1(n5428), .IN2(n9376), .IN3(n9064), .Q(n14813) );
  AND2X1 U15830 ( .IN1(n12549), .IN2(test_so33), .Q(n9376) );
  INVX0 U15831 ( .INP(n843), .ZN(n12549) );
  OR2X1 U15832 ( .IN1(n5564), .IN2(n5387), .Q(n843) );
  OR2X1 U15833 ( .IN1(n14816), .IN2(n14817), .Q(g25678) );
  AND3X1 U15834 ( .IN1(n8317), .IN2(n14818), .IN3(n9065), .Q(n14817) );
  OR2X1 U15835 ( .IN1(n14819), .IN2(g3752), .Q(n14818) );
  AND2X1 U15836 ( .IN1(n8318), .IN2(g8344), .Q(n14819) );
  AND2X1 U15837 ( .IN1(n9148), .IN2(g3802), .Q(n14816) );
  OR2X1 U15838 ( .IN1(n14820), .IN2(n14821), .Q(g25677) );
  AND2X1 U15839 ( .IN1(n9148), .IN2(g3752), .Q(n14821) );
  AND2X1 U15840 ( .IN1(n9041), .IN2(g4040), .Q(n14820) );
  AND2X1 U15841 ( .IN1(g3881), .IN2(n9028), .Q(g25676) );
  OR2X1 U15842 ( .IN1(n14822), .IN2(n14823), .Q(g25670) );
  AND2X1 U15843 ( .IN1(n14824), .IN2(g3498), .Q(n14823) );
  AND2X1 U15844 ( .IN1(n12616), .IN2(g3462), .Q(n14822) );
  OR3X1 U15845 ( .IN1(n14825), .IN2(n14826), .IN3(n14827), .Q(g25669) );
  AND2X1 U15846 ( .IN1(n12616), .IN2(g3494), .Q(n14827) );
  AND4X1 U15847 ( .IN1(n10982), .IN2(n9081), .IN3(n5668), .IN4(n5454), .Q(
        n14826) );
  AND2X1 U15848 ( .IN1(n14828), .IN2(g3490), .Q(n14825) );
  OR2X1 U15849 ( .IN1(n9126), .IN2(n14829), .Q(n14828) );
  AND2X1 U15850 ( .IN1(n10982), .IN2(g3484), .Q(n14829) );
  OR2X1 U15851 ( .IN1(n14830), .IN2(n14831), .Q(g25668) );
  AND2X1 U15852 ( .IN1(n14824), .IN2(g3484), .Q(n14831) );
  AND2X1 U15853 ( .IN1(n12616), .IN2(g3490), .Q(n14830) );
  OR3X1 U15854 ( .IN1(n14832), .IN2(n14833), .IN3(n14834), .Q(g25667) );
  AND2X1 U15855 ( .IN1(n12616), .IN2(g3470), .Q(n14834) );
  INVX0 U15856 ( .INP(n14824), .ZN(n12616) );
  OR2X1 U15857 ( .IN1(n9125), .IN2(n10982), .Q(n14824) );
  INVX0 U15858 ( .INP(n14835), .ZN(n14833) );
  OR2X1 U15859 ( .IN1(n9008), .IN2(n8760), .Q(n14835) );
  AND3X1 U15860 ( .IN1(n5424), .IN2(n10982), .IN3(n9065), .Q(n14832) );
  AND2X1 U15861 ( .IN1(g3518), .IN2(n12634), .Q(n10982) );
  INVX0 U15862 ( .INP(n470), .ZN(n12634) );
  OR2X1 U15863 ( .IN1(n5569), .IN2(n5383), .Q(n470) );
  OR2X1 U15864 ( .IN1(n14836), .IN2(n14837), .Q(g25664) );
  AND3X1 U15865 ( .IN1(n8301), .IN2(n14838), .IN3(n9065), .Q(n14837) );
  OR2X1 U15866 ( .IN1(n14839), .IN2(g3401), .Q(n14838) );
  AND2X1 U15867 ( .IN1(n8302), .IN2(g8279), .Q(n14839) );
  AND2X1 U15868 ( .IN1(n9148), .IN2(g3451), .Q(n14836) );
  OR2X1 U15869 ( .IN1(n14840), .IN2(n14841), .Q(g25663) );
  AND2X1 U15870 ( .IN1(n9148), .IN2(g3401), .Q(n14841) );
  AND2X1 U15871 ( .IN1(n9041), .IN2(g3689), .Q(n14840) );
  AND2X1 U15872 ( .IN1(g3530), .IN2(n9028), .Q(g25662) );
  OR2X1 U15873 ( .IN1(n14842), .IN2(n14843), .Q(g25656) );
  AND2X1 U15874 ( .IN1(n14844), .IN2(g3147), .Q(n14843) );
  AND2X1 U15875 ( .IN1(n12701), .IN2(g3111), .Q(n14842) );
  OR3X1 U15876 ( .IN1(n14845), .IN2(n14846), .IN3(n14847), .Q(g25655) );
  INVX0 U15877 ( .INP(n14848), .ZN(n14847) );
  OR2X1 U15878 ( .IN1(n14844), .IN2(n5882), .Q(n14848) );
  AND4X1 U15879 ( .IN1(n10977), .IN2(n9080), .IN3(n5661), .IN4(n5447), .Q(
        n14846) );
  AND2X1 U15880 ( .IN1(n14849), .IN2(g3139), .Q(n14845) );
  OR2X1 U15881 ( .IN1(n9125), .IN2(n14850), .Q(n14849) );
  AND2X1 U15882 ( .IN1(n10977), .IN2(g3133), .Q(n14850) );
  OR2X1 U15883 ( .IN1(n14851), .IN2(n14852), .Q(g25654) );
  AND2X1 U15884 ( .IN1(n14844), .IN2(g3133), .Q(n14852) );
  AND2X1 U15885 ( .IN1(n12701), .IN2(g3139), .Q(n14851) );
  OR3X1 U15886 ( .IN1(n14853), .IN2(n14854), .IN3(n14855), .Q(g25653) );
  AND2X1 U15887 ( .IN1(n12701), .IN2(g3119), .Q(n14855) );
  INVX0 U15888 ( .INP(n14844), .ZN(n12701) );
  OR2X1 U15889 ( .IN1(n9125), .IN2(n10977), .Q(n14844) );
  AND2X1 U15890 ( .IN1(n9148), .IN2(g3115), .Q(n14854) );
  AND3X1 U15891 ( .IN1(n5423), .IN2(n10977), .IN3(n9065), .Q(n14853) );
  AND2X1 U15892 ( .IN1(g3167), .IN2(n12719), .Q(n10977) );
  INVX0 U15893 ( .INP(n563), .ZN(n12719) );
  OR2X1 U15894 ( .IN1(n5603), .IN2(n5390), .Q(n563) );
  OR2X1 U15895 ( .IN1(n14856), .IN2(n14857), .Q(g25650) );
  AND3X1 U15896 ( .IN1(n8323), .IN2(n14858), .IN3(n9065), .Q(n14857) );
  OR2X1 U15897 ( .IN1(n14859), .IN2(g3050), .Q(n14858) );
  AND2X1 U15898 ( .IN1(n8324), .IN2(g8215), .Q(n14859) );
  AND2X1 U15899 ( .IN1(n9148), .IN2(g3100), .Q(n14856) );
  OR2X1 U15900 ( .IN1(n14860), .IN2(n14861), .Q(g25649) );
  AND2X1 U15901 ( .IN1(n9148), .IN2(g3050), .Q(n14861) );
  AND2X1 U15902 ( .IN1(n9041), .IN2(g3338), .Q(n14860) );
  AND2X1 U15903 ( .IN1(g3179), .IN2(n9027), .Q(g25648) );
  OR3X1 U15904 ( .IN1(n14862), .IN2(n14863), .IN3(n5045), .Q(g25639) );
  AND2X1 U15905 ( .IN1(n13558), .IN2(n9027), .Q(n14863) );
  AND2X1 U15906 ( .IN1(g2719), .IN2(n5299), .Q(n13558) );
  AND2X1 U15907 ( .IN1(n9148), .IN2(g2715), .Q(n14862) );
  OR2X1 U15908 ( .IN1(n14864), .IN2(n14865), .Q(g25638) );
  AND2X1 U15909 ( .IN1(n14866), .IN2(n9027), .Q(n14865) );
  OR2X1 U15910 ( .IN1(n14867), .IN2(n14868), .Q(n14866) );
  AND3X1 U15911 ( .IN1(n14869), .IN2(n5768), .IN3(n5441), .Q(n14868) );
  AND2X1 U15912 ( .IN1(n14870), .IN2(g1559), .Q(n14867) );
  AND2X1 U15913 ( .IN1(n9148), .IN2(g1564), .Q(n14864) );
  OR2X1 U15914 ( .IN1(n14871), .IN2(n14872), .Q(g25637) );
  AND2X1 U15915 ( .IN1(n14873), .IN2(g1559), .Q(n14872) );
  OR2X1 U15916 ( .IN1(n9124), .IN2(n14874), .Q(n14873) );
  AND2X1 U15917 ( .IN1(n14869), .IN2(n5768), .Q(n14874) );
  INVX0 U15918 ( .INP(n14870), .ZN(n14869) );
  AND3X1 U15919 ( .IN1(n9055), .IN2(g1554), .IN3(n14870), .Q(n14871) );
  OR2X1 U15920 ( .IN1(n14875), .IN2(n14876), .Q(g25636) );
  AND2X1 U15921 ( .IN1(n14877), .IN2(n9027), .Q(n14876) );
  OR2X1 U15922 ( .IN1(n14878), .IN2(n14879), .Q(n14877) );
  AND2X1 U15923 ( .IN1(n14880), .IN2(g1306), .Q(n14879) );
  INVX0 U15924 ( .INP(n14881), .ZN(n14880) );
  AND2X1 U15925 ( .IN1(n14881), .IN2(g1339), .Q(n14878) );
  AND2X1 U15926 ( .IN1(g7946), .IN2(n11216), .Q(n14881) );
  INVX0 U15927 ( .INP(n13627), .ZN(n11216) );
  OR2X1 U15928 ( .IN1(n5364), .IN2(n8819), .Q(n13627) );
  AND2X1 U15929 ( .IN1(n9148), .IN2(g1521), .Q(n14875) );
  OR2X1 U15930 ( .IN1(n14882), .IN2(n14883), .Q(g25635) );
  AND2X1 U15931 ( .IN1(n14884), .IN2(g1300), .Q(n14883) );
  OR2X1 U15932 ( .IN1(n14885), .IN2(n13616), .Q(n14884) );
  AND2X1 U15933 ( .IN1(n14886), .IN2(n9027), .Q(n14885) );
  OR2X1 U15934 ( .IN1(n5865), .IN2(n14500), .Q(n14886) );
  AND2X1 U15935 ( .IN1(n14887), .IN2(g1484), .Q(n14882) );
  OR2X1 U15936 ( .IN1(n9125), .IN2(n14888), .Q(n14887) );
  AND3X1 U15937 ( .IN1(n13621), .IN2(n5483), .IN3(n14889), .Q(n14888) );
  INVX0 U15938 ( .INP(n14500), .ZN(n14889) );
  OR2X1 U15939 ( .IN1(n8551), .IN2(test_so12), .Q(n14500) );
  AND3X1 U15940 ( .IN1(n14506), .IN2(n8824), .IN3(n14890), .Q(g25634) );
  OR2X1 U15941 ( .IN1(n14891), .IN2(n14892), .Q(n14890) );
  AND2X1 U15942 ( .IN1(n9042), .IN2(g1395), .Q(n14892) );
  AND2X1 U15943 ( .IN1(n11485), .IN2(n14893), .Q(n14891) );
  INVX0 U15944 ( .INP(n14505), .ZN(n14506) );
  AND3X1 U15945 ( .IN1(g1395), .IN2(g12923), .IN3(n14893), .Q(n14505) );
  INVX0 U15946 ( .INP(n14894), .ZN(n14893) );
  OR3X1 U15947 ( .IN1(n14895), .IN2(n14896), .IN3(n14897), .Q(g25633) );
  AND3X1 U15948 ( .IN1(n14898), .IN2(n8764), .IN3(n14510), .Q(n14897) );
  AND2X1 U15949 ( .IN1(n9148), .IN2(g1379), .Q(n14896) );
  AND3X1 U15950 ( .IN1(n14512), .IN2(g1384), .IN3(n9058), .Q(n14895) );
  OR2X1 U15951 ( .IN1(n14899), .IN2(n14900), .Q(g25632) );
  AND3X1 U15952 ( .IN1(n14901), .IN2(n14902), .IN3(n14510), .Q(n14900) );
  AND2X1 U15953 ( .IN1(g1351), .IN2(n9027), .Q(n14510) );
  OR2X1 U15954 ( .IN1(n13089), .IN2(n14903), .Q(n14902) );
  OR2X1 U15955 ( .IN1(n8655), .IN2(n14512), .Q(n14901) );
  AND2X1 U15956 ( .IN1(n14904), .IN2(g1312), .Q(n14899) );
  OR2X1 U15957 ( .IN1(n9125), .IN2(n14898), .Q(n14904) );
  AND2X1 U15958 ( .IN1(n14905), .IN2(n9027), .Q(g25631) );
  OR2X1 U15959 ( .IN1(n14906), .IN2(n14907), .Q(n14905) );
  AND2X1 U15960 ( .IN1(n14512), .IN2(g1312), .Q(n14907) );
  AND3X1 U15961 ( .IN1(n14908), .IN2(n14909), .IN3(n14228), .Q(n14906) );
  INVX0 U15962 ( .INP(n13089), .ZN(n14228) );
  OR2X1 U15963 ( .IN1(n9380), .IN2(g1351), .Q(n14909) );
  AND4X1 U15964 ( .IN1(g1379), .IN2(n14234), .IN3(g1345), .IN4(g1367), .Q(
        n9380) );
  OR2X1 U15965 ( .IN1(n5322), .IN2(n14910), .Q(n14908) );
  AND2X1 U15966 ( .IN1(n14233), .IN2(n14229), .Q(n14910) );
  OR2X1 U15967 ( .IN1(n8655), .IN2(n14234), .Q(n14229) );
  INVX0 U15968 ( .INP(n14903), .ZN(n14233) );
  OR2X1 U15969 ( .IN1(n8657), .IN2(n8654), .Q(n14903) );
  OR2X1 U15970 ( .IN1(n14911), .IN2(n14912), .Q(g25630) );
  AND2X1 U15971 ( .IN1(g24247), .IN2(g1266), .Q(n14912) );
  AND2X1 U15972 ( .IN1(n14913), .IN2(g1249), .Q(n14911) );
  OR2X1 U15973 ( .IN1(n9124), .IN2(n14914), .Q(n14913) );
  AND2X1 U15974 ( .IN1(n8369), .IN2(g12923), .Q(n14914) );
  OR2X1 U15975 ( .IN1(n14915), .IN2(n14916), .Q(g25629) );
  AND2X1 U15976 ( .IN1(n14917), .IN2(n9026), .Q(n14916) );
  OR2X1 U15977 ( .IN1(n14918), .IN2(n14919), .Q(n14917) );
  AND3X1 U15978 ( .IN1(n14920), .IN2(n8839), .IN3(n5442), .Q(n14919) );
  AND2X1 U15979 ( .IN1(n14921), .IN2(g1216), .Q(n14918) );
  AND2X1 U15980 ( .IN1(n9149), .IN2(g1221), .Q(n14915) );
  OR2X1 U15981 ( .IN1(n14922), .IN2(n14923), .Q(g25628) );
  AND2X1 U15982 ( .IN1(n14924), .IN2(g1216), .Q(n14923) );
  OR2X1 U15983 ( .IN1(n9124), .IN2(n14925), .Q(n14924) );
  AND2X1 U15984 ( .IN1(n14920), .IN2(n8839), .Q(n14925) );
  AND3X1 U15985 ( .IN1(n14921), .IN2(n9053), .IN3(test_so76), .Q(n14922) );
  OR2X1 U15986 ( .IN1(n14926), .IN2(n14927), .Q(g25627) );
  AND2X1 U15987 ( .IN1(n14928), .IN2(n9026), .Q(n14927) );
  OR2X1 U15988 ( .IN1(n14929), .IN2(n14930), .Q(n14928) );
  AND2X1 U15989 ( .IN1(n14931), .IN2(g962), .Q(n14930) );
  INVX0 U15990 ( .INP(n14932), .ZN(n14931) );
  AND2X1 U15991 ( .IN1(n14932), .IN2(g996), .Q(n14929) );
  AND2X1 U15992 ( .IN1(g7916), .IN2(n11387), .Q(n14932) );
  AND2X1 U15993 ( .IN1(g1183), .IN2(g1171), .Q(n11387) );
  AND2X1 U15994 ( .IN1(n9149), .IN2(g1178), .Q(n14926) );
  OR2X1 U15995 ( .IN1(n14933), .IN2(n14934), .Q(g25626) );
  AND2X1 U15996 ( .IN1(n14935), .IN2(g956), .Q(n14934) );
  OR2X1 U15997 ( .IN1(n14936), .IN2(n13659), .Q(n14935) );
  AND2X1 U15998 ( .IN1(n14937), .IN2(n9026), .Q(n14936) );
  OR2X1 U15999 ( .IN1(n5691), .IN2(n14532), .Q(n14937) );
  AND2X1 U16000 ( .IN1(n14938), .IN2(g1141), .Q(n14933) );
  OR2X1 U16001 ( .IN1(n9124), .IN2(n14939), .Q(n14938) );
  AND3X1 U16002 ( .IN1(n13664), .IN2(n5341), .IN3(n14538), .Q(n14939) );
  INVX0 U16003 ( .INP(n14532), .ZN(n14538) );
  OR2X1 U16004 ( .IN1(n8820), .IN2(g1152), .Q(n14532) );
  AND3X1 U16005 ( .IN1(n14940), .IN2(n14544), .IN3(n5320), .Q(g25625) );
  INVX0 U16006 ( .INP(n14543), .ZN(n14544) );
  AND3X1 U16007 ( .IN1(g1052), .IN2(g12919), .IN3(n14941), .Q(n14543) );
  OR2X1 U16008 ( .IN1(n14942), .IN2(n14943), .Q(n14940) );
  AND2X1 U16009 ( .IN1(n9042), .IN2(g1052), .Q(n14943) );
  AND2X1 U16010 ( .IN1(n11500), .IN2(n14941), .Q(n14942) );
  INVX0 U16011 ( .INP(n14944), .ZN(n14941) );
  OR3X1 U16012 ( .IN1(n14945), .IN2(n14946), .IN3(n14947), .Q(g25624) );
  AND3X1 U16013 ( .IN1(n14948), .IN2(n8765), .IN3(n14548), .Q(n14947) );
  AND2X1 U16014 ( .IN1(n9149), .IN2(g1036), .Q(n14946) );
  AND3X1 U16015 ( .IN1(n14550), .IN2(g1041), .IN3(n9065), .Q(n14945) );
  OR2X1 U16016 ( .IN1(n14949), .IN2(n14950), .Q(g25623) );
  AND3X1 U16017 ( .IN1(n14951), .IN2(n14952), .IN3(n14548), .Q(n14950) );
  AND2X1 U16018 ( .IN1(g1008), .IN2(n9026), .Q(n14548) );
  OR2X1 U16019 ( .IN1(n13124), .IN2(n14953), .Q(n14952) );
  OR2X1 U16020 ( .IN1(n8572), .IN2(n14550), .Q(n14951) );
  AND2X1 U16021 ( .IN1(test_so20), .IN2(n14954), .Q(n14949) );
  OR2X1 U16022 ( .IN1(n9124), .IN2(n14948), .Q(n14954) );
  INVX0 U16023 ( .INP(n14550), .ZN(n14948) );
  AND2X1 U16024 ( .IN1(n14955), .IN2(n9026), .Q(g25622) );
  OR2X1 U16025 ( .IN1(n14956), .IN2(n14957), .Q(n14955) );
  AND2X1 U16026 ( .IN1(test_so20), .IN2(n14550), .Q(n14957) );
  AND3X1 U16027 ( .IN1(n14958), .IN2(n14959), .IN3(n14242), .Q(n14956) );
  INVX0 U16028 ( .INP(n13124), .ZN(n14242) );
  OR2X1 U16029 ( .IN1(n9379), .IN2(g1008), .Q(n14959) );
  AND4X1 U16030 ( .IN1(g1036), .IN2(n14249), .IN3(g1002), .IN4(g1024), .Q(
        n9379) );
  OR2X1 U16031 ( .IN1(n5321), .IN2(n14960), .Q(n14958) );
  AND2X1 U16032 ( .IN1(n14248), .IN2(n14250), .Q(n14960) );
  OR2X1 U16033 ( .IN1(n8572), .IN2(n14249), .Q(n14250) );
  INVX0 U16034 ( .INP(n14953), .ZN(n14248) );
  OR2X1 U16035 ( .IN1(n8656), .IN2(n8653), .Q(n14953) );
  OR2X1 U16036 ( .IN1(n14961), .IN2(n14962), .Q(g25621) );
  AND2X1 U16037 ( .IN1(g24231), .IN2(g921), .Q(n14962) );
  AND2X1 U16038 ( .IN1(n14963), .IN2(g904), .Q(n14961) );
  OR2X1 U16039 ( .IN1(n9124), .IN2(n14964), .Q(n14963) );
  AND2X1 U16040 ( .IN1(n8368), .IN2(g12919), .Q(n14964) );
  AND2X1 U16041 ( .IN1(n14965), .IN2(g837), .Q(g25619) );
  OR2X1 U16042 ( .IN1(n9125), .IN2(n14966), .Q(n14965) );
  AND2X1 U16043 ( .IN1(n14967), .IN2(n14968), .Q(n14966) );
  OR2X1 U16044 ( .IN1(n14599), .IN2(g843), .Q(n14968) );
  OR2X1 U16045 ( .IN1(n8356), .IN2(n14969), .Q(n14967) );
  INVX0 U16046 ( .INP(n14599), .ZN(n14969) );
  OR2X1 U16047 ( .IN1(n14970), .IN2(n14971), .Q(g25618) );
  AND2X1 U16048 ( .IN1(n14972), .IN2(g832), .Q(n14971) );
  OR2X1 U16049 ( .IN1(n14973), .IN2(n14974), .Q(n14972) );
  AND2X1 U16050 ( .IN1(n5822), .IN2(n4518), .Q(n14974) );
  AND2X1 U16051 ( .IN1(n9043), .IN2(n13689), .Q(n4518) );
  AND2X1 U16052 ( .IN1(n13727), .IN2(n13689), .Q(n14973) );
  AND2X1 U16053 ( .IN1(n14975), .IN2(g817), .Q(n14970) );
  OR2X1 U16054 ( .IN1(n9124), .IN2(n14976), .Q(n14975) );
  AND3X1 U16055 ( .IN1(n4948), .IN2(n13689), .IN3(n8545), .Q(n14976) );
  OR2X1 U16056 ( .IN1(n14977), .IN2(n14978), .Q(g25617) );
  AND2X1 U16057 ( .IN1(n9149), .IN2(g812), .Q(n14978) );
  AND3X1 U16058 ( .IN1(n14979), .IN2(n14980), .IN3(n13689), .Q(n14977) );
  OR2X1 U16059 ( .IN1(n14981), .IN2(n5709), .Q(n13689) );
  AND2X1 U16060 ( .IN1(n5733), .IN2(g837), .Q(n14981) );
  OR2X1 U16061 ( .IN1(n13728), .IN2(g817), .Q(n14980) );
  OR2X1 U16062 ( .IN1(n5822), .IN2(n13727), .Q(n14979) );
  AND2X1 U16063 ( .IN1(n14982), .IN2(n9026), .Q(g25616) );
  OR3X1 U16064 ( .IN1(n14983), .IN2(n14984), .IN3(n14985), .Q(n14982) );
  AND2X1 U16065 ( .IN1(n14986), .IN2(n14987), .Q(n14985) );
  INVX0 U16066 ( .INP(n14317), .ZN(n14986) );
  AND2X1 U16067 ( .IN1(n14987), .IN2(n5732), .Q(n14984) );
  AND3X1 U16068 ( .IN1(n14988), .IN2(n14317), .IN3(g732), .Q(n14983) );
  OR4X1 U16069 ( .IN1(n14297), .IN2(n14295), .IN3(g528), .IN4(n14989), .Q(
        n14317) );
  OR2X1 U16070 ( .IN1(g490), .IN2(g482), .Q(n14989) );
  OR2X1 U16071 ( .IN1(test_so54), .IN2(g518), .Q(n14297) );
  INVX0 U16072 ( .INP(n14987), .ZN(n14988) );
  OR2X1 U16073 ( .IN1(n14990), .IN2(n14991), .Q(n14987) );
  INVX0 U16074 ( .INP(n14992), .ZN(n14991) );
  OR2X1 U16075 ( .IN1(n14993), .IN2(n14994), .Q(n14992) );
  AND2X1 U16076 ( .IN1(n14994), .IN2(n14993), .Q(n14990) );
  AND2X1 U16077 ( .IN1(n14995), .IN2(n14996), .Q(n14993) );
  OR2X1 U16078 ( .IN1(n14997), .IN2(n5597), .Q(n14996) );
  OR2X1 U16079 ( .IN1(g225), .IN2(n14998), .Q(n14995) );
  INVX0 U16080 ( .INP(n14997), .ZN(n14998) );
  OR2X1 U16081 ( .IN1(n14999), .IN2(n15000), .Q(n14997) );
  AND3X1 U16082 ( .IN1(n15001), .IN2(n15002), .IN3(n15003), .Q(n15000) );
  OR2X1 U16083 ( .IN1(n15004), .IN2(n15005), .Q(n15003) );
  AND2X1 U16084 ( .IN1(n8658), .IN2(g239), .Q(n15005) );
  AND2X1 U16085 ( .IN1(n8659), .IN2(g232), .Q(n15004) );
  OR2X1 U16086 ( .IN1(n8660), .IN2(g255), .Q(n15002) );
  OR2X1 U16087 ( .IN1(n8661), .IN2(g269), .Q(n15001) );
  AND3X1 U16088 ( .IN1(n15006), .IN2(n15007), .IN3(n15008), .Q(n14999) );
  OR2X1 U16089 ( .IN1(n15009), .IN2(n15010), .Q(n15008) );
  AND2X1 U16090 ( .IN1(n8660), .IN2(g255), .Q(n15010) );
  AND2X1 U16091 ( .IN1(n8661), .IN2(g269), .Q(n15009) );
  OR2X1 U16092 ( .IN1(n8658), .IN2(g239), .Q(n15007) );
  OR2X1 U16093 ( .IN1(n8659), .IN2(g232), .Q(n15006) );
  OR2X1 U16094 ( .IN1(n15011), .IN2(n15012), .Q(n14994) );
  AND2X1 U16095 ( .IN1(n6008), .IN2(g262), .Q(n15012) );
  AND2X1 U16096 ( .IN1(n8662), .IN2(g246), .Q(n15011) );
  OR2X1 U16097 ( .IN1(n15013), .IN2(n15014), .Q(g25615) );
  AND2X1 U16098 ( .IN1(n15015), .IN2(g686), .Q(n15014) );
  AND2X1 U16099 ( .IN1(n14280), .IN2(g667), .Q(n15013) );
  OR3X1 U16100 ( .IN1(n15016), .IN2(n15017), .IN3(n15018), .Q(g25614) );
  AND2X1 U16101 ( .IN1(n9149), .IN2(g691), .Q(n15018) );
  AND2X1 U16102 ( .IN1(n5111), .IN2(n14281), .Q(n15017) );
  AND2X1 U16103 ( .IN1(n14280), .IN2(g686), .Q(n15016) );
  OR2X1 U16104 ( .IN1(n15019), .IN2(n15020), .Q(g25613) );
  AND2X1 U16105 ( .IN1(n9149), .IN2(g559), .Q(n15020) );
  AND4X1 U16106 ( .IN1(n2421), .IN2(n15021), .IN3(n15022), .IN4(n14617), .Q(
        n15019) );
  OR2X1 U16107 ( .IN1(n8281), .IN2(n15023), .Q(n14617) );
  OR2X1 U16108 ( .IN1(n15024), .IN2(g562), .Q(n15022) );
  INVX0 U16109 ( .INP(n15023), .ZN(n15024) );
  OR2X1 U16110 ( .IN1(n15025), .IN2(n8688), .Q(n15023) );
  AND2X1 U16111 ( .IN1(n8272), .IN2(g12368), .Q(n15025) );
  OR2X1 U16112 ( .IN1(n5288), .IN2(n15421), .Q(n15021) );
  OR2X1 U16113 ( .IN1(n15026), .IN2(n15027), .Q(g25612) );
  AND2X1 U16114 ( .IN1(n14280), .IN2(g518), .Q(n15027) );
  AND2X1 U16115 ( .IN1(n15028), .IN2(g513), .Q(n15026) );
  OR2X1 U16116 ( .IN1(n15029), .IN2(n15030), .Q(g25611) );
  AND2X1 U16117 ( .IN1(n14280), .IN2(g513), .Q(n15030) );
  AND2X1 U16118 ( .IN1(n15028), .IN2(g504), .Q(n15029) );
  OR2X1 U16119 ( .IN1(n9136), .IN2(n15031), .Q(n15028) );
  AND2X1 U16120 ( .IN1(n14281), .IN2(n14623), .Q(n15031) );
  INVX0 U16121 ( .INP(n4962), .ZN(n14623) );
  OR3X1 U16122 ( .IN1(n15032), .IN2(n15033), .IN3(n15034), .Q(g25610) );
  AND2X1 U16123 ( .IN1(test_so54), .IN2(n15015), .Q(n15033) );
  AND2X1 U16124 ( .IN1(n14280), .IN2(g504), .Q(n15032) );
  OR3X1 U16125 ( .IN1(n15034), .IN2(n15035), .IN3(n15036), .Q(g25609) );
  AND2X1 U16126 ( .IN1(test_so54), .IN2(n15037), .Q(n15036) );
  OR2X1 U16127 ( .IN1(n15038), .IN2(n14280), .Q(n15037) );
  INVX0 U16128 ( .INP(n15015), .ZN(n14280) );
  OR2X1 U16129 ( .IN1(n9136), .IN2(n14281), .Q(n15015) );
  AND2X1 U16130 ( .IN1(n5548), .IN2(n9025), .Q(n15038) );
  AND3X1 U16131 ( .IN1(n5287), .IN2(n9053), .IN3(n14281), .Q(n15035) );
  AND2X1 U16132 ( .IN1(n14281), .IN2(n13718), .Q(n15034) );
  AND2X1 U16133 ( .IN1(n9043), .IN2(n4962), .Q(n13718) );
  AND3X1 U16134 ( .IN1(g358), .IN2(g385), .IN3(n5633), .Q(n14281) );
  OR3X1 U16135 ( .IN1(n15039), .IN2(n15040), .IN3(n15041), .Q(g25605) );
  AND2X1 U16136 ( .IN1(n15042), .IN2(g460), .Q(n15041) );
  AND3X1 U16137 ( .IN1(n15043), .IN2(g246), .IN3(n9064), .Q(n15040) );
  AND2X1 U16138 ( .IN1(n9149), .IN2(g168), .Q(n15039) );
  OR2X1 U16139 ( .IN1(n15044), .IN2(n15045), .Q(g25604) );
  AND2X1 U16140 ( .IN1(n15046), .IN2(g460), .Q(n15045) );
  AND2X1 U16141 ( .IN1(n15042), .IN2(g452), .Q(n15044) );
  OR3X1 U16142 ( .IN1(n15047), .IN2(n15048), .IN3(n15049), .Q(g25602) );
  AND2X1 U16143 ( .IN1(n15042), .IN2(test_so72), .Q(n15049) );
  AND3X1 U16144 ( .IN1(n15043), .IN2(g446), .IN3(n9064), .Q(n15048) );
  AND2X1 U16145 ( .IN1(n9149), .IN2(g405), .Q(n15047) );
  OR2X1 U16146 ( .IN1(n15050), .IN2(n15051), .Q(g25601) );
  AND2X1 U16147 ( .IN1(test_so72), .IN2(n15046), .Q(n15051) );
  AND2X1 U16148 ( .IN1(n15042), .IN2(g174), .Q(n15050) );
  OR2X1 U16149 ( .IN1(n15052), .IN2(n15053), .Q(g25600) );
  AND2X1 U16150 ( .IN1(n15046), .IN2(g174), .Q(n15053) );
  AND2X1 U16151 ( .IN1(n15042), .IN2(g168), .Q(n15052) );
  INVX0 U16152 ( .INP(n15046), .ZN(n15042) );
  OR2X1 U16153 ( .IN1(n9136), .IN2(n15043), .Q(n15046) );
  INVX0 U16154 ( .INP(n14295), .ZN(n15043) );
  OR2X1 U16155 ( .IN1(n5121), .IN2(g370), .Q(n14295) );
  OR2X1 U16156 ( .IN1(n15054), .IN2(n15055), .Q(g25599) );
  AND2X1 U16157 ( .IN1(n9149), .IN2(g385), .Q(n15054) );
  OR2X1 U16158 ( .IN1(n15056), .IN2(n15057), .Q(g25598) );
  AND2X1 U16159 ( .IN1(n15058), .IN2(g376), .Q(n15057) );
  OR2X1 U16160 ( .IN1(n9135), .IN2(n15059), .Q(n15058) );
  AND2X1 U16161 ( .IN1(n5121), .IN2(g358), .Q(n15059) );
  AND3X1 U16162 ( .IN1(n9054), .IN2(g385), .IN3(n5121), .Q(n15056) );
  OR3X1 U16163 ( .IN1(n8788), .IN2(n5633), .IN3(n5632), .Q(n5121) );
  OR2X1 U16164 ( .IN1(n15060), .IN2(n15061), .Q(g25597) );
  AND3X1 U16165 ( .IN1(n15062), .IN2(n15063), .IN3(n9064), .Q(n15061) );
  OR2X1 U16166 ( .IN1(n15055), .IN2(g370), .Q(n15063) );
  INVX0 U16167 ( .INP(n10206), .ZN(n15055) );
  OR2X1 U16168 ( .IN1(n8636), .IN2(n10206), .Q(n15062) );
  OR3X1 U16169 ( .IN1(n8690), .IN2(n5633), .IN3(n5632), .Q(n10206) );
  AND2X1 U16170 ( .IN1(n9149), .IN2(g358), .Q(n15060) );
  OR2X1 U16171 ( .IN1(n15064), .IN2(n15065), .Q(g25596) );
  AND2X1 U16172 ( .IN1(n15066), .IN2(n9025), .Q(n15065) );
  OR2X1 U16173 ( .IN1(n15067), .IN2(n15068), .Q(n15066) );
  AND2X1 U16174 ( .IN1(n5633), .IN2(g358), .Q(n15068) );
  AND2X1 U16175 ( .IN1(n8788), .IN2(g376), .Q(n15067) );
  AND2X1 U16176 ( .IN1(n9149), .IN2(g370), .Q(n15064) );
  AND3X1 U16177 ( .IN1(n8788), .IN2(n9052), .IN3(n8690), .Q(g25595) );
  AND3X1 U16178 ( .IN1(n14315), .IN2(n9053), .IN3(n14313), .Q(g25594) );
  OR2X1 U16179 ( .IN1(n15069), .IN2(g278), .Q(n14313) );
  AND4X1 U16180 ( .IN1(n6008), .IN2(n8658), .IN3(n8659), .IN4(n15070), .Q(
        n15069) );
  AND4X1 U16181 ( .IN1(g269), .IN2(n5597), .IN3(g262), .IN4(g255), .Q(n15070)
         );
  OR4X1 U16182 ( .IN1(g269), .IN2(g255), .IN3(g262), .IN4(n15071), .Q(n14315)
         );
  OR4X1 U16183 ( .IN1(n6008), .IN2(n5597), .IN3(n8659), .IN4(n8658), .Q(n15071) );
  OR2X1 U16184 ( .IN1(n15072), .IN2(n15073), .Q(g25593) );
  AND2X1 U16185 ( .IN1(n15074), .IN2(n9025), .Q(n15073) );
  OR2X1 U16186 ( .IN1(n15075), .IN2(n15076), .Q(n15074) );
  AND2X1 U16187 ( .IN1(n15077), .IN2(n15078), .Q(n15076) );
  INVX0 U16188 ( .INP(n15079), .ZN(n15078) );
  AND2X1 U16189 ( .IN1(n15079), .IN2(g209), .Q(n15075) );
  AND2X1 U16190 ( .IN1(n9149), .IN2(g191), .Q(n15072) );
  OR2X1 U16191 ( .IN1(n15080), .IN2(n15081), .Q(g25592) );
  AND3X1 U16192 ( .IN1(n15082), .IN2(n15083), .IN3(n9064), .Q(n15081) );
  INVX0 U16193 ( .INP(n15084), .ZN(n15083) );
  AND2X1 U16194 ( .IN1(n15085), .IN2(n8374), .Q(n15084) );
  OR2X1 U16195 ( .IN1(n8374), .IN2(n15085), .Q(n15082) );
  OR2X1 U16196 ( .IN1(n15079), .IN2(n15077), .Q(n15085) );
  OR2X1 U16197 ( .IN1(n15086), .IN2(n15087), .Q(n15077) );
  AND2X1 U16198 ( .IN1(n8374), .IN2(g191), .Q(n15087) );
  AND2X1 U16199 ( .IN1(n8375), .IN2(g8358), .Q(n15086) );
  OR2X1 U16200 ( .IN1(n8548), .IN2(n8547), .Q(n15079) );
  AND2X1 U16201 ( .IN1(n9149), .IN2(g222), .Q(n15080) );
  OR2X1 U16202 ( .IN1(n15088), .IN2(n15089), .Q(g25591) );
  AND2X1 U16203 ( .IN1(n9149), .IN2(g209), .Q(n15089) );
  AND2X1 U16204 ( .IN1(n8548), .IN2(n9025), .Q(n15088) );
  AND2X1 U16205 ( .IN1(test_so94), .IN2(n5525), .Q(g25167) );
  AND2X1 U16206 ( .IN1(n15090), .IN2(g6732), .Q(g24355) );
  OR2X1 U16207 ( .IN1(n9135), .IN2(n15091), .Q(n15090) );
  OR2X1 U16208 ( .IN1(n15092), .IN2(n15093), .Q(g24354) );
  AND3X1 U16209 ( .IN1(n8753), .IN2(n15091), .IN3(n9063), .Q(n15093) );
  AND2X1 U16210 ( .IN1(n9150), .IN2(g6727), .Q(n15092) );
  OR2X1 U16211 ( .IN1(n15094), .IN2(n15095), .Q(g24353) );
  AND3X1 U16212 ( .IN1(n15091), .IN2(n15096), .IN3(n9063), .Q(n15095) );
  OR2X1 U16213 ( .IN1(n15097), .IN2(g6727), .Q(n15096) );
  OR2X1 U16214 ( .IN1(n5531), .IN2(n15098), .Q(n15091) );
  INVX0 U16215 ( .INP(n15097), .ZN(n15098) );
  AND4X1 U16216 ( .IN1(g14828), .IN2(test_so80), .IN3(g17688), .IN4(g17778), 
        .Q(n15097) );
  AND2X1 U16217 ( .IN1(n9150), .IN2(g6723), .Q(n15094) );
  AND4X1 U16218 ( .IN1(n15099), .IN2(n15100), .IN3(n8717), .IN4(n15101), .Q(
        g24352) );
  AND3X1 U16219 ( .IN1(n8715), .IN2(n9052), .IN3(n8716), .Q(n15101) );
  OR2X1 U16220 ( .IN1(n8668), .IN2(g14828), .Q(n15100) );
  OR2X1 U16221 ( .IN1(test_so80), .IN2(n5700), .Q(n15099) );
  AND2X1 U16222 ( .IN1(n15102), .IN2(g6386), .Q(g24351) );
  OR2X1 U16223 ( .IN1(n9134), .IN2(n15103), .Q(n15102) );
  OR2X1 U16224 ( .IN1(n15104), .IN2(n15105), .Q(g24350) );
  AND3X1 U16225 ( .IN1(n8744), .IN2(n15103), .IN3(n9062), .Q(n15105) );
  OR2X1 U16226 ( .IN1(n8829), .IN2(n15106), .Q(n15103) );
  AND2X1 U16227 ( .IN1(test_so69), .IN2(n9138), .Q(n15104) );
  OR2X1 U16228 ( .IN1(n15107), .IN2(n15108), .Q(g24349) );
  AND2X1 U16229 ( .IN1(n15109), .IN2(n9025), .Q(n15108) );
  OR2X1 U16230 ( .IN1(n15110), .IN2(n15111), .Q(n15109) );
  AND2X1 U16231 ( .IN1(n15112), .IN2(n8829), .Q(n15111) );
  AND2X1 U16232 ( .IN1(test_so69), .IN2(n15106), .Q(n15110) );
  INVX0 U16233 ( .INP(n15112), .ZN(n15106) );
  AND4X1 U16234 ( .IN1(g14779), .IN2(g12422), .IN3(g17649), .IN4(g17760), .Q(
        n15112) );
  AND2X1 U16235 ( .IN1(n9150), .IN2(g6377), .Q(n15107) );
  AND4X1 U16236 ( .IN1(n15113), .IN2(n15114), .IN3(n8708), .IN4(n15115), .Q(
        g24348) );
  AND3X1 U16237 ( .IN1(n8706), .IN2(n9051), .IN3(n8707), .Q(n15115) );
  OR2X1 U16238 ( .IN1(n8665), .IN2(g14779), .Q(n15114) );
  OR2X1 U16239 ( .IN1(n5703), .IN2(g12422), .Q(n15113) );
  AND2X1 U16240 ( .IN1(n15116), .IN2(g6040), .Q(g24347) );
  OR2X1 U16241 ( .IN1(n9134), .IN2(n15117), .Q(n15116) );
  OR2X1 U16242 ( .IN1(n15118), .IN2(n15119), .Q(g24346) );
  AND3X1 U16243 ( .IN1(n15117), .IN2(n8844), .IN3(n9062), .Q(n15119) );
  AND2X1 U16244 ( .IN1(n9150), .IN2(g6035), .Q(n15118) );
  OR2X1 U16245 ( .IN1(n15120), .IN2(n15121), .Q(g24345) );
  AND3X1 U16246 ( .IN1(n15117), .IN2(n15122), .IN3(n9062), .Q(n15121) );
  OR2X1 U16247 ( .IN1(n15123), .IN2(g6035), .Q(n15122) );
  OR2X1 U16248 ( .IN1(n5528), .IN2(n15124), .Q(n15117) );
  INVX0 U16249 ( .INP(n15123), .ZN(n15124) );
  AND4X1 U16250 ( .IN1(g14738), .IN2(g12350), .IN3(g17607), .IN4(g17739), .Q(
        n15123) );
  AND2X1 U16251 ( .IN1(n9151), .IN2(g6031), .Q(n15120) );
  AND4X1 U16252 ( .IN1(n15125), .IN2(n15126), .IN3(n8763), .IN4(n15127), .Q(
        g24344) );
  AND3X1 U16253 ( .IN1(n8761), .IN2(n9052), .IN3(n8762), .Q(n15127) );
  OR2X1 U16254 ( .IN1(n8667), .IN2(g14738), .Q(n15126) );
  OR2X1 U16255 ( .IN1(n5698), .IN2(g12350), .Q(n15125) );
  AND2X1 U16256 ( .IN1(n15128), .IN2(g5694), .Q(g24343) );
  OR2X1 U16257 ( .IN1(n9134), .IN2(n15129), .Q(n15128) );
  OR2X1 U16258 ( .IN1(n15130), .IN2(n15131), .Q(g24342) );
  AND3X1 U16259 ( .IN1(n8754), .IN2(n15129), .IN3(n9062), .Q(n15131) );
  AND2X1 U16260 ( .IN1(n9151), .IN2(g5689), .Q(n15130) );
  OR2X1 U16261 ( .IN1(n15132), .IN2(n15133), .Q(g24341) );
  AND3X1 U16262 ( .IN1(n15129), .IN2(n15134), .IN3(n9062), .Q(n15133) );
  OR2X1 U16263 ( .IN1(n15135), .IN2(g5689), .Q(n15134) );
  OR2X1 U16264 ( .IN1(n5529), .IN2(n15136), .Q(n15129) );
  INVX0 U16265 ( .INP(n15135), .ZN(n15136) );
  AND4X1 U16266 ( .IN1(g14694), .IN2(g12300), .IN3(g17580), .IN4(g17711), .Q(
        n15135) );
  AND2X1 U16267 ( .IN1(n9151), .IN2(g5685), .Q(n15132) );
  AND4X1 U16268 ( .IN1(n15137), .IN2(n15138), .IN3(n8702), .IN4(n15139), .Q(
        g24340) );
  AND3X1 U16269 ( .IN1(n8700), .IN2(n9052), .IN3(n8701), .Q(n15139) );
  OR2X1 U16270 ( .IN1(n8669), .IN2(g14694), .Q(n15138) );
  OR2X1 U16271 ( .IN1(n5705), .IN2(g12300), .Q(n15137) );
  AND2X1 U16272 ( .IN1(n15140), .IN2(g5348), .Q(g24339) );
  OR2X1 U16273 ( .IN1(n9134), .IN2(n15141), .Q(n15140) );
  OR2X1 U16274 ( .IN1(n15142), .IN2(n15143), .Q(g24338) );
  AND3X1 U16275 ( .IN1(n8774), .IN2(n15141), .IN3(n9062), .Q(n15143) );
  OR2X1 U16276 ( .IN1(n8828), .IN2(n15144), .Q(n15141) );
  AND2X1 U16277 ( .IN1(test_so10), .IN2(n9139), .Q(n15142) );
  OR2X1 U16278 ( .IN1(n15145), .IN2(n15146), .Q(g24337) );
  AND2X1 U16279 ( .IN1(n15147), .IN2(n9025), .Q(n15146) );
  OR2X1 U16280 ( .IN1(n15148), .IN2(n15149), .Q(n15147) );
  AND2X1 U16281 ( .IN1(n15150), .IN2(n8828), .Q(n15149) );
  AND2X1 U16282 ( .IN1(test_so10), .IN2(n15144), .Q(n15148) );
  INVX0 U16283 ( .INP(n15150), .ZN(n15144) );
  AND4X1 U16284 ( .IN1(g14662), .IN2(g12238), .IN3(g17519), .IN4(g17674), .Q(
        n15150) );
  AND2X1 U16285 ( .IN1(n9151), .IN2(g5339), .Q(n15145) );
  AND4X1 U16286 ( .IN1(n15151), .IN2(n15152), .IN3(n8705), .IN4(n15153), .Q(
        g24336) );
  AND3X1 U16287 ( .IN1(n8703), .IN2(n9051), .IN3(n8704), .Q(n15153) );
  OR2X1 U16288 ( .IN1(n8670), .IN2(g14662), .Q(n15152) );
  OR2X1 U16289 ( .IN1(n5704), .IN2(g12238), .Q(n15151) );
  OR2X1 U16290 ( .IN1(n15154), .IN2(n15155), .Q(g24335) );
  AND2X1 U16291 ( .IN1(n9151), .IN2(g18881), .Q(n15155) );
  AND3X1 U16292 ( .IN1(n5653), .IN2(g4643), .IN3(n15156), .Q(n15154) );
  OR2X1 U16293 ( .IN1(n15157), .IN2(n15158), .Q(g24334) );
  AND2X1 U16294 ( .IN1(n9151), .IN2(g4358), .Q(n15158) );
  AND4X1 U16295 ( .IN1(n14427), .IN2(n5608), .IN3(n15156), .IN4(n15159), .Q(
        n15157) );
  AND4X1 U16296 ( .IN1(n5274), .IN2(n5539), .IN3(n5303), .IN4(n5365), .Q(
        n15159) );
  AND4X1 U16297 ( .IN1(n8822), .IN2(n9082), .IN3(n5506), .IN4(n15160), .Q(
        n15156) );
  AND3X1 U16298 ( .IN1(n5540), .IN2(n5323), .IN3(n5348), .Q(n15160) );
  AND4X1 U16299 ( .IN1(n5727), .IN2(test_so3), .IN3(g4633), .IN4(g4340), .Q(
        n14427) );
  AND2X1 U16300 ( .IN1(n9141), .IN2(g4392), .Q(g24298) );
  OR2X1 U16301 ( .IN1(n15161), .IN2(n15162), .Q(g24282) );
  AND2X1 U16302 ( .IN1(g24281), .IN2(g9251), .Q(n15162) );
  AND2X1 U16303 ( .IN1(n15163), .IN2(g4308), .Q(n15161) );
  OR2X1 U16304 ( .IN1(n8511), .IN2(n9123), .Q(n15163) );
  AND2X1 U16305 ( .IN1(n9045), .IN2(n8542), .Q(g24281) );
  OR2X1 U16306 ( .IN1(n15164), .IN2(n15165), .Q(g24280) );
  AND2X1 U16307 ( .IN1(n15166), .IN2(g4273), .Q(n15165) );
  OR2X1 U16308 ( .IN1(n15167), .IN2(n15168), .Q(n15166) );
  AND2X1 U16309 ( .IN1(n5763), .IN2(n9025), .Q(n15167) );
  AND2X1 U16310 ( .IN1(n15169), .IN2(g4269), .Q(n15164) );
  OR2X1 U16311 ( .IN1(n9133), .IN2(n15170), .Q(n15169) );
  AND3X1 U16312 ( .IN1(g4264), .IN2(g4258), .IN3(n5764), .Q(n15170) );
  OR2X1 U16313 ( .IN1(n15171), .IN2(n15172), .Q(g24279) );
  AND3X1 U16314 ( .IN1(n15173), .IN2(n15174), .IN3(n9062), .Q(n15172) );
  OR2X1 U16315 ( .IN1(n15175), .IN2(n15176), .Q(n15174) );
  INVX0 U16316 ( .INP(n15177), .ZN(n15173) );
  AND2X1 U16317 ( .IN1(n15176), .IN2(n15175), .Q(n15177) );
  AND2X1 U16318 ( .IN1(n15178), .IN2(n15179), .Q(n15176) );
  INVX0 U16319 ( .INP(n15180), .ZN(n15179) );
  AND3X1 U16320 ( .IN1(n5726), .IN2(n15181), .IN3(n8620), .Q(n15180) );
  OR4X1 U16321 ( .IN1(g11770), .IN2(g8916), .IN3(g8915), .IN4(n15182), .Q(
        n15181) );
  OR4X1 U16322 ( .IN1(g8920), .IN2(g8919), .IN3(g8918), .IN4(g8917), .Q(n15182) );
  OR2X1 U16323 ( .IN1(n5726), .IN2(n8620), .Q(n15178) );
  INVX0 U16324 ( .INP(n15183), .ZN(n15171) );
  OR2X1 U16325 ( .IN1(n9008), .IN2(n8620), .Q(n15183) );
  AND2X1 U16326 ( .IN1(n15184), .IN2(g4045), .Q(g24278) );
  OR2X1 U16327 ( .IN1(n9133), .IN2(n15185), .Q(n15184) );
  OR2X1 U16328 ( .IN1(n15186), .IN2(n15187), .Q(g24277) );
  AND3X1 U16329 ( .IN1(n8746), .IN2(n15185), .IN3(n9061), .Q(n15187) );
  AND2X1 U16330 ( .IN1(n9140), .IN2(g4040), .Q(n15186) );
  OR2X1 U16331 ( .IN1(n15188), .IN2(n15189), .Q(g24276) );
  AND3X1 U16332 ( .IN1(n15185), .IN2(n15190), .IN3(n9061), .Q(n15189) );
  OR2X1 U16333 ( .IN1(n15191), .IN2(g4040), .Q(n15190) );
  OR2X1 U16334 ( .IN1(n5530), .IN2(n15192), .Q(n15185) );
  INVX0 U16335 ( .INP(n15191), .ZN(n15192) );
  AND4X1 U16336 ( .IN1(g13966), .IN2(g11418), .IN3(g16659), .IN4(g16775), .Q(
        n15191) );
  AND2X1 U16337 ( .IN1(n9141), .IN2(g4031), .Q(n15188) );
  AND4X1 U16338 ( .IN1(n15193), .IN2(n15194), .IN3(n8714), .IN4(n15195), .Q(
        g24275) );
  AND3X1 U16339 ( .IN1(n8712), .IN2(n9051), .IN3(n8713), .Q(n15195) );
  OR2X1 U16340 ( .IN1(n8666), .IN2(g13966), .Q(n15194) );
  OR2X1 U16341 ( .IN1(n5701), .IN2(g11418), .Q(n15193) );
  AND2X1 U16342 ( .IN1(n15196), .IN2(g3694), .Q(g24274) );
  OR2X1 U16343 ( .IN1(n9133), .IN2(n15197), .Q(n15196) );
  OR2X1 U16344 ( .IN1(n15198), .IN2(n15199), .Q(g24273) );
  AND3X1 U16345 ( .IN1(n8755), .IN2(n15197), .IN3(n9061), .Q(n15199) );
  AND2X1 U16346 ( .IN1(n9140), .IN2(g3689), .Q(n15198) );
  OR2X1 U16347 ( .IN1(n15200), .IN2(n15201), .Q(g24272) );
  AND3X1 U16348 ( .IN1(n15197), .IN2(n15202), .IN3(n9061), .Q(n15201) );
  OR2X1 U16349 ( .IN1(n15203), .IN2(g3689), .Q(n15202) );
  OR2X1 U16350 ( .IN1(n5532), .IN2(n15204), .Q(n15197) );
  INVX0 U16351 ( .INP(n15203), .ZN(n15204) );
  AND4X1 U16352 ( .IN1(g13926), .IN2(g11388), .IN3(g16627), .IN4(g16744), .Q(
        n15203) );
  AND2X1 U16353 ( .IN1(n9140), .IN2(g3680), .Q(n15200) );
  AND4X1 U16354 ( .IN1(n15205), .IN2(n15206), .IN3(n8720), .IN4(n15207), .Q(
        g24271) );
  AND3X1 U16355 ( .IN1(n8718), .IN2(n9051), .IN3(n8719), .Q(n15207) );
  OR2X1 U16356 ( .IN1(n8663), .IN2(g13926), .Q(n15206) );
  OR2X1 U16357 ( .IN1(n5699), .IN2(g11388), .Q(n15205) );
  AND2X1 U16358 ( .IN1(n15208), .IN2(g3343), .Q(g24270) );
  OR2X1 U16359 ( .IN1(n9133), .IN2(n15209), .Q(n15208) );
  OR2X1 U16360 ( .IN1(n15210), .IN2(n15211), .Q(g24269) );
  AND3X1 U16361 ( .IN1(n8743), .IN2(n15209), .IN3(n9060), .Q(n15211) );
  AND2X1 U16362 ( .IN1(n9140), .IN2(g3338), .Q(n15210) );
  OR2X1 U16363 ( .IN1(n15212), .IN2(n15213), .Q(g24268) );
  AND3X1 U16364 ( .IN1(n15209), .IN2(n15214), .IN3(n9060), .Q(n15213) );
  OR2X1 U16365 ( .IN1(n15215), .IN2(g3338), .Q(n15214) );
  OR2X1 U16366 ( .IN1(n5527), .IN2(n15216), .Q(n15209) );
  INVX0 U16367 ( .INP(n15215), .ZN(n15216) );
  AND4X1 U16368 ( .IN1(g13895), .IN2(g11349), .IN3(g16603), .IN4(g16718), .Q(
        n15215) );
  AND2X1 U16369 ( .IN1(test_so91), .IN2(n9138), .Q(n15212) );
  AND4X1 U16370 ( .IN1(n15217), .IN2(n15218), .IN3(n8711), .IN4(n15219), .Q(
        g24267) );
  AND3X1 U16371 ( .IN1(n8709), .IN2(n9050), .IN3(n8710), .Q(n15219) );
  OR2X1 U16372 ( .IN1(n8664), .IN2(g13895), .Q(n15218) );
  OR2X1 U16373 ( .IN1(n5702), .IN2(g11349), .Q(n15217) );
  OR2X1 U16374 ( .IN1(n15220), .IN2(n15221), .Q(g24266) );
  AND3X1 U16375 ( .IN1(test_so9), .IN2(n8751), .IN3(n9060), .Q(n15221) );
  AND2X1 U16376 ( .IN1(n9140), .IN2(g2841), .Q(n15220) );
  OR3X1 U16377 ( .IN1(n15222), .IN2(n15223), .IN3(n2787), .Q(g24263) );
  AND2X1 U16378 ( .IN1(n9046), .IN2(n5963), .Q(n2787) );
  AND2X1 U16379 ( .IN1(n9140), .IN2(g2712), .Q(n15223) );
  AND2X1 U16380 ( .IN1(n5299), .IN2(n9025), .Q(n15222) );
  OR2X1 U16381 ( .IN1(n15224), .IN2(n11485), .Q(g24261) );
  AND2X1 U16382 ( .IN1(n9140), .IN2(g1585), .Q(n15224) );
  AND2X1 U16383 ( .IN1(n15225), .IN2(n15226), .Q(g24260) );
  OR2X1 U16384 ( .IN1(n15227), .IN2(g1430), .Q(n15226) );
  AND2X1 U16385 ( .IN1(n9047), .IN2(g1548), .Q(n15227) );
  OR2X1 U16386 ( .IN1(n9132), .IN2(n9350), .Q(n15225) );
  OR2X1 U16387 ( .IN1(n15228), .IN2(n11485), .Q(g24259) );
  AND2X1 U16388 ( .IN1(n9140), .IN2(g1579), .Q(n15228) );
  OR2X1 U16389 ( .IN1(n15229), .IN2(n15230), .Q(g24258) );
  AND2X1 U16390 ( .IN1(n9140), .IN2(g1554), .Q(n15230) );
  AND2X1 U16391 ( .IN1(n9045), .IN2(g496), .Q(n15229) );
  AND2X1 U16392 ( .IN1(n15231), .IN2(n15232), .Q(g24257) );
  INVX0 U16393 ( .INP(n15233), .ZN(n15232) );
  AND2X1 U16394 ( .IN1(n15234), .IN2(n5616), .Q(n15233) );
  OR2X1 U16395 ( .IN1(n5616), .IN2(n15234), .Q(n15231) );
  OR2X1 U16396 ( .IN1(n9132), .IN2(n15235), .Q(n15234) );
  OR2X1 U16397 ( .IN1(n15236), .IN2(n15237), .Q(g24256) );
  AND2X1 U16398 ( .IN1(n15238), .IN2(n9025), .Q(n15237) );
  OR2X1 U16399 ( .IN1(n15239), .IN2(n15240), .Q(n15238) );
  AND4X1 U16400 ( .IN1(n8740), .IN2(n14894), .IN3(n8741), .IN4(n15235), .Q(
        n15240) );
  INVX0 U16401 ( .INP(n15241), .ZN(n15239) );
  OR2X1 U16402 ( .IN1(n15235), .IN2(n15242), .Q(n15241) );
  AND3X1 U16403 ( .IN1(n14894), .IN2(n8740), .IN3(n8741), .Q(n15242) );
  AND3X1 U16404 ( .IN1(n5616), .IN2(n5302), .IN3(n5401), .Q(n14894) );
  OR4X1 U16405 ( .IN1(n1392), .IN2(n14512), .IN3(n15243), .IN4(n15244), .Q(
        n15235) );
  AND2X1 U16406 ( .IN1(n8360), .IN2(n8824), .Q(n15244) );
  AND2X1 U16407 ( .IN1(test_so68), .IN2(g1579), .Q(n15243) );
  AND2X1 U16408 ( .IN1(n9141), .IN2(g1339), .Q(n15236) );
  OR3X1 U16409 ( .IN1(n15245), .IN2(n15246), .IN3(n15247), .Q(g24255) );
  AND2X1 U16410 ( .IN1(n11485), .IN2(g17423), .Q(n15247) );
  AND2X1 U16411 ( .IN1(n9141), .IN2(g1589), .Q(n15246) );
  AND3X1 U16412 ( .IN1(n8734), .IN2(g10527), .IN3(n9061), .Q(n15245) );
  AND3X1 U16413 ( .IN1(n8735), .IN2(n8733), .IN3(n15248), .Q(g24254) );
  AND3X1 U16414 ( .IN1(n15249), .IN2(n9051), .IN3(n8734), .Q(n15248) );
  OR3X1 U16415 ( .IN1(n5768), .IN2(n15250), .IN3(n14870), .Q(n15249) );
  OR2X1 U16416 ( .IN1(n8729), .IN2(n9350), .Q(n14870) );
  OR2X1 U16417 ( .IN1(n5546), .IN2(n8544), .Q(n9350) );
  AND2X1 U16418 ( .IN1(n14898), .IN2(n14320), .Q(n15250) );
  INVX0 U16419 ( .INP(n1392), .ZN(n14320) );
  OR2X1 U16420 ( .IN1(g1351), .IN2(g1312), .Q(n1392) );
  INVX0 U16421 ( .INP(n14512), .ZN(n14898) );
  OR2X1 U16422 ( .IN1(n13089), .IN2(n14234), .Q(n14512) );
  OR2X1 U16423 ( .IN1(n15251), .IN2(n15252), .Q(n14234) );
  AND2X1 U16424 ( .IN1(n5381), .IN2(n8824), .Q(n15252) );
  AND2X1 U16425 ( .IN1(test_so68), .IN2(g1339), .Q(n15251) );
  AND2X1 U16426 ( .IN1(n8824), .IN2(n5616), .Q(n13089) );
  OR2X1 U16427 ( .IN1(n15253), .IN2(n15254), .Q(g24253) );
  AND2X1 U16428 ( .IN1(n15255), .IN2(n9025), .Q(n15254) );
  OR2X1 U16429 ( .IN1(n15256), .IN2(n15257), .Q(n15255) );
  AND2X1 U16430 ( .IN1(g7946), .IN2(g1521), .Q(n15257) );
  AND2X1 U16431 ( .IN1(n5302), .IN2(g1532), .Q(n15256) );
  AND2X1 U16432 ( .IN1(n9141), .IN2(g1306), .Q(n15253) );
  OR2X1 U16433 ( .IN1(n15258), .IN2(n15259), .Q(g24252) );
  AND2X1 U16434 ( .IN1(n15260), .IN2(n9024), .Q(n15259) );
  OR2X1 U16435 ( .IN1(n15261), .IN2(n15262), .Q(n15260) );
  AND2X1 U16436 ( .IN1(g7946), .IN2(g1339), .Q(n15262) );
  AND2X1 U16437 ( .IN1(n5302), .IN2(g1521), .Q(n15261) );
  AND2X1 U16438 ( .IN1(test_so49), .IN2(n9139), .Q(n15258) );
  OR2X1 U16439 ( .IN1(n15263), .IN2(n15264), .Q(g24251) );
  AND2X1 U16440 ( .IN1(test_so12), .IN2(n15265), .Q(n15264) );
  AND2X1 U16441 ( .IN1(n13616), .IN2(g1442), .Q(n15263) );
  OR2X1 U16442 ( .IN1(n15266), .IN2(n15267), .Q(g24250) );
  AND2X1 U16443 ( .IN1(n15265), .IN2(g1489), .Q(n15267) );
  AND2X1 U16444 ( .IN1(test_so12), .IN2(n13616), .Q(n15266) );
  INVX0 U16445 ( .INP(n15265), .ZN(n13616) );
  OR2X1 U16446 ( .IN1(n15268), .IN2(n15269), .Q(g24249) );
  AND2X1 U16447 ( .IN1(n15270), .IN2(g1489), .Q(n15269) );
  INVX0 U16448 ( .INP(n15271), .ZN(n15270) );
  AND2X1 U16449 ( .IN1(n15272), .IN2(n15265), .Q(n15271) );
  OR2X1 U16450 ( .IN1(n9132), .IN2(n13621), .Q(n15265) );
  OR2X1 U16451 ( .IN1(n9132), .IN2(test_so12), .Q(n15272) );
  AND3X1 U16452 ( .IN1(n8551), .IN2(n9051), .IN3(n13621), .Q(n15268) );
  AND3X1 U16453 ( .IN1(n8819), .IN2(g13272), .IN3(n5364), .Q(n13621) );
  OR3X1 U16454 ( .IN1(n15273), .IN2(n15274), .IN3(n15275), .Q(g24248) );
  AND2X1 U16455 ( .IN1(n11485), .IN2(g1395), .Q(n15275) );
  AND2X1 U16456 ( .IN1(n15276), .IN2(g1404), .Q(n15274) );
  AND2X1 U16457 ( .IN1(n15277), .IN2(n9024), .Q(n15273) );
  OR2X1 U16458 ( .IN1(n15278), .IN2(n5401), .Q(n15277) );
  AND2X1 U16459 ( .IN1(n5655), .IN2(n15276), .Q(n15278) );
  OR3X1 U16460 ( .IN1(n8757), .IN2(n9121), .IN3(g12923), .Q(n15276) );
  AND2X1 U16461 ( .IN1(n11485), .IN2(n8770), .Q(g24247) );
  AND2X1 U16462 ( .IN1(g12923), .IN2(n9029), .Q(n11485) );
  OR2X1 U16463 ( .IN1(n15279), .IN2(n11500), .Q(g24245) );
  AND2X1 U16464 ( .IN1(n9141), .IN2(g30332), .Q(n15279) );
  AND2X1 U16465 ( .IN1(n15280), .IN2(n15281), .Q(g24244) );
  OR2X1 U16466 ( .IN1(n15282), .IN2(g1087), .Q(n15281) );
  AND2X1 U16467 ( .IN1(n9045), .IN2(g1205), .Q(n15282) );
  OR2X1 U16468 ( .IN1(n9132), .IN2(n9483), .Q(n15280) );
  OR2X1 U16469 ( .IN1(n15283), .IN2(n11500), .Q(g24243) );
  AND2X1 U16470 ( .IN1(n9141), .IN2(g1236), .Q(n15283) );
  OR2X1 U16471 ( .IN1(n15284), .IN2(n15285), .Q(g24242) );
  AND2X1 U16472 ( .IN1(test_so76), .IN2(n9137), .Q(n15285) );
  AND2X1 U16473 ( .IN1(n9047), .IN2(g29215), .Q(n15284) );
  AND2X1 U16474 ( .IN1(n15286), .IN2(n15287), .Q(g24241) );
  INVX0 U16475 ( .INP(n15288), .ZN(n15287) );
  AND2X1 U16476 ( .IN1(n15289), .IN2(n5622), .Q(n15288) );
  OR2X1 U16477 ( .IN1(n5622), .IN2(n15289), .Q(n15286) );
  OR2X1 U16478 ( .IN1(n9132), .IN2(n15290), .Q(n15289) );
  OR2X1 U16479 ( .IN1(n15291), .IN2(n15292), .Q(g24240) );
  AND2X1 U16480 ( .IN1(n15293), .IN2(n9024), .Q(n15292) );
  OR2X1 U16481 ( .IN1(n15294), .IN2(n15295), .Q(n15293) );
  AND4X1 U16482 ( .IN1(n8747), .IN2(n14944), .IN3(n8748), .IN4(n15290), .Q(
        n15295) );
  INVX0 U16483 ( .INP(n15296), .ZN(n15294) );
  OR2X1 U16484 ( .IN1(n15290), .IN2(n15297), .Q(n15296) );
  AND3X1 U16485 ( .IN1(n14944), .IN2(n8747), .IN3(n8748), .Q(n15297) );
  AND3X1 U16486 ( .IN1(n5622), .IN2(n5304), .IN3(n5392), .Q(n14944) );
  OR3X1 U16487 ( .IN1(n4837), .IN2(n15298), .IN3(n14550), .Q(n15290) );
  AND2X1 U16488 ( .IN1(n15299), .IN2(n15300), .Q(n15298) );
  OR2X1 U16489 ( .IN1(n5320), .IN2(g1236), .Q(n15300) );
  OR2X1 U16490 ( .IN1(n8359), .IN2(g979), .Q(n15299) );
  AND2X1 U16491 ( .IN1(n9142), .IN2(g996), .Q(n15291) );
  OR3X1 U16492 ( .IN1(n15301), .IN2(n15302), .IN3(n15303), .Q(g24239) );
  AND2X1 U16493 ( .IN1(n11500), .IN2(g17400), .Q(n15303) );
  AND2X1 U16494 ( .IN1(n9142), .IN2(g1246), .Q(n15302) );
  AND3X1 U16495 ( .IN1(n8698), .IN2(g10500), .IN3(n9059), .Q(n15301) );
  AND3X1 U16496 ( .IN1(n8699), .IN2(n8698), .IN3(n15304), .Q(g24238) );
  AND3X1 U16497 ( .IN1(n9053), .IN2(n8841), .IN3(n15305), .Q(n15304) );
  INVX0 U16498 ( .INP(n15306), .ZN(n15305) );
  AND3X1 U16499 ( .IN1(n15307), .IN2(n14920), .IN3(test_so76), .Q(n15306) );
  INVX0 U16500 ( .INP(n14921), .ZN(n14920) );
  OR2X1 U16501 ( .IN1(n8730), .IN2(n9483), .Q(n14921) );
  OR2X1 U16502 ( .IN1(n5547), .IN2(n8543), .Q(n9483) );
  OR2X1 U16503 ( .IN1(n14550), .IN2(n4837), .Q(n15307) );
  OR2X1 U16504 ( .IN1(test_so20), .IN2(g1008), .Q(n4837) );
  OR2X1 U16505 ( .IN1(n13124), .IN2(n14249), .Q(n14550) );
  INVX0 U16506 ( .INP(n14247), .ZN(n14249) );
  OR2X1 U16507 ( .IN1(n15308), .IN2(n15309), .Q(n14247) );
  AND2X1 U16508 ( .IN1(n5320), .IN2(g996), .Q(n15309) );
  AND2X1 U16509 ( .IN1(n8373), .IN2(g979), .Q(n15308) );
  AND2X1 U16510 ( .IN1(n5320), .IN2(n5622), .Q(n13124) );
  OR2X1 U16511 ( .IN1(n15310), .IN2(n15311), .Q(g24237) );
  AND2X1 U16512 ( .IN1(n15312), .IN2(n9024), .Q(n15311) );
  OR2X1 U16513 ( .IN1(n15313), .IN2(n15314), .Q(n15312) );
  AND2X1 U16514 ( .IN1(g7916), .IN2(g1178), .Q(n15314) );
  AND2X1 U16515 ( .IN1(n5304), .IN2(g1189), .Q(n15313) );
  AND2X1 U16516 ( .IN1(n9142), .IN2(g962), .Q(n15310) );
  OR2X1 U16517 ( .IN1(n15315), .IN2(n15316), .Q(g24236) );
  AND2X1 U16518 ( .IN1(n15317), .IN2(n9024), .Q(n15316) );
  OR2X1 U16519 ( .IN1(n15318), .IN2(n15319), .Q(n15317) );
  AND2X1 U16520 ( .IN1(g7916), .IN2(g996), .Q(n15319) );
  AND2X1 U16521 ( .IN1(n5304), .IN2(g1178), .Q(n15318) );
  AND2X1 U16522 ( .IN1(n9142), .IN2(g1183), .Q(n15315) );
  OR2X1 U16523 ( .IN1(n15320), .IN2(n15321), .Q(g24235) );
  AND2X1 U16524 ( .IN1(n15322), .IN2(g1152), .Q(n15321) );
  AND2X1 U16525 ( .IN1(test_so7), .IN2(n13659), .Q(n15320) );
  OR2X1 U16526 ( .IN1(n15323), .IN2(n15324), .Q(g24234) );
  AND2X1 U16527 ( .IN1(n15322), .IN2(g1146), .Q(n15324) );
  AND2X1 U16528 ( .IN1(n13659), .IN2(g1152), .Q(n15323) );
  OR2X1 U16529 ( .IN1(n15325), .IN2(n15326), .Q(g24233) );
  AND2X1 U16530 ( .IN1(n15327), .IN2(g1146), .Q(n15326) );
  OR2X1 U16531 ( .IN1(n15328), .IN2(n13659), .Q(n15327) );
  INVX0 U16532 ( .INP(n15322), .ZN(n13659) );
  OR2X1 U16533 ( .IN1(n9131), .IN2(n13664), .Q(n15322) );
  AND2X1 U16534 ( .IN1(n5618), .IN2(n9024), .Q(n15328) );
  AND3X1 U16535 ( .IN1(n9053), .IN2(n8820), .IN3(n13664), .Q(n15325) );
  AND3X1 U16536 ( .IN1(g13259), .IN2(n5363), .IN3(n5599), .Q(n13664) );
  OR3X1 U16537 ( .IN1(n15329), .IN2(n15330), .IN3(n15331), .Q(g24232) );
  AND2X1 U16538 ( .IN1(n11500), .IN2(g1052), .Q(n15331) );
  AND2X1 U16539 ( .IN1(n15332), .IN2(g1061), .Q(n15330) );
  AND2X1 U16540 ( .IN1(n15333), .IN2(n9024), .Q(n15329) );
  OR2X1 U16541 ( .IN1(n15334), .IN2(n5392), .Q(n15333) );
  AND2X1 U16542 ( .IN1(n5654), .IN2(n15332), .Q(n15334) );
  OR3X1 U16543 ( .IN1(n8756), .IN2(n9121), .IN3(g12919), .Q(n15332) );
  AND2X1 U16544 ( .IN1(n11500), .IN2(n8771), .Q(g24231) );
  AND2X1 U16545 ( .IN1(g12919), .IN2(n9024), .Q(n11500) );
  OR2X1 U16546 ( .IN1(n15335), .IN2(n15336), .Q(g24216) );
  AND2X1 U16547 ( .IN1(n15337), .IN2(g854), .Q(n15336) );
  AND2X1 U16548 ( .IN1(n13727), .IN2(g847), .Q(n15335) );
  OR2X1 U16549 ( .IN1(n15338), .IN2(n15339), .Q(g24215) );
  AND2X1 U16550 ( .IN1(n15340), .IN2(g703), .Q(n15339) );
  OR2X1 U16551 ( .IN1(n9131), .IN2(n15341), .Q(n15340) );
  AND2X1 U16552 ( .IN1(n5562), .IN2(n14599), .Q(n15341) );
  AND2X1 U16553 ( .IN1(g847), .IN2(n4948), .Q(n14599) );
  AND2X1 U16554 ( .IN1(n15342), .IN2(g837), .Q(n15338) );
  OR2X1 U16555 ( .IN1(n15343), .IN2(n13727), .Q(n15342) );
  AND3X1 U16556 ( .IN1(n15344), .IN2(n9050), .IN3(n15345), .Q(n15343) );
  OR2X1 U16557 ( .IN1(n5728), .IN2(n8545), .Q(n15345) );
  OR3X1 U16558 ( .IN1(n15346), .IN2(n15347), .IN3(n15348), .Q(g24214) );
  AND2X1 U16559 ( .IN1(n15349), .IN2(g703), .Q(n15348) );
  OR2X1 U16560 ( .IN1(n15350), .IN2(n13727), .Q(n15349) );
  AND2X1 U16561 ( .IN1(n15351), .IN2(n9024), .Q(n15350) );
  OR2X1 U16562 ( .IN1(n5562), .IN2(n15344), .Q(n15351) );
  OR2X1 U16563 ( .IN1(n5709), .IN2(n5733), .Q(n15344) );
  AND4X1 U16564 ( .IN1(n13728), .IN2(g822), .IN3(n15352), .IN4(n5709), .Q(
        n15347) );
  AND2X1 U16565 ( .IN1(g817), .IN2(g723), .Q(n15352) );
  AND2X1 U16566 ( .IN1(n9142), .IN2(g847), .Q(n15346) );
  OR2X1 U16567 ( .IN1(n15353), .IN2(g24212), .Q(g24213) );
  AND2X1 U16568 ( .IN1(n9142), .IN2(g753), .Q(n15353) );
  OR2X1 U16569 ( .IN1(n15354), .IN2(n15355), .Q(g24211) );
  AND2X1 U16570 ( .IN1(n9142), .IN2(g546), .Q(n15355) );
  AND2X1 U16571 ( .IN1(n2404), .IN2(n15356), .Q(n15354) );
  OR2X1 U16572 ( .IN1(n5520), .IN2(test_so41), .Q(n15356) );
  AND3X1 U16573 ( .IN1(n15357), .IN2(n9051), .IN3(n12052), .Q(g24210) );
  INVX0 U16574 ( .INP(n13144), .ZN(n12052) );
  OR3X1 U16575 ( .IN1(n8672), .IN2(n5287), .IN3(g513), .Q(n13144) );
  OR2X1 U16576 ( .IN1(n15358), .IN2(n15359), .Q(n15357) );
  AND2X1 U16577 ( .IN1(g174), .IN2(g168), .Q(n15359) );
  AND2X1 U16578 ( .IN1(test_so72), .IN2(n15360), .Q(n15358) );
  OR2X1 U16579 ( .IN1(g174), .IN2(g168), .Q(n15360) );
  OR2X1 U16580 ( .IN1(n15361), .IN2(n15362), .Q(g24209) );
  AND2X1 U16581 ( .IN1(n13728), .IN2(g446), .Q(n15362) );
  AND2X1 U16582 ( .IN1(n13727), .IN2(g417), .Q(n15361) );
  OR3X1 U16583 ( .IN1(n15363), .IN2(n15364), .IN3(n15365), .Q(g24208) );
  AND2X1 U16584 ( .IN1(n9142), .IN2(g424), .Q(n15365) );
  AND2X1 U16585 ( .IN1(n13728), .IN2(g246), .Q(n15364) );
  AND2X1 U16586 ( .IN1(n13727), .IN2(g475), .Q(n15363) );
  OR2X1 U16587 ( .IN1(n15366), .IN2(n15367), .Q(g24207) );
  AND2X1 U16588 ( .IN1(n15337), .IN2(g475), .Q(n15367) );
  AND2X1 U16589 ( .IN1(n13727), .IN2(g441), .Q(n15366) );
  OR2X1 U16590 ( .IN1(n15368), .IN2(n15369), .Q(g24206) );
  AND2X1 U16591 ( .IN1(n15337), .IN2(g441), .Q(n15369) );
  AND2X1 U16592 ( .IN1(n13727), .IN2(g437), .Q(n15368) );
  OR3X1 U16593 ( .IN1(n15370), .IN2(n15371), .IN3(n15372), .Q(g24205) );
  AND2X1 U16594 ( .IN1(n9142), .IN2(g437), .Q(n15372) );
  AND2X1 U16595 ( .IN1(n13728), .IN2(g269), .Q(n15371) );
  AND2X1 U16596 ( .IN1(test_so23), .IN2(n13727), .Q(n15370) );
  OR2X1 U16597 ( .IN1(n15373), .IN2(n15374), .Q(g24204) );
  AND2X1 U16598 ( .IN1(test_so23), .IN2(n15337), .Q(n15374) );
  AND2X1 U16599 ( .IN1(n13727), .IN2(g429), .Q(n15373) );
  OR2X1 U16600 ( .IN1(n15375), .IN2(n15376), .Q(g24203) );
  AND2X1 U16601 ( .IN1(n15337), .IN2(g429), .Q(n15376) );
  AND2X1 U16602 ( .IN1(n13727), .IN2(g401), .Q(n15375) );
  OR2X1 U16603 ( .IN1(n15377), .IN2(n15378), .Q(g24202) );
  AND2X1 U16604 ( .IN1(n15337), .IN2(g411), .Q(n15378) );
  AND2X1 U16605 ( .IN1(n13727), .IN2(g424), .Q(n15377) );
  OR2X1 U16606 ( .IN1(n15379), .IN2(n15380), .Q(g24201) );
  AND2X1 U16607 ( .IN1(n15337), .IN2(g392), .Q(n15380) );
  AND2X1 U16608 ( .IN1(n13727), .IN2(g405), .Q(n15379) );
  OR3X1 U16609 ( .IN1(n15381), .IN2(n15382), .IN3(n15383), .Q(g24200) );
  AND2X1 U16610 ( .IN1(n9142), .IN2(g401), .Q(n15383) );
  AND2X1 U16611 ( .IN1(n13727), .IN2(g392), .Q(n15382) );
  INVX0 U16612 ( .INP(n15337), .ZN(n13727) );
  OR2X1 U16613 ( .IN1(n4948), .IN2(n9123), .Q(n15337) );
  AND3X1 U16614 ( .IN1(n5821), .IN2(g854), .IN3(n13728), .Q(n15381) );
  AND2X1 U16615 ( .IN1(n9046), .IN2(n4948), .Q(n13728) );
  AND2X1 U16616 ( .IN1(n8789), .IN2(n8679), .Q(g23190) );
  OR2X1 U16617 ( .IN1(n15384), .IN2(n15385), .Q(g21901) );
  AND2X1 U16618 ( .IN1(n15386), .IN2(n9023), .Q(n15385) );
  OR2X1 U16619 ( .IN1(n15387), .IN2(n15388), .Q(n15386) );
  AND2X1 U16620 ( .IN1(n5380), .IN2(n15389), .Q(n15388) );
  OR2X1 U16621 ( .IN1(n15390), .IN2(g8786), .Q(n15389) );
  AND4X1 U16622 ( .IN1(n8651), .IN2(n8650), .IN3(n8652), .IN4(n15391), .Q(
        n15390) );
  AND4X1 U16623 ( .IN1(DFF_480_n1), .IN2(DFF_909_n1), .IN3(n8649), .IN4(
        DFF_1234_n1), .Q(n15391) );
  AND2X1 U16624 ( .IN1(n5694), .IN2(g4180), .Q(n15387) );
  AND2X1 U16625 ( .IN1(n9142), .IN2(g2946), .Q(n15384) );
  OR2X1 U16626 ( .IN1(n15392), .IN2(n15393), .Q(g21900) );
  AND3X1 U16627 ( .IN1(n8750), .IN2(n8749), .IN3(n9066), .Q(n15393) );
  AND2X1 U16628 ( .IN1(n9142), .IN2(g4239), .Q(n15392) );
  AND2X1 U16629 ( .IN1(n15394), .IN2(n15395), .Q(g21899) );
  INVX0 U16630 ( .INP(n15396), .ZN(n15395) );
  AND2X1 U16631 ( .IN1(n15397), .IN2(n8540), .Q(n15396) );
  OR2X1 U16632 ( .IN1(n8540), .IN2(n15397), .Q(n15394) );
  OR2X1 U16633 ( .IN1(n8512), .IN2(n9122), .Q(n15397) );
  OR2X1 U16634 ( .IN1(n15398), .IN2(n15399), .Q(g21898) );
  INVX0 U16635 ( .INP(n15400), .ZN(n15399) );
  OR2X1 U16636 ( .IN1(n9008), .IN2(n8361), .Q(n15400) );
  AND2X1 U16637 ( .IN1(n8540), .IN2(n9023), .Q(n15398) );
  AND2X1 U16638 ( .IN1(n15401), .IN2(n15402), .Q(g21897) );
  INVX0 U16639 ( .INP(n15403), .ZN(n15402) );
  AND2X1 U16640 ( .IN1(n15404), .IN2(n8541), .Q(n15403) );
  OR2X1 U16641 ( .IN1(n8541), .IN2(n15404), .Q(n15401) );
  OR2X1 U16642 ( .IN1(n8513), .IN2(n9123), .Q(n15404) );
  OR2X1 U16643 ( .IN1(n15405), .IN2(n15406), .Q(g21896) );
  AND2X1 U16644 ( .IN1(n9142), .IN2(g4245), .Q(n15406) );
  AND2X1 U16645 ( .IN1(n8541), .IN2(n9023), .Q(n15405) );
  OR2X1 U16646 ( .IN1(n15407), .IN2(n15408), .Q(g21895) );
  AND2X1 U16647 ( .IN1(n15168), .IN2(g4269), .Q(n15408) );
  OR2X1 U16648 ( .IN1(n15409), .IN2(g21893), .Q(n15168) );
  AND2X1 U16649 ( .IN1(n5823), .IN2(n9023), .Q(n15409) );
  AND2X1 U16650 ( .IN1(n15410), .IN2(g4264), .Q(n15407) );
  OR2X1 U16651 ( .IN1(n9131), .IN2(n15411), .Q(n15410) );
  AND2X1 U16652 ( .IN1(n5763), .IN2(g4258), .Q(n15411) );
  OR2X1 U16653 ( .IN1(n15412), .IN2(n15413), .Q(g21894) );
  AND2X1 U16654 ( .IN1(g21893), .IN2(g4264), .Q(n15413) );
  AND2X1 U16655 ( .IN1(n15414), .IN2(g4258), .Q(n15412) );
  OR2X1 U16656 ( .IN1(n5823), .IN2(n9122), .Q(n15414) );
  AND2X1 U16657 ( .IN1(n9032), .IN2(n8758), .Q(g21893) );
  OR2X1 U16658 ( .IN1(n15415), .IN2(n15416), .Q(g21892) );
  AND2X1 U16659 ( .IN1(n9142), .IN2(g4273), .Q(n15416) );
  AND2X1 U16660 ( .IN1(n8354), .IN2(n9024), .Q(n15415) );
  OR2X1 U16661 ( .IN1(n15417), .IN2(n15418), .Q(g21891) );
  AND2X1 U16662 ( .IN1(n15175), .IN2(n9023), .Q(n15418) );
  OR2X1 U16663 ( .IN1(n15419), .IN2(n15420), .Q(n15175) );
  AND2X1 U16664 ( .IN1(n8515), .IN2(n5484), .Q(n15420) );
  AND2X1 U16665 ( .IN1(n8516), .IN2(g4253), .Q(n15419) );
  AND2X1 U16666 ( .IN1(n9143), .IN2(g4180), .Q(n15417) );
  AND2X1 U16667 ( .IN1(n9143), .IN2(n9240), .Q(g21727) );
  AND2X1 U16668 ( .IN1(n9155), .IN2(g2975), .Q(g18597) );
  INVX0 U16669 ( .INP(g5), .ZN(g12833) );
  OR2X1 U5116_U1 ( .IN1(g34783), .IN2(n338), .Q(g34221) );
  OR2X1 U5126_U1 ( .IN1(n1392), .IN2(n4896), .Q(n4895) );
  OR2X1 U5127_U1 ( .IN1(n4837), .IN2(n4921), .Q(n4920) );
  OR2X1 U5128_U1 ( .IN1(n2787), .IN2(n1256), .Q(n5045) );
  OR2X1 U5129_U1 ( .IN1(g559), .IN2(g9048), .Q(n4959) );
  INVX0 U5353_U2 ( .INP(n8809), .ZN(U5353_n1) );
  AND2X1 U5353_U1 ( .IN1(n5960), .IN2(U5353_n1), .Q(n4689) );
  INVX0 U5355_U2 ( .INP(n8804), .ZN(U5355_n1) );
  AND2X1 U5355_U1 ( .IN1(n5961), .IN2(U5355_n1), .Q(n4708) );
  INVX0 U5961_U2 ( .INP(n791), .ZN(U5961_n1) );
  AND2X1 U5961_U1 ( .IN1(n3593), .IN2(U5961_n1), .Q(n3595) );
  INVX0 U5962_U2 ( .INP(n1369), .ZN(U5962_n1) );
  AND2X1 U5962_U1 ( .IN1(n3574), .IN2(U5962_n1), .Q(n3576) );
  INVX0 U5963_U2 ( .INP(n1371), .ZN(U5963_n1) );
  AND2X1 U5963_U1 ( .IN1(n3517), .IN2(U5963_n1), .Q(n3519) );
  INVX0 U5964_U2 ( .INP(n1731), .ZN(U5964_n1) );
  AND2X1 U5964_U1 ( .IN1(n3628), .IN2(U5964_n1), .Q(n3630) );
  INVX0 U5965_U2 ( .INP(n1367), .ZN(U5965_n1) );
  AND2X1 U5965_U1 ( .IN1(n3555), .IN2(U5965_n1), .Q(n3557) );
  INVX0 U5966_U2 ( .INP(n795), .ZN(U5966_n1) );
  AND2X1 U5966_U1 ( .IN1(n3646), .IN2(U5966_n1), .Q(n3648) );
  INVX0 U5967_U2 ( .INP(n1373), .ZN(U5967_n1) );
  AND2X1 U5967_U1 ( .IN1(n3536), .IN2(U5967_n1), .Q(n3538) );
  INVX0 U5968_U2 ( .INP(n789), .ZN(U5968_n1) );
  AND2X1 U5968_U1 ( .IN1(n3611), .IN2(U5968_n1), .Q(n3613) );
  AND2X1 U6100_U2 ( .IN1(n3635), .IN2(U6100_n1), .Q(n4888) );
  INVX0 U6100_U1 ( .INP(n9136), .ZN(U6100_n1) );
  INVX0 U6211_U2 ( .INP(n1733), .ZN(U6211_n1) );
  AND2X1 U6211_U1 ( .IN1(n3623), .IN2(U6211_n1), .Q(n3622) );
  INVX0 U6212_U2 ( .INP(n790), .ZN(U6212_n1) );
  AND2X1 U6212_U1 ( .IN1(n3587), .IN2(U6212_n1), .Q(n3586) );
  INVX0 U6213_U2 ( .INP(n788), .ZN(U6213_n1) );
  AND2X1 U6213_U1 ( .IN1(n3605), .IN2(U6213_n1), .Q(n3604) );
  INVX0 U6214_U2 ( .INP(n1368), .ZN(U6214_n1) );
  AND2X1 U6214_U1 ( .IN1(n3568), .IN2(U6214_n1), .Q(n3567) );
  INVX0 U6215_U2 ( .INP(n1366), .ZN(U6215_n1) );
  AND2X1 U6215_U1 ( .IN1(n3549), .IN2(U6215_n1), .Q(n3548) );
  INVX0 U6216_U2 ( .INP(n1370), .ZN(U6216_n1) );
  AND2X1 U6216_U1 ( .IN1(n3512), .IN2(U6216_n1), .Q(n3511) );
  INVX0 U6217_U2 ( .INP(n1372), .ZN(U6217_n1) );
  AND2X1 U6217_U1 ( .IN1(n3531), .IN2(U6217_n1), .Q(n3530) );
  INVX0 U6218_U2 ( .INP(n794), .ZN(U6218_n1) );
  AND2X1 U6218_U1 ( .IN1(n3641), .IN2(U6218_n1), .Q(n3640) );
  INVX0 U6279_U2 ( .INP(n5337), .ZN(U6279_n1) );
  AND2X1 U6279_U1 ( .IN1(n4537), .IN2(U6279_n1), .Q(n4201) );
  INVX0 U6280_U2 ( .INP(n5336), .ZN(U6280_n1) );
  AND2X1 U6280_U1 ( .IN1(n4201), .IN2(U6280_n1), .Q(n3745) );
  INVX0 U6281_U2 ( .INP(n5294), .ZN(U6281_n1) );
  AND2X1 U6281_U1 ( .IN1(n3745), .IN2(U6281_n1), .Q(n3684) );
  INVX0 U6282_U2 ( .INP(n5552), .ZN(U6282_n1) );
  AND2X1 U6282_U1 ( .IN1(n3684), .IN2(U6282_n1), .Q(n3274) );
  INVX0 U6283_U2 ( .INP(n5472), .ZN(U6283_n1) );
  AND2X1 U6283_U1 ( .IN1(n3274), .IN2(U6283_n1), .Q(n2982) );
  INVX0 U6284_U2 ( .INP(n5476), .ZN(U6284_n1) );
  AND2X1 U6284_U1 ( .IN1(n2982), .IN2(U6284_n1), .Q(n2706) );
  INVX0 U6285_U2 ( .INP(n5550), .ZN(U6285_n1) );
  AND2X1 U6285_U1 ( .IN1(n2706), .IN2(U6285_n1), .Q(n2649) );
  INVX0 U6286_U2 ( .INP(n5473), .ZN(U6286_n1) );
  AND2X1 U6286_U1 ( .IN1(n2649), .IN2(U6286_n1), .Q(n2556) );
  INVX0 U6287_U2 ( .INP(n5475), .ZN(U6287_n1) );
  AND2X1 U6287_U1 ( .IN1(n2556), .IN2(U6287_n1), .Q(n2509) );
  INVX0 U6288_U2 ( .INP(n5474), .ZN(U6288_n1) );
  AND2X1 U6288_U1 ( .IN1(n2509), .IN2(U6288_n1), .Q(n2487) );
  INVX0 U6289_U2 ( .INP(n5339), .ZN(U6289_n1) );
  AND2X1 U6289_U1 ( .IN1(n2487), .IN2(U6289_n1), .Q(n2427) );
  INVX0 U6290_U2 ( .INP(n5672), .ZN(U6290_n1) );
  AND2X1 U6290_U1 ( .IN1(n2427), .IN2(U6290_n1), .Q(n2423) );
  INVX0 U6291_U2 ( .INP(n5335), .ZN(U6291_n1) );
  AND2X1 U6291_U1 ( .IN1(n4826), .IN2(U6291_n1), .Q(n4537) );
  AND2X1 U6292_U2 ( .IN1(n4959), .IN2(U6292_n1), .Q(n2421) );
  INVX0 U6292_U1 ( .INP(n9136), .ZN(U6292_n1) );
  AND2X1 U6338_U2 ( .IN1(n4210), .IN2(U6338_n1), .Q(n3765) );
  INVX0 U6338_U1 ( .INP(n9137), .ZN(U6338_n1) );
  INVX0 U6341_U2 ( .INP(n1151), .ZN(U6341_n1) );
  AND2X1 U6341_U1 ( .IN1(n3765), .IN2(U6341_n1), .Q(n3951) );
  INVX0 U6342_U2 ( .INP(n769), .ZN(U6342_n1) );
  AND2X1 U6342_U1 ( .IN1(n3765), .IN2(U6342_n1), .Q(n3774) );
  INVX0 U6343_U2 ( .INP(n1084), .ZN(U6343_n1) );
  AND2X1 U6343_U1 ( .IN1(n3765), .IN2(U6343_n1), .Q(n3842) );
  INVX0 U6344_U2 ( .INP(n1022), .ZN(U6344_n1) );
  AND2X1 U6344_U1 ( .IN1(n3765), .IN2(U6344_n1), .Q(n3808) );
  INVX0 U6345_U2 ( .INP(n764), .ZN(U6345_n1) );
  AND2X1 U6345_U1 ( .IN1(n3765), .IN2(U6345_n1), .Q(n3908) );
  INVX0 U6346_U2 ( .INP(n115), .ZN(U6346_n1) );
  AND2X1 U6346_U1 ( .IN1(n3765), .IN2(U6346_n1), .Q(n3984) );
  INVX0 U6347_U2 ( .INP(n528), .ZN(U6347_n1) );
  AND2X1 U6347_U1 ( .IN1(n3765), .IN2(U6347_n1), .Q(n3875) );
  INVX0 U6348_U2 ( .INP(n130), .ZN(U6348_n1) );
  AND2X1 U6348_U1 ( .IN1(n3765), .IN2(U6348_n1), .Q(n4015) );
  INVX0 U6349_U2 ( .INP(n3446), .ZN(U6349_n1) );
  AND2X1 U6349_U1 ( .IN1(n3765), .IN2(U6349_n1), .Q(n3914) );
  INVX0 U6350_U2 ( .INP(n3406), .ZN(U6350_n1) );
  AND2X1 U6350_U1 ( .IN1(n3765), .IN2(U6350_n1), .Q(n3780) );
  INVX0 U6351_U2 ( .INP(n3481), .ZN(U6351_n1) );
  AND2X1 U6351_U1 ( .IN1(n3765), .IN2(U6351_n1), .Q(n3957) );
  INVX0 U6352_U2 ( .INP(n3426), .ZN(U6352_n1) );
  AND2X1 U6352_U1 ( .IN1(n3765), .IN2(U6352_n1), .Q(n3848) );
  INVX0 U6353_U2 ( .INP(n3491), .ZN(U6353_n1) );
  AND2X1 U6353_U1 ( .IN1(n3765), .IN2(U6353_n1), .Q(n3990) );
  INVX0 U6354_U2 ( .INP(n3416), .ZN(U6354_n1) );
  AND2X1 U6354_U1 ( .IN1(n3765), .IN2(U6354_n1), .Q(n3814) );
  INVX0 U6355_U2 ( .INP(n3436), .ZN(U6355_n1) );
  AND2X1 U6355_U1 ( .IN1(n3765), .IN2(U6355_n1), .Q(n3881) );
  INVX0 U6356_U2 ( .INP(n3502), .ZN(U6356_n1) );
  AND2X1 U6356_U1 ( .IN1(n3765), .IN2(U6356_n1), .Q(n4022) );
  INVX0 U6357_U2 ( .INP(n3501), .ZN(U6357_n1) );
  AND2X1 U6357_U1 ( .IN1(n3765), .IN2(U6357_n1), .Q(n4027) );
  INVX0 U6358_U2 ( .INP(n3407), .ZN(U6358_n1) );
  AND2X1 U6358_U1 ( .IN1(n3765), .IN2(U6358_n1), .Q(n3785) );
  INVX0 U6359_U2 ( .INP(n3482), .ZN(U6359_n1) );
  AND2X1 U6359_U1 ( .IN1(n3765), .IN2(U6359_n1), .Q(n3962) );
  INVX0 U6360_U2 ( .INP(n3427), .ZN(U6360_n1) );
  AND2X1 U6360_U1 ( .IN1(n3765), .IN2(U6360_n1), .Q(n3853) );
  INVX0 U6361_U2 ( .INP(n3437), .ZN(U6361_n1) );
  AND2X1 U6361_U1 ( .IN1(n3765), .IN2(U6361_n1), .Q(n3886) );
  INVX0 U6362_U2 ( .INP(n3417), .ZN(U6362_n1) );
  AND2X1 U6362_U1 ( .IN1(n3765), .IN2(U6362_n1), .Q(n3819) );
  INVX0 U6363_U2 ( .INP(n3492), .ZN(U6363_n1) );
  AND2X1 U6363_U1 ( .IN1(n3765), .IN2(U6363_n1), .Q(n3995) );
  INVX0 U6364_U2 ( .INP(n3447), .ZN(U6364_n1) );
  AND2X1 U6364_U1 ( .IN1(n3765), .IN2(U6364_n1), .Q(n3919) );
  INVX0 U6365_U2 ( .INP(n5471), .ZN(U6365_n1) );
  AND2X1 U6365_U1 ( .IN1(n3682), .IN2(U6365_n1), .Q(n3272) );
  INVX0 U6366_U2 ( .INP(n5331), .ZN(U6366_n1) );
  AND2X1 U6366_U1 ( .IN1(n3272), .IN2(U6366_n1), .Q(n2980) );
  INVX0 U6367_U2 ( .INP(n5332), .ZN(U6367_n1) );
  AND2X1 U6367_U1 ( .IN1(n2980), .IN2(U6367_n1), .Q(n2704) );
  INVX0 U6368_U2 ( .INP(n5333), .ZN(U6368_n1) );
  AND2X1 U6368_U1 ( .IN1(n2704), .IN2(U6368_n1), .Q(n2647) );
  INVX0 U6369_U2 ( .INP(n5334), .ZN(U6369_n1) );
  AND2X1 U6369_U1 ( .IN1(n2647), .IN2(U6369_n1), .Q(n2554) );
  INVX0 U6370_U2 ( .INP(n5330), .ZN(U6370_n1) );
  AND2X1 U6370_U1 ( .IN1(n2554), .IN2(U6370_n1), .Q(n2507) );
  INVX0 U6371_U2 ( .INP(n5551), .ZN(U6371_n1) );
  AND2X1 U6371_U1 ( .IN1(n2507), .IN2(U6371_n1), .Q(n2485) );
  INVX0 U6372_U2 ( .INP(n5293), .ZN(U6372_n1) );
  AND2X1 U6372_U1 ( .IN1(n2485), .IN2(U6372_n1), .Q(n2425) );
  INVX0 U6373_U2 ( .INP(n5292), .ZN(U6373_n1) );
  AND2X1 U6373_U1 ( .IN1(n2425), .IN2(U6373_n1), .Q(n2419) );
  INVX0 U6374_U2 ( .INP(n5470), .ZN(U6374_n1) );
  AND2X1 U6374_U1 ( .IN1(n3743), .IN2(U6374_n1), .Q(n3682) );
  INVX0 U6375_U2 ( .INP(n5291), .ZN(U6375_n1) );
  AND2X1 U6375_U1 ( .IN1(n2419), .IN2(U6375_n1), .Q(n2405) );
  AND2X1 U6417_U2 ( .IN1(n4198), .IN2(U6417_n1), .Q(n2404) );
  INVX0 U6417_U1 ( .INP(n9136), .ZN(U6417_n1) );
  INVX0 U6446_U2 ( .INP(n1795), .ZN(U6446_n1) );
  AND2X1 U6446_U1 ( .IN1(g110), .IN2(U6446_n1), .Q(n3524) );
  INVX0 U6465_U2 ( .INP(n5600), .ZN(U6465_n1) );
  AND2X1 U6465_U1 ( .IN1(n797), .IN2(U6465_n1), .Q(n4388) );
  INVX0 U6497_U2 ( .INP(n3635), .ZN(U6497_n1) );
  AND2X1 U6497_U1 ( .IN1(n822), .IN2(U6497_n1), .Q(n3005) );
  AND2X1 U6523_U2 ( .IN1(n1039), .IN2(U6523_n1), .Q(n4945) );
  INVX0 U6523_U1 ( .INP(n9137), .ZN(U6523_n1) );
  INVX0 U6542_U2 ( .INP(n5300), .ZN(U6542_n1) );
  AND2X1 U6542_U1 ( .IN1(n822), .IN2(U6542_n1), .Q(n3525) );
  INVX0 U6552_U2 ( .INP(n5676), .ZN(U6552_n1) );
  AND2X1 U6552_U1 ( .IN1(n3281), .IN2(U6552_n1), .Q(n3277) );
  INVX0 U6553_U2 ( .INP(n5680), .ZN(U6553_n1) );
  AND2X1 U6553_U1 ( .IN1(n3276), .IN2(U6553_n1), .Q(n2989) );
  INVX0 U6554_U2 ( .INP(n5677), .ZN(U6554_n1) );
  AND2X1 U6554_U1 ( .IN1(n3277), .IN2(U6554_n1), .Q(n2991) );
  INVX0 U6555_U2 ( .INP(n5561), .ZN(U6555_n1) );
  AND2X1 U6555_U1 ( .IN1(n3687), .IN2(U6555_n1), .Q(n3281) );
  INVX0 U6556_U2 ( .INP(n5679), .ZN(U6556_n1) );
  AND2X1 U6556_U1 ( .IN1(n3279), .IN2(U6556_n1), .Q(n3276) );
  INVX0 U6559_U2 ( .INP(n5678), .ZN(U6559_n1) );
  AND2X1 U6559_U1 ( .IN1(n2991), .IN2(U6559_n1), .Q(n2710) );
  INVX0 U6560_U2 ( .INP(n5675), .ZN(U6560_n1) );
  AND2X1 U6560_U1 ( .IN1(n2989), .IN2(U6560_n1), .Q(n2707) );
  INVX0 U6561_U2 ( .INP(n5327), .ZN(U6561_n1) );
  AND2X1 U6561_U1 ( .IN1(n3174), .IN2(U6561_n1), .Q(n3116) );
  INVX0 U6570_U2 ( .INP(n5477), .ZN(U6570_n1) );
  AND2X1 U6570_U1 ( .IN1(n3362), .IN2(U6570_n1), .Q(n2527) );
  INVX0 U6911_U2 ( .INP(n985), .ZN(U6911_n1) );
  AND2X1 U6911_U1 ( .IN1(n3115), .IN2(U6911_n1), .Q(n3111) );
  INVX0 U6912_U2 ( .INP(n998), .ZN(U6912_n1) );
  AND2X1 U6912_U1 ( .IN1(n3115), .IN2(U6912_n1), .Q(n3131) );
  INVX0 U6917_U2 ( .INP(n5350), .ZN(U6917_n1) );
  AND2X1 U6917_U1 ( .IN1(n3933), .IN2(U6917_n1), .Q(n3799) );
  INVX0 U6926_U2 ( .INP(n5674), .ZN(U6926_n1) );
  AND2X1 U6926_U1 ( .IN1(n3664), .IN2(U6926_n1), .Q(n3662) );
  INVX0 U6927_U2 ( .INP(n5673), .ZN(U6927_n1) );
  AND2X1 U6927_U1 ( .IN1(n3673), .IN2(U6927_n1), .Q(n3671) );
  INVX0 U6929_U2 ( .INP(n1122), .ZN(U6929_n1) );
  AND2X1 U6929_U1 ( .IN1(n3505), .IN2(U6929_n1), .Q(n2790) );
  INVX0 U6931_U2 ( .INP(n5554), .ZN(U6931_n1) );
  AND2X1 U6931_U1 ( .IN1(n4490), .IN2(U6931_n1), .Q(n4178) );
  INVX0 U6932_U2 ( .INP(n5555), .ZN(U6932_n1) );
  AND2X1 U6932_U1 ( .IN1(n4514), .IN2(U6932_n1), .Q(n4196) );
  INVX0 U6933_U2 ( .INP(n5558), .ZN(U6933_n1) );
  AND2X1 U6933_U1 ( .IN1(n4178), .IN2(U6933_n1), .Q(n3736) );
  INVX0 U6934_U2 ( .INP(n5559), .ZN(U6934_n1) );
  AND2X1 U6934_U1 ( .IN1(n4196), .IN2(U6934_n1), .Q(n3741) );
  INVX0 U6935_U2 ( .INP(n5553), .ZN(U6935_n1) );
  AND2X1 U6935_U1 ( .IN1(n3736), .IN2(U6935_n1), .Q(n3664) );
  INVX0 U6936_U2 ( .INP(n5560), .ZN(U6936_n1) );
  AND2X1 U6936_U1 ( .IN1(n3741), .IN2(U6936_n1), .Q(n3673) );
  INVX0 U6937_U2 ( .INP(n5303), .ZN(U6937_n1) );
  AND2X1 U6937_U1 ( .IN1(n141), .IN2(U6937_n1), .Q(n2598) );
  INVX0 U6938_U2 ( .INP(n5556), .ZN(U6938_n1) );
  AND2X1 U6938_U1 ( .IN1(n4804), .IN2(U6938_n1), .Q(n4490) );
  INVX0 U6939_U2 ( .INP(n5557), .ZN(U6939_n1) );
  AND2X1 U6939_U1 ( .IN1(n4811), .IN2(U6939_n1), .Q(n4514) );
  INVX0 U6940_U2 ( .INP(n5422), .ZN(U6940_n1) );
  AND2X1 U6940_U1 ( .IN1(n4814), .IN2(U6940_n1), .Q(n4519) );
  INVX0 U6941_U2 ( .INP(n5323), .ZN(U6941_n1) );
  AND2X1 U6941_U1 ( .IN1(n2607), .IN2(U6941_n1), .Q(n2594) );
  INVX0 U6944_U2 ( .INP(n5348), .ZN(U6944_n1) );
  AND2X1 U6944_U1 ( .IN1(n3084), .IN2(U6944_n1), .Q(n3033) );
  INVX0 U6950_U2 ( .INP(n5365), .ZN(U6950_n1) );
  AND2X1 U6950_U1 ( .IN1(n2598), .IN2(U6950_n1), .Q(n2590) );
  INVX0 U6954_U2 ( .INP(n998), .ZN(U6954_n1) );
  AND2X1 U6954_U1 ( .IN1(n724), .IN2(U6954_n1), .Q(n3125) );
  INVX0 U6955_U2 ( .INP(n985), .ZN(U6955_n1) );
  AND2X1 U6955_U1 ( .IN1(n705), .IN2(U6955_n1), .Q(n3105) );
  INVX0 U6956_U2 ( .INP(n997), .ZN(U6956_n1) );
  AND2X1 U6956_U1 ( .IN1(n388), .IN2(U6956_n1), .Q(n3145) );
  INVX0 U6957_U2 ( .INP(n987), .ZN(U6957_n1) );
  AND2X1 U6957_U1 ( .IN1(n719), .IN2(U6957_n1), .Q(n3164) );
  INVX0 U7174_U2 ( .INP(n5288), .ZN(U7174_n1) );
  AND2X1 U7174_U1 ( .IN1(n2423), .IN2(U7174_n1), .Q(n2422) );
  INVX0 U7248_U2 ( .INP(g1536), .ZN(U7248_n1) );
  AND2X1 U7248_U1 ( .IN1(n4172), .IN2(U7248_n1), .Q(n4173) );
  INVX0 U7249_U2 ( .INP(g1193), .ZN(U7249_n1) );
  AND2X1 U7249_U1 ( .IN1(n4190), .IN2(U7249_n1), .Q(n4191) );
  INVX0 U7402_U2 ( .INP(n561), .ZN(U7402_n1) );
  AND2X1 U7402_U1 ( .IN1(n4034), .IN2(U7402_n1), .Q(n4037) );
  INVX0 U7405_U2 ( .INP(n562), .ZN(U7405_n1) );
  AND2X1 U7405_U1 ( .IN1(n4034), .IN2(U7405_n1), .Q(n4039) );
  INVX0 U7413_U2 ( .INP(n844), .ZN(U7413_n1) );
  AND2X1 U7413_U1 ( .IN1(n3969), .IN2(U7413_n1), .Q(n3972) );
  INVX0 U7416_U2 ( .INP(n232), .ZN(U7416_n1) );
  AND2X1 U7416_U1 ( .IN1(n3926), .IN2(U7416_n1), .Q(n3929) );
  INVX0 U7427_U2 ( .INP(n736), .ZN(U7427_n1) );
  AND2X1 U7427_U1 ( .IN1(n3860), .IN2(U7427_n1), .Q(n3863) );
  INVX0 U7438_U2 ( .INP(n471), .ZN(U7438_n1) );
  AND2X1 U7438_U1 ( .IN1(n4002), .IN2(U7438_n1), .Q(n4003) );
  INVX0 U7449_U2 ( .INP(n563), .ZN(U7449_n1) );
  AND2X1 U7449_U1 ( .IN1(n4034), .IN2(U7449_n1), .Q(n4032) );
  INVX0 U7455_U2 ( .INP(n564), .ZN(U7455_n1) );
  AND2X1 U7455_U1 ( .IN1(n4034), .IN2(U7455_n1), .Q(n4035) );
  INVX0 U7464_U2 ( .INP(n1418), .ZN(U7464_n1) );
  AND2X1 U7464_U1 ( .IN1(n3792), .IN2(U7464_n1), .Q(n3797) );
  INVX0 U7467_U2 ( .INP(n1422), .ZN(U7467_n1) );
  AND2X1 U7467_U1 ( .IN1(n3792), .IN2(U7467_n1), .Q(n3790) );
  INVX0 U7482_U2 ( .INP(n1416), .ZN(U7482_n1) );
  AND2X1 U7482_U1 ( .IN1(n3792), .IN2(U7482_n1), .Q(n3795) );
  INVX0 U7492_U2 ( .INP(n945), .ZN(U7492_n1) );
  AND2X1 U7492_U1 ( .IN1(n3893), .IN2(U7492_n1), .Q(n3891) );
  INVX0 U7513_U2 ( .INP(n55), .ZN(U7513_n1) );
  AND2X1 U7513_U1 ( .IN1(n3826), .IN2(U7513_n1), .Q(n3827) );
  INVX0 U7516_U2 ( .INP(n943), .ZN(U7516_n1) );
  AND2X1 U7516_U1 ( .IN1(n3893), .IN2(U7516_n1), .Q(n3896) );
  INVX0 U7549_U2 ( .INP(n465), .ZN(U7549_n1) );
  AND2X1 U7549_U1 ( .IN1(n4002), .IN2(U7549_n1), .Q(n4007) );
  INVX0 U7561_U2 ( .INP(n225), .ZN(U7561_n1) );
  AND2X1 U7561_U1 ( .IN1(n3926), .IN2(U7561_n1), .Q(n3931) );
  INVX0 U7574_U2 ( .INP(n1423), .ZN(U7574_n1) );
  AND2X1 U7574_U1 ( .IN1(n3792), .IN2(U7574_n1), .Q(n3793) );
  INVX0 U7577_U2 ( .INP(n231), .ZN(U7577_n1) );
  AND2X1 U7577_U1 ( .IN1(n3926), .IN2(U7577_n1), .Q(n3924) );
  INVX0 U7585_U2 ( .INP(n57), .ZN(U7585_n1) );
  AND2X1 U7585_U1 ( .IN1(n3826), .IN2(U7585_n1), .Q(n3831) );
  INVX0 U7595_U2 ( .INP(n93), .ZN(U7595_n1) );
  AND2X1 U7595_U1 ( .IN1(n3826), .IN2(U7595_n1), .Q(n3829) );
  INVX0 U7614_U2 ( .INP(n223), .ZN(U7614_n1) );
  AND2X1 U7614_U1 ( .IN1(n3926), .IN2(U7614_n1), .Q(n3927) );
  INVX0 U7621_U2 ( .INP(n839), .ZN(U7621_n1) );
  AND2X1 U7621_U1 ( .IN1(n3969), .IN2(U7621_n1), .Q(n3974) );
  INVX0 U7629_U2 ( .INP(n944), .ZN(U7629_n1) );
  AND2X1 U7629_U1 ( .IN1(n3893), .IN2(U7629_n1), .Q(n3898) );
  INVX0 U7636_U2 ( .INP(n837), .ZN(U7636_n1) );
  AND2X1 U7636_U1 ( .IN1(n3969), .IN2(U7636_n1), .Q(n3970) );
  INVX0 U7639_U2 ( .INP(n470), .ZN(U7639_n1) );
  AND2X1 U7639_U1 ( .IN1(n4002), .IN2(U7639_n1), .Q(n4000) );
  INVX0 U7649_U2 ( .INP(n731), .ZN(U7649_n1) );
  AND2X1 U7649_U1 ( .IN1(n3860), .IN2(U7649_n1), .Q(n3865) );
  INVX0 U7652_U2 ( .INP(n729), .ZN(U7652_n1) );
  AND2X1 U7652_U1 ( .IN1(n3860), .IN2(U7652_n1), .Q(n3861) );
  INVX0 U7668_U2 ( .INP(n92), .ZN(U7668_n1) );
  AND2X1 U7668_U1 ( .IN1(n3826), .IN2(U7668_n1), .Q(n3824) );
  INVX0 U7673_U2 ( .INP(n946), .ZN(U7673_n1) );
  AND2X1 U7673_U1 ( .IN1(n3893), .IN2(U7673_n1), .Q(n3894) );
  INVX0 U7690_U2 ( .INP(n843), .ZN(U7690_n1) );
  AND2X1 U7690_U1 ( .IN1(n3969), .IN2(U7690_n1), .Q(n3967) );
  INVX0 U7707_U2 ( .INP(n735), .ZN(U7707_n1) );
  AND2X1 U7707_U1 ( .IN1(n3860), .IN2(U7707_n1), .Q(n3858) );
  INVX0 U7712_U2 ( .INP(n463), .ZN(U7712_n1) );
  AND2X1 U7712_U1 ( .IN1(n4002), .IN2(U7712_n1), .Q(n4005) );
  AND2X1 U7792_U2 ( .IN1(g952), .IN2(U7792_n1), .Q(n2505) );
  INVX0 U7792_U1 ( .INP(n9137), .ZN(U7792_n1) );
  AND2X1 U7794_U2 ( .IN1(g1296), .IN2(U7794_n1), .Q(n2499) );
  INVX0 U7794_U1 ( .INP(n9136), .ZN(U7794_n1) );
  INVX0 U7895_U2 ( .INP(g113), .ZN(U7895_n1) );
  AND2X1 U7895_U1 ( .IN1(n2668), .IN2(U7895_n1), .Q(n2760) );
  INVX0 U7897_U2 ( .INP(g31), .ZN(U7897_n1) );
  AND2X1 U7897_U1 ( .IN1(g6), .IN2(U7897_n1), .Q(n3395) );
  AND2X1 U7977_U2 ( .IN1(g661), .IN2(U7977_n1), .Q(n4956) );
  INVX0 U7977_U1 ( .INP(n9136), .ZN(U7977_n1) );
  INVX0 U8034_U2 ( .INP(n5612), .ZN(U8034_n1) );
  AND2X1 U8034_U1 ( .IN1(n1253), .IN2(U8034_n1), .Q(n5026) );
  INVX0 U8036_U2 ( .INP(n5340), .ZN(U8036_n1) );
  AND2X1 U8036_U1 ( .IN1(n3729), .IN2(U8036_n1), .Q(n3941) );
  INVX0 U8050_U2 ( .INP(g1367), .ZN(U8050_n1) );
  AND2X1 U8050_U1 ( .IN1(n217), .IN2(U8050_n1), .Q(n3733) );
  AND2X1 U8055_U2 ( .IN1(g1345), .IN2(U8055_n1), .Q(n4798) );
  INVX0 U8055_U1 ( .INP(n9137), .ZN(U8055_n1) );
  AND2X1 U8060_U2 ( .IN1(g1002), .IN2(U8060_n1), .Q(n4805) );
  INVX0 U8060_U1 ( .INP(n9136), .ZN(U8060_n1) );
  INVX0 U8070_U2 ( .INP(g1361), .ZN(U8070_n1) );
  AND2X1 U8070_U1 ( .IN1(n218), .IN2(U8070_n1), .Q(n4175) );
  INVX0 U8074_U2 ( .INP(g1018), .ZN(U8074_n1) );
  AND2X1 U8074_U1 ( .IN1(n581), .IN2(U8074_n1), .Q(n4193) );
  INVX0 U8088_U2 ( .INP(g1024), .ZN(U8088_n1) );
  AND2X1 U8088_U1 ( .IN1(n580), .IN2(U8088_n1), .Q(n3738) );
  INVX0 U8112_U2 ( .INP(n4523), .ZN(U8112_n1) );
  AND2X1 U8112_U1 ( .IN1(n4525), .IN2(U8112_n1), .Q(n4524) );
  INVX0 U8113_U2 ( .INP(n5751), .ZN(U8113_n1) );
  AND2X1 U8113_U1 ( .IN1(n4526), .IN2(U8113_n1), .Q(n4523) );
  INVX0 U8147_U2 ( .INP(n2573), .ZN(U8147_n1) );
  AND2X1 U8147_U1 ( .IN1(g4659), .IN2(U8147_n1), .Q(n2577) );
  INVX0 U8165_U2 ( .INP(n2563), .ZN(U8165_n1) );
  AND2X1 U8165_U1 ( .IN1(g4849), .IN2(U8165_n1), .Q(n2567) );
  INVX0 U8185_U2 ( .INP(g1046), .ZN(U8185_n1) );
  AND2X1 U8185_U1 ( .IN1(n865), .IN2(U8185_n1), .Q(n4938) );
  INVX0 U8192_U2 ( .INP(g1389), .ZN(U8192_n1) );
  AND2X1 U8192_U1 ( .IN1(n209), .IN2(U8192_n1), .Q(n4913) );
  INVX0 U8210_U2 ( .INP(n1253), .ZN(U8210_n1) );
  AND2X1 U8210_U1 ( .IN1(n4722), .IN2(U8210_n1), .Q(n4714) );
  INVX0 U8223_U2 ( .INP(n4516), .ZN(U8223_n1) );
  AND2X1 U8223_U1 ( .IN1(n4518), .IN2(U8223_n1), .Q(n4517) );
  INVX0 U8224_U2 ( .INP(n5728), .ZN(U8224_n1) );
  AND2X1 U8224_U1 ( .IN1(n4519), .IN2(U8224_n1), .Q(n4516) );
  AND2X1 U8281_U2 ( .IN1(n939), .IN2(U8281_n1), .Q(n5111) );
  INVX0 U8281_U1 ( .INP(n9137), .ZN(U8281_n1) );
  AND2X1 U8307_U2 ( .IN1(g29216), .IN2(U8307_n1), .Q(g26900) );
  INVX0 U8307_U1 ( .INP(n9137), .ZN(U8307_n1) );
  INVX0 U8974_U2 ( .INP(test_so25), .ZN(U8974_n1) );
  AND2X1 U8974_U1 ( .IN1(n3362), .IN2(U8974_n1), .Q(n2552) );
  INVX0 U8975_U2 ( .INP(g528), .ZN(U8975_n1) );
  AND2X1 U8975_U1 ( .IN1(n3174), .IN2(U8975_n1), .Q(n3195) );
  AND2X1 U9065_U2 ( .IN1(g4145), .IN2(U9065_n1), .Q(n4721) );
  INVX0 U9065_U1 ( .INP(n9137), .ZN(U9065_n1) );
  AND2X1 U9070_U2 ( .IN1(g2841), .IN2(U9070_n1), .Q(n3730) );
  INVX0 U9070_U1 ( .INP(n9137), .ZN(U9070_n1) );
  INVX0 U9075_U2 ( .INP(g9), .ZN(U9075_n1) );
  AND2X1 U9075_U1 ( .IN1(g19), .IN2(U9075_n1), .Q(n3362) );
  AND2X1 U9076_U2 ( .IN1(g113), .IN2(U9076_n1), .Q(g25694) );
  INVX0 U9076_U1 ( .INP(n9136), .ZN(U9076_n1) );
  AND2X1 U9080_U2 ( .IN1(n4305), .IN2(U9080_n1), .Q(g29277) );
  INVX0 U9080_U1 ( .INP(n9137), .ZN(U9080_n1) );
  AND2X1 U9084_U2 ( .IN1(g4423), .IN2(U9084_n1), .Q(g26953) );
  INVX0 U9084_U1 ( .INP(n9137), .ZN(U9084_n1) );
  AND2X1 U9085_U2 ( .IN1(g64), .IN2(U9085_n1), .Q(g24212) );
  INVX0 U9085_U1 ( .INP(n9137), .ZN(U9085_n1) );
  AND2X1 U9086_U2 ( .IN1(n4283), .IN2(U9086_n1), .Q(g29279) );
  INVX0 U9086_U1 ( .INP(n9136), .ZN(U9086_n1) );
  AND2X1 U9090_U2 ( .IN1(g125), .IN2(U9090_n1), .Q(g25688) );
  INVX0 U9090_U1 ( .INP(n9136), .ZN(U9090_n1) );
  INVX0 U9098_U2 ( .INP(n342), .ZN(U9098_n1) );
  AND2X1 U9098_U1 ( .IN1(g4681), .IN2(U9098_n1), .Q(g34028) );
  INVX0 U9099_U2 ( .INP(n2608), .ZN(U9099_n1) );
  AND2X1 U9099_U1 ( .IN1(n2595), .IN2(U9099_n1), .Q(g34449) );
  AND2X1 U9101_U2 ( .IN1(g6745), .IN2(U9101_n1), .Q(g26880) );
  INVX0 U9101_U1 ( .INP(n9137), .ZN(U9101_n1) );
  INVX0 U9107_U2 ( .INP(n8813), .ZN(U9107_n1) );
  AND2X1 U9107_U1 ( .IN1(n4448), .IN2(U9107_n1), .Q(n4447) );
  INVX0 U9111_U2 ( .INP(n8810), .ZN(U9111_n1) );
  AND2X1 U9111_U1 ( .IN1(n4403), .IN2(U9111_n1), .Q(n4402) );
  INVX0 U9116_U2 ( .INP(n8818), .ZN(U9116_n1) );
  AND2X1 U9116_U1 ( .IN1(n4426), .IN2(U9116_n1), .Q(n4425) );
  INVX0 U9120_U2 ( .INP(n8807), .ZN(U9120_n1) );
  AND2X1 U9120_U1 ( .IN1(n4437), .IN2(U9120_n1), .Q(n4436) );
  INVX0 U9124_U2 ( .INP(n8815), .ZN(U9124_n1) );
  AND2X1 U9124_U1 ( .IN1(n4392), .IN2(U9124_n1), .Q(n4391) );
  INVX0 U9128_U2 ( .INP(n8808), .ZN(U9128_n1) );
  AND2X1 U9128_U1 ( .IN1(n4380), .IN2(U9128_n1), .Q(n4379) );
  INVX0 U9132_U2 ( .INP(n8816), .ZN(U9132_n1) );
  AND2X1 U9132_U1 ( .IN1(n4415), .IN2(U9132_n1), .Q(n4414) );
  INVX0 U9136_U2 ( .INP(n8817), .ZN(U9136_n1) );
  AND2X1 U9136_U1 ( .IN1(n4459), .IN2(U9136_n1), .Q(n4458) );
  INVX0 U9315_U2 ( .INP(n5753), .ZN(U9315_n1) );
  AND2X1 U9315_U1 ( .IN1(n5016), .IN2(U9315_n1), .Q(n5014) );
  INVX0 U9453_U2 ( .INP(n8811), .ZN(U9453_n1) );
  AND2X1 U9453_U1 ( .IN1(n3065), .IN2(U9453_n1), .Q(n3064) );
  INVX0 U9825_U2 ( .INP(n1795), .ZN(U9825_n1) );
  AND2X1 U9825_U1 ( .IN1(g112), .IN2(U9825_n1), .Q(n3115) );
  INVX0 U9886_U2 ( .INP(n5121), .ZN(U9886_n1) );
  AND2X1 U9886_U1 ( .IN1(g370), .IN2(U9886_n1), .Q(n4948) );
  INVX0 U9927_U2 ( .INP(g4098), .ZN(U9927_n1) );
  AND2X1 U9927_U1 ( .IN1(n3933), .IN2(U9927_n1), .Q(n3833) );
  INVX0 U9953_U2 ( .INP(n158), .ZN(U9953_n1) );
  AND2X1 U9953_U1 ( .IN1(g671), .IN2(U9953_n1), .Q(n4526) );
  INVX0 U9957_U2 ( .INP(n5283), .ZN(U9957_n1) );
  AND2X1 U9957_U1 ( .IN1(g4843), .IN2(U9957_n1), .Q(n2563) );
  INVX0 U9958_U2 ( .INP(n5656), .ZN(U9958_n1) );
  AND2X1 U9958_U1 ( .IN1(test_so19), .IN2(U9958_n1), .Q(n2573) );
  INVX0 U9968_U2 ( .INP(g4358), .ZN(U9968_n1) );
  AND2X1 U9968_U1 ( .IN1(n3084), .IN2(U9968_n1), .Q(n3023) );
  INVX0 U9972_U2 ( .INP(n4535), .ZN(U9972_n1) );
  AND2X1 U9972_U1 ( .IN1(g681), .IN2(U9972_n1), .Q(n5112) );
  INVX0 U9992_U2 ( .INP(n517), .ZN(U9992_n1) );
  AND2X1 U9992_U1 ( .IN1(n3675), .IN2(U9992_n1), .Q(n2644) );
  INVX0 U10314_U2 ( .INP(g686), .ZN(U10314_n1) );
  AND2X1 U10314_U1 ( .IN1(g667), .IN2(U10314_n1), .Q(n4962) );
  INVX0 U10318_U2 ( .INP(n5681), .ZN(U10318_n1) );
  AND2X1 U10318_U1 ( .IN1(g5092), .IN2(U10318_n1), .Q(n5016) );
endmodule

