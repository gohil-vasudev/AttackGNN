module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n639_, new_n484_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n883_, new_n1005_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n676_, new_n970_, new_n466_, new_n262_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n932_, new_n878_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n493_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n407_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n933_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n765_, new_n405_;

not g000 ( new_n202_, keyIn_0_55 );
xnor g001 ( new_n203_, N65, N69 );
xnor g002 ( new_n204_, new_n203_, keyIn_0_8 );
not g003 ( new_n205_, keyIn_0_9 );
xnor g004 ( new_n206_, N73, N77 );
xnor g005 ( new_n207_, new_n206_, new_n205_ );
xnor g006 ( new_n208_, new_n204_, new_n207_ );
xnor g007 ( new_n209_, new_n208_, keyIn_0_32 );
xor g008 ( new_n210_, N81, N85 );
xnor g009 ( new_n211_, new_n210_, keyIn_0_10 );
xnor g010 ( new_n212_, N89, N93 );
xnor g011 ( new_n213_, new_n212_, keyIn_0_11 );
xnor g012 ( new_n214_, new_n211_, new_n213_ );
xnor g013 ( new_n215_, new_n214_, keyIn_0_33 );
xnor g014 ( new_n216_, new_n215_, new_n209_ );
xnor g015 ( new_n217_, new_n216_, keyIn_0_43 );
nand g016 ( new_n218_, N129, N137 );
xnor g017 ( new_n219_, new_n217_, new_n218_ );
xnor g018 ( new_n220_, new_n219_, keyIn_0_47 );
xnor g019 ( new_n221_, N33, N49 );
xnor g020 ( new_n222_, N1, N17 );
xnor g021 ( new_n223_, new_n221_, new_n222_ );
xnor g022 ( new_n224_, new_n220_, new_n223_ );
xnor g023 ( new_n225_, new_n224_, new_n202_ );
xnor g024 ( new_n226_, N97, N101 );
xnor g025 ( new_n227_, new_n226_, keyIn_0_12 );
xnor g026 ( new_n228_, N105, N109 );
xnor g027 ( new_n229_, new_n228_, keyIn_0_13 );
xnor g028 ( new_n230_, new_n227_, new_n229_ );
xnor g029 ( new_n231_, new_n230_, keyIn_0_34 );
xnor g030 ( new_n232_, new_n209_, new_n231_ );
xnor g031 ( new_n233_, new_n232_, keyIn_0_45 );
xnor g032 ( new_n234_, new_n233_, keyIn_0_16 );
nand g033 ( new_n235_, N131, N137 );
not g034 ( new_n236_, new_n235_ );
xnor g035 ( new_n237_, new_n234_, new_n236_ );
nand g036 ( new_n238_, new_n237_, keyIn_0_49 );
not g037 ( new_n239_, keyIn_0_49 );
xnor g038 ( new_n240_, new_n234_, new_n235_ );
nand g039 ( new_n241_, new_n240_, new_n239_ );
nand g040 ( new_n242_, new_n238_, new_n241_ );
xnor g041 ( new_n243_, N41, N57 );
xnor g042 ( new_n244_, new_n243_, keyIn_0_22 );
xnor g043 ( new_n245_, N9, N25 );
xnor g044 ( new_n246_, new_n245_, keyIn_0_21 );
xnor g045 ( new_n247_, new_n244_, new_n246_ );
xor g046 ( new_n248_, new_n247_, keyIn_0_36 );
not g047 ( new_n249_, new_n248_ );
xnor g048 ( new_n250_, new_n242_, new_n249_ );
nand g049 ( new_n251_, new_n250_, keyIn_0_57 );
not g050 ( new_n252_, keyIn_0_57 );
xnor g051 ( new_n253_, new_n242_, new_n248_ );
nand g052 ( new_n254_, new_n253_, new_n252_ );
nand g053 ( new_n255_, new_n251_, new_n254_ );
not g054 ( new_n256_, keyIn_0_56 );
not g055 ( new_n257_, keyIn_0_35 );
not g056 ( new_n258_, keyIn_0_15 );
xnor g057 ( new_n259_, N121, N125 );
xnor g058 ( new_n260_, new_n259_, new_n258_ );
xnor g059 ( new_n261_, N113, N117 );
xnor g060 ( new_n262_, new_n261_, keyIn_0_14 );
xnor g061 ( new_n263_, new_n260_, new_n262_ );
xnor g062 ( new_n264_, new_n263_, new_n257_ );
xnor g063 ( new_n265_, new_n231_, new_n264_ );
xnor g064 ( new_n266_, new_n265_, keyIn_0_44 );
nand g065 ( new_n267_, N130, N137 );
xor g066 ( new_n268_, new_n266_, new_n267_ );
xnor g067 ( new_n269_, new_n268_, keyIn_0_48 );
xnor g068 ( new_n270_, N37, N53 );
xnor g069 ( new_n271_, N5, N21 );
xnor g070 ( new_n272_, new_n270_, new_n271_ );
not g071 ( new_n273_, new_n272_ );
nand g072 ( new_n274_, new_n269_, new_n273_ );
not g073 ( new_n275_, keyIn_0_48 );
xnor g074 ( new_n276_, new_n268_, new_n275_ );
nand g075 ( new_n277_, new_n276_, new_n272_ );
nand g076 ( new_n278_, new_n274_, new_n277_ );
xnor g077 ( new_n279_, new_n278_, new_n256_ );
xnor g078 ( new_n280_, new_n215_, new_n264_ );
xnor g079 ( new_n281_, new_n280_, keyIn_0_46 );
nand g080 ( new_n282_, N132, N137 );
xnor g081 ( new_n283_, new_n281_, new_n282_ );
xnor g082 ( new_n284_, new_n283_, keyIn_0_50 );
xor g083 ( new_n285_, N13, N29 );
xnor g084 ( new_n286_, new_n285_, keyIn_0_23 );
xnor g085 ( new_n287_, N45, N61 );
xnor g086 ( new_n288_, new_n286_, new_n287_ );
xnor g087 ( new_n289_, new_n284_, new_n288_ );
xnor g088 ( new_n290_, new_n289_, keyIn_0_58 );
nor g089 ( new_n291_, new_n279_, new_n290_ );
nand g090 ( new_n292_, new_n255_, new_n291_ );
nor g091 ( new_n293_, new_n255_, new_n291_ );
not g092 ( new_n294_, new_n225_ );
nand g093 ( new_n295_, new_n279_, new_n290_ );
nand g094 ( new_n296_, new_n295_, new_n294_ );
nor g095 ( new_n297_, new_n293_, new_n296_ );
nand g096 ( new_n298_, new_n297_, new_n292_ );
not g097 ( new_n299_, new_n255_ );
nand g098 ( new_n300_, new_n299_, keyIn_0_63 );
not g099 ( new_n301_, keyIn_0_63 );
nand g100 ( new_n302_, new_n255_, new_n301_ );
xnor g101 ( new_n303_, new_n278_, keyIn_0_56 );
nand g102 ( new_n304_, new_n303_, new_n225_ );
nor g103 ( new_n305_, new_n304_, new_n290_ );
and g104 ( new_n306_, new_n302_, new_n305_ );
nand g105 ( new_n307_, new_n306_, new_n300_ );
nand g106 ( new_n308_, new_n307_, new_n298_ );
not g107 ( new_n309_, keyIn_0_59 );
not g108 ( new_n310_, keyIn_0_29 );
not g109 ( new_n311_, N29 );
nand g110 ( new_n312_, new_n311_, N25 );
not g111 ( new_n313_, N25 );
nand g112 ( new_n314_, new_n313_, N29 );
nand g113 ( new_n315_, new_n312_, new_n314_ );
nand g114 ( new_n316_, new_n315_, keyIn_0_3 );
not g115 ( new_n317_, keyIn_0_3 );
xnor g116 ( new_n318_, N25, N29 );
nand g117 ( new_n319_, new_n318_, new_n317_ );
nand g118 ( new_n320_, new_n316_, new_n319_ );
xnor g119 ( new_n321_, N17, N21 );
nand g120 ( new_n322_, new_n321_, keyIn_0_2 );
not g121 ( new_n323_, keyIn_0_2 );
and g122 ( new_n324_, N17, N21 );
nor g123 ( new_n325_, N17, N21 );
nor g124 ( new_n326_, new_n324_, new_n325_ );
nand g125 ( new_n327_, new_n326_, new_n323_ );
nand g126 ( new_n328_, new_n327_, new_n322_ );
nand g127 ( new_n329_, new_n320_, new_n328_ );
and g128 ( new_n330_, new_n316_, new_n319_ );
and g129 ( new_n331_, new_n327_, new_n322_ );
nand g130 ( new_n332_, new_n330_, new_n331_ );
nand g131 ( new_n333_, new_n332_, new_n329_ );
nand g132 ( new_n334_, new_n333_, new_n310_ );
and g133 ( new_n335_, new_n320_, new_n328_ );
nor g134 ( new_n336_, new_n320_, new_n328_ );
nor g135 ( new_n337_, new_n335_, new_n336_ );
nand g136 ( new_n338_, new_n337_, keyIn_0_29 );
nand g137 ( new_n339_, new_n338_, new_n334_ );
xnor g138 ( new_n340_, N9, N13 );
nand g139 ( new_n341_, new_n340_, keyIn_0_1 );
not g140 ( new_n342_, keyIn_0_1 );
and g141 ( new_n343_, N9, N13 );
nor g142 ( new_n344_, N9, N13 );
nor g143 ( new_n345_, new_n343_, new_n344_ );
nand g144 ( new_n346_, new_n345_, new_n342_ );
nand g145 ( new_n347_, new_n346_, new_n341_ );
xnor g146 ( new_n348_, N1, N5 );
nand g147 ( new_n349_, new_n348_, keyIn_0_0 );
not g148 ( new_n350_, keyIn_0_0 );
and g149 ( new_n351_, N1, N5 );
nor g150 ( new_n352_, N1, N5 );
nor g151 ( new_n353_, new_n351_, new_n352_ );
nand g152 ( new_n354_, new_n353_, new_n350_ );
nand g153 ( new_n355_, new_n354_, new_n349_ );
nand g154 ( new_n356_, new_n347_, new_n355_ );
and g155 ( new_n357_, new_n346_, new_n341_ );
and g156 ( new_n358_, new_n354_, new_n349_ );
nand g157 ( new_n359_, new_n357_, new_n358_ );
nand g158 ( new_n360_, new_n359_, new_n356_ );
xnor g159 ( new_n361_, new_n360_, keyIn_0_28 );
nand g160 ( new_n362_, new_n361_, new_n339_ );
xnor g161 ( new_n363_, new_n333_, keyIn_0_29 );
not g162 ( new_n364_, keyIn_0_28 );
xnor g163 ( new_n365_, new_n360_, new_n364_ );
nand g164 ( new_n366_, new_n363_, new_n365_ );
nand g165 ( new_n367_, new_n366_, new_n362_ );
nand g166 ( new_n368_, new_n367_, keyIn_0_39 );
not g167 ( new_n369_, keyIn_0_39 );
xnor g168 ( new_n370_, new_n365_, new_n339_ );
nand g169 ( new_n371_, new_n370_, new_n369_ );
nand g170 ( new_n372_, new_n371_, new_n368_ );
nand g171 ( new_n373_, N133, N137 );
xnor g172 ( new_n374_, new_n373_, keyIn_0_17 );
not g173 ( new_n375_, new_n374_ );
nand g174 ( new_n376_, new_n372_, new_n375_ );
xnor g175 ( new_n377_, new_n367_, new_n369_ );
nand g176 ( new_n378_, new_n377_, new_n374_ );
nand g177 ( new_n379_, new_n378_, new_n376_ );
nand g178 ( new_n380_, new_n379_, keyIn_0_51 );
not g179 ( new_n381_, keyIn_0_51 );
xnor g180 ( new_n382_, new_n372_, new_n374_ );
nand g181 ( new_n383_, new_n382_, new_n381_ );
nand g182 ( new_n384_, new_n383_, new_n380_ );
xor g183 ( new_n385_, N97, N113 );
xnor g184 ( new_n386_, N65, N81 );
xnor g185 ( new_n387_, new_n385_, new_n386_ );
not g186 ( new_n388_, new_n387_ );
nand g187 ( new_n389_, new_n384_, new_n388_ );
xnor g188 ( new_n390_, new_n379_, new_n381_ );
nand g189 ( new_n391_, new_n390_, new_n387_ );
nand g190 ( new_n392_, new_n391_, new_n389_ );
xnor g191 ( new_n393_, new_n392_, new_n309_ );
not g192 ( new_n394_, keyIn_0_60 );
xnor g193 ( new_n395_, N49, N53 );
nand g194 ( new_n396_, new_n395_, keyIn_0_6 );
not g195 ( new_n397_, keyIn_0_6 );
and g196 ( new_n398_, N49, N53 );
nor g197 ( new_n399_, N49, N53 );
nor g198 ( new_n400_, new_n398_, new_n399_ );
nand g199 ( new_n401_, new_n400_, new_n397_ );
nand g200 ( new_n402_, new_n401_, new_n396_ );
xnor g201 ( new_n403_, N57, N61 );
nand g202 ( new_n404_, new_n403_, keyIn_0_7 );
not g203 ( new_n405_, keyIn_0_7 );
and g204 ( new_n406_, N57, N61 );
nor g205 ( new_n407_, N57, N61 );
nor g206 ( new_n408_, new_n406_, new_n407_ );
nand g207 ( new_n409_, new_n408_, new_n405_ );
nand g208 ( new_n410_, new_n409_, new_n404_ );
nand g209 ( new_n411_, new_n402_, new_n410_ );
and g210 ( new_n412_, new_n401_, new_n396_ );
xnor g211 ( new_n413_, new_n403_, new_n405_ );
nand g212 ( new_n414_, new_n412_, new_n413_ );
nand g213 ( new_n415_, new_n414_, new_n411_ );
xnor g214 ( new_n416_, new_n415_, keyIn_0_31 );
not g215 ( new_n417_, keyIn_0_30 );
not g216 ( new_n418_, keyIn_0_4 );
xnor g217 ( new_n419_, N33, N37 );
nand g218 ( new_n420_, new_n419_, new_n418_ );
and g219 ( new_n421_, N33, N37 );
nor g220 ( new_n422_, N33, N37 );
nor g221 ( new_n423_, new_n421_, new_n422_ );
nand g222 ( new_n424_, new_n423_, keyIn_0_4 );
nand g223 ( new_n425_, new_n424_, new_n420_ );
xnor g224 ( new_n426_, N41, N45 );
nand g225 ( new_n427_, new_n426_, keyIn_0_5 );
not g226 ( new_n428_, keyIn_0_5 );
and g227 ( new_n429_, N41, N45 );
nor g228 ( new_n430_, N41, N45 );
nor g229 ( new_n431_, new_n429_, new_n430_ );
nand g230 ( new_n432_, new_n431_, new_n428_ );
nand g231 ( new_n433_, new_n432_, new_n427_ );
xnor g232 ( new_n434_, new_n425_, new_n433_ );
nand g233 ( new_n435_, new_n434_, new_n417_ );
and g234 ( new_n436_, new_n425_, new_n433_ );
nor g235 ( new_n437_, new_n425_, new_n433_ );
nor g236 ( new_n438_, new_n436_, new_n437_ );
nand g237 ( new_n439_, new_n438_, keyIn_0_30 );
nand g238 ( new_n440_, new_n439_, new_n435_ );
nand g239 ( new_n441_, new_n416_, new_n440_ );
not g240 ( new_n442_, keyIn_0_31 );
xnor g241 ( new_n443_, new_n415_, new_n442_ );
and g242 ( new_n444_, new_n439_, new_n435_ );
nand g243 ( new_n445_, new_n444_, new_n443_ );
nand g244 ( new_n446_, new_n445_, new_n441_ );
xnor g245 ( new_n447_, new_n446_, keyIn_0_40 );
nand g246 ( new_n448_, N134, N137 );
xor g247 ( new_n449_, new_n448_, keyIn_0_18 );
not g248 ( new_n450_, new_n449_ );
nand g249 ( new_n451_, new_n447_, new_n450_ );
not g250 ( new_n452_, keyIn_0_40 );
xnor g251 ( new_n453_, new_n446_, new_n452_ );
nand g252 ( new_n454_, new_n453_, new_n449_ );
nand g253 ( new_n455_, new_n451_, new_n454_ );
nand g254 ( new_n456_, new_n455_, keyIn_0_52 );
not g255 ( new_n457_, keyIn_0_52 );
xnor g256 ( new_n458_, new_n447_, new_n449_ );
nand g257 ( new_n459_, new_n458_, new_n457_ );
nand g258 ( new_n460_, new_n459_, new_n456_ );
xor g259 ( new_n461_, N69, N85 );
xnor g260 ( new_n462_, new_n461_, keyIn_0_24 );
xnor g261 ( new_n463_, N101, N117 );
xnor g262 ( new_n464_, new_n463_, keyIn_0_25 );
xnor g263 ( new_n465_, new_n462_, new_n464_ );
xnor g264 ( new_n466_, new_n465_, keyIn_0_37 );
not g265 ( new_n467_, new_n466_ );
nand g266 ( new_n468_, new_n460_, new_n467_ );
xnor g267 ( new_n469_, new_n455_, new_n457_ );
nand g268 ( new_n470_, new_n469_, new_n466_ );
nand g269 ( new_n471_, new_n470_, new_n468_ );
nand g270 ( new_n472_, new_n471_, new_n394_ );
xnor g271 ( new_n473_, new_n460_, new_n466_ );
nand g272 ( new_n474_, new_n473_, keyIn_0_60 );
nand g273 ( new_n475_, new_n474_, new_n472_ );
nand g274 ( new_n476_, new_n475_, new_n393_ );
nand g275 ( new_n477_, new_n416_, new_n339_ );
nand g276 ( new_n478_, new_n363_, new_n443_ );
nand g277 ( new_n479_, new_n478_, new_n477_ );
nand g278 ( new_n480_, new_n479_, keyIn_0_42 );
not g279 ( new_n481_, keyIn_0_42 );
xnor g280 ( new_n482_, new_n443_, new_n339_ );
nand g281 ( new_n483_, new_n482_, new_n481_ );
nand g282 ( new_n484_, new_n483_, new_n480_ );
nand g283 ( new_n485_, N136, N137 );
xor g284 ( new_n486_, new_n485_, keyIn_0_20 );
not g285 ( new_n487_, new_n486_ );
nand g286 ( new_n488_, new_n484_, new_n487_ );
xnor g287 ( new_n489_, new_n479_, new_n481_ );
nand g288 ( new_n490_, new_n489_, new_n486_ );
nand g289 ( new_n491_, new_n490_, new_n488_ );
nand g290 ( new_n492_, new_n491_, keyIn_0_54 );
not g291 ( new_n493_, keyIn_0_54 );
xnor g292 ( new_n494_, new_n484_, new_n486_ );
nand g293 ( new_n495_, new_n494_, new_n493_ );
nand g294 ( new_n496_, new_n495_, new_n492_ );
xor g295 ( new_n497_, N109, N125 );
xnor g296 ( new_n498_, N77, N93 );
xnor g297 ( new_n499_, new_n497_, new_n498_ );
not g298 ( new_n500_, new_n499_ );
nand g299 ( new_n501_, new_n496_, new_n500_ );
xnor g300 ( new_n502_, new_n491_, new_n493_ );
nand g301 ( new_n503_, new_n502_, new_n499_ );
nand g302 ( new_n504_, new_n503_, new_n501_ );
xnor g303 ( new_n505_, new_n504_, keyIn_0_62 );
nand g304 ( new_n506_, new_n361_, new_n440_ );
nand g305 ( new_n507_, new_n444_, new_n365_ );
nand g306 ( new_n508_, new_n507_, new_n506_ );
nand g307 ( new_n509_, new_n508_, keyIn_0_41 );
not g308 ( new_n510_, keyIn_0_41 );
xnor g309 ( new_n511_, new_n365_, new_n440_ );
nand g310 ( new_n512_, new_n511_, new_n510_ );
nand g311 ( new_n513_, new_n512_, new_n509_ );
nand g312 ( new_n514_, N135, N137 );
xor g313 ( new_n515_, new_n514_, keyIn_0_19 );
not g314 ( new_n516_, new_n515_ );
nand g315 ( new_n517_, new_n513_, new_n516_ );
xnor g316 ( new_n518_, new_n508_, new_n510_ );
nand g317 ( new_n519_, new_n518_, new_n515_ );
nand g318 ( new_n520_, new_n519_, new_n517_ );
nand g319 ( new_n521_, new_n520_, keyIn_0_53 );
not g320 ( new_n522_, keyIn_0_53 );
xnor g321 ( new_n523_, new_n513_, new_n515_ );
nand g322 ( new_n524_, new_n523_, new_n522_ );
nand g323 ( new_n525_, new_n524_, new_n521_ );
xor g324 ( new_n526_, N105, N121 );
xnor g325 ( new_n527_, new_n526_, keyIn_0_27 );
xnor g326 ( new_n528_, N73, N89 );
xnor g327 ( new_n529_, new_n528_, keyIn_0_26 );
xnor g328 ( new_n530_, new_n527_, new_n529_ );
xnor g329 ( new_n531_, new_n530_, keyIn_0_38 );
not g330 ( new_n532_, new_n531_ );
nand g331 ( new_n533_, new_n525_, new_n532_ );
xnor g332 ( new_n534_, new_n520_, new_n522_ );
nand g333 ( new_n535_, new_n534_, new_n531_ );
nand g334 ( new_n536_, new_n535_, new_n533_ );
xnor g335 ( new_n537_, new_n536_, keyIn_0_61 );
nand g336 ( new_n538_, new_n537_, new_n505_ );
nor g337 ( new_n539_, new_n476_, new_n538_ );
nand g338 ( new_n540_, new_n308_, new_n539_ );
not g339 ( new_n541_, new_n540_ );
nand g340 ( new_n542_, new_n541_, new_n225_ );
xnor g341 ( N724, new_n542_, N1 );
nand g342 ( new_n544_, new_n541_, new_n279_ );
xnor g343 ( N725, new_n544_, N5 );
nand g344 ( new_n546_, new_n541_, new_n299_ );
xnor g345 ( N726, new_n546_, N9 );
nand g346 ( new_n548_, new_n541_, new_n290_ );
xnor g347 ( N727, new_n548_, N13 );
not g348 ( new_n550_, N17 );
not g349 ( new_n551_, keyIn_0_76 );
not g350 ( new_n552_, keyIn_0_62 );
nand g351 ( new_n553_, new_n504_, new_n552_ );
xnor g352 ( new_n554_, new_n496_, new_n499_ );
nand g353 ( new_n555_, new_n554_, keyIn_0_62 );
nand g354 ( new_n556_, new_n555_, new_n553_ );
not g355 ( new_n557_, keyIn_0_61 );
nand g356 ( new_n558_, new_n536_, new_n557_ );
xnor g357 ( new_n559_, new_n525_, new_n531_ );
nand g358 ( new_n560_, new_n559_, keyIn_0_61 );
nand g359 ( new_n561_, new_n560_, new_n558_ );
nand g360 ( new_n562_, new_n561_, new_n556_ );
nor g361 ( new_n563_, new_n476_, new_n562_ );
nand g362 ( new_n564_, new_n308_, new_n563_ );
xnor g363 ( new_n565_, new_n564_, new_n551_ );
nand g364 ( new_n566_, new_n565_, new_n225_ );
xor g365 ( new_n567_, new_n566_, keyIn_0_82 );
xnor g366 ( new_n568_, new_n567_, new_n550_ );
nand g367 ( new_n569_, new_n568_, keyIn_0_105 );
not g368 ( new_n570_, keyIn_0_105 );
xnor g369 ( new_n571_, new_n567_, N17 );
nand g370 ( new_n572_, new_n571_, new_n570_ );
nand g371 ( N728, new_n569_, new_n572_ );
not g372 ( new_n574_, N21 );
nand g373 ( new_n575_, new_n565_, new_n279_ );
xnor g374 ( new_n576_, new_n575_, keyIn_0_83 );
xnor g375 ( new_n577_, new_n576_, new_n574_ );
xnor g376 ( N729, new_n577_, keyIn_0_106 );
nand g377 ( new_n579_, new_n565_, new_n299_ );
xnor g378 ( N730, new_n579_, N25 );
nand g379 ( new_n581_, new_n565_, new_n290_ );
xnor g380 ( new_n582_, new_n581_, keyIn_0_84 );
xnor g381 ( new_n583_, new_n582_, N29 );
xnor g382 ( N731, new_n583_, keyIn_0_107 );
not g383 ( new_n585_, keyIn_0_85 );
not g384 ( new_n586_, keyIn_0_77 );
nor g385 ( new_n587_, new_n393_, new_n556_ );
nand g386 ( new_n588_, new_n587_, new_n537_ );
not g387 ( new_n589_, new_n475_ );
nand g388 ( new_n590_, new_n308_, new_n589_ );
nor g389 ( new_n591_, new_n590_, new_n588_ );
xnor g390 ( new_n592_, new_n591_, new_n586_ );
nor g391 ( new_n593_, new_n592_, new_n294_ );
nand g392 ( new_n594_, new_n593_, new_n585_ );
xnor g393 ( new_n595_, new_n591_, keyIn_0_77 );
nand g394 ( new_n596_, new_n595_, new_n225_ );
nand g395 ( new_n597_, new_n596_, keyIn_0_85 );
nand g396 ( new_n598_, new_n594_, new_n597_ );
nand g397 ( new_n599_, new_n598_, N33 );
not g398 ( new_n600_, N33 );
xnor g399 ( new_n601_, new_n596_, new_n585_ );
nand g400 ( new_n602_, new_n601_, new_n600_ );
nand g401 ( new_n603_, new_n602_, new_n599_ );
nand g402 ( new_n604_, new_n603_, keyIn_0_108 );
not g403 ( new_n605_, keyIn_0_108 );
xnor g404 ( new_n606_, new_n598_, new_n600_ );
nand g405 ( new_n607_, new_n606_, new_n605_ );
nand g406 ( N732, new_n607_, new_n604_ );
not g407 ( new_n609_, keyIn_0_109 );
nor g408 ( new_n610_, new_n592_, new_n303_ );
nand g409 ( new_n611_, new_n610_, keyIn_0_86 );
not g410 ( new_n612_, keyIn_0_86 );
nand g411 ( new_n613_, new_n595_, new_n279_ );
nand g412 ( new_n614_, new_n613_, new_n612_ );
nand g413 ( new_n615_, new_n611_, new_n614_ );
nand g414 ( new_n616_, new_n615_, N37 );
not g415 ( new_n617_, N37 );
xnor g416 ( new_n618_, new_n613_, keyIn_0_86 );
nand g417 ( new_n619_, new_n618_, new_n617_ );
nand g418 ( new_n620_, new_n619_, new_n616_ );
nand g419 ( new_n621_, new_n620_, new_n609_ );
xnor g420 ( new_n622_, new_n615_, new_n617_ );
nand g421 ( new_n623_, new_n622_, keyIn_0_109 );
nand g422 ( N733, new_n623_, new_n621_ );
not g423 ( new_n625_, N41 );
nor g424 ( new_n626_, new_n592_, new_n255_ );
nand g425 ( new_n627_, new_n626_, keyIn_0_87 );
not g426 ( new_n628_, keyIn_0_87 );
nand g427 ( new_n629_, new_n595_, new_n299_ );
nand g428 ( new_n630_, new_n629_, new_n628_ );
nand g429 ( new_n631_, new_n627_, new_n630_ );
nand g430 ( new_n632_, new_n631_, new_n625_ );
xnor g431 ( new_n633_, new_n629_, keyIn_0_87 );
nand g432 ( new_n634_, new_n633_, N41 );
nand g433 ( new_n635_, new_n634_, new_n632_ );
nand g434 ( new_n636_, new_n635_, keyIn_0_110 );
not g435 ( new_n637_, keyIn_0_110 );
xnor g436 ( new_n638_, new_n631_, N41 );
nand g437 ( new_n639_, new_n638_, new_n637_ );
nand g438 ( N734, new_n639_, new_n636_ );
not g439 ( new_n641_, N45 );
not g440 ( new_n642_, new_n290_ );
nor g441 ( new_n643_, new_n592_, new_n642_ );
nand g442 ( new_n644_, new_n643_, keyIn_0_88 );
not g443 ( new_n645_, keyIn_0_88 );
nand g444 ( new_n646_, new_n595_, new_n290_ );
nand g445 ( new_n647_, new_n646_, new_n645_ );
nand g446 ( new_n648_, new_n644_, new_n647_ );
nand g447 ( new_n649_, new_n648_, new_n641_ );
xnor g448 ( new_n650_, new_n646_, keyIn_0_88 );
nand g449 ( new_n651_, new_n650_, N45 );
nand g450 ( new_n652_, new_n651_, new_n649_ );
nand g451 ( new_n653_, new_n652_, keyIn_0_111 );
not g452 ( new_n654_, keyIn_0_111 );
xnor g453 ( new_n655_, new_n648_, N45 );
nand g454 ( new_n656_, new_n655_, new_n654_ );
nand g455 ( N735, new_n656_, new_n653_ );
nor g456 ( new_n658_, new_n393_, new_n505_ );
nand g457 ( new_n659_, new_n658_, new_n561_ );
nor g458 ( new_n660_, new_n590_, new_n659_ );
nand g459 ( new_n661_, new_n660_, new_n225_ );
xnor g460 ( N736, new_n661_, N49 );
nand g461 ( new_n663_, new_n660_, new_n279_ );
xnor g462 ( N737, new_n663_, N53 );
nand g463 ( new_n665_, new_n660_, new_n299_ );
xnor g464 ( N738, new_n665_, N57 );
nand g465 ( new_n667_, new_n660_, new_n290_ );
xnor g466 ( N739, new_n667_, N61 );
not g467 ( new_n669_, N65 );
not g468 ( new_n670_, keyIn_0_71 );
nand g469 ( new_n671_, new_n658_, new_n475_ );
not g470 ( new_n672_, keyIn_0_64 );
nand g471 ( new_n673_, new_n561_, new_n672_ );
nand g472 ( new_n674_, new_n537_, keyIn_0_64 );
nand g473 ( new_n675_, new_n674_, new_n673_ );
nor g474 ( new_n676_, new_n671_, new_n675_ );
nand g475 ( new_n677_, new_n676_, new_n670_ );
nand g476 ( new_n678_, new_n392_, keyIn_0_59 );
xnor g477 ( new_n679_, new_n384_, new_n387_ );
nand g478 ( new_n680_, new_n679_, new_n309_ );
nand g479 ( new_n681_, new_n680_, new_n678_ );
nand g480 ( new_n682_, new_n681_, new_n556_ );
nor g481 ( new_n683_, new_n682_, new_n589_ );
xnor g482 ( new_n684_, new_n561_, keyIn_0_64 );
nand g483 ( new_n685_, new_n684_, new_n683_ );
nand g484 ( new_n686_, new_n685_, keyIn_0_71 );
nand g485 ( new_n687_, new_n677_, new_n686_ );
not g486 ( new_n688_, keyIn_0_72 );
nor g487 ( new_n689_, new_n588_, new_n589_ );
nand g488 ( new_n690_, new_n689_, new_n688_ );
nand g489 ( new_n691_, new_n505_, new_n681_ );
nor g490 ( new_n692_, new_n691_, new_n561_ );
nand g491 ( new_n693_, new_n692_, new_n475_ );
nand g492 ( new_n694_, new_n693_, keyIn_0_72 );
nand g493 ( new_n695_, new_n690_, new_n694_ );
nand g494 ( new_n696_, new_n687_, new_n695_ );
nand g495 ( new_n697_, new_n561_, keyIn_0_66 );
not g496 ( new_n698_, keyIn_0_66 );
nand g497 ( new_n699_, new_n537_, new_n698_ );
nand g498 ( new_n700_, new_n699_, new_n697_ );
nor g499 ( new_n701_, new_n476_, new_n556_ );
nand g500 ( new_n702_, new_n701_, new_n700_ );
xnor g501 ( new_n703_, new_n702_, keyIn_0_74 );
not g502 ( new_n704_, keyIn_0_73 );
nand g503 ( new_n705_, new_n561_, keyIn_0_65 );
not g504 ( new_n706_, keyIn_0_65 );
nand g505 ( new_n707_, new_n537_, new_n706_ );
nand g506 ( new_n708_, new_n707_, new_n705_ );
nor g507 ( new_n709_, new_n691_, new_n475_ );
nand g508 ( new_n710_, new_n709_, new_n708_ );
xnor g509 ( new_n711_, new_n710_, new_n704_ );
nand g510 ( new_n712_, new_n703_, new_n711_ );
nor g511 ( new_n713_, new_n712_, new_n696_ );
nand g512 ( new_n714_, new_n713_, keyIn_0_75 );
not g513 ( new_n715_, keyIn_0_75 );
and g514 ( new_n716_, new_n687_, new_n695_ );
not g515 ( new_n717_, keyIn_0_74 );
xnor g516 ( new_n718_, new_n702_, new_n717_ );
xnor g517 ( new_n719_, new_n710_, keyIn_0_73 );
nor g518 ( new_n720_, new_n718_, new_n719_ );
nand g519 ( new_n721_, new_n720_, new_n716_ );
nand g520 ( new_n722_, new_n721_, new_n715_ );
nand g521 ( new_n723_, new_n722_, new_n714_ );
nor g522 ( new_n724_, new_n279_, keyIn_0_67 );
nand g523 ( new_n725_, new_n279_, keyIn_0_67 );
nor g524 ( new_n726_, new_n294_, new_n290_ );
nand g525 ( new_n727_, new_n726_, new_n725_ );
nor g526 ( new_n728_, new_n727_, new_n724_ );
and g527 ( new_n729_, new_n728_, new_n299_ );
nand g528 ( new_n730_, new_n723_, new_n729_ );
nor g529 ( new_n731_, new_n730_, keyIn_0_78 );
nand g530 ( new_n732_, new_n730_, keyIn_0_78 );
nand g531 ( new_n733_, new_n732_, new_n393_ );
nor g532 ( new_n734_, new_n733_, new_n731_ );
nand g533 ( new_n735_, new_n734_, keyIn_0_89 );
not g534 ( new_n736_, keyIn_0_89 );
not g535 ( new_n737_, new_n731_ );
and g536 ( new_n738_, new_n732_, new_n393_ );
nand g537 ( new_n739_, new_n738_, new_n737_ );
nand g538 ( new_n740_, new_n739_, new_n736_ );
nand g539 ( new_n741_, new_n740_, new_n735_ );
nand g540 ( new_n742_, new_n741_, new_n669_ );
xnor g541 ( new_n743_, new_n734_, new_n736_ );
nand g542 ( new_n744_, new_n743_, N65 );
nand g543 ( new_n745_, new_n744_, new_n742_ );
nand g544 ( new_n746_, new_n745_, keyIn_0_112 );
not g545 ( new_n747_, keyIn_0_112 );
xnor g546 ( new_n748_, new_n741_, N65 );
nand g547 ( new_n749_, new_n748_, new_n747_ );
nand g548 ( N740, new_n749_, new_n746_ );
not g549 ( new_n751_, keyIn_0_113 );
nand g550 ( new_n752_, new_n732_, new_n589_ );
nor g551 ( new_n753_, new_n752_, new_n731_ );
nand g552 ( new_n754_, new_n753_, keyIn_0_90 );
not g553 ( new_n755_, keyIn_0_90 );
and g554 ( new_n756_, new_n732_, new_n589_ );
nand g555 ( new_n757_, new_n756_, new_n737_ );
nand g556 ( new_n758_, new_n757_, new_n755_ );
nand g557 ( new_n759_, new_n758_, new_n754_ );
nand g558 ( new_n760_, new_n759_, N69 );
not g559 ( new_n761_, N69 );
xnor g560 ( new_n762_, new_n753_, new_n755_ );
nand g561 ( new_n763_, new_n762_, new_n761_ );
nand g562 ( new_n764_, new_n763_, new_n760_ );
nand g563 ( new_n765_, new_n764_, new_n751_ );
xnor g564 ( new_n766_, new_n759_, new_n761_ );
nand g565 ( new_n767_, new_n766_, keyIn_0_113 );
nand g566 ( N741, new_n767_, new_n765_ );
not g567 ( new_n769_, keyIn_0_114 );
nand g568 ( new_n770_, new_n732_, new_n537_ );
nor g569 ( new_n771_, new_n770_, new_n731_ );
nand g570 ( new_n772_, new_n771_, keyIn_0_91 );
not g571 ( new_n773_, keyIn_0_91 );
and g572 ( new_n774_, new_n732_, new_n537_ );
nand g573 ( new_n775_, new_n774_, new_n737_ );
nand g574 ( new_n776_, new_n775_, new_n773_ );
nand g575 ( new_n777_, new_n776_, new_n772_ );
nand g576 ( new_n778_, new_n777_, N73 );
not g577 ( new_n779_, N73 );
xnor g578 ( new_n780_, new_n771_, new_n773_ );
nand g579 ( new_n781_, new_n780_, new_n779_ );
nand g580 ( new_n782_, new_n781_, new_n778_ );
nand g581 ( new_n783_, new_n782_, new_n769_ );
xnor g582 ( new_n784_, new_n777_, new_n779_ );
nand g583 ( new_n785_, new_n784_, keyIn_0_114 );
nand g584 ( N742, new_n785_, new_n783_ );
nand g585 ( new_n787_, new_n732_, new_n556_ );
nor g586 ( new_n788_, new_n787_, new_n731_ );
nand g587 ( new_n789_, new_n788_, keyIn_0_92 );
not g588 ( new_n790_, keyIn_0_92 );
and g589 ( new_n791_, new_n732_, new_n556_ );
nand g590 ( new_n792_, new_n791_, new_n737_ );
nand g591 ( new_n793_, new_n792_, new_n790_ );
nand g592 ( new_n794_, new_n793_, new_n789_ );
nand g593 ( new_n795_, new_n794_, N77 );
not g594 ( new_n796_, N77 );
xnor g595 ( new_n797_, new_n788_, new_n790_ );
nand g596 ( new_n798_, new_n797_, new_n796_ );
nand g597 ( new_n799_, new_n798_, new_n795_ );
nand g598 ( new_n800_, new_n799_, keyIn_0_115 );
not g599 ( new_n801_, keyIn_0_115 );
xnor g600 ( new_n802_, new_n794_, new_n796_ );
nand g601 ( new_n803_, new_n802_, new_n801_ );
nand g602 ( N743, new_n803_, new_n800_ );
not g603 ( new_n805_, keyIn_0_116 );
not g604 ( new_n806_, keyIn_0_79 );
not g605 ( new_n807_, keyIn_0_68 );
nor g606 ( new_n808_, new_n299_, new_n807_ );
nand g607 ( new_n809_, new_n299_, new_n807_ );
nor g608 ( new_n810_, new_n304_, new_n642_ );
nand g609 ( new_n811_, new_n809_, new_n810_ );
nor g610 ( new_n812_, new_n811_, new_n808_ );
nand g611 ( new_n813_, new_n723_, new_n812_ );
nor g612 ( new_n814_, new_n813_, new_n806_ );
nand g613 ( new_n815_, new_n813_, new_n806_ );
nand g614 ( new_n816_, new_n815_, new_n393_ );
nor g615 ( new_n817_, new_n816_, new_n814_ );
nand g616 ( new_n818_, new_n817_, keyIn_0_93 );
not g617 ( new_n819_, keyIn_0_93 );
not g618 ( new_n820_, new_n814_ );
and g619 ( new_n821_, new_n815_, new_n393_ );
nand g620 ( new_n822_, new_n821_, new_n820_ );
nand g621 ( new_n823_, new_n822_, new_n819_ );
nand g622 ( new_n824_, new_n823_, new_n818_ );
nand g623 ( new_n825_, new_n824_, N81 );
not g624 ( new_n826_, N81 );
xnor g625 ( new_n827_, new_n817_, new_n819_ );
nand g626 ( new_n828_, new_n827_, new_n826_ );
nand g627 ( new_n829_, new_n828_, new_n825_ );
nand g628 ( new_n830_, new_n829_, new_n805_ );
xnor g629 ( new_n831_, new_n824_, new_n826_ );
nand g630 ( new_n832_, new_n831_, keyIn_0_116 );
nand g631 ( N744, new_n832_, new_n830_ );
nand g632 ( new_n834_, new_n815_, new_n589_ );
nor g633 ( new_n835_, new_n834_, new_n814_ );
nand g634 ( new_n836_, new_n835_, keyIn_0_94 );
not g635 ( new_n837_, keyIn_0_94 );
and g636 ( new_n838_, new_n815_, new_n589_ );
nand g637 ( new_n839_, new_n838_, new_n820_ );
nand g638 ( new_n840_, new_n839_, new_n837_ );
nand g639 ( new_n841_, new_n840_, new_n836_ );
nand g640 ( new_n842_, new_n841_, N85 );
not g641 ( new_n843_, N85 );
xnor g642 ( new_n844_, new_n835_, new_n837_ );
nand g643 ( new_n845_, new_n844_, new_n843_ );
nand g644 ( new_n846_, new_n845_, new_n842_ );
nand g645 ( new_n847_, new_n846_, keyIn_0_117 );
not g646 ( new_n848_, keyIn_0_117 );
xnor g647 ( new_n849_, new_n841_, new_n843_ );
nand g648 ( new_n850_, new_n849_, new_n848_ );
nand g649 ( N745, new_n850_, new_n847_ );
not g650 ( new_n852_, keyIn_0_118 );
nand g651 ( new_n853_, new_n815_, new_n537_ );
nor g652 ( new_n854_, new_n853_, new_n814_ );
nand g653 ( new_n855_, new_n854_, keyIn_0_95 );
not g654 ( new_n856_, keyIn_0_95 );
and g655 ( new_n857_, new_n815_, new_n537_ );
nand g656 ( new_n858_, new_n857_, new_n820_ );
nand g657 ( new_n859_, new_n858_, new_n856_ );
nand g658 ( new_n860_, new_n859_, new_n855_ );
nand g659 ( new_n861_, new_n860_, N89 );
not g660 ( new_n862_, N89 );
xnor g661 ( new_n863_, new_n854_, new_n856_ );
nand g662 ( new_n864_, new_n863_, new_n862_ );
nand g663 ( new_n865_, new_n864_, new_n861_ );
nand g664 ( new_n866_, new_n865_, new_n852_ );
xnor g665 ( new_n867_, new_n860_, new_n862_ );
nand g666 ( new_n868_, new_n867_, keyIn_0_118 );
nand g667 ( N746, new_n868_, new_n866_ );
not g668 ( new_n870_, keyIn_0_119 );
nand g669 ( new_n871_, new_n815_, new_n556_ );
nor g670 ( new_n872_, new_n871_, new_n814_ );
nand g671 ( new_n873_, new_n872_, keyIn_0_96 );
not g672 ( new_n874_, keyIn_0_96 );
and g673 ( new_n875_, new_n815_, new_n556_ );
nand g674 ( new_n876_, new_n875_, new_n820_ );
nand g675 ( new_n877_, new_n876_, new_n874_ );
nand g676 ( new_n878_, new_n877_, new_n873_ );
nand g677 ( new_n879_, new_n878_, N93 );
not g678 ( new_n880_, N93 );
xnor g679 ( new_n881_, new_n872_, new_n874_ );
nand g680 ( new_n882_, new_n881_, new_n880_ );
nand g681 ( new_n883_, new_n882_, new_n879_ );
nand g682 ( new_n884_, new_n883_, new_n870_ );
xnor g683 ( new_n885_, new_n878_, new_n880_ );
nand g684 ( new_n886_, new_n885_, keyIn_0_119 );
nand g685 ( N747, new_n886_, new_n884_ );
not g686 ( new_n888_, keyIn_0_120 );
not g687 ( new_n889_, keyIn_0_97 );
nand g688 ( new_n890_, new_n294_, new_n279_ );
nor g689 ( new_n891_, new_n890_, new_n290_ );
nand g690 ( new_n892_, new_n891_, new_n299_ );
not g691 ( new_n893_, new_n892_ );
nand g692 ( new_n894_, new_n723_, new_n893_ );
nor g693 ( new_n895_, new_n894_, keyIn_0_80 );
nand g694 ( new_n896_, new_n894_, keyIn_0_80 );
nand g695 ( new_n897_, new_n896_, new_n393_ );
nor g696 ( new_n898_, new_n897_, new_n895_ );
nand g697 ( new_n899_, new_n898_, new_n889_ );
not g698 ( new_n900_, new_n895_ );
and g699 ( new_n901_, new_n896_, new_n393_ );
nand g700 ( new_n902_, new_n901_, new_n900_ );
nand g701 ( new_n903_, new_n902_, keyIn_0_97 );
nand g702 ( new_n904_, new_n903_, new_n899_ );
nand g703 ( new_n905_, new_n904_, N97 );
not g704 ( new_n906_, N97 );
xnor g705 ( new_n907_, new_n898_, keyIn_0_97 );
nand g706 ( new_n908_, new_n907_, new_n906_ );
nand g707 ( new_n909_, new_n908_, new_n905_ );
nand g708 ( new_n910_, new_n909_, new_n888_ );
xnor g709 ( new_n911_, new_n904_, new_n906_ );
nand g710 ( new_n912_, new_n911_, keyIn_0_120 );
nand g711 ( N748, new_n912_, new_n910_ );
nand g712 ( new_n914_, new_n896_, new_n589_ );
nor g713 ( new_n915_, new_n914_, new_n895_ );
nand g714 ( new_n916_, new_n915_, keyIn_0_98 );
not g715 ( new_n917_, keyIn_0_98 );
and g716 ( new_n918_, new_n896_, new_n589_ );
nand g717 ( new_n919_, new_n918_, new_n900_ );
nand g718 ( new_n920_, new_n919_, new_n917_ );
nand g719 ( new_n921_, new_n920_, new_n916_ );
nand g720 ( new_n922_, new_n921_, N101 );
not g721 ( new_n923_, N101 );
xnor g722 ( new_n924_, new_n915_, new_n917_ );
nand g723 ( new_n925_, new_n924_, new_n923_ );
nand g724 ( new_n926_, new_n925_, new_n922_ );
nand g725 ( new_n927_, new_n926_, keyIn_0_121 );
not g726 ( new_n928_, keyIn_0_121 );
xnor g727 ( new_n929_, new_n921_, new_n923_ );
nand g728 ( new_n930_, new_n929_, new_n928_ );
nand g729 ( N749, new_n930_, new_n927_ );
not g730 ( new_n932_, keyIn_0_99 );
nand g731 ( new_n933_, new_n896_, new_n537_ );
nor g732 ( new_n934_, new_n933_, new_n895_ );
nand g733 ( new_n935_, new_n934_, new_n932_ );
and g734 ( new_n936_, new_n896_, new_n537_ );
nand g735 ( new_n937_, new_n936_, new_n900_ );
nand g736 ( new_n938_, new_n937_, keyIn_0_99 );
nand g737 ( new_n939_, new_n938_, new_n935_ );
nand g738 ( new_n940_, new_n939_, N105 );
not g739 ( new_n941_, N105 );
xnor g740 ( new_n942_, new_n934_, keyIn_0_99 );
nand g741 ( new_n943_, new_n942_, new_n941_ );
nand g742 ( new_n944_, new_n943_, new_n940_ );
nand g743 ( new_n945_, new_n944_, keyIn_0_122 );
not g744 ( new_n946_, keyIn_0_122 );
xnor g745 ( new_n947_, new_n939_, new_n941_ );
nand g746 ( new_n948_, new_n947_, new_n946_ );
nand g747 ( N750, new_n948_, new_n945_ );
not g748 ( new_n950_, keyIn_0_123 );
not g749 ( new_n951_, keyIn_0_100 );
nand g750 ( new_n952_, new_n896_, new_n556_ );
nor g751 ( new_n953_, new_n952_, new_n895_ );
nand g752 ( new_n954_, new_n953_, new_n951_ );
and g753 ( new_n955_, new_n896_, new_n556_ );
nand g754 ( new_n956_, new_n955_, new_n900_ );
nand g755 ( new_n957_, new_n956_, keyIn_0_100 );
nand g756 ( new_n958_, new_n957_, new_n954_ );
nand g757 ( new_n959_, new_n958_, N109 );
not g758 ( new_n960_, N109 );
xnor g759 ( new_n961_, new_n953_, keyIn_0_100 );
nand g760 ( new_n962_, new_n961_, new_n960_ );
nand g761 ( new_n963_, new_n962_, new_n959_ );
nand g762 ( new_n964_, new_n963_, new_n950_ );
xnor g763 ( new_n965_, new_n958_, new_n960_ );
nand g764 ( new_n966_, new_n965_, keyIn_0_123 );
nand g765 ( N751, new_n966_, new_n964_ );
not g766 ( new_n968_, keyIn_0_70 );
nand g767 ( new_n969_, new_n299_, new_n968_ );
nor g768 ( new_n970_, new_n299_, new_n968_ );
not g769 ( new_n971_, keyIn_0_69 );
nand g770 ( new_n972_, new_n294_, new_n971_ );
nor g771 ( new_n973_, new_n294_, new_n971_ );
nor g772 ( new_n974_, new_n973_, new_n295_ );
nand g773 ( new_n975_, new_n974_, new_n972_ );
nor g774 ( new_n976_, new_n975_, new_n970_ );
and g775 ( new_n977_, new_n976_, new_n969_ );
nand g776 ( new_n978_, new_n723_, new_n977_ );
nor g777 ( new_n979_, new_n978_, keyIn_0_81 );
nand g778 ( new_n980_, new_n978_, keyIn_0_81 );
nand g779 ( new_n981_, new_n980_, new_n393_ );
nor g780 ( new_n982_, new_n981_, new_n979_ );
nand g781 ( new_n983_, new_n982_, keyIn_0_101 );
not g782 ( new_n984_, keyIn_0_101 );
not g783 ( new_n985_, new_n979_ );
and g784 ( new_n986_, new_n980_, new_n393_ );
nand g785 ( new_n987_, new_n986_, new_n985_ );
nand g786 ( new_n988_, new_n987_, new_n984_ );
nand g787 ( new_n989_, new_n988_, new_n983_ );
nand g788 ( new_n990_, new_n989_, N113 );
not g789 ( new_n991_, N113 );
xnor g790 ( new_n992_, new_n982_, new_n984_ );
nand g791 ( new_n993_, new_n992_, new_n991_ );
nand g792 ( new_n994_, new_n993_, new_n990_ );
nand g793 ( new_n995_, new_n994_, keyIn_0_124 );
not g794 ( new_n996_, keyIn_0_124 );
xnor g795 ( new_n997_, new_n989_, new_n991_ );
nand g796 ( new_n998_, new_n997_, new_n996_ );
nand g797 ( N752, new_n998_, new_n995_ );
not g798 ( new_n1000_, keyIn_0_125 );
nand g799 ( new_n1001_, new_n980_, new_n589_ );
nor g800 ( new_n1002_, new_n1001_, new_n979_ );
nand g801 ( new_n1003_, new_n1002_, keyIn_0_102 );
not g802 ( new_n1004_, keyIn_0_102 );
and g803 ( new_n1005_, new_n980_, new_n589_ );
nand g804 ( new_n1006_, new_n1005_, new_n985_ );
nand g805 ( new_n1007_, new_n1006_, new_n1004_ );
nand g806 ( new_n1008_, new_n1007_, new_n1003_ );
nand g807 ( new_n1009_, new_n1008_, N117 );
not g808 ( new_n1010_, N117 );
xnor g809 ( new_n1011_, new_n1002_, new_n1004_ );
nand g810 ( new_n1012_, new_n1011_, new_n1010_ );
nand g811 ( new_n1013_, new_n1012_, new_n1009_ );
nand g812 ( new_n1014_, new_n1013_, new_n1000_ );
xnor g813 ( new_n1015_, new_n1008_, new_n1010_ );
nand g814 ( new_n1016_, new_n1015_, keyIn_0_125 );
nand g815 ( N753, new_n1016_, new_n1014_ );
not g816 ( new_n1018_, N121 );
nand g817 ( new_n1019_, new_n980_, new_n537_ );
nor g818 ( new_n1020_, new_n1019_, new_n979_ );
nand g819 ( new_n1021_, new_n1020_, keyIn_0_103 );
not g820 ( new_n1022_, keyIn_0_103 );
and g821 ( new_n1023_, new_n980_, new_n537_ );
nand g822 ( new_n1024_, new_n1023_, new_n985_ );
nand g823 ( new_n1025_, new_n1024_, new_n1022_ );
nand g824 ( new_n1026_, new_n1025_, new_n1021_ );
nand g825 ( new_n1027_, new_n1026_, new_n1018_ );
xnor g826 ( new_n1028_, new_n1020_, new_n1022_ );
nand g827 ( new_n1029_, new_n1028_, N121 );
nand g828 ( new_n1030_, new_n1029_, new_n1027_ );
nand g829 ( new_n1031_, new_n1030_, keyIn_0_126 );
not g830 ( new_n1032_, keyIn_0_126 );
xnor g831 ( new_n1033_, new_n1026_, N121 );
nand g832 ( new_n1034_, new_n1033_, new_n1032_ );
nand g833 ( N754, new_n1034_, new_n1031_ );
not g834 ( new_n1036_, keyIn_0_127 );
nand g835 ( new_n1037_, new_n980_, new_n556_ );
nor g836 ( new_n1038_, new_n1037_, new_n979_ );
nand g837 ( new_n1039_, new_n1038_, keyIn_0_104 );
not g838 ( new_n1040_, keyIn_0_104 );
and g839 ( new_n1041_, new_n980_, new_n556_ );
nand g840 ( new_n1042_, new_n1041_, new_n985_ );
nand g841 ( new_n1043_, new_n1042_, new_n1040_ );
nand g842 ( new_n1044_, new_n1043_, new_n1039_ );
nand g843 ( new_n1045_, new_n1044_, N125 );
not g844 ( new_n1046_, N125 );
xnor g845 ( new_n1047_, new_n1038_, new_n1040_ );
nand g846 ( new_n1048_, new_n1047_, new_n1046_ );
nand g847 ( new_n1049_, new_n1048_, new_n1045_ );
nand g848 ( new_n1050_, new_n1049_, new_n1036_ );
xnor g849 ( new_n1051_, new_n1044_, new_n1046_ );
nand g850 ( new_n1052_, new_n1051_, keyIn_0_127 );
nand g851 ( N755, new_n1052_, new_n1050_ );
endmodule