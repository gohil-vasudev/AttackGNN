module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n256_, new_n452_, new_n381_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n126_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n813_, new_n830_, new_n480_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n837_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n765_, new_n405_;

not g000 ( new_n106_, N65 );
or g001 ( new_n107_, new_n106_, N69 );
not g002 ( new_n108_, N69 );
or g003 ( new_n109_, new_n108_, N65 );
and g004 ( new_n110_, new_n107_, new_n109_ );
and g005 ( new_n111_, N73, N77 );
not g006 ( new_n112_, new_n111_ );
or g007 ( new_n113_, N73, N77 );
and g008 ( new_n114_, new_n112_, new_n113_ );
or g009 ( new_n115_, new_n110_, new_n114_ );
and g010 ( new_n116_, new_n110_, new_n114_ );
not g011 ( new_n117_, new_n116_ );
and g012 ( new_n118_, new_n117_, new_n115_ );
not g013 ( new_n119_, new_n118_ );
not g014 ( new_n120_, N81 );
or g015 ( new_n121_, new_n120_, N85 );
not g016 ( new_n122_, N85 );
or g017 ( new_n123_, new_n122_, N81 );
and g018 ( new_n124_, new_n121_, new_n123_ );
and g019 ( new_n125_, N89, N93 );
not g020 ( new_n126_, new_n125_ );
or g021 ( new_n127_, N89, N93 );
and g022 ( new_n128_, new_n126_, new_n127_ );
or g023 ( new_n129_, new_n124_, new_n128_ );
and g024 ( new_n130_, new_n124_, new_n128_ );
not g025 ( new_n131_, new_n130_ );
and g026 ( new_n132_, new_n131_, new_n129_ );
not g027 ( new_n133_, new_n132_ );
and g028 ( new_n134_, new_n119_, new_n133_ );
and g029 ( new_n135_, new_n118_, new_n132_ );
or g030 ( new_n136_, new_n134_, new_n135_ );
and g031 ( new_n137_, N129, N137 );
and g032 ( new_n138_, new_n136_, new_n137_ );
not g033 ( new_n139_, new_n134_ );
not g034 ( new_n140_, new_n135_ );
not g035 ( new_n141_, new_n137_ );
and g036 ( new_n142_, new_n139_, new_n140_, new_n141_ );
or g037 ( new_n143_, new_n138_, new_n142_ );
not g038 ( new_n144_, keyIn_0_9 );
not g039 ( new_n145_, N17 );
and g040 ( new_n146_, new_n145_, N1 );
not g041 ( new_n147_, N1 );
and g042 ( new_n148_, new_n147_, N17 );
or g043 ( new_n149_, new_n146_, new_n148_ );
and g044 ( new_n150_, N33, N49 );
not g045 ( new_n151_, N33 );
not g046 ( new_n152_, N49 );
and g047 ( new_n153_, new_n151_, new_n152_ );
or g048 ( new_n154_, new_n153_, new_n150_ );
and g049 ( new_n155_, new_n149_, new_n154_ );
not g050 ( new_n156_, new_n149_ );
not g051 ( new_n157_, new_n154_ );
and g052 ( new_n158_, new_n156_, new_n157_ );
or g053 ( new_n159_, new_n158_, new_n155_ );
and g054 ( new_n160_, new_n159_, new_n144_ );
not g055 ( new_n161_, new_n160_ );
or g056 ( new_n162_, new_n159_, new_n144_ );
and g057 ( new_n163_, new_n161_, new_n162_ );
not g058 ( new_n164_, new_n163_ );
and g059 ( new_n165_, new_n143_, new_n164_ );
not g060 ( new_n166_, new_n138_ );
not g061 ( new_n167_, new_n142_ );
and g062 ( new_n168_, new_n166_, new_n167_, new_n163_ );
or g063 ( new_n169_, new_n165_, new_n168_ );
not g064 ( new_n170_, keyIn_0_24 );
not g065 ( new_n171_, keyIn_0_5 );
and g066 ( new_n172_, N1, N5 );
not g067 ( new_n173_, N5 );
and g068 ( new_n174_, new_n147_, new_n173_ );
or g069 ( new_n175_, new_n174_, new_n172_ );
and g070 ( new_n176_, N9, N13 );
not g071 ( new_n177_, N9 );
not g072 ( new_n178_, N13 );
and g073 ( new_n179_, new_n177_, new_n178_ );
or g074 ( new_n180_, new_n179_, new_n176_ );
and g075 ( new_n181_, new_n175_, new_n180_ );
not g076 ( new_n182_, new_n175_ );
not g077 ( new_n183_, new_n180_ );
and g078 ( new_n184_, new_n182_, new_n183_ );
or g079 ( new_n185_, new_n184_, new_n181_ );
not g080 ( new_n186_, new_n185_ );
not g081 ( new_n187_, keyIn_0_8 );
or g082 ( new_n188_, N41, N45 );
and g083 ( new_n189_, N41, N45 );
not g084 ( new_n190_, new_n189_ );
and g085 ( new_n191_, new_n190_, new_n188_ );
or g086 ( new_n192_, new_n191_, keyIn_0_2 );
and g087 ( new_n193_, new_n190_, keyIn_0_2, new_n188_ );
not g088 ( new_n194_, new_n193_ );
and g089 ( new_n195_, new_n192_, new_n194_ );
not g090 ( new_n196_, keyIn_0_1 );
and g091 ( new_n197_, N33, N37 );
not g092 ( new_n198_, new_n197_ );
or g093 ( new_n199_, N33, N37 );
and g094 ( new_n200_, new_n198_, new_n199_ );
or g095 ( new_n201_, new_n200_, new_n196_ );
and g096 ( new_n202_, new_n198_, new_n196_, new_n199_ );
not g097 ( new_n203_, new_n202_ );
and g098 ( new_n204_, new_n201_, new_n203_ );
or g099 ( new_n205_, new_n195_, new_n204_ );
and g100 ( new_n206_, new_n192_, new_n201_, new_n194_, new_n203_ );
not g101 ( new_n207_, new_n206_ );
and g102 ( new_n208_, new_n205_, new_n207_ );
or g103 ( new_n209_, new_n208_, new_n187_ );
and g104 ( new_n210_, new_n205_, new_n187_, new_n207_ );
not g105 ( new_n211_, new_n210_ );
and g106 ( new_n212_, new_n209_, new_n211_ );
or g107 ( new_n213_, new_n212_, new_n186_ );
and g108 ( new_n214_, new_n209_, new_n186_, new_n211_ );
not g109 ( new_n215_, new_n214_ );
and g110 ( new_n216_, new_n213_, new_n215_ );
or g111 ( new_n217_, new_n216_, new_n171_ );
and g112 ( new_n218_, new_n213_, new_n171_, new_n215_ );
not g113 ( new_n219_, new_n218_ );
and g114 ( new_n220_, new_n217_, new_n219_ );
and g115 ( new_n221_, N135, N137 );
or g116 ( new_n222_, new_n220_, new_n221_ );
and g117 ( new_n223_, new_n217_, new_n219_, new_n221_ );
not g118 ( new_n224_, new_n223_ );
and g119 ( new_n225_, new_n222_, new_n224_ );
and g120 ( new_n226_, N105, N121 );
not g121 ( new_n227_, N105 );
not g122 ( new_n228_, N121 );
and g123 ( new_n229_, new_n227_, new_n228_ );
or g124 ( new_n230_, new_n229_, new_n226_ );
and g125 ( new_n231_, new_n230_, keyIn_0_7 );
not g126 ( new_n232_, new_n231_ );
or g127 ( new_n233_, new_n230_, keyIn_0_7 );
and g128 ( new_n234_, new_n232_, new_n233_ );
not g129 ( new_n235_, new_n234_ );
and g130 ( new_n236_, N73, N89 );
not g131 ( new_n237_, N73 );
not g132 ( new_n238_, N89 );
and g133 ( new_n239_, new_n237_, new_n238_ );
or g134 ( new_n240_, new_n239_, new_n236_ );
and g135 ( new_n241_, new_n235_, new_n240_ );
not g136 ( new_n242_, new_n241_ );
or g137 ( new_n243_, new_n235_, new_n240_ );
and g138 ( new_n244_, new_n242_, new_n243_ );
or g139 ( new_n245_, new_n225_, new_n244_ );
and g140 ( new_n246_, new_n222_, new_n224_, new_n244_ );
not g141 ( new_n247_, new_n246_ );
and g142 ( new_n248_, new_n245_, new_n247_ );
not g143 ( new_n249_, keyIn_0_2 );
not g144 ( new_n250_, N41 );
not g145 ( new_n251_, N45 );
and g146 ( new_n252_, new_n250_, new_n251_ );
or g147 ( new_n253_, new_n252_, new_n189_ );
and g148 ( new_n254_, new_n253_, new_n249_ );
or g149 ( new_n255_, new_n254_, new_n193_ );
not g150 ( new_n256_, N37 );
and g151 ( new_n257_, new_n151_, new_n256_ );
or g152 ( new_n258_, new_n257_, new_n197_ );
and g153 ( new_n259_, new_n258_, keyIn_0_1 );
or g154 ( new_n260_, new_n259_, new_n202_ );
and g155 ( new_n261_, new_n255_, new_n260_ );
or g156 ( new_n262_, new_n261_, new_n206_ );
and g157 ( new_n263_, new_n262_, keyIn_0_8 );
or g158 ( new_n264_, new_n263_, new_n210_ );
and g159 ( new_n265_, N49, N53 );
not g160 ( new_n266_, new_n265_ );
or g161 ( new_n267_, N49, N53 );
and g162 ( new_n268_, new_n266_, new_n267_ );
and g163 ( new_n269_, N57, N61 );
not g164 ( new_n270_, new_n269_ );
or g165 ( new_n271_, N57, N61 );
and g166 ( new_n272_, new_n270_, new_n271_ );
or g167 ( new_n273_, new_n268_, new_n272_ );
and g168 ( new_n274_, new_n268_, new_n272_ );
not g169 ( new_n275_, new_n274_ );
and g170 ( new_n276_, new_n275_, new_n273_ );
and g171 ( new_n277_, new_n264_, new_n276_ );
not g172 ( new_n278_, new_n276_ );
and g173 ( new_n279_, new_n212_, new_n278_ );
or g174 ( new_n280_, new_n277_, new_n279_ );
and g175 ( new_n281_, N134, N137 );
and g176 ( new_n282_, new_n280_, new_n281_ );
or g177 ( new_n283_, new_n212_, new_n278_ );
or g178 ( new_n284_, new_n264_, new_n276_ );
and g179 ( new_n285_, new_n284_, new_n283_ );
not g180 ( new_n286_, new_n281_ );
and g181 ( new_n287_, new_n285_, new_n286_ );
or g182 ( new_n288_, new_n282_, new_n287_ );
and g183 ( new_n289_, N101, N117 );
not g184 ( new_n290_, N101 );
not g185 ( new_n291_, N117 );
and g186 ( new_n292_, new_n290_, new_n291_ );
or g187 ( new_n293_, new_n292_, new_n289_ );
and g188 ( new_n294_, N69, N85 );
and g189 ( new_n295_, new_n108_, new_n122_ );
or g190 ( new_n296_, new_n295_, new_n294_ );
and g191 ( new_n297_, new_n293_, new_n296_ );
not g192 ( new_n298_, new_n293_ );
not g193 ( new_n299_, new_n296_ );
and g194 ( new_n300_, new_n298_, new_n299_ );
or g195 ( new_n301_, new_n300_, new_n297_ );
not g196 ( new_n302_, new_n301_ );
and g197 ( new_n303_, new_n288_, new_n302_ );
or g198 ( new_n304_, new_n285_, new_n286_ );
or g199 ( new_n305_, new_n280_, new_n281_ );
and g200 ( new_n306_, new_n305_, new_n304_, new_n301_ );
or g201 ( new_n307_, new_n303_, new_n306_ );
not g202 ( new_n308_, new_n307_ );
or g203 ( new_n309_, new_n308_, keyIn_0_14 );
not g204 ( new_n310_, keyIn_0_0 );
or g205 ( new_n311_, N17, N21 );
not g206 ( new_n312_, new_n311_ );
and g207 ( new_n313_, N17, N21 );
or g208 ( new_n314_, new_n312_, new_n313_ );
and g209 ( new_n315_, new_n314_, new_n310_ );
not g210 ( new_n316_, new_n313_ );
and g211 ( new_n317_, new_n316_, keyIn_0_0, new_n311_ );
or g212 ( new_n318_, new_n315_, new_n317_ );
and g213 ( new_n319_, N25, N29 );
not g214 ( new_n320_, N25 );
not g215 ( new_n321_, N29 );
and g216 ( new_n322_, new_n320_, new_n321_ );
or g217 ( new_n323_, new_n322_, new_n319_ );
not g218 ( new_n324_, new_n323_ );
and g219 ( new_n325_, new_n318_, new_n324_ );
and g220 ( new_n326_, new_n316_, new_n311_ );
or g221 ( new_n327_, new_n326_, keyIn_0_0 );
not g222 ( new_n328_, new_n317_ );
and g223 ( new_n329_, new_n327_, new_n328_ );
and g224 ( new_n330_, new_n329_, new_n323_ );
or g225 ( new_n331_, new_n325_, new_n330_ );
and g226 ( new_n332_, new_n331_, new_n185_ );
or g227 ( new_n333_, new_n329_, new_n323_ );
or g228 ( new_n334_, new_n318_, new_n324_ );
and g229 ( new_n335_, new_n334_, new_n333_ );
and g230 ( new_n336_, new_n335_, new_n186_ );
or g231 ( new_n337_, new_n332_, new_n336_ );
and g232 ( new_n338_, N133, N137 );
and g233 ( new_n339_, new_n337_, new_n338_ );
not g234 ( new_n340_, new_n339_ );
or g235 ( new_n341_, new_n337_, new_n338_ );
and g236 ( new_n342_, new_n340_, new_n341_ );
and g237 ( new_n343_, N65, N81 );
and g238 ( new_n344_, new_n106_, new_n120_ );
or g239 ( new_n345_, new_n344_, new_n343_ );
and g240 ( new_n346_, N97, N113 );
not g241 ( new_n347_, N97 );
not g242 ( new_n348_, N113 );
and g243 ( new_n349_, new_n347_, new_n348_ );
or g244 ( new_n350_, new_n349_, new_n346_ );
and g245 ( new_n351_, new_n345_, new_n350_ );
not g246 ( new_n352_, new_n345_ );
not g247 ( new_n353_, new_n350_ );
and g248 ( new_n354_, new_n352_, new_n353_ );
or g249 ( new_n355_, new_n354_, new_n351_ );
not g250 ( new_n356_, new_n355_ );
or g251 ( new_n357_, new_n342_, new_n356_ );
and g252 ( new_n358_, new_n342_, new_n356_ );
not g253 ( new_n359_, new_n358_ );
and g254 ( new_n360_, new_n359_, new_n357_ );
not g255 ( new_n361_, new_n360_ );
not g256 ( new_n362_, keyIn_0_14 );
or g257 ( new_n363_, new_n307_, new_n362_ );
and g258 ( new_n364_, new_n248_, new_n309_, new_n361_, new_n363_ );
not g259 ( new_n365_, keyIn_0_15 );
not g260 ( new_n366_, keyIn_0_10 );
or g261 ( new_n367_, new_n335_, new_n276_ );
or g262 ( new_n368_, new_n331_, new_n278_ );
and g263 ( new_n369_, new_n368_, new_n367_ );
and g264 ( new_n370_, N136, N137 );
not g265 ( new_n371_, new_n370_ );
and g266 ( new_n372_, new_n369_, new_n371_ );
and g267 ( new_n373_, new_n331_, new_n278_ );
and g268 ( new_n374_, new_n335_, new_n276_ );
or g269 ( new_n375_, new_n373_, new_n374_ );
and g270 ( new_n376_, new_n375_, new_n370_ );
or g271 ( new_n377_, new_n376_, new_n372_ );
and g272 ( new_n378_, new_n377_, new_n366_ );
or g273 ( new_n379_, new_n375_, new_n370_ );
or g274 ( new_n380_, new_n369_, new_n371_ );
and g275 ( new_n381_, new_n379_, new_n380_ );
and g276 ( new_n382_, new_n381_, keyIn_0_10 );
or g277 ( new_n383_, new_n378_, new_n382_ );
and g278 ( new_n384_, N109, N125 );
not g279 ( new_n385_, N109 );
not g280 ( new_n386_, N125 );
and g281 ( new_n387_, new_n385_, new_n386_ );
or g282 ( new_n388_, new_n387_, new_n384_ );
and g283 ( new_n389_, N77, N93 );
not g284 ( new_n390_, N77 );
not g285 ( new_n391_, N93 );
and g286 ( new_n392_, new_n390_, new_n391_ );
or g287 ( new_n393_, new_n392_, new_n389_ );
and g288 ( new_n394_, new_n388_, new_n393_ );
not g289 ( new_n395_, new_n388_ );
not g290 ( new_n396_, new_n393_ );
and g291 ( new_n397_, new_n395_, new_n396_ );
or g292 ( new_n398_, new_n397_, new_n394_ );
and g293 ( new_n399_, new_n383_, new_n398_ );
or g294 ( new_n400_, new_n381_, keyIn_0_10 );
or g295 ( new_n401_, new_n377_, new_n366_ );
and g296 ( new_n402_, new_n401_, new_n400_ );
not g297 ( new_n403_, new_n398_ );
and g298 ( new_n404_, new_n402_, new_n403_ );
or g299 ( new_n405_, new_n399_, new_n404_ );
and g300 ( new_n406_, new_n405_, new_n365_ );
or g301 ( new_n407_, new_n402_, new_n403_ );
or g302 ( new_n408_, new_n383_, new_n398_ );
and g303 ( new_n409_, new_n408_, new_n407_ );
and g304 ( new_n410_, new_n409_, keyIn_0_15 );
or g305 ( new_n411_, new_n406_, new_n410_ );
and g306 ( new_n412_, N97, N101 );
and g307 ( new_n413_, new_n347_, new_n290_ );
or g308 ( new_n414_, new_n413_, new_n412_ );
and g309 ( new_n415_, new_n414_, keyIn_0_3 );
not g310 ( new_n416_, new_n415_ );
or g311 ( new_n417_, new_n414_, keyIn_0_3 );
and g312 ( new_n418_, new_n416_, new_n417_ );
not g313 ( new_n419_, new_n418_ );
and g314 ( new_n420_, N105, N109 );
and g315 ( new_n421_, new_n227_, new_n385_ );
or g316 ( new_n422_, new_n421_, new_n420_ );
and g317 ( new_n423_, new_n419_, new_n422_ );
not g318 ( new_n424_, new_n423_ );
or g319 ( new_n425_, new_n419_, new_n422_ );
and g320 ( new_n426_, new_n424_, new_n425_ );
and g321 ( new_n427_, N121, N125 );
and g322 ( new_n428_, new_n228_, new_n386_ );
or g323 ( new_n429_, new_n428_, new_n427_ );
and g324 ( new_n430_, new_n429_, keyIn_0_4 );
not g325 ( new_n431_, new_n430_ );
or g326 ( new_n432_, new_n429_, keyIn_0_4 );
and g327 ( new_n433_, new_n431_, new_n432_ );
not g328 ( new_n434_, new_n433_ );
and g329 ( new_n435_, N113, N117 );
and g330 ( new_n436_, new_n348_, new_n291_ );
or g331 ( new_n437_, new_n436_, new_n435_ );
and g332 ( new_n438_, new_n434_, new_n437_ );
not g333 ( new_n439_, new_n438_ );
or g334 ( new_n440_, new_n434_, new_n437_ );
and g335 ( new_n441_, new_n439_, new_n440_ );
or g336 ( new_n442_, new_n426_, new_n441_ );
and g337 ( new_n443_, new_n426_, new_n441_ );
not g338 ( new_n444_, new_n443_ );
and g339 ( new_n445_, new_n444_, new_n442_ );
and g340 ( new_n446_, N130, N137 );
or g341 ( new_n447_, new_n445_, new_n446_ );
not g342 ( new_n448_, new_n425_ );
or g343 ( new_n449_, new_n448_, new_n423_ );
not g344 ( new_n450_, new_n441_ );
and g345 ( new_n451_, new_n450_, new_n449_ );
not g346 ( new_n452_, new_n446_ );
or g347 ( new_n453_, new_n451_, new_n443_, new_n452_ );
and g348 ( new_n454_, new_n447_, new_n453_ );
and g349 ( new_n455_, N37, N53 );
not g350 ( new_n456_, N53 );
and g351 ( new_n457_, new_n256_, new_n456_ );
or g352 ( new_n458_, new_n457_, new_n455_ );
and g353 ( new_n459_, N5, N21 );
not g354 ( new_n460_, N21 );
and g355 ( new_n461_, new_n173_, new_n460_ );
or g356 ( new_n462_, new_n461_, new_n459_ );
and g357 ( new_n463_, new_n458_, new_n462_ );
not g358 ( new_n464_, new_n458_ );
not g359 ( new_n465_, new_n462_ );
and g360 ( new_n466_, new_n464_, new_n465_ );
or g361 ( new_n467_, new_n466_, new_n463_ );
not g362 ( new_n468_, new_n467_ );
or g363 ( new_n469_, new_n454_, new_n468_ );
not g364 ( new_n470_, new_n447_ );
not g365 ( new_n471_, new_n453_ );
or g366 ( new_n472_, new_n470_, new_n471_, new_n467_ );
and g367 ( new_n473_, new_n469_, new_n472_ );
not g368 ( new_n474_, new_n473_ );
and g369 ( new_n475_, new_n449_, new_n119_ );
and g370 ( new_n476_, new_n426_, new_n118_ );
or g371 ( new_n477_, new_n475_, new_n476_ );
and g372 ( new_n478_, N131, N137 );
and g373 ( new_n479_, new_n477_, new_n478_ );
or g374 ( new_n480_, new_n426_, new_n118_ );
not g375 ( new_n481_, new_n476_ );
and g376 ( new_n482_, new_n481_, new_n480_ );
not g377 ( new_n483_, new_n478_ );
and g378 ( new_n484_, new_n482_, new_n483_ );
or g379 ( new_n485_, new_n484_, new_n479_ );
and g380 ( new_n486_, N41, N57 );
not g381 ( new_n487_, N57 );
and g382 ( new_n488_, new_n250_, new_n487_ );
or g383 ( new_n489_, new_n488_, new_n486_ );
and g384 ( new_n490_, new_n489_, keyIn_0_6 );
not g385 ( new_n491_, new_n490_ );
or g386 ( new_n492_, new_n489_, keyIn_0_6 );
and g387 ( new_n493_, new_n491_, new_n492_ );
not g388 ( new_n494_, new_n493_ );
and g389 ( new_n495_, new_n320_, N9 );
and g390 ( new_n496_, new_n177_, N25 );
or g391 ( new_n497_, new_n495_, new_n496_ );
and g392 ( new_n498_, new_n494_, new_n497_ );
not g393 ( new_n499_, new_n498_ );
or g394 ( new_n500_, new_n494_, new_n497_ );
and g395 ( new_n501_, new_n499_, new_n500_ );
not g396 ( new_n502_, new_n501_ );
and g397 ( new_n503_, new_n485_, new_n502_ );
or g398 ( new_n504_, new_n482_, new_n483_ );
or g399 ( new_n505_, new_n477_, new_n478_ );
and g400 ( new_n506_, new_n504_, new_n505_ );
and g401 ( new_n507_, new_n506_, new_n501_ );
or g402 ( new_n508_, new_n503_, new_n507_ );
and g403 ( new_n509_, new_n508_, keyIn_0_12 );
or g404 ( new_n510_, new_n509_, new_n474_ );
not g405 ( new_n511_, keyIn_0_12 );
or g406 ( new_n512_, new_n506_, new_n501_ );
or g407 ( new_n513_, new_n485_, new_n502_ );
and g408 ( new_n514_, new_n513_, new_n512_ );
or g409 ( new_n515_, new_n473_, new_n514_, new_n511_ );
not g410 ( new_n516_, new_n169_ );
or g411 ( new_n517_, new_n441_, new_n132_ );
not g412 ( new_n518_, new_n517_ );
and g413 ( new_n519_, new_n441_, new_n132_ );
or g414 ( new_n520_, new_n518_, new_n519_ );
and g415 ( new_n521_, N132, N137 );
and g416 ( new_n522_, new_n520_, new_n521_ );
not g417 ( new_n523_, new_n519_ );
not g418 ( new_n524_, new_n521_ );
and g419 ( new_n525_, new_n523_, new_n517_, new_n524_ );
or g420 ( new_n526_, new_n522_, new_n525_ );
and g421 ( new_n527_, N45, N61 );
not g422 ( new_n528_, N61 );
and g423 ( new_n529_, new_n251_, new_n528_ );
or g424 ( new_n530_, new_n529_, new_n527_ );
and g425 ( new_n531_, N13, N29 );
and g426 ( new_n532_, new_n178_, new_n321_ );
or g427 ( new_n533_, new_n532_, new_n531_ );
and g428 ( new_n534_, new_n530_, new_n533_ );
not g429 ( new_n535_, new_n530_ );
not g430 ( new_n536_, new_n533_ );
and g431 ( new_n537_, new_n535_, new_n536_ );
or g432 ( new_n538_, new_n537_, new_n534_ );
and g433 ( new_n539_, new_n526_, new_n538_ );
not g434 ( new_n540_, new_n522_ );
not g435 ( new_n541_, new_n525_ );
not g436 ( new_n542_, new_n538_ );
and g437 ( new_n543_, new_n540_, new_n541_, new_n542_ );
or g438 ( new_n544_, new_n539_, new_n543_ );
not g439 ( new_n545_, new_n544_ );
and g440 ( new_n546_, new_n545_, new_n516_ );
and g441 ( new_n547_, new_n510_, new_n515_, new_n546_ );
and g442 ( new_n548_, new_n544_, new_n514_ );
not g443 ( new_n549_, keyIn_0_11 );
and g444 ( new_n550_, new_n169_, new_n549_ );
and g445 ( new_n551_, new_n516_, keyIn_0_11 );
or g446 ( new_n552_, new_n551_, new_n550_ );
and g447 ( new_n553_, new_n548_, new_n552_, new_n473_ );
and g448 ( new_n554_, new_n553_, keyIn_0_19 );
or g449 ( new_n555_, new_n553_, keyIn_0_19 );
not g450 ( new_n556_, new_n555_ );
and g451 ( new_n557_, new_n514_, new_n169_ );
or g452 ( new_n558_, new_n473_, keyIn_0_13 );
and g453 ( new_n559_, new_n473_, keyIn_0_13 );
not g454 ( new_n560_, new_n559_ );
and g455 ( new_n561_, new_n560_, new_n545_, new_n557_, new_n558_ );
or g456 ( new_n562_, new_n556_, new_n547_, new_n554_, new_n561_ );
and g457 ( new_n563_, new_n562_, new_n364_, new_n411_ );
or g458 ( new_n564_, new_n563_, new_n170_ );
and g459 ( new_n565_, new_n563_, new_n170_ );
not g460 ( new_n566_, new_n565_ );
and g461 ( new_n567_, new_n566_, new_n564_ );
not g462 ( new_n568_, new_n567_ );
and g463 ( new_n569_, new_n568_, new_n169_ );
not g464 ( new_n570_, new_n569_ );
and g465 ( new_n571_, new_n570_, N1 );
and g466 ( new_n572_, new_n569_, new_n147_ );
or g467 ( N724, new_n571_, new_n572_ );
and g468 ( new_n574_, new_n568_, new_n474_ );
not g469 ( new_n575_, new_n574_ );
and g470 ( new_n576_, new_n575_, N5 );
and g471 ( new_n577_, new_n574_, new_n173_ );
or g472 ( N725, new_n576_, new_n577_ );
or g473 ( new_n579_, new_n567_, new_n514_ );
and g474 ( new_n580_, new_n579_, N9 );
or g475 ( new_n581_, new_n364_, new_n170_ );
and g476 ( new_n582_, new_n567_, new_n581_ );
not g477 ( new_n583_, new_n582_ );
and g478 ( new_n584_, new_n583_, new_n177_, new_n508_ );
or g479 ( new_n585_, new_n584_, new_n580_ );
and g480 ( new_n586_, new_n585_, keyIn_0_30 );
not g481 ( new_n587_, keyIn_0_30 );
not g482 ( new_n588_, new_n580_ );
not g483 ( new_n589_, new_n584_ );
and g484 ( new_n590_, new_n589_, new_n587_, new_n588_ );
or g485 ( N726, new_n586_, new_n590_ );
or g486 ( new_n592_, new_n567_, new_n545_ );
and g487 ( new_n593_, new_n592_, N13 );
and g488 ( new_n594_, new_n568_, new_n178_, new_n544_ );
or g489 ( new_n595_, new_n593_, new_n594_ );
and g490 ( new_n596_, new_n595_, keyIn_0_31 );
not g491 ( new_n597_, keyIn_0_31 );
not g492 ( new_n598_, new_n593_ );
not g493 ( new_n599_, new_n594_ );
and g494 ( new_n600_, new_n598_, new_n597_, new_n599_ );
or g495 ( N727, new_n596_, new_n600_ );
and g496 ( new_n602_, new_n264_, new_n185_ );
or g497 ( new_n603_, new_n602_, new_n214_ );
and g498 ( new_n604_, new_n603_, keyIn_0_5 );
or g499 ( new_n605_, new_n604_, new_n218_ );
not g500 ( new_n606_, new_n221_ );
and g501 ( new_n607_, new_n605_, new_n606_ );
or g502 ( new_n608_, new_n607_, new_n223_ );
not g503 ( new_n609_, new_n244_ );
and g504 ( new_n610_, new_n608_, new_n609_ );
or g505 ( new_n611_, new_n610_, new_n246_ );
and g506 ( new_n612_, new_n611_, new_n405_ );
or g507 ( new_n613_, new_n308_, new_n360_ );
not g508 ( new_n614_, new_n613_ );
and g509 ( new_n615_, new_n562_, new_n612_, new_n614_ );
and g510 ( new_n616_, new_n615_, new_n169_ );
not g511 ( new_n617_, new_n616_ );
and g512 ( new_n618_, new_n617_, N17 );
and g513 ( new_n619_, new_n616_, new_n145_ );
or g514 ( N728, new_n618_, new_n619_ );
and g515 ( new_n621_, new_n615_, new_n474_ );
not g516 ( new_n622_, new_n621_ );
and g517 ( new_n623_, new_n622_, N21 );
and g518 ( new_n624_, new_n621_, new_n460_ );
or g519 ( N729, new_n623_, new_n624_ );
not g520 ( new_n626_, keyIn_0_25 );
and g521 ( new_n627_, new_n615_, new_n508_ );
or g522 ( new_n628_, new_n627_, new_n626_ );
and g523 ( new_n629_, new_n627_, new_n626_ );
not g524 ( new_n630_, new_n629_ );
and g525 ( new_n631_, new_n630_, new_n628_ );
not g526 ( new_n632_, new_n631_ );
and g527 ( new_n633_, new_n632_, new_n320_ );
and g528 ( new_n634_, new_n631_, N25 );
or g529 ( N730, new_n633_, new_n634_ );
not g530 ( new_n636_, keyIn_0_26 );
and g531 ( new_n637_, new_n615_, new_n544_ );
or g532 ( new_n638_, new_n637_, new_n636_ );
and g533 ( new_n639_, new_n637_, new_n636_ );
not g534 ( new_n640_, new_n639_ );
and g535 ( new_n641_, new_n640_, new_n638_ );
not g536 ( new_n642_, new_n641_ );
and g537 ( new_n643_, new_n642_, N29 );
and g538 ( new_n644_, new_n641_, new_n321_ );
or g539 ( N731, new_n643_, new_n644_ );
and g540 ( new_n646_, new_n562_, new_n308_ );
not g541 ( new_n647_, keyIn_0_16 );
or g542 ( new_n648_, new_n360_, new_n647_ );
or g543 ( new_n649_, new_n361_, keyIn_0_16 );
and g544 ( new_n650_, new_n248_, new_n409_, new_n648_, new_n649_ );
and g545 ( new_n651_, new_n646_, new_n650_ );
and g546 ( new_n652_, new_n651_, new_n169_ );
not g547 ( new_n653_, new_n652_ );
and g548 ( new_n654_, new_n653_, N33 );
and g549 ( new_n655_, new_n652_, new_n151_ );
or g550 ( N732, new_n654_, new_n655_ );
and g551 ( new_n657_, new_n651_, new_n474_ );
not g552 ( new_n658_, new_n657_ );
and g553 ( new_n659_, new_n658_, N37 );
and g554 ( new_n660_, new_n657_, new_n256_ );
or g555 ( N733, new_n659_, new_n660_ );
and g556 ( new_n662_, new_n651_, new_n508_ );
not g557 ( new_n663_, new_n662_ );
and g558 ( new_n664_, new_n663_, N41 );
and g559 ( new_n665_, new_n662_, new_n250_ );
or g560 ( N734, new_n664_, new_n665_ );
and g561 ( new_n667_, new_n651_, new_n544_ );
not g562 ( new_n668_, new_n667_ );
and g563 ( new_n669_, new_n668_, N45 );
and g564 ( new_n670_, new_n667_, new_n251_ );
or g565 ( N735, new_n669_, new_n670_ );
not g566 ( new_n672_, keyIn_0_17 );
or g567 ( new_n673_, new_n361_, new_n672_ );
or g568 ( new_n674_, new_n360_, keyIn_0_17 );
and g569 ( new_n675_, new_n646_, new_n612_, new_n673_, new_n674_ );
and g570 ( new_n676_, new_n675_, new_n169_ );
not g571 ( new_n677_, new_n676_ );
and g572 ( new_n678_, new_n677_, N49 );
and g573 ( new_n679_, new_n676_, new_n152_ );
or g574 ( N736, new_n678_, new_n679_ );
and g575 ( new_n681_, new_n675_, new_n474_ );
not g576 ( new_n682_, new_n681_ );
and g577 ( new_n683_, new_n682_, N53 );
and g578 ( new_n684_, new_n681_, new_n456_ );
or g579 ( N737, new_n683_, new_n684_ );
and g580 ( new_n686_, new_n675_, new_n508_ );
not g581 ( new_n687_, new_n686_ );
and g582 ( new_n688_, new_n687_, N57 );
and g583 ( new_n689_, new_n686_, new_n487_ );
or g584 ( N738, new_n688_, new_n689_ );
and g585 ( new_n691_, new_n675_, new_n544_ );
not g586 ( new_n692_, new_n691_ );
and g587 ( new_n693_, new_n692_, N61 );
and g588 ( new_n694_, new_n691_, new_n528_ );
or g589 ( N739, new_n693_, new_n694_ );
and g590 ( new_n696_, new_n473_, new_n169_ );
and g591 ( new_n697_, new_n696_, new_n508_, new_n545_ );
not g592 ( new_n698_, new_n697_ );
not g593 ( new_n699_, keyIn_0_23 );
or g594 ( new_n700_, new_n405_, new_n307_, new_n361_ );
or g595 ( new_n701_, new_n248_, new_n700_ );
and g596 ( new_n702_, new_n701_, keyIn_0_22 );
not g597 ( new_n703_, keyIn_0_22 );
and g598 ( new_n704_, new_n308_, new_n360_, new_n409_ );
and g599 ( new_n705_, new_n611_, new_n704_ );
and g600 ( new_n706_, new_n705_, new_n703_ );
or g601 ( new_n707_, new_n702_, new_n706_ );
not g602 ( new_n708_, keyIn_0_18 );
or g603 ( new_n709_, new_n248_, new_n708_ );
and g604 ( new_n710_, new_n245_, new_n708_, new_n247_ );
not g605 ( new_n711_, new_n710_ );
and g606 ( new_n712_, new_n709_, new_n711_ );
and g607 ( new_n713_, new_n614_, new_n409_ );
not g608 ( new_n714_, new_n713_ );
or g609 ( new_n715_, new_n712_, new_n714_ );
not g610 ( new_n716_, keyIn_0_21 );
and g611 ( new_n717_, new_n409_, new_n307_, new_n360_ );
and g612 ( new_n718_, new_n717_, new_n245_, new_n247_ );
or g613 ( new_n719_, new_n718_, new_n716_ );
not g614 ( new_n720_, new_n719_ );
and g615 ( new_n721_, new_n718_, new_n716_ );
or g616 ( new_n722_, new_n720_, new_n721_ );
and g617 ( new_n723_, new_n307_, new_n360_ );
not g618 ( new_n724_, new_n723_ );
or g619 ( new_n725_, new_n248_, new_n409_, new_n724_ );
and g620 ( new_n726_, new_n725_, keyIn_0_20 );
or g621 ( new_n727_, new_n248_, new_n724_, keyIn_0_20, new_n409_ );
not g622 ( new_n728_, new_n727_ );
or g623 ( new_n729_, new_n726_, new_n728_ );
and g624 ( new_n730_, new_n729_, new_n707_, new_n715_, new_n722_ );
or g625 ( new_n731_, new_n730_, new_n699_ );
not g626 ( new_n732_, new_n721_ );
and g627 ( new_n733_, new_n732_, new_n719_ );
not g628 ( new_n734_, keyIn_0_20 );
and g629 ( new_n735_, new_n611_, new_n405_, new_n723_ );
or g630 ( new_n736_, new_n735_, new_n734_ );
and g631 ( new_n737_, new_n736_, new_n727_ );
or g632 ( new_n738_, new_n737_, new_n733_ );
or g633 ( new_n739_, new_n705_, new_n703_ );
or g634 ( new_n740_, new_n701_, keyIn_0_22 );
and g635 ( new_n741_, new_n740_, new_n739_ );
and g636 ( new_n742_, new_n611_, keyIn_0_18 );
or g637 ( new_n743_, new_n742_, new_n710_ );
and g638 ( new_n744_, new_n743_, new_n713_ );
or g639 ( new_n745_, new_n741_, new_n744_, keyIn_0_23 );
or g640 ( new_n746_, new_n745_, new_n738_ );
and g641 ( new_n747_, new_n731_, new_n746_ );
not g642 ( new_n748_, new_n747_ );
and g643 ( new_n749_, new_n748_, new_n361_ );
not g644 ( new_n750_, new_n749_ );
or g645 ( new_n751_, new_n750_, new_n698_ );
and g646 ( new_n752_, new_n751_, N65 );
and g647 ( new_n753_, new_n749_, new_n106_, new_n697_ );
or g648 ( N740, new_n752_, new_n753_ );
and g649 ( new_n755_, new_n748_, new_n308_ );
not g650 ( new_n756_, new_n755_ );
or g651 ( new_n757_, new_n756_, new_n698_ );
and g652 ( new_n758_, new_n757_, N69 );
and g653 ( new_n759_, new_n755_, new_n108_, new_n697_ );
or g654 ( N741, new_n758_, new_n759_ );
and g655 ( new_n761_, new_n748_, new_n248_ );
not g656 ( new_n762_, new_n761_ );
or g657 ( new_n763_, new_n762_, new_n698_ );
and g658 ( new_n764_, new_n763_, N73 );
and g659 ( new_n765_, new_n761_, new_n237_, new_n697_ );
or g660 ( N742, new_n764_, new_n765_ );
and g661 ( new_n767_, new_n748_, new_n405_ );
not g662 ( new_n768_, new_n767_ );
or g663 ( new_n769_, new_n768_, new_n698_ );
and g664 ( new_n770_, new_n769_, N77 );
and g665 ( new_n771_, new_n767_, new_n390_, new_n697_ );
or g666 ( N743, new_n770_, new_n771_ );
and g667 ( new_n773_, new_n548_, new_n696_ );
not g668 ( new_n774_, new_n773_ );
or g669 ( new_n775_, new_n750_, new_n774_ );
and g670 ( new_n776_, new_n775_, N81 );
and g671 ( new_n777_, new_n749_, new_n120_, new_n773_ );
or g672 ( N744, new_n776_, new_n777_ );
not g673 ( new_n779_, keyIn_0_27 );
or g674 ( new_n780_, new_n747_, new_n307_, new_n774_ );
and g675 ( new_n781_, new_n780_, new_n779_ );
and g676 ( new_n782_, new_n748_, keyIn_0_27, new_n308_, new_n773_ );
or g677 ( new_n783_, new_n781_, new_n782_ );
and g678 ( new_n784_, new_n783_, new_n122_ );
not g679 ( new_n785_, new_n781_ );
not g680 ( new_n786_, new_n782_ );
and g681 ( new_n787_, new_n785_, N85, new_n786_ );
or g682 ( N745, new_n784_, new_n787_ );
or g683 ( new_n789_, new_n762_, new_n774_ );
and g684 ( new_n790_, new_n789_, N89 );
and g685 ( new_n791_, new_n761_, new_n238_, new_n773_ );
or g686 ( N746, new_n790_, new_n791_ );
or g687 ( new_n793_, new_n768_, new_n774_ );
and g688 ( new_n794_, new_n793_, N93 );
and g689 ( new_n795_, new_n767_, new_n391_, new_n773_ );
or g690 ( N747, new_n794_, new_n795_ );
and g691 ( new_n797_, new_n546_, new_n474_, new_n508_ );
not g692 ( new_n798_, new_n797_ );
or g693 ( new_n799_, new_n750_, new_n798_ );
and g694 ( new_n800_, new_n799_, N97 );
and g695 ( new_n801_, new_n749_, new_n347_, new_n797_ );
or g696 ( N748, new_n800_, new_n801_ );
or g697 ( new_n803_, new_n756_, new_n798_ );
and g698 ( new_n804_, new_n803_, N101 );
and g699 ( new_n805_, new_n755_, new_n290_, new_n797_ );
or g700 ( N749, new_n804_, new_n805_ );
or g701 ( new_n807_, new_n762_, new_n798_ );
and g702 ( new_n808_, new_n807_, N105 );
and g703 ( new_n809_, new_n761_, new_n227_, new_n797_ );
or g704 ( N750, new_n808_, new_n809_ );
or g705 ( new_n811_, new_n747_, new_n409_, new_n798_ );
and g706 ( new_n812_, new_n811_, keyIn_0_28 );
not g707 ( new_n813_, keyIn_0_28 );
and g708 ( new_n814_, new_n748_, new_n813_, new_n405_, new_n797_ );
or g709 ( new_n815_, new_n812_, new_n814_ );
and g710 ( new_n816_, new_n815_, new_n385_ );
not g711 ( new_n817_, new_n812_ );
not g712 ( new_n818_, new_n814_ );
and g713 ( new_n819_, new_n817_, N109, new_n818_ );
or g714 ( N751, new_n816_, new_n819_ );
and g715 ( new_n821_, new_n548_, new_n516_, new_n474_ );
not g716 ( new_n822_, new_n821_ );
or g717 ( new_n823_, new_n750_, new_n822_ );
and g718 ( new_n824_, new_n823_, N113 );
and g719 ( new_n825_, new_n749_, new_n348_, new_n821_ );
or g720 ( N752, new_n824_, new_n825_ );
or g721 ( new_n827_, new_n747_, new_n307_, new_n822_ );
and g722 ( new_n828_, new_n827_, keyIn_0_29 );
not g723 ( new_n829_, keyIn_0_29 );
and g724 ( new_n830_, new_n748_, new_n829_, new_n308_, new_n821_ );
or g725 ( new_n831_, new_n828_, new_n830_ );
and g726 ( new_n832_, new_n831_, N117 );
not g727 ( new_n833_, new_n828_ );
not g728 ( new_n834_, new_n830_ );
and g729 ( new_n835_, new_n833_, new_n291_, new_n834_ );
or g730 ( N753, new_n832_, new_n835_ );
or g731 ( new_n837_, new_n762_, new_n822_ );
and g732 ( new_n838_, new_n837_, N121 );
and g733 ( new_n839_, new_n761_, new_n228_, new_n821_ );
or g734 ( N754, new_n838_, new_n839_ );
or g735 ( new_n841_, new_n768_, new_n822_ );
and g736 ( new_n842_, new_n841_, N125 );
and g737 ( new_n843_, new_n767_, new_n386_, new_n821_ );
or g738 ( N755, new_n842_, new_n843_ );
endmodule