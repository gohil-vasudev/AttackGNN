module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n1233_, new_n479_, new_n1105_, new_n1215_, new_n1249_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n1157_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n566_, new_n641_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n1207_, new_n1211_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1237_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n1210_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n1213_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n1188_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n1221_, new_n1167_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n1238_, new_n792_, new_n1058_, new_n953_, new_n1162_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n449_, new_n580_, new_n639_, new_n484_, new_n832_, new_n766_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n1250_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n1151_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1203_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n1257_, new_n988_, new_n478_, new_n694_, new_n461_, new_n1228_, new_n710_, new_n971_, new_n565_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1196_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1216_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n1214_, new_n1005_, new_n883_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n1170_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n1182_, new_n1200_, new_n650_, new_n708_, new_n750_, new_n1217_, new_n887_, new_n355_, new_n926_, new_n353_, new_n1222_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1226_, new_n778_, new_n452_, new_n1198_, new_n1219_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n1168_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n1007_, new_n935_, new_n1241_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1159_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n398_, new_n1177_, new_n646_, new_n395_, new_n538_, new_n1026_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1106_, new_n1132_, new_n473_, new_n1147_, new_n1229_, new_n790_, new_n1081_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n1234_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n1245_, new_n402_, new_n663_, new_n579_, new_n1209_, new_n659_, new_n1254_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n1201_, new_n948_, new_n1231_, new_n762_, new_n1055_, new_n1193_, new_n838_, new_n923_, new_n1187_, new_n469_, new_n1205_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n1253_, new_n1256_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n1171_, new_n688_, new_n1255_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n1160_, new_n1166_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1175_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n380_, new_n1251_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n1252_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n1191_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1224_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n1186_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1261_, new_n1040_, new_n1246_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n1179_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n1240_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n1195_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n1227_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n1248_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n1244_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n769_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n1220_, new_n989_, new_n1204_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n1206_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n905_, new_n539_, new_n1258_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n1197_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1194_, new_n1077_, new_n1243_, new_n490_, new_n560_, new_n1100_, new_n1230_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n1165_, new_n1259_, new_n425_, new_n896_, new_n802_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n1236_, new_n709_, new_n866_, new_n1235_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1225_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n1192_, new_n573_, new_n765_, new_n405_, new_n1103_;

and g000 ( new_n343_, N29, N42 );
and g001 ( N388, new_n343_, N75 );
not g002 ( new_n345_, N80 );
nand g003 ( new_n346_, N29, N36 );
nor g004 ( N389, new_n346_, new_n345_ );
not g005 ( new_n348_, N42 );
nor g006 ( N390, new_n346_, new_n348_ );
and g007 ( N391, N85, N86 );
not g008 ( new_n351_, N13 );
nand g009 ( new_n352_, N1, N8 );
nor g010 ( new_n353_, new_n352_, new_n351_ );
and g011 ( N418, new_n353_, N17 );
not g012 ( new_n355_, N390 );
nand g013 ( new_n356_, N1, N26 );
nand g014 ( new_n357_, N13, N17 );
nor g015 ( new_n358_, new_n356_, new_n357_ );
nand g016 ( new_n359_, new_n355_, new_n358_ );
xnor g017 ( N419, new_n359_, keyIn_0_8 );
nand g018 ( new_n361_, N59, N75 );
or g019 ( N420, new_n361_, new_n345_ );
and g020 ( new_n363_, N36, N59 );
nand g021 ( N421, new_n363_, N80 );
nand g022 ( N422, new_n363_, N42 );
not g023 ( new_n366_, N90 );
nor g024 ( new_n367_, N87, N88 );
nor g025 ( N423, new_n367_, new_n366_ );
nand g026 ( new_n369_, new_n358_, N390 );
xnor g027 ( N446, new_n369_, keyIn_0_25 );
not g028 ( new_n371_, N51 );
nor g029 ( new_n372_, new_n356_, new_n371_ );
xnor g030 ( N447, new_n372_, keyIn_0_0 );
nand g031 ( new_n374_, new_n353_, N55 );
nand g032 ( new_n375_, N29, N68 );
nor g033 ( new_n376_, new_n374_, new_n375_ );
xor g034 ( N448, new_n376_, keyIn_0_12 );
and g035 ( new_n378_, N59, N68 );
nand g036 ( new_n379_, new_n378_, N74 );
nor g037 ( new_n380_, new_n374_, new_n379_ );
xor g038 ( N449, new_n380_, keyIn_0_13 );
not g039 ( new_n382_, N89 );
nor g040 ( N450, new_n367_, new_n382_ );
xor g041 ( new_n384_, N111, N116 );
xnor g042 ( new_n385_, new_n384_, keyIn_0_17 );
xor g043 ( new_n386_, new_n385_, keyIn_0_31 );
xnor g044 ( new_n387_, N121, N126 );
xnor g045 ( new_n388_, new_n387_, keyIn_0_18 );
xor g046 ( new_n389_, new_n388_, keyIn_0_32 );
nand g047 ( new_n390_, new_n386_, new_n389_ );
xor g048 ( new_n391_, new_n390_, keyIn_0_43 );
nand g049 ( new_n392_, new_n385_, new_n388_ );
xor g050 ( new_n393_, new_n392_, keyIn_0_33 );
nand g051 ( new_n394_, new_n391_, new_n393_ );
xnor g052 ( new_n395_, new_n394_, keyIn_0_53 );
not g053 ( new_n396_, new_n395_ );
nor g054 ( new_n397_, new_n396_, N135 );
xor g055 ( new_n398_, new_n397_, keyIn_0_73 );
nand g056 ( new_n399_, new_n396_, N135 );
xnor g057 ( new_n400_, new_n399_, keyIn_0_72 );
nand g058 ( new_n401_, new_n398_, new_n400_ );
xnor g059 ( new_n402_, new_n401_, keyIn_0_95 );
not g060 ( new_n403_, N130 );
xor g061 ( new_n404_, N101, N106 );
xnor g062 ( new_n405_, new_n404_, keyIn_0_16 );
xor g063 ( new_n406_, new_n405_, keyIn_0_29 );
xnor g064 ( new_n407_, N91, N96 );
xnor g065 ( new_n408_, new_n407_, keyIn_0_15 );
xor g066 ( new_n409_, new_n408_, keyIn_0_28 );
nand g067 ( new_n410_, new_n406_, new_n409_ );
nand g068 ( new_n411_, new_n410_, keyIn_0_42 );
nand g069 ( new_n412_, new_n405_, new_n408_ );
xor g070 ( new_n413_, new_n412_, keyIn_0_30 );
nor g071 ( new_n414_, new_n410_, keyIn_0_42 );
nor g072 ( new_n415_, new_n414_, new_n413_ );
nand g073 ( new_n416_, new_n415_, new_n411_ );
xor g074 ( new_n417_, new_n416_, keyIn_0_52 );
nor g075 ( new_n418_, new_n417_, new_n403_ );
xnor g076 ( new_n419_, new_n418_, keyIn_0_70 );
nand g077 ( new_n420_, new_n417_, new_n403_ );
xnor g078 ( new_n421_, new_n420_, keyIn_0_71 );
nand g079 ( new_n422_, new_n419_, new_n421_ );
xor g080 ( new_n423_, new_n422_, keyIn_0_94 );
nand g081 ( new_n424_, new_n402_, new_n423_ );
xnor g082 ( new_n425_, new_n424_, keyIn_0_116 );
nor g083 ( new_n426_, new_n402_, new_n423_ );
xnor g084 ( new_n427_, new_n426_, keyIn_0_106 );
nand g085 ( new_n428_, new_n427_, new_n425_ );
xnor g086 ( N767, new_n428_, keyIn_0_139 );
not g087 ( new_n430_, N207 );
xor g088 ( new_n431_, N195, N201 );
xnor g089 ( new_n432_, new_n431_, keyIn_0_24 );
xnor g090 ( new_n433_, new_n432_, keyIn_0_39 );
xor g091 ( new_n434_, N183, N189 );
xnor g092 ( new_n435_, new_n434_, keyIn_0_23 );
xnor g093 ( new_n436_, new_n435_, keyIn_0_38 );
nand g094 ( new_n437_, new_n433_, new_n436_ );
nand g095 ( new_n438_, new_n437_, keyIn_0_50 );
nand g096 ( new_n439_, new_n432_, new_n435_ );
xor g097 ( new_n440_, new_n439_, keyIn_0_40 );
nor g098 ( new_n441_, new_n437_, keyIn_0_50 );
nor g099 ( new_n442_, new_n441_, new_n440_ );
nand g100 ( new_n443_, new_n442_, new_n438_ );
xor g101 ( new_n444_, new_n443_, keyIn_0_69 );
nor g102 ( new_n445_, new_n444_, new_n430_ );
xor g103 ( new_n446_, new_n445_, keyIn_0_92 );
nand g104 ( new_n447_, new_n444_, new_n430_ );
xor g105 ( new_n448_, new_n447_, keyIn_0_93 );
nand g106 ( new_n449_, new_n446_, new_n448_ );
xnor g107 ( new_n450_, new_n449_, keyIn_0_105 );
not g108 ( new_n451_, keyIn_0_49 );
xor g109 ( new_n452_, N159, N165 );
xnor g110 ( new_n453_, new_n452_, keyIn_0_21 );
xor g111 ( new_n454_, new_n453_, keyIn_0_35 );
xnor g112 ( new_n455_, N171, N177 );
xnor g113 ( new_n456_, new_n455_, keyIn_0_22 );
xor g114 ( new_n457_, new_n456_, keyIn_0_36 );
nand g115 ( new_n458_, new_n454_, new_n457_ );
nor g116 ( new_n459_, new_n458_, new_n451_ );
nand g117 ( new_n460_, new_n453_, new_n456_ );
xor g118 ( new_n461_, new_n460_, keyIn_0_37 );
nand g119 ( new_n462_, new_n458_, new_n451_ );
nand g120 ( new_n463_, new_n462_, new_n461_ );
nor g121 ( new_n464_, new_n463_, new_n459_ );
xor g122 ( new_n465_, new_n464_, keyIn_0_68 );
nor g123 ( new_n466_, new_n465_, N130 );
xor g124 ( new_n467_, new_n466_, keyIn_0_91 );
nand g125 ( new_n468_, new_n465_, N130 );
xnor g126 ( new_n469_, new_n468_, keyIn_0_90 );
nand g127 ( new_n470_, new_n467_, new_n469_ );
xor g128 ( new_n471_, new_n470_, keyIn_0_104 );
nand g129 ( new_n472_, new_n471_, new_n450_ );
xnor g130 ( new_n473_, new_n472_, keyIn_0_117 );
nor g131 ( new_n474_, new_n471_, new_n450_ );
xor g132 ( new_n475_, new_n474_, keyIn_0_115 );
nand g133 ( new_n476_, new_n475_, new_n473_ );
xnor g134 ( N768, new_n476_, keyIn_0_140 );
not g135 ( new_n478_, keyIn_0_210 );
not g136 ( new_n479_, keyIn_0_202 );
not g137 ( new_n480_, N261 );
not g138 ( new_n481_, N201 );
not g139 ( new_n482_, keyIn_0_103 );
not g140 ( new_n483_, keyIn_0_63 );
not g141 ( new_n484_, keyIn_0_9 );
and g142 ( new_n485_, N1, N26 );
nand g143 ( new_n486_, new_n485_, N51 );
nand g144 ( new_n487_, new_n486_, keyIn_0_0 );
not g145 ( new_n488_, keyIn_0_0 );
nand g146 ( new_n489_, new_n372_, new_n488_ );
nand g147 ( new_n490_, new_n487_, new_n489_ );
nand g148 ( new_n491_, new_n490_, new_n484_ );
nand g149 ( new_n492_, N447, keyIn_0_9 );
nand g150 ( new_n493_, new_n492_, new_n491_ );
xnor g151 ( new_n494_, new_n493_, keyIn_0_26 );
not g152 ( new_n495_, N17 );
nand g153 ( new_n496_, N59, N156 );
xnor g154 ( new_n497_, new_n496_, keyIn_0_5 );
not g155 ( new_n498_, new_n497_ );
nor g156 ( new_n499_, new_n498_, new_n495_ );
nand g157 ( new_n500_, new_n494_, new_n499_ );
nand g158 ( new_n501_, new_n500_, keyIn_0_48 );
not g159 ( new_n502_, keyIn_0_48 );
not g160 ( new_n503_, keyIn_0_26 );
nand g161 ( new_n504_, new_n493_, new_n503_ );
xnor g162 ( new_n505_, new_n490_, keyIn_0_9 );
nand g163 ( new_n506_, new_n505_, keyIn_0_26 );
nand g164 ( new_n507_, new_n506_, new_n504_ );
not g165 ( new_n508_, new_n499_ );
nor g166 ( new_n509_, new_n507_, new_n508_ );
nand g167 ( new_n510_, new_n509_, new_n502_ );
nand g168 ( new_n511_, new_n501_, new_n510_ );
nand g169 ( new_n512_, new_n511_, N1 );
xnor g170 ( new_n513_, new_n512_, new_n483_ );
nand g171 ( new_n514_, new_n513_, N153 );
nand g172 ( new_n515_, new_n514_, keyIn_0_88 );
not g173 ( new_n516_, keyIn_0_88 );
not g174 ( new_n517_, N153 );
xnor g175 ( new_n518_, new_n512_, keyIn_0_63 );
nor g176 ( new_n519_, new_n518_, new_n517_ );
nand g177 ( new_n520_, new_n519_, new_n516_ );
nand g178 ( new_n521_, new_n520_, new_n515_ );
not g179 ( new_n522_, keyIn_0_89 );
not g180 ( new_n523_, keyIn_0_54 );
not g181 ( new_n524_, keyIn_0_20 );
nand g182 ( new_n525_, N17, N42 );
xor g183 ( new_n526_, new_n525_, keyIn_0_7 );
not g184 ( new_n527_, keyIn_0_6 );
nor g185 ( new_n528_, N17, N42 );
xnor g186 ( new_n529_, new_n528_, new_n527_ );
nand g187 ( new_n530_, new_n526_, new_n529_ );
nand g188 ( new_n531_, new_n530_, new_n524_ );
nor g189 ( new_n532_, new_n530_, new_n524_ );
nor g190 ( new_n533_, new_n532_, new_n496_ );
and g191 ( new_n534_, new_n533_, new_n531_ );
nand g192 ( new_n535_, new_n494_, new_n534_ );
nor g193 ( new_n536_, new_n535_, keyIn_0_47 );
not g194 ( new_n537_, new_n536_ );
not g195 ( new_n538_, keyIn_0_34 );
nand g196 ( new_n539_, N17, N51 );
nor g197 ( new_n540_, new_n352_, new_n539_ );
xnor g198 ( new_n541_, new_n540_, keyIn_0_1 );
xnor g199 ( new_n542_, new_n541_, keyIn_0_10 );
nor g200 ( new_n543_, new_n361_, new_n348_ );
xnor g201 ( new_n544_, new_n543_, keyIn_0_3 );
xnor g202 ( new_n545_, new_n544_, keyIn_0_14 );
nand g203 ( new_n546_, new_n542_, new_n545_ );
xnor g204 ( new_n547_, new_n546_, new_n538_ );
not g205 ( new_n548_, keyIn_0_47 );
nand g206 ( new_n549_, new_n533_, new_n531_ );
nor g207 ( new_n550_, new_n507_, new_n549_ );
nor g208 ( new_n551_, new_n550_, new_n548_ );
nor g209 ( new_n552_, new_n551_, new_n547_ );
nand g210 ( new_n553_, new_n552_, new_n537_ );
nand g211 ( new_n554_, new_n553_, new_n523_ );
xnor g212 ( new_n555_, new_n546_, keyIn_0_34 );
nand g213 ( new_n556_, new_n535_, keyIn_0_47 );
nand g214 ( new_n557_, new_n556_, new_n555_ );
nor g215 ( new_n558_, new_n557_, new_n536_ );
nand g216 ( new_n559_, new_n558_, keyIn_0_54 );
nand g217 ( new_n560_, new_n554_, new_n559_ );
nand g218 ( new_n561_, new_n560_, N126 );
xnor g219 ( new_n562_, new_n561_, new_n522_ );
nand g220 ( new_n563_, new_n562_, new_n521_ );
nor g221 ( new_n564_, new_n563_, new_n482_ );
not g222 ( new_n565_, new_n564_ );
nand g223 ( new_n566_, N29, N75 );
nor g224 ( new_n567_, new_n566_, new_n345_ );
xor g225 ( new_n568_, new_n567_, keyIn_0_2 );
nor g226 ( new_n569_, new_n507_, new_n568_ );
nand g227 ( new_n570_, new_n569_, N55 );
nor g228 ( new_n571_, new_n570_, keyIn_0_46 );
xnor g229 ( new_n572_, keyIn_0_4, N268 );
xor g230 ( new_n573_, new_n572_, keyIn_0_19 );
and g231 ( new_n574_, new_n570_, keyIn_0_46 );
or g232 ( new_n575_, new_n574_, new_n573_ );
nor g233 ( new_n576_, new_n575_, new_n571_ );
xor g234 ( new_n577_, new_n576_, keyIn_0_67 );
nand g235 ( new_n578_, new_n563_, new_n482_ );
and g236 ( new_n579_, new_n578_, new_n577_ );
nand g237 ( new_n580_, new_n579_, new_n565_ );
nand g238 ( new_n581_, new_n580_, keyIn_0_114 );
not g239 ( new_n582_, keyIn_0_114 );
nand g240 ( new_n583_, new_n578_, new_n577_ );
nor g241 ( new_n584_, new_n583_, new_n564_ );
nand g242 ( new_n585_, new_n584_, new_n582_ );
nand g243 ( new_n586_, new_n581_, new_n585_ );
nand g244 ( new_n587_, new_n586_, new_n481_ );
xnor g245 ( new_n588_, new_n587_, keyIn_0_138 );
not g246 ( new_n589_, keyIn_0_137 );
xnor g247 ( new_n590_, new_n584_, keyIn_0_114 );
nand g248 ( new_n591_, new_n590_, N201 );
nand g249 ( new_n592_, new_n591_, new_n589_ );
nor g250 ( new_n593_, new_n586_, new_n481_ );
nand g251 ( new_n594_, new_n593_, keyIn_0_137 );
nand g252 ( new_n595_, new_n592_, new_n594_ );
nor g253 ( new_n596_, new_n588_, new_n595_ );
xor g254 ( new_n597_, new_n596_, keyIn_0_163 );
nor g255 ( new_n598_, new_n597_, new_n480_ );
xnor g256 ( new_n599_, new_n598_, keyIn_0_185 );
nand g257 ( new_n600_, new_n597_, new_n480_ );
xnor g258 ( new_n601_, new_n600_, keyIn_0_184 );
nand g259 ( new_n602_, new_n599_, new_n601_ );
nand g260 ( new_n603_, new_n602_, new_n479_ );
not g261 ( new_n604_, N219 );
nor g262 ( new_n605_, new_n602_, new_n479_ );
nor g263 ( new_n606_, new_n605_, new_n604_ );
nand g264 ( new_n607_, new_n606_, new_n603_ );
nand g265 ( new_n608_, new_n607_, new_n478_ );
and g266 ( new_n609_, N121, N210 );
nor g267 ( new_n610_, new_n607_, new_n478_ );
nor g268 ( new_n611_, new_n610_, new_n609_ );
nand g269 ( new_n612_, new_n611_, new_n608_ );
nand g270 ( new_n613_, new_n612_, keyIn_0_216 );
nor g271 ( new_n614_, new_n612_, keyIn_0_216 );
not g272 ( new_n615_, N228 );
nor g273 ( new_n616_, new_n597_, new_n615_ );
xnor g274 ( new_n617_, new_n595_, keyIn_0_162 );
and g275 ( new_n618_, new_n617_, N237 );
nor g276 ( new_n619_, new_n616_, new_n618_ );
nor g277 ( new_n620_, new_n619_, keyIn_0_203 );
nand g278 ( new_n621_, new_n619_, keyIn_0_203 );
not g279 ( new_n622_, keyIn_0_164 );
nand g280 ( new_n623_, N255, N267 );
nand g281 ( new_n624_, new_n590_, N246 );
nand g282 ( new_n625_, new_n624_, new_n623_ );
nor g283 ( new_n626_, new_n625_, new_n622_ );
and g284 ( new_n627_, N42, N72 );
nand g285 ( new_n628_, new_n378_, new_n627_ );
nor g286 ( new_n629_, new_n374_, new_n628_ );
xnor g287 ( new_n630_, new_n629_, keyIn_0_11 );
nand g288 ( new_n631_, new_n630_, N73 );
xor g289 ( new_n632_, new_n631_, keyIn_0_27 );
xnor g290 ( new_n633_, new_n632_, keyIn_0_41 );
xnor g291 ( new_n634_, new_n633_, keyIn_0_51 );
not g292 ( new_n635_, new_n634_ );
nand g293 ( new_n636_, new_n635_, N201 );
nand g294 ( new_n637_, new_n625_, new_n622_ );
nand g295 ( new_n638_, new_n637_, new_n636_ );
nor g296 ( new_n639_, new_n638_, new_n626_ );
nand g297 ( new_n640_, new_n621_, new_n639_ );
or g298 ( new_n641_, new_n640_, new_n620_ );
nor g299 ( new_n642_, new_n614_, new_n641_ );
nand g300 ( new_n643_, new_n642_, new_n613_ );
xnor g301 ( N850, new_n643_, keyIn_0_222 );
not g302 ( new_n645_, keyIn_0_230 );
not g303 ( new_n646_, keyIn_0_219 );
nand g304 ( new_n647_, new_n513_, N143 );
xor g305 ( new_n648_, new_n647_, keyIn_0_82 );
nand g306 ( new_n649_, new_n560_, N111 );
xor g307 ( new_n650_, new_n649_, keyIn_0_83 );
nand g308 ( new_n651_, new_n648_, new_n650_ );
xor g309 ( new_n652_, new_n651_, keyIn_0_100 );
xor g310 ( new_n653_, new_n576_, keyIn_0_64 );
nand g311 ( new_n654_, new_n652_, new_n653_ );
xnor g312 ( new_n655_, new_n654_, keyIn_0_111 );
nand g313 ( new_n656_, new_n655_, N183 );
xnor g314 ( new_n657_, new_n656_, keyIn_0_130 );
nor g315 ( new_n658_, new_n655_, N183 );
xnor g316 ( new_n659_, new_n658_, keyIn_0_131 );
nand g317 ( new_n660_, new_n659_, new_n657_ );
xnor g318 ( new_n661_, new_n660_, keyIn_0_154 );
not g319 ( new_n662_, keyIn_0_196 );
not g320 ( new_n663_, keyIn_0_167 );
nor g321 ( new_n664_, new_n588_, new_n480_ );
not g322 ( new_n665_, N189 );
not g323 ( new_n666_, keyIn_0_112 );
nand g324 ( new_n667_, new_n513_, N146 );
nand g325 ( new_n668_, new_n667_, keyIn_0_84 );
not g326 ( new_n669_, keyIn_0_84 );
not g327 ( new_n670_, N146 );
nor g328 ( new_n671_, new_n518_, new_n670_ );
nand g329 ( new_n672_, new_n671_, new_n669_ );
nand g330 ( new_n673_, new_n672_, new_n668_ );
not g331 ( new_n674_, keyIn_0_85 );
nand g332 ( new_n675_, new_n560_, N116 );
xnor g333 ( new_n676_, new_n675_, new_n674_ );
nand g334 ( new_n677_, new_n676_, new_n673_ );
nor g335 ( new_n678_, new_n677_, keyIn_0_101 );
xor g336 ( new_n679_, new_n576_, keyIn_0_65 );
nand g337 ( new_n680_, new_n677_, keyIn_0_101 );
nand g338 ( new_n681_, new_n680_, new_n679_ );
nor g339 ( new_n682_, new_n681_, new_n678_ );
xnor g340 ( new_n683_, new_n682_, new_n666_ );
nand g341 ( new_n684_, new_n683_, new_n665_ );
nand g342 ( new_n685_, new_n684_, keyIn_0_134 );
not g343 ( new_n686_, keyIn_0_134 );
not g344 ( new_n687_, new_n678_ );
and g345 ( new_n688_, new_n680_, new_n679_ );
nand g346 ( new_n689_, new_n688_, new_n687_ );
nand g347 ( new_n690_, new_n689_, new_n666_ );
nand g348 ( new_n691_, new_n682_, keyIn_0_112 );
nand g349 ( new_n692_, new_n690_, new_n691_ );
nor g350 ( new_n693_, new_n692_, N189 );
nand g351 ( new_n694_, new_n693_, new_n686_ );
nand g352 ( new_n695_, new_n685_, new_n694_ );
not g353 ( new_n696_, N195 );
not g354 ( new_n697_, keyIn_0_113 );
not g355 ( new_n698_, keyIn_0_102 );
not g356 ( new_n699_, keyIn_0_86 );
nand g357 ( new_n700_, new_n513_, N149 );
nand g358 ( new_n701_, new_n700_, new_n699_ );
not g359 ( new_n702_, N149 );
nor g360 ( new_n703_, new_n518_, new_n702_ );
nand g361 ( new_n704_, new_n703_, keyIn_0_86 );
nand g362 ( new_n705_, new_n704_, new_n701_ );
not g363 ( new_n706_, keyIn_0_87 );
nand g364 ( new_n707_, new_n560_, N121 );
xnor g365 ( new_n708_, new_n707_, new_n706_ );
nand g366 ( new_n709_, new_n708_, new_n705_ );
nor g367 ( new_n710_, new_n709_, new_n698_ );
xor g368 ( new_n711_, new_n576_, keyIn_0_66 );
nand g369 ( new_n712_, new_n709_, new_n698_ );
nand g370 ( new_n713_, new_n712_, new_n711_ );
nor g371 ( new_n714_, new_n713_, new_n710_ );
xnor g372 ( new_n715_, new_n714_, new_n697_ );
nand g373 ( new_n716_, new_n715_, new_n696_ );
nand g374 ( new_n717_, new_n716_, keyIn_0_136 );
not g375 ( new_n718_, keyIn_0_136 );
not g376 ( new_n719_, new_n710_ );
and g377 ( new_n720_, new_n712_, new_n711_ );
nand g378 ( new_n721_, new_n720_, new_n719_ );
nand g379 ( new_n722_, new_n721_, new_n697_ );
nand g380 ( new_n723_, new_n714_, keyIn_0_113 );
nand g381 ( new_n724_, new_n722_, new_n723_ );
nor g382 ( new_n725_, new_n724_, N195 );
nand g383 ( new_n726_, new_n725_, new_n718_ );
nand g384 ( new_n727_, new_n717_, new_n726_ );
and g385 ( new_n728_, new_n695_, new_n727_ );
nand g386 ( new_n729_, new_n728_, new_n664_ );
nand g387 ( new_n730_, new_n729_, new_n663_ );
not g388 ( new_n731_, keyIn_0_138 );
nand g389 ( new_n732_, new_n587_, new_n731_ );
nor g390 ( new_n733_, new_n590_, N201 );
nand g391 ( new_n734_, new_n733_, keyIn_0_138 );
nand g392 ( new_n735_, new_n734_, new_n732_ );
nand g393 ( new_n736_, new_n735_, N261 );
nand g394 ( new_n737_, new_n695_, new_n727_ );
nor g395 ( new_n738_, new_n737_, new_n736_ );
nand g396 ( new_n739_, new_n738_, keyIn_0_167 );
nand g397 ( new_n740_, new_n730_, new_n739_ );
not g398 ( new_n741_, keyIn_0_177 );
not g399 ( new_n742_, keyIn_0_133 );
nand g400 ( new_n743_, new_n692_, N189 );
nand g401 ( new_n744_, new_n743_, new_n742_ );
nor g402 ( new_n745_, new_n683_, new_n665_ );
nand g403 ( new_n746_, new_n745_, keyIn_0_133 );
nand g404 ( new_n747_, new_n746_, new_n744_ );
nand g405 ( new_n748_, new_n747_, keyIn_0_156 );
not g406 ( new_n749_, keyIn_0_156 );
xnor g407 ( new_n750_, new_n743_, keyIn_0_133 );
nand g408 ( new_n751_, new_n750_, new_n749_ );
nand g409 ( new_n752_, new_n751_, new_n748_ );
nand g410 ( new_n753_, new_n752_, new_n741_ );
xnor g411 ( new_n754_, new_n747_, new_n749_ );
nand g412 ( new_n755_, new_n754_, keyIn_0_177 );
nand g413 ( new_n756_, new_n755_, new_n753_ );
and g414 ( new_n757_, new_n756_, new_n740_ );
not g415 ( new_n758_, keyIn_0_187 );
not g416 ( new_n759_, keyIn_0_135 );
nand g417 ( new_n760_, new_n724_, N195 );
xnor g418 ( new_n761_, new_n760_, new_n759_ );
nand g419 ( new_n762_, new_n761_, keyIn_0_159 );
not g420 ( new_n763_, keyIn_0_159 );
xnor g421 ( new_n764_, new_n760_, keyIn_0_135 );
nand g422 ( new_n765_, new_n764_, new_n763_ );
nand g423 ( new_n766_, new_n762_, new_n765_ );
nand g424 ( new_n767_, new_n766_, new_n695_ );
xnor g425 ( new_n768_, new_n767_, new_n758_ );
nand g426 ( new_n769_, new_n757_, new_n768_ );
not g427 ( new_n770_, keyIn_0_162 );
xnor g428 ( new_n771_, new_n595_, new_n770_ );
not g429 ( new_n772_, new_n727_ );
nor g430 ( new_n773_, new_n771_, new_n772_ );
nand g431 ( new_n774_, new_n773_, new_n695_ );
nand g432 ( new_n775_, new_n774_, keyIn_0_188 );
not g433 ( new_n776_, keyIn_0_188 );
not g434 ( new_n777_, new_n695_ );
nand g435 ( new_n778_, new_n617_, new_n727_ );
nor g436 ( new_n779_, new_n778_, new_n777_ );
nand g437 ( new_n780_, new_n779_, new_n776_ );
nand g438 ( new_n781_, new_n775_, new_n780_ );
nor g439 ( new_n782_, new_n769_, new_n781_ );
nand g440 ( new_n783_, new_n782_, new_n662_ );
nand g441 ( new_n784_, new_n756_, new_n740_ );
xnor g442 ( new_n785_, new_n767_, keyIn_0_187 );
nor g443 ( new_n786_, new_n785_, new_n784_ );
xnor g444 ( new_n787_, new_n779_, keyIn_0_188 );
nand g445 ( new_n788_, new_n787_, new_n786_ );
nand g446 ( new_n789_, new_n788_, keyIn_0_196 );
nand g447 ( new_n790_, new_n783_, new_n789_ );
not g448 ( new_n791_, new_n790_ );
nand g449 ( new_n792_, new_n791_, new_n661_ );
xnor g450 ( new_n793_, new_n792_, keyIn_0_204 );
nor g451 ( new_n794_, new_n791_, new_n661_ );
xnor g452 ( new_n795_, new_n794_, keyIn_0_205 );
nand g453 ( new_n796_, new_n795_, new_n793_ );
xnor g454 ( new_n797_, new_n796_, keyIn_0_213 );
nand g455 ( new_n798_, new_n797_, N219 );
nor g456 ( new_n799_, new_n798_, new_n646_ );
nand g457 ( new_n800_, N106, N210 );
nand g458 ( new_n801_, new_n798_, new_n646_ );
nand g459 ( new_n802_, new_n801_, new_n800_ );
nor g460 ( new_n803_, new_n802_, new_n799_ );
nor g461 ( new_n804_, new_n803_, new_n645_ );
nand g462 ( new_n805_, new_n803_, new_n645_ );
not g463 ( new_n806_, keyIn_0_197 );
nor g464 ( new_n807_, new_n661_, new_n615_ );
nand g465 ( new_n808_, new_n807_, keyIn_0_175 );
xor g466 ( new_n809_, new_n657_, keyIn_0_153 );
nand g467 ( new_n810_, new_n809_, N237 );
xor g468 ( new_n811_, new_n810_, keyIn_0_176 );
nor g469 ( new_n812_, new_n807_, keyIn_0_175 );
nor g470 ( new_n813_, new_n811_, new_n812_ );
nand g471 ( new_n814_, new_n813_, new_n808_ );
nor g472 ( new_n815_, new_n814_, new_n806_ );
nand g473 ( new_n816_, new_n814_, new_n806_ );
not g474 ( new_n817_, keyIn_0_132 );
nand g475 ( new_n818_, new_n655_, N246 );
nor g476 ( new_n819_, new_n818_, new_n817_ );
nand g477 ( new_n820_, new_n635_, N183 );
nand g478 ( new_n821_, new_n818_, new_n817_ );
nand g479 ( new_n822_, new_n821_, new_n820_ );
nor g480 ( new_n823_, new_n822_, new_n819_ );
xnor g481 ( new_n824_, new_n823_, keyIn_0_155 );
nand g482 ( new_n825_, new_n816_, new_n824_ );
nor g483 ( new_n826_, new_n825_, new_n815_ );
nand g484 ( new_n827_, new_n805_, new_n826_ );
nor g485 ( new_n828_, new_n827_, new_n804_ );
xnor g486 ( N863, new_n828_, keyIn_0_240 );
not g487 ( new_n830_, keyIn_0_231 );
not g488 ( new_n831_, keyIn_0_220 );
nand g489 ( new_n832_, new_n747_, new_n695_ );
xnor g490 ( new_n833_, new_n832_, keyIn_0_157 );
xnor g491 ( new_n834_, new_n773_, keyIn_0_186 );
nand g492 ( new_n835_, new_n664_, new_n727_ );
xnor g493 ( new_n836_, new_n835_, keyIn_0_166 );
xnor g494 ( new_n837_, new_n766_, keyIn_0_180 );
nor g495 ( new_n838_, new_n836_, new_n837_ );
nand g496 ( new_n839_, new_n834_, new_n838_ );
xor g497 ( new_n840_, new_n839_, keyIn_0_198 );
nor g498 ( new_n841_, new_n840_, new_n833_ );
xnor g499 ( new_n842_, new_n841_, keyIn_0_206 );
nand g500 ( new_n843_, new_n840_, new_n833_ );
xnor g501 ( new_n844_, new_n843_, keyIn_0_207 );
nand g502 ( new_n845_, new_n842_, new_n844_ );
xor g503 ( new_n846_, new_n845_, keyIn_0_214 );
nand g504 ( new_n847_, new_n846_, N219 );
nor g505 ( new_n848_, new_n847_, new_n831_ );
nand g506 ( new_n849_, N111, N210 );
nand g507 ( new_n850_, new_n847_, new_n831_ );
nand g508 ( new_n851_, new_n850_, new_n849_ );
nor g509 ( new_n852_, new_n851_, new_n848_ );
nor g510 ( new_n853_, new_n852_, new_n830_ );
nand g511 ( new_n854_, new_n852_, new_n830_ );
not g512 ( new_n855_, keyIn_0_199 );
nand g513 ( new_n856_, new_n752_, N237 );
xor g514 ( new_n857_, new_n856_, keyIn_0_179 );
nand g515 ( new_n858_, new_n833_, N228 );
xor g516 ( new_n859_, new_n858_, keyIn_0_178 );
nand g517 ( new_n860_, new_n859_, new_n857_ );
nor g518 ( new_n861_, new_n860_, new_n855_ );
nand g519 ( new_n862_, new_n860_, new_n855_ );
not g520 ( new_n863_, keyIn_0_158 );
nand g521 ( new_n864_, new_n692_, N246 );
nand g522 ( new_n865_, N255, N259 );
and g523 ( new_n866_, new_n864_, new_n865_ );
nor g524 ( new_n867_, new_n866_, new_n863_ );
nand g525 ( new_n868_, new_n866_, new_n863_ );
nand g526 ( new_n869_, new_n635_, N189 );
nand g527 ( new_n870_, new_n868_, new_n869_ );
nor g528 ( new_n871_, new_n870_, new_n867_ );
nand g529 ( new_n872_, new_n862_, new_n871_ );
nor g530 ( new_n873_, new_n872_, new_n861_ );
nand g531 ( new_n874_, new_n854_, new_n873_ );
nor g532 ( new_n875_, new_n874_, new_n853_ );
xnor g533 ( N864, new_n875_, keyIn_0_241 );
not g534 ( new_n877_, keyIn_0_215 );
nand g535 ( new_n878_, new_n764_, new_n727_ );
xor g536 ( new_n879_, new_n878_, keyIn_0_160 );
xnor g537 ( new_n880_, new_n617_, keyIn_0_183 );
xnor g538 ( new_n881_, new_n736_, keyIn_0_165 );
nand g539 ( new_n882_, new_n880_, new_n881_ );
xor g540 ( new_n883_, new_n882_, keyIn_0_200 );
nand g541 ( new_n884_, new_n883_, new_n879_ );
xor g542 ( new_n885_, new_n884_, keyIn_0_209 );
nor g543 ( new_n886_, new_n883_, new_n879_ );
xnor g544 ( new_n887_, new_n886_, keyIn_0_208 );
nand g545 ( new_n888_, new_n885_, new_n887_ );
nand g546 ( new_n889_, new_n888_, new_n877_ );
nor g547 ( new_n890_, new_n888_, new_n877_ );
nor g548 ( new_n891_, new_n890_, new_n604_ );
nand g549 ( new_n892_, new_n891_, new_n889_ );
nand g550 ( new_n893_, new_n892_, keyIn_0_221 );
and g551 ( new_n894_, N116, N210 );
nor g552 ( new_n895_, new_n892_, keyIn_0_221 );
nor g553 ( new_n896_, new_n895_, new_n894_ );
nand g554 ( new_n897_, new_n896_, new_n893_ );
xnor g555 ( new_n898_, new_n897_, keyIn_0_232 );
not g556 ( new_n899_, keyIn_0_201 );
nand g557 ( new_n900_, new_n879_, N228 );
nand g558 ( new_n901_, new_n900_, keyIn_0_181 );
nand g559 ( new_n902_, new_n766_, N237 );
xnor g560 ( new_n903_, new_n902_, keyIn_0_182 );
nor g561 ( new_n904_, new_n900_, keyIn_0_181 );
nor g562 ( new_n905_, new_n904_, new_n903_ );
nand g563 ( new_n906_, new_n905_, new_n901_ );
nor g564 ( new_n907_, new_n906_, new_n899_ );
nand g565 ( new_n908_, new_n906_, new_n899_ );
nand g566 ( new_n909_, new_n724_, N246 );
nand g567 ( new_n910_, N255, N260 );
nand g568 ( new_n911_, new_n909_, new_n910_ );
nor g569 ( new_n912_, new_n911_, keyIn_0_161 );
nand g570 ( new_n913_, new_n635_, N195 );
nand g571 ( new_n914_, new_n911_, keyIn_0_161 );
nand g572 ( new_n915_, new_n914_, new_n913_ );
nor g573 ( new_n916_, new_n915_, new_n912_ );
nand g574 ( new_n917_, new_n908_, new_n916_ );
nor g575 ( new_n918_, new_n917_, new_n907_ );
nand g576 ( new_n919_, new_n898_, new_n918_ );
xor g577 ( N865, new_n919_, keyIn_0_242 );
not g578 ( new_n921_, keyIn_0_226 );
nand g579 ( new_n922_, new_n560_, N96 );
nand g580 ( new_n923_, new_n922_, keyIn_0_76 );
not g581 ( new_n924_, N138 );
nor g582 ( new_n925_, new_n371_, new_n924_ );
nor g583 ( new_n926_, new_n922_, keyIn_0_76 );
nor g584 ( new_n927_, new_n926_, new_n925_ );
nand g585 ( new_n928_, new_n927_, new_n923_ );
nor g586 ( new_n929_, new_n928_, keyIn_0_97 );
nand g587 ( new_n930_, new_n928_, keyIn_0_97 );
nand g588 ( new_n931_, new_n569_, N17 );
nor g589 ( new_n932_, new_n931_, keyIn_0_45 );
and g590 ( new_n933_, new_n931_, keyIn_0_45 );
or g591 ( new_n934_, new_n933_, new_n572_ );
nor g592 ( new_n935_, new_n934_, new_n932_ );
xnor g593 ( new_n936_, new_n935_, keyIn_0_58 );
and g594 ( new_n937_, new_n497_, N55 );
nand g595 ( new_n938_, new_n494_, new_n937_ );
xor g596 ( new_n939_, new_n938_, keyIn_0_44 );
nand g597 ( new_n940_, new_n939_, N146 );
xor g598 ( new_n941_, new_n940_, keyIn_0_57 );
nand g599 ( new_n942_, new_n936_, new_n941_ );
xor g600 ( new_n943_, new_n942_, keyIn_0_77 );
nand g601 ( new_n944_, new_n943_, new_n930_ );
nor g602 ( new_n945_, new_n944_, new_n929_ );
xor g603 ( new_n946_, new_n945_, keyIn_0_108 );
nor g604 ( new_n947_, new_n946_, N165 );
xor g605 ( new_n948_, new_n947_, keyIn_0_122 );
xnor g606 ( new_n949_, new_n935_, keyIn_0_60 );
nand g607 ( new_n950_, new_n939_, N149 );
xnor g608 ( new_n951_, new_n950_, keyIn_0_59 );
nand g609 ( new_n952_, new_n949_, new_n951_ );
xor g610 ( new_n953_, new_n952_, keyIn_0_79 );
nand g611 ( new_n954_, new_n560_, N101 );
nand g612 ( new_n955_, new_n954_, keyIn_0_78 );
nor g613 ( new_n956_, new_n495_, new_n924_ );
nor g614 ( new_n957_, new_n954_, keyIn_0_78 );
nor g615 ( new_n958_, new_n957_, new_n956_ );
nand g616 ( new_n959_, new_n958_, new_n955_ );
xnor g617 ( new_n960_, new_n959_, keyIn_0_98 );
nand g618 ( new_n961_, new_n960_, new_n953_ );
xor g619 ( new_n962_, new_n961_, keyIn_0_109 );
or g620 ( new_n963_, new_n962_, N171 );
xnor g621 ( new_n964_, new_n963_, keyIn_0_125 );
not g622 ( new_n965_, new_n964_ );
nand g623 ( new_n966_, new_n948_, new_n965_ );
not g624 ( new_n967_, new_n966_ );
not g625 ( new_n968_, keyIn_0_212 );
nand g626 ( new_n969_, new_n790_, new_n659_ );
nand g627 ( new_n970_, new_n969_, keyIn_0_211 );
not g628 ( new_n971_, keyIn_0_211 );
and g629 ( new_n972_, new_n790_, new_n659_ );
nand g630 ( new_n973_, new_n972_, new_n971_ );
nand g631 ( new_n974_, new_n973_, new_n970_ );
xnor g632 ( new_n975_, new_n809_, keyIn_0_174 );
not g633 ( new_n976_, new_n975_ );
nand g634 ( new_n977_, new_n974_, new_n976_ );
xnor g635 ( new_n978_, new_n977_, new_n968_ );
not g636 ( new_n979_, keyIn_0_99 );
nand g637 ( new_n980_, new_n560_, N106 );
nand g638 ( new_n981_, new_n980_, keyIn_0_80 );
and g639 ( new_n982_, N138, N152 );
nor g640 ( new_n983_, new_n980_, keyIn_0_80 );
nor g641 ( new_n984_, new_n983_, new_n982_ );
nand g642 ( new_n985_, new_n984_, new_n981_ );
nand g643 ( new_n986_, new_n985_, new_n979_ );
nor g644 ( new_n987_, new_n985_, new_n979_ );
xnor g645 ( new_n988_, new_n935_, keyIn_0_62 );
nand g646 ( new_n989_, new_n939_, N153 );
xnor g647 ( new_n990_, new_n989_, keyIn_0_61 );
nand g648 ( new_n991_, new_n988_, new_n990_ );
xor g649 ( new_n992_, new_n991_, keyIn_0_81 );
nor g650 ( new_n993_, new_n992_, new_n987_ );
nand g651 ( new_n994_, new_n993_, new_n986_ );
xnor g652 ( new_n995_, new_n994_, keyIn_0_110 );
nor g653 ( new_n996_, new_n995_, N177 );
xor g654 ( new_n997_, new_n996_, keyIn_0_128 );
nor g655 ( new_n998_, new_n978_, new_n997_ );
nand g656 ( new_n999_, new_n998_, new_n967_ );
nor g657 ( new_n1000_, new_n999_, keyIn_0_225 );
not g658 ( new_n1001_, new_n1000_ );
not g659 ( new_n1002_, keyIn_0_225 );
nand g660 ( new_n1003_, new_n977_, keyIn_0_212 );
xnor g661 ( new_n1004_, new_n969_, new_n971_ );
nor g662 ( new_n1005_, new_n1004_, new_n975_ );
nand g663 ( new_n1006_, new_n1005_, new_n968_ );
nand g664 ( new_n1007_, new_n1006_, new_n1003_ );
not g665 ( new_n1008_, new_n997_ );
nand g666 ( new_n1009_, new_n1007_, new_n1008_ );
nor g667 ( new_n1010_, new_n1009_, new_n966_ );
nor g668 ( new_n1011_, new_n1010_, new_n1002_ );
not g669 ( new_n1012_, keyIn_0_190 );
nand g670 ( new_n1013_, new_n962_, N171 );
xor g671 ( new_n1014_, new_n1013_, keyIn_0_124 );
xnor g672 ( new_n1015_, new_n1014_, keyIn_0_147 );
nand g673 ( new_n1016_, new_n1015_, new_n948_ );
nor g674 ( new_n1017_, new_n1016_, new_n1012_ );
not g675 ( new_n1018_, keyIn_0_191 );
nand g676 ( new_n1019_, new_n995_, N177 );
xor g677 ( new_n1020_, new_n1019_, keyIn_0_127 );
xor g678 ( new_n1021_, new_n1020_, keyIn_0_150 );
nand g679 ( new_n1022_, new_n1021_, new_n967_ );
nor g680 ( new_n1023_, new_n1022_, new_n1018_ );
nor g681 ( new_n1024_, new_n1023_, new_n1017_ );
not g682 ( new_n1025_, new_n1024_ );
nand g683 ( new_n1026_, new_n1016_, new_n1012_ );
nand g684 ( new_n1027_, new_n946_, N165 );
xnor g685 ( new_n1028_, new_n1027_, keyIn_0_121 );
xor g686 ( new_n1029_, new_n1028_, keyIn_0_144 );
xnor g687 ( new_n1030_, new_n1029_, keyIn_0_168 );
nand g688 ( new_n1031_, new_n1022_, new_n1018_ );
not g689 ( new_n1032_, new_n1031_ );
nor g690 ( new_n1033_, new_n1032_, new_n1030_ );
nand g691 ( new_n1034_, new_n1033_, new_n1026_ );
nor g692 ( new_n1035_, new_n1034_, new_n1025_ );
not g693 ( new_n1036_, new_n1035_ );
nor g694 ( new_n1037_, new_n1011_, new_n1036_ );
nand g695 ( new_n1038_, new_n1037_, new_n1001_ );
nand g696 ( new_n1039_, new_n1038_, new_n921_ );
nand g697 ( new_n1040_, new_n999_, keyIn_0_225 );
nand g698 ( new_n1041_, new_n1040_, new_n1035_ );
nor g699 ( new_n1042_, new_n1041_, new_n1000_ );
nand g700 ( new_n1043_, new_n1042_, keyIn_0_226 );
nand g701 ( new_n1044_, new_n1043_, new_n1039_ );
nand g702 ( new_n1045_, new_n560_, N91 );
nand g703 ( new_n1046_, new_n1045_, keyIn_0_74 );
and g704 ( new_n1047_, N8, N138 );
nor g705 ( new_n1048_, new_n1045_, keyIn_0_74 );
nor g706 ( new_n1049_, new_n1048_, new_n1047_ );
nand g707 ( new_n1050_, new_n1049_, new_n1046_ );
nor g708 ( new_n1051_, new_n1050_, keyIn_0_96 );
nand g709 ( new_n1052_, new_n1050_, keyIn_0_96 );
xnor g710 ( new_n1053_, new_n935_, keyIn_0_56 );
nand g711 ( new_n1054_, new_n939_, N143 );
xor g712 ( new_n1055_, new_n1054_, keyIn_0_55 );
nand g713 ( new_n1056_, new_n1053_, new_n1055_ );
xor g714 ( new_n1057_, new_n1056_, keyIn_0_75 );
nand g715 ( new_n1058_, new_n1057_, new_n1052_ );
nor g716 ( new_n1059_, new_n1058_, new_n1051_ );
xor g717 ( new_n1060_, new_n1059_, keyIn_0_107 );
nor g718 ( new_n1061_, new_n1060_, N159 );
xor g719 ( new_n1062_, new_n1061_, keyIn_0_119 );
not g720 ( new_n1063_, new_n1062_ );
nand g721 ( new_n1064_, new_n1044_, new_n1063_ );
nand g722 ( new_n1065_, new_n1064_, keyIn_0_243 );
nand g723 ( new_n1066_, new_n1060_, N159 );
xnor g724 ( new_n1067_, new_n1066_, keyIn_0_118 );
xnor g725 ( new_n1068_, new_n1067_, keyIn_0_141 );
nor g726 ( new_n1069_, new_n1064_, keyIn_0_243 );
nor g727 ( new_n1070_, new_n1069_, new_n1068_ );
nand g728 ( new_n1071_, new_n1070_, new_n1065_ );
xor g729 ( N866, new_n1071_, keyIn_0_248 );
not g730 ( new_n1073_, keyIn_0_247 );
nand g731 ( new_n1074_, new_n1008_, new_n1020_ );
xnor g732 ( new_n1075_, new_n1074_, keyIn_0_151 );
nor g733 ( new_n1076_, new_n1007_, new_n1075_ );
xor g734 ( new_n1077_, new_n1076_, keyIn_0_217 );
nand g735 ( new_n1078_, new_n1007_, new_n1075_ );
xnor g736 ( new_n1079_, new_n1078_, keyIn_0_218 );
nand g737 ( new_n1080_, new_n1077_, new_n1079_ );
nor g738 ( new_n1081_, new_n1080_, keyIn_0_229 );
nand g739 ( new_n1082_, new_n1080_, keyIn_0_229 );
nand g740 ( new_n1083_, new_n1082_, N219 );
nor g741 ( new_n1084_, new_n1083_, new_n1081_ );
nor g742 ( new_n1085_, new_n1084_, keyIn_0_239 );
nand g743 ( new_n1086_, N101, N210 );
nand g744 ( new_n1087_, new_n1084_, keyIn_0_239 );
nand g745 ( new_n1088_, new_n1087_, new_n1086_ );
nor g746 ( new_n1089_, new_n1088_, new_n1085_ );
nor g747 ( new_n1090_, new_n1089_, new_n1073_ );
nand g748 ( new_n1091_, new_n1089_, new_n1073_ );
not g749 ( new_n1092_, keyIn_0_172 );
nand g750 ( new_n1093_, new_n1075_, N228 );
nand g751 ( new_n1094_, new_n1093_, new_n1092_ );
nor g752 ( new_n1095_, new_n1093_, new_n1092_ );
nand g753 ( new_n1096_, new_n1021_, N237 );
xnor g754 ( new_n1097_, new_n1096_, keyIn_0_173 );
nor g755 ( new_n1098_, new_n1095_, new_n1097_ );
nand g756 ( new_n1099_, new_n1098_, new_n1094_ );
nor g757 ( new_n1100_, new_n1099_, keyIn_0_195 );
nand g758 ( new_n1101_, new_n1099_, keyIn_0_195 );
nand g759 ( new_n1102_, new_n995_, N246 );
nand g760 ( new_n1103_, new_n1102_, keyIn_0_129 );
and g761 ( new_n1104_, new_n635_, N177 );
nor g762 ( new_n1105_, new_n1102_, keyIn_0_129 );
nor g763 ( new_n1106_, new_n1105_, new_n1104_ );
nand g764 ( new_n1107_, new_n1106_, new_n1103_ );
xnor g765 ( new_n1108_, new_n1107_, keyIn_0_152 );
nand g766 ( new_n1109_, new_n1101_, new_n1108_ );
nor g767 ( new_n1110_, new_n1109_, new_n1100_ );
nand g768 ( new_n1111_, new_n1091_, new_n1110_ );
nor g769 ( new_n1112_, new_n1111_, new_n1090_ );
xor g770 ( N874, new_n1112_, keyIn_0_249 );
not g771 ( new_n1114_, keyIn_0_253 );
not g772 ( new_n1115_, keyIn_0_250 );
not g773 ( new_n1116_, keyIn_0_244 );
not g774 ( new_n1117_, keyIn_0_233 );
nand g775 ( new_n1118_, new_n1063_, new_n1067_ );
xnor g776 ( new_n1119_, new_n1118_, keyIn_0_142 );
not g777 ( new_n1120_, new_n1119_ );
nor g778 ( new_n1121_, new_n1044_, new_n1120_ );
nand g779 ( new_n1122_, new_n1121_, new_n1117_ );
xnor g780 ( new_n1123_, new_n1038_, keyIn_0_226 );
nand g781 ( new_n1124_, new_n1123_, new_n1119_ );
nand g782 ( new_n1125_, new_n1124_, keyIn_0_233 );
nand g783 ( new_n1126_, new_n1125_, new_n1122_ );
nand g784 ( new_n1127_, new_n1044_, new_n1120_ );
xnor g785 ( new_n1128_, new_n1127_, keyIn_0_234 );
nand g786 ( new_n1129_, new_n1128_, new_n1126_ );
nand g787 ( new_n1130_, new_n1129_, new_n1116_ );
nor g788 ( new_n1131_, new_n1129_, new_n1116_ );
nor g789 ( new_n1132_, new_n1131_, new_n604_ );
nand g790 ( new_n1133_, new_n1132_, new_n1130_ );
nand g791 ( new_n1134_, new_n573_, N210 );
nand g792 ( new_n1135_, new_n1133_, new_n1134_ );
nor g793 ( new_n1136_, new_n1135_, new_n1115_ );
nand g794 ( new_n1137_, new_n1135_, new_n1115_ );
nand g795 ( new_n1138_, new_n1120_, N228 );
nand g796 ( new_n1139_, new_n1068_, N237 );
nand g797 ( new_n1140_, new_n1138_, new_n1139_ );
nor g798 ( new_n1141_, new_n1140_, keyIn_0_192 );
nand g799 ( new_n1142_, new_n1140_, keyIn_0_192 );
nand g800 ( new_n1143_, new_n1060_, N246 );
xor g801 ( new_n1144_, new_n1143_, keyIn_0_120 );
nand g802 ( new_n1145_, new_n635_, N159 );
nand g803 ( new_n1146_, new_n1144_, new_n1145_ );
xor g804 ( new_n1147_, new_n1146_, keyIn_0_143 );
nand g805 ( new_n1148_, new_n1142_, new_n1147_ );
nor g806 ( new_n1149_, new_n1148_, new_n1141_ );
nand g807 ( new_n1150_, new_n1137_, new_n1149_ );
nor g808 ( new_n1151_, new_n1150_, new_n1136_ );
xnor g809 ( N878, new_n1151_, new_n1114_ );
not g810 ( new_n1153_, keyIn_0_254 );
not g811 ( new_n1154_, keyIn_0_251 );
not g812 ( new_n1155_, keyIn_0_227 );
not g813 ( new_n1156_, keyIn_0_224 );
nand g814 ( new_n1157_, new_n998_, new_n965_ );
nand g815 ( new_n1158_, new_n1157_, new_n1156_ );
nor g816 ( new_n1159_, new_n1009_, new_n964_ );
nand g817 ( new_n1160_, new_n1159_, keyIn_0_224 );
nand g818 ( new_n1161_, new_n1158_, new_n1160_ );
not g819 ( new_n1162_, keyIn_0_189 );
nand g820 ( new_n1163_, new_n1021_, new_n965_ );
nand g821 ( new_n1164_, new_n1163_, new_n1162_ );
nor g822 ( new_n1165_, new_n1163_, new_n1162_ );
xor g823 ( new_n1166_, new_n1015_, keyIn_0_169 );
nor g824 ( new_n1167_, new_n1165_, new_n1166_ );
nand g825 ( new_n1168_, new_n1167_, new_n1164_ );
not g826 ( new_n1169_, new_n1168_ );
nand g827 ( new_n1170_, new_n1161_, new_n1169_ );
nand g828 ( new_n1171_, new_n1170_, new_n1155_ );
xnor g829 ( new_n1172_, new_n1159_, new_n1156_ );
nor g830 ( new_n1173_, new_n1172_, new_n1168_ );
nand g831 ( new_n1174_, new_n1173_, keyIn_0_227 );
nand g832 ( new_n1175_, new_n1174_, new_n1171_ );
nand g833 ( new_n1176_, new_n948_, new_n1028_ );
xnor g834 ( new_n1177_, new_n1176_, keyIn_0_145 );
nand g835 ( new_n1178_, new_n1175_, new_n1177_ );
nand g836 ( new_n1179_, new_n1178_, keyIn_0_235 );
not g837 ( new_n1180_, keyIn_0_235 );
xnor g838 ( new_n1181_, new_n1170_, keyIn_0_227 );
not g839 ( new_n1182_, new_n1177_ );
nor g840 ( new_n1183_, new_n1181_, new_n1182_ );
nand g841 ( new_n1184_, new_n1183_, new_n1180_ );
nand g842 ( new_n1185_, new_n1184_, new_n1179_ );
not g843 ( new_n1186_, keyIn_0_236 );
nand g844 ( new_n1187_, new_n1181_, new_n1182_ );
nand g845 ( new_n1188_, new_n1187_, new_n1186_ );
nor g846 ( new_n1189_, new_n1175_, new_n1177_ );
nand g847 ( new_n1190_, new_n1189_, keyIn_0_236 );
nand g848 ( new_n1191_, new_n1190_, new_n1188_ );
nand g849 ( new_n1192_, new_n1185_, new_n1191_ );
nand g850 ( new_n1193_, new_n1192_, keyIn_0_245 );
nor g851 ( new_n1194_, new_n1192_, keyIn_0_245 );
nor g852 ( new_n1195_, new_n1194_, new_n604_ );
nand g853 ( new_n1196_, new_n1195_, new_n1193_ );
nand g854 ( new_n1197_, N91, N210 );
nand g855 ( new_n1198_, new_n1196_, new_n1197_ );
xnor g856 ( new_n1199_, new_n1198_, new_n1154_ );
nand g857 ( new_n1200_, new_n1182_, N228 );
nand g858 ( new_n1201_, new_n1029_, N237 );
nand g859 ( new_n1202_, new_n1200_, new_n1201_ );
nor g860 ( new_n1203_, new_n1202_, keyIn_0_193 );
nand g861 ( new_n1204_, new_n1202_, keyIn_0_193 );
nand g862 ( new_n1205_, new_n946_, N246 );
xnor g863 ( new_n1206_, new_n1205_, keyIn_0_123 );
nand g864 ( new_n1207_, new_n635_, N165 );
nand g865 ( new_n1208_, new_n1206_, new_n1207_ );
xnor g866 ( new_n1209_, new_n1208_, keyIn_0_146 );
nand g867 ( new_n1210_, new_n1204_, new_n1209_ );
nor g868 ( new_n1211_, new_n1210_, new_n1203_ );
nand g869 ( new_n1212_, new_n1199_, new_n1211_ );
nand g870 ( new_n1213_, new_n1212_, new_n1153_ );
xnor g871 ( new_n1214_, new_n1198_, keyIn_0_251 );
not g872 ( new_n1215_, new_n1211_ );
nor g873 ( new_n1216_, new_n1214_, new_n1215_ );
nand g874 ( new_n1217_, new_n1216_, keyIn_0_254 );
nand g875 ( N879, new_n1217_, new_n1213_ );
not g876 ( new_n1219_, keyIn_0_252 );
nand g877 ( new_n1220_, new_n965_, new_n1014_ );
xor g878 ( new_n1221_, new_n1220_, keyIn_0_148 );
not g879 ( new_n1222_, new_n1221_ );
nand g880 ( new_n1223_, new_n1009_, keyIn_0_223 );
xnor g881 ( new_n1224_, new_n1021_, keyIn_0_171 );
nor g882 ( new_n1225_, new_n1009_, keyIn_0_223 );
nor g883 ( new_n1226_, new_n1225_, new_n1224_ );
nand g884 ( new_n1227_, new_n1226_, new_n1223_ );
xnor g885 ( new_n1228_, new_n1227_, keyIn_0_228 );
nor g886 ( new_n1229_, new_n1228_, new_n1222_ );
xor g887 ( new_n1230_, new_n1229_, keyIn_0_237 );
nand g888 ( new_n1231_, new_n1228_, new_n1222_ );
xor g889 ( new_n1232_, new_n1231_, keyIn_0_238 );
nand g890 ( new_n1233_, new_n1230_, new_n1232_ );
nand g891 ( new_n1234_, new_n1233_, keyIn_0_246 );
nor g892 ( new_n1235_, new_n1233_, keyIn_0_246 );
nor g893 ( new_n1236_, new_n1235_, new_n604_ );
nand g894 ( new_n1237_, new_n1236_, new_n1234_ );
nand g895 ( new_n1238_, N96, N210 );
nand g896 ( new_n1239_, new_n1237_, new_n1238_ );
nor g897 ( new_n1240_, new_n1239_, new_n1219_ );
nand g898 ( new_n1241_, new_n1239_, new_n1219_ );
nand g899 ( new_n1242_, new_n1015_, N237 );
xnor g900 ( new_n1243_, new_n1242_, keyIn_0_170 );
nand g901 ( new_n1244_, new_n1222_, N228 );
nand g902 ( new_n1245_, new_n1244_, new_n1243_ );
nor g903 ( new_n1246_, new_n1245_, keyIn_0_194 );
nand g904 ( new_n1247_, new_n1245_, keyIn_0_194 );
not g905 ( new_n1248_, keyIn_0_126 );
nand g906 ( new_n1249_, new_n962_, N246 );
nor g907 ( new_n1250_, new_n1249_, new_n1248_ );
nand g908 ( new_n1251_, new_n635_, N171 );
nand g909 ( new_n1252_, new_n1249_, new_n1248_ );
nand g910 ( new_n1253_, new_n1252_, new_n1251_ );
nor g911 ( new_n1254_, new_n1253_, new_n1250_ );
xnor g912 ( new_n1255_, new_n1254_, keyIn_0_149 );
nand g913 ( new_n1256_, new_n1247_, new_n1255_ );
nor g914 ( new_n1257_, new_n1256_, new_n1246_ );
nand g915 ( new_n1258_, new_n1241_, new_n1257_ );
or g916 ( new_n1259_, new_n1258_, new_n1240_ );
nand g917 ( new_n1260_, new_n1259_, keyIn_0_255 );
not g918 ( new_n1261_, keyIn_0_255 );
nor g919 ( new_n1262_, new_n1258_, new_n1240_ );
nand g920 ( new_n1263_, new_n1262_, new_n1261_ );
nand g921 ( N880, new_n1260_, new_n1263_ );
endmodule