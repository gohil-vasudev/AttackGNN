module add_mul_comp_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, 
        a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, 
        a_27_, a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, 
        b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, 
        b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, 
        b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   Result_9_, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_31_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_28_ = Result_9_;
  assign Result_26_ = Result_9_;
  assign Result_24_ = Result_9_;
  assign Result_22_ = Result_9_;
  assign Result_20_ = Result_9_;
  assign Result_19_ = Result_9_;
  assign Result_17_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_16_ = Result_9_;
  assign Result_18_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_21_ = Result_9_;
  assign Result_23_ = Result_9_;
  assign Result_25_ = Result_9_;
  assign Result_27_ = Result_9_;
  assign Result_29_ = Result_9_;
  assign Result_30_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  OR2_X2 U729 ( .A1(n1229), .A2(n1230), .ZN(Result_9_) );
  INV_X1 U730 ( .A(n696), .ZN(Result_63_) );
  AND2_X1 U731 ( .A1(n697), .A2(n698), .ZN(n696) );
  OR2_X1 U732 ( .A1(n699), .A2(n700), .ZN(Result_62_) );
  AND2_X1 U733 ( .A1(n701), .A2(n702), .ZN(n700) );
  OR2_X1 U734 ( .A1(n703), .A2(n704), .ZN(n702) );
  AND2_X1 U735 ( .A1(Result_9_), .A2(n697), .ZN(n704) );
  INV_X1 U736 ( .A(n705), .ZN(n697) );
  INV_X1 U737 ( .A(n706), .ZN(n703) );
  OR2_X1 U738 ( .A1(n707), .A2(n708), .ZN(n706) );
  AND2_X1 U739 ( .A1(a_31_), .A2(b_31_), .ZN(n708) );
  INV_X1 U740 ( .A(n709), .ZN(n701) );
  AND2_X1 U741 ( .A1(n709), .A2(n710), .ZN(n699) );
  OR2_X1 U742 ( .A1(n711), .A2(n712), .ZN(n710) );
  AND2_X1 U743 ( .A1(n705), .A2(Result_9_), .ZN(n712) );
  AND3_X1 U744 ( .A1(b_31_), .A2(a_31_), .A3(n713), .ZN(n711) );
  AND2_X1 U745 ( .A1(n714), .A2(n715), .ZN(n709) );
  INV_X1 U746 ( .A(n716), .ZN(n714) );
  OR2_X1 U747 ( .A1(n717), .A2(n718), .ZN(Result_61_) );
  AND2_X1 U748 ( .A1(n719), .A2(Result_9_), .ZN(n718) );
  OR2_X1 U749 ( .A1(n720), .A2(n721), .ZN(n719) );
  INV_X1 U750 ( .A(n722), .ZN(n721) );
  OR2_X1 U751 ( .A1(n723), .A2(n724), .ZN(n722) );
  AND2_X1 U752 ( .A1(n724), .A2(n723), .ZN(n720) );
  AND2_X1 U753 ( .A1(n713), .A2(n725), .ZN(n717) );
  OR2_X1 U754 ( .A1(n726), .A2(n727), .ZN(n725) );
  INV_X1 U755 ( .A(n728), .ZN(n727) );
  OR2_X1 U756 ( .A1(n729), .A2(n724), .ZN(n728) );
  AND2_X1 U757 ( .A1(n724), .A2(n729), .ZN(n726) );
  AND2_X1 U758 ( .A1(n730), .A2(n731), .ZN(n724) );
  OR2_X1 U759 ( .A1(n732), .A2(b_29_), .ZN(n731) );
  OR2_X1 U760 ( .A1(n733), .A2(n734), .ZN(Result_60_) );
  AND2_X1 U761 ( .A1(n735), .A2(Result_9_), .ZN(n734) );
  OR2_X1 U762 ( .A1(n736), .A2(n737), .ZN(n735) );
  INV_X1 U763 ( .A(n738), .ZN(n737) );
  OR2_X1 U764 ( .A1(n739), .A2(n740), .ZN(n738) );
  AND2_X1 U765 ( .A1(n740), .A2(n739), .ZN(n736) );
  AND3_X1 U766 ( .A1(n741), .A2(n742), .A3(n713), .ZN(n733) );
  INV_X1 U767 ( .A(n743), .ZN(n742) );
  AND2_X1 U768 ( .A1(n744), .A2(n740), .ZN(n743) );
  OR2_X1 U769 ( .A1(n740), .A2(n744), .ZN(n741) );
  AND2_X1 U770 ( .A1(n745), .A2(n746), .ZN(n740) );
  OR2_X1 U771 ( .A1(n747), .A2(b_28_), .ZN(n746) );
  OR2_X1 U772 ( .A1(n748), .A2(n749), .ZN(Result_59_) );
  AND2_X1 U773 ( .A1(n750), .A2(Result_9_), .ZN(n749) );
  OR2_X1 U774 ( .A1(n751), .A2(n752), .ZN(n750) );
  INV_X1 U775 ( .A(n753), .ZN(n752) );
  OR2_X1 U776 ( .A1(n754), .A2(n755), .ZN(n753) );
  AND2_X1 U777 ( .A1(n755), .A2(n754), .ZN(n751) );
  AND3_X1 U778 ( .A1(n756), .A2(n757), .A3(n713), .ZN(n748) );
  INV_X1 U779 ( .A(n758), .ZN(n757) );
  AND2_X1 U780 ( .A1(n759), .A2(n755), .ZN(n758) );
  OR2_X1 U781 ( .A1(n755), .A2(n759), .ZN(n756) );
  AND2_X1 U782 ( .A1(n760), .A2(n761), .ZN(n755) );
  OR2_X1 U783 ( .A1(n762), .A2(b_27_), .ZN(n761) );
  OR2_X1 U784 ( .A1(n763), .A2(n764), .ZN(Result_58_) );
  AND2_X1 U785 ( .A1(n765), .A2(Result_9_), .ZN(n764) );
  OR2_X1 U786 ( .A1(n766), .A2(n767), .ZN(n765) );
  INV_X1 U787 ( .A(n768), .ZN(n767) );
  OR2_X1 U788 ( .A1(n769), .A2(n770), .ZN(n768) );
  AND2_X1 U789 ( .A1(n770), .A2(n769), .ZN(n766) );
  AND3_X1 U790 ( .A1(n771), .A2(n772), .A3(n713), .ZN(n763) );
  INV_X1 U791 ( .A(n773), .ZN(n772) );
  AND2_X1 U792 ( .A1(n774), .A2(n770), .ZN(n773) );
  OR2_X1 U793 ( .A1(n770), .A2(n774), .ZN(n771) );
  AND2_X1 U794 ( .A1(n775), .A2(n776), .ZN(n770) );
  OR2_X1 U795 ( .A1(n777), .A2(b_26_), .ZN(n776) );
  OR2_X1 U796 ( .A1(n778), .A2(n779), .ZN(Result_57_) );
  AND2_X1 U797 ( .A1(n780), .A2(Result_9_), .ZN(n779) );
  OR2_X1 U798 ( .A1(n781), .A2(n782), .ZN(n780) );
  INV_X1 U799 ( .A(n783), .ZN(n782) );
  OR2_X1 U800 ( .A1(n784), .A2(n785), .ZN(n783) );
  AND2_X1 U801 ( .A1(n785), .A2(n784), .ZN(n781) );
  AND3_X1 U802 ( .A1(n786), .A2(n787), .A3(n713), .ZN(n778) );
  INV_X1 U803 ( .A(n788), .ZN(n787) );
  AND2_X1 U804 ( .A1(n789), .A2(n785), .ZN(n788) );
  OR2_X1 U805 ( .A1(n785), .A2(n789), .ZN(n786) );
  AND2_X1 U806 ( .A1(n790), .A2(n791), .ZN(n785) );
  OR2_X1 U807 ( .A1(n792), .A2(b_25_), .ZN(n791) );
  OR2_X1 U808 ( .A1(n793), .A2(n794), .ZN(Result_56_) );
  AND2_X1 U809 ( .A1(n795), .A2(Result_9_), .ZN(n794) );
  OR2_X1 U810 ( .A1(n796), .A2(n797), .ZN(n795) );
  INV_X1 U811 ( .A(n798), .ZN(n797) );
  OR2_X1 U812 ( .A1(n799), .A2(n800), .ZN(n798) );
  AND2_X1 U813 ( .A1(n800), .A2(n799), .ZN(n796) );
  AND3_X1 U814 ( .A1(n801), .A2(n802), .A3(n713), .ZN(n793) );
  INV_X1 U815 ( .A(n803), .ZN(n802) );
  AND2_X1 U816 ( .A1(n804), .A2(n800), .ZN(n803) );
  OR2_X1 U817 ( .A1(n800), .A2(n804), .ZN(n801) );
  AND2_X1 U818 ( .A1(n805), .A2(n806), .ZN(n800) );
  OR2_X1 U819 ( .A1(n807), .A2(b_24_), .ZN(n806) );
  OR2_X1 U820 ( .A1(n808), .A2(n809), .ZN(Result_55_) );
  AND2_X1 U821 ( .A1(n810), .A2(Result_9_), .ZN(n809) );
  OR2_X1 U822 ( .A1(n811), .A2(n812), .ZN(n810) );
  INV_X1 U823 ( .A(n813), .ZN(n812) );
  OR2_X1 U824 ( .A1(n814), .A2(n815), .ZN(n813) );
  AND2_X1 U825 ( .A1(n815), .A2(n814), .ZN(n811) );
  AND3_X1 U826 ( .A1(n816), .A2(n817), .A3(n713), .ZN(n808) );
  INV_X1 U827 ( .A(n818), .ZN(n817) );
  AND2_X1 U828 ( .A1(n819), .A2(n815), .ZN(n818) );
  OR2_X1 U829 ( .A1(n815), .A2(n819), .ZN(n816) );
  AND2_X1 U830 ( .A1(n820), .A2(n821), .ZN(n815) );
  OR2_X1 U831 ( .A1(n822), .A2(b_23_), .ZN(n821) );
  OR2_X1 U832 ( .A1(n823), .A2(n824), .ZN(Result_54_) );
  AND2_X1 U833 ( .A1(n825), .A2(Result_9_), .ZN(n824) );
  OR2_X1 U834 ( .A1(n826), .A2(n827), .ZN(n825) );
  INV_X1 U835 ( .A(n828), .ZN(n827) );
  OR2_X1 U836 ( .A1(n829), .A2(n830), .ZN(n828) );
  AND2_X1 U837 ( .A1(n830), .A2(n829), .ZN(n826) );
  AND3_X1 U838 ( .A1(n831), .A2(n832), .A3(n713), .ZN(n823) );
  INV_X1 U839 ( .A(n833), .ZN(n832) );
  AND2_X1 U840 ( .A1(n834), .A2(n830), .ZN(n833) );
  OR2_X1 U841 ( .A1(n830), .A2(n834), .ZN(n831) );
  AND2_X1 U842 ( .A1(n835), .A2(n836), .ZN(n830) );
  OR2_X1 U843 ( .A1(n837), .A2(b_22_), .ZN(n836) );
  OR2_X1 U844 ( .A1(n838), .A2(n839), .ZN(Result_53_) );
  AND2_X1 U845 ( .A1(n840), .A2(Result_9_), .ZN(n839) );
  OR2_X1 U846 ( .A1(n841), .A2(n842), .ZN(n840) );
  INV_X1 U847 ( .A(n843), .ZN(n842) );
  OR2_X1 U848 ( .A1(n844), .A2(n845), .ZN(n843) );
  AND2_X1 U849 ( .A1(n845), .A2(n844), .ZN(n841) );
  AND3_X1 U850 ( .A1(n846), .A2(n847), .A3(n713), .ZN(n838) );
  INV_X1 U851 ( .A(n848), .ZN(n847) );
  AND2_X1 U852 ( .A1(n849), .A2(n845), .ZN(n848) );
  OR2_X1 U853 ( .A1(n845), .A2(n849), .ZN(n846) );
  AND2_X1 U854 ( .A1(n850), .A2(n851), .ZN(n845) );
  OR2_X1 U855 ( .A1(n852), .A2(b_21_), .ZN(n851) );
  OR2_X1 U856 ( .A1(n853), .A2(n854), .ZN(Result_52_) );
  AND2_X1 U857 ( .A1(n855), .A2(Result_9_), .ZN(n854) );
  OR2_X1 U858 ( .A1(n856), .A2(n857), .ZN(n855) );
  INV_X1 U859 ( .A(n858), .ZN(n857) );
  OR2_X1 U860 ( .A1(n859), .A2(n860), .ZN(n858) );
  AND2_X1 U861 ( .A1(n860), .A2(n859), .ZN(n856) );
  AND3_X1 U862 ( .A1(n861), .A2(n862), .A3(n713), .ZN(n853) );
  INV_X1 U863 ( .A(n863), .ZN(n862) );
  AND2_X1 U864 ( .A1(n864), .A2(n860), .ZN(n863) );
  OR2_X1 U865 ( .A1(n860), .A2(n864), .ZN(n861) );
  AND2_X1 U866 ( .A1(n865), .A2(n866), .ZN(n860) );
  OR2_X1 U867 ( .A1(n867), .A2(b_20_), .ZN(n866) );
  OR2_X1 U868 ( .A1(n868), .A2(n869), .ZN(Result_51_) );
  AND2_X1 U869 ( .A1(n870), .A2(Result_9_), .ZN(n869) );
  OR2_X1 U870 ( .A1(n871), .A2(n872), .ZN(n870) );
  INV_X1 U871 ( .A(n873), .ZN(n872) );
  OR2_X1 U872 ( .A1(n874), .A2(n875), .ZN(n873) );
  AND2_X1 U873 ( .A1(n875), .A2(n874), .ZN(n871) );
  AND3_X1 U874 ( .A1(n876), .A2(n877), .A3(n713), .ZN(n868) );
  INV_X1 U875 ( .A(n878), .ZN(n877) );
  AND2_X1 U876 ( .A1(n879), .A2(n875), .ZN(n878) );
  OR2_X1 U877 ( .A1(n875), .A2(n879), .ZN(n876) );
  AND2_X1 U878 ( .A1(n880), .A2(n881), .ZN(n875) );
  OR2_X1 U879 ( .A1(n882), .A2(b_19_), .ZN(n881) );
  OR2_X1 U880 ( .A1(n883), .A2(n884), .ZN(Result_50_) );
  AND2_X1 U881 ( .A1(n885), .A2(Result_9_), .ZN(n884) );
  OR2_X1 U882 ( .A1(n886), .A2(n887), .ZN(n885) );
  INV_X1 U883 ( .A(n888), .ZN(n887) );
  OR2_X1 U884 ( .A1(n889), .A2(n890), .ZN(n888) );
  AND2_X1 U885 ( .A1(n890), .A2(n889), .ZN(n886) );
  AND3_X1 U886 ( .A1(n891), .A2(n892), .A3(n713), .ZN(n883) );
  INV_X1 U887 ( .A(n893), .ZN(n892) );
  AND2_X1 U888 ( .A1(n894), .A2(n890), .ZN(n893) );
  OR2_X1 U889 ( .A1(n890), .A2(n894), .ZN(n891) );
  AND2_X1 U890 ( .A1(n895), .A2(n896), .ZN(n890) );
  OR2_X1 U891 ( .A1(n897), .A2(b_18_), .ZN(n896) );
  OR2_X1 U892 ( .A1(n898), .A2(n899), .ZN(Result_49_) );
  AND2_X1 U893 ( .A1(n900), .A2(Result_9_), .ZN(n899) );
  OR2_X1 U894 ( .A1(n901), .A2(n902), .ZN(n900) );
  INV_X1 U895 ( .A(n903), .ZN(n902) );
  OR2_X1 U896 ( .A1(n904), .A2(n905), .ZN(n903) );
  AND2_X1 U897 ( .A1(n905), .A2(n904), .ZN(n901) );
  AND3_X1 U898 ( .A1(n906), .A2(n907), .A3(n713), .ZN(n898) );
  INV_X1 U899 ( .A(n908), .ZN(n907) );
  AND2_X1 U900 ( .A1(n909), .A2(n905), .ZN(n908) );
  OR2_X1 U901 ( .A1(n905), .A2(n909), .ZN(n906) );
  AND2_X1 U902 ( .A1(n910), .A2(n911), .ZN(n905) );
  OR2_X1 U903 ( .A1(n912), .A2(b_17_), .ZN(n911) );
  OR2_X1 U904 ( .A1(n913), .A2(n914), .ZN(Result_48_) );
  AND2_X1 U905 ( .A1(n915), .A2(Result_9_), .ZN(n914) );
  OR2_X1 U906 ( .A1(n916), .A2(n917), .ZN(n915) );
  INV_X1 U907 ( .A(n918), .ZN(n917) );
  OR2_X1 U908 ( .A1(n919), .A2(n920), .ZN(n918) );
  AND2_X1 U909 ( .A1(n920), .A2(n919), .ZN(n916) );
  AND3_X1 U910 ( .A1(n921), .A2(n922), .A3(n713), .ZN(n913) );
  INV_X1 U911 ( .A(n923), .ZN(n922) );
  AND2_X1 U912 ( .A1(n924), .A2(n920), .ZN(n923) );
  OR2_X1 U913 ( .A1(n920), .A2(n924), .ZN(n921) );
  AND2_X1 U914 ( .A1(n925), .A2(n926), .ZN(n920) );
  OR2_X1 U915 ( .A1(n927), .A2(b_16_), .ZN(n926) );
  OR2_X1 U916 ( .A1(n928), .A2(n929), .ZN(Result_47_) );
  AND2_X1 U917 ( .A1(n930), .A2(Result_9_), .ZN(n929) );
  OR2_X1 U918 ( .A1(n931), .A2(n932), .ZN(n930) );
  INV_X1 U919 ( .A(n933), .ZN(n932) );
  OR2_X1 U920 ( .A1(n934), .A2(n935), .ZN(n933) );
  AND2_X1 U921 ( .A1(n935), .A2(n934), .ZN(n931) );
  AND3_X1 U922 ( .A1(n936), .A2(n937), .A3(n713), .ZN(n928) );
  INV_X1 U923 ( .A(n938), .ZN(n937) );
  AND2_X1 U924 ( .A1(n939), .A2(n935), .ZN(n938) );
  OR2_X1 U925 ( .A1(n935), .A2(n939), .ZN(n936) );
  AND2_X1 U926 ( .A1(n940), .A2(n941), .ZN(n935) );
  OR2_X1 U927 ( .A1(n942), .A2(b_15_), .ZN(n941) );
  OR2_X1 U928 ( .A1(n943), .A2(n944), .ZN(Result_46_) );
  AND2_X1 U929 ( .A1(n945), .A2(Result_9_), .ZN(n944) );
  OR2_X1 U930 ( .A1(n946), .A2(n947), .ZN(n945) );
  INV_X1 U931 ( .A(n948), .ZN(n947) );
  OR2_X1 U932 ( .A1(n949), .A2(n950), .ZN(n948) );
  AND2_X1 U933 ( .A1(n950), .A2(n949), .ZN(n946) );
  AND3_X1 U934 ( .A1(n951), .A2(n952), .A3(n713), .ZN(n943) );
  INV_X1 U935 ( .A(n953), .ZN(n952) );
  AND2_X1 U936 ( .A1(n954), .A2(n950), .ZN(n953) );
  OR2_X1 U937 ( .A1(n950), .A2(n954), .ZN(n951) );
  AND2_X1 U938 ( .A1(n955), .A2(n956), .ZN(n950) );
  OR2_X1 U939 ( .A1(n957), .A2(b_14_), .ZN(n956) );
  OR2_X1 U940 ( .A1(n958), .A2(n959), .ZN(Result_45_) );
  AND2_X1 U941 ( .A1(n960), .A2(Result_9_), .ZN(n959) );
  OR2_X1 U942 ( .A1(n961), .A2(n962), .ZN(n960) );
  INV_X1 U943 ( .A(n963), .ZN(n962) );
  OR2_X1 U944 ( .A1(n964), .A2(n965), .ZN(n963) );
  AND2_X1 U945 ( .A1(n965), .A2(n964), .ZN(n961) );
  AND3_X1 U946 ( .A1(n966), .A2(n967), .A3(n713), .ZN(n958) );
  INV_X1 U947 ( .A(n968), .ZN(n967) );
  AND2_X1 U948 ( .A1(n969), .A2(n965), .ZN(n968) );
  OR2_X1 U949 ( .A1(n965), .A2(n969), .ZN(n966) );
  AND2_X1 U950 ( .A1(n970), .A2(n971), .ZN(n965) );
  OR2_X1 U951 ( .A1(n972), .A2(b_13_), .ZN(n971) );
  OR2_X1 U952 ( .A1(n973), .A2(n974), .ZN(Result_44_) );
  AND2_X1 U953 ( .A1(n975), .A2(Result_9_), .ZN(n974) );
  OR2_X1 U954 ( .A1(n976), .A2(n977), .ZN(n975) );
  INV_X1 U955 ( .A(n978), .ZN(n977) );
  OR2_X1 U956 ( .A1(n979), .A2(n980), .ZN(n978) );
  AND2_X1 U957 ( .A1(n980), .A2(n979), .ZN(n976) );
  AND3_X1 U958 ( .A1(n981), .A2(n982), .A3(n713), .ZN(n973) );
  INV_X1 U959 ( .A(n983), .ZN(n982) );
  AND2_X1 U960 ( .A1(n984), .A2(n980), .ZN(n983) );
  OR2_X1 U961 ( .A1(n980), .A2(n984), .ZN(n981) );
  AND2_X1 U962 ( .A1(n985), .A2(n986), .ZN(n980) );
  OR2_X1 U963 ( .A1(n987), .A2(b_12_), .ZN(n986) );
  OR2_X1 U964 ( .A1(n988), .A2(n989), .ZN(Result_43_) );
  AND2_X1 U965 ( .A1(n990), .A2(Result_9_), .ZN(n989) );
  OR2_X1 U966 ( .A1(n991), .A2(n992), .ZN(n990) );
  INV_X1 U967 ( .A(n993), .ZN(n992) );
  OR2_X1 U968 ( .A1(n994), .A2(n995), .ZN(n993) );
  AND2_X1 U969 ( .A1(n995), .A2(n994), .ZN(n991) );
  AND3_X1 U970 ( .A1(n996), .A2(n997), .A3(n713), .ZN(n988) );
  INV_X1 U971 ( .A(n998), .ZN(n997) );
  AND2_X1 U972 ( .A1(n999), .A2(n995), .ZN(n998) );
  OR2_X1 U973 ( .A1(n995), .A2(n999), .ZN(n996) );
  AND2_X1 U974 ( .A1(n1000), .A2(n1001), .ZN(n995) );
  OR2_X1 U975 ( .A1(n1002), .A2(b_11_), .ZN(n1001) );
  OR2_X1 U976 ( .A1(n1003), .A2(n1004), .ZN(Result_42_) );
  AND2_X1 U977 ( .A1(n1005), .A2(Result_9_), .ZN(n1004) );
  OR2_X1 U978 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
  INV_X1 U979 ( .A(n1008), .ZN(n1007) );
  OR2_X1 U980 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
  AND2_X1 U981 ( .A1(n1010), .A2(n1009), .ZN(n1006) );
  AND3_X1 U982 ( .A1(n1011), .A2(n1012), .A3(n713), .ZN(n1003) );
  INV_X1 U983 ( .A(n1013), .ZN(n1012) );
  AND2_X1 U984 ( .A1(n1014), .A2(n1010), .ZN(n1013) );
  OR2_X1 U985 ( .A1(n1010), .A2(n1014), .ZN(n1011) );
  AND2_X1 U986 ( .A1(n1015), .A2(n1016), .ZN(n1010) );
  OR2_X1 U987 ( .A1(n1017), .A2(b_10_), .ZN(n1016) );
  OR2_X1 U988 ( .A1(n1018), .A2(n1019), .ZN(Result_41_) );
  AND2_X1 U989 ( .A1(n1020), .A2(Result_9_), .ZN(n1019) );
  OR2_X1 U990 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
  INV_X1 U991 ( .A(n1023), .ZN(n1022) );
  OR2_X1 U992 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
  AND2_X1 U993 ( .A1(n1025), .A2(n1024), .ZN(n1021) );
  AND3_X1 U994 ( .A1(n1026), .A2(n1027), .A3(n713), .ZN(n1018) );
  INV_X1 U995 ( .A(n1028), .ZN(n1027) );
  AND2_X1 U996 ( .A1(n1029), .A2(n1025), .ZN(n1028) );
  OR2_X1 U997 ( .A1(n1025), .A2(n1029), .ZN(n1026) );
  AND2_X1 U998 ( .A1(n1030), .A2(n1031), .ZN(n1025) );
  OR2_X1 U999 ( .A1(n1032), .A2(b_9_), .ZN(n1031) );
  OR2_X1 U1000 ( .A1(n1033), .A2(n1034), .ZN(Result_40_) );
  AND2_X1 U1001 ( .A1(n1035), .A2(Result_9_), .ZN(n1034) );
  OR2_X1 U1002 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
  INV_X1 U1003 ( .A(n1038), .ZN(n1037) );
  OR2_X1 U1004 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
  AND2_X1 U1005 ( .A1(n1040), .A2(n1039), .ZN(n1036) );
  AND3_X1 U1006 ( .A1(n1041), .A2(n1042), .A3(n713), .ZN(n1033) );
  INV_X1 U1007 ( .A(n1043), .ZN(n1042) );
  AND2_X1 U1008 ( .A1(n1044), .A2(n1040), .ZN(n1043) );
  OR2_X1 U1009 ( .A1(n1040), .A2(n1044), .ZN(n1041) );
  AND2_X1 U1010 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
  OR2_X1 U1011 ( .A1(n1047), .A2(b_8_), .ZN(n1046) );
  OR2_X1 U1012 ( .A1(n1048), .A2(n1049), .ZN(Result_39_) );
  AND2_X1 U1013 ( .A1(n1050), .A2(Result_9_), .ZN(n1049) );
  OR2_X1 U1014 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
  INV_X1 U1015 ( .A(n1053), .ZN(n1052) );
  OR2_X1 U1016 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
  AND2_X1 U1017 ( .A1(n1055), .A2(n1054), .ZN(n1051) );
  AND3_X1 U1018 ( .A1(n1056), .A2(n1057), .A3(n713), .ZN(n1048) );
  INV_X1 U1019 ( .A(n1058), .ZN(n1057) );
  AND2_X1 U1020 ( .A1(n1059), .A2(n1055), .ZN(n1058) );
  OR2_X1 U1021 ( .A1(n1055), .A2(n1059), .ZN(n1056) );
  AND2_X1 U1022 ( .A1(n1060), .A2(n1061), .ZN(n1055) );
  OR2_X1 U1023 ( .A1(n1062), .A2(b_7_), .ZN(n1061) );
  OR2_X1 U1024 ( .A1(n1063), .A2(n1064), .ZN(Result_38_) );
  AND2_X1 U1025 ( .A1(n1065), .A2(Result_9_), .ZN(n1064) );
  OR2_X1 U1026 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
  INV_X1 U1027 ( .A(n1068), .ZN(n1067) );
  OR2_X1 U1028 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
  AND2_X1 U1029 ( .A1(n1070), .A2(n1069), .ZN(n1066) );
  AND3_X1 U1030 ( .A1(n1071), .A2(n1072), .A3(n713), .ZN(n1063) );
  INV_X1 U1031 ( .A(n1073), .ZN(n1072) );
  AND2_X1 U1032 ( .A1(n1074), .A2(n1070), .ZN(n1073) );
  OR2_X1 U1033 ( .A1(n1070), .A2(n1074), .ZN(n1071) );
  AND2_X1 U1034 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
  OR2_X1 U1035 ( .A1(n1077), .A2(b_6_), .ZN(n1076) );
  OR2_X1 U1036 ( .A1(n1078), .A2(n1079), .ZN(Result_37_) );
  AND2_X1 U1037 ( .A1(n1080), .A2(Result_9_), .ZN(n1079) );
  OR2_X1 U1038 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
  INV_X1 U1039 ( .A(n1083), .ZN(n1082) );
  OR2_X1 U1040 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
  AND2_X1 U1041 ( .A1(n1085), .A2(n1084), .ZN(n1081) );
  AND3_X1 U1042 ( .A1(n1086), .A2(n1087), .A3(n713), .ZN(n1078) );
  INV_X1 U1043 ( .A(n1088), .ZN(n1087) );
  AND2_X1 U1044 ( .A1(n1089), .A2(n1085), .ZN(n1088) );
  OR2_X1 U1045 ( .A1(n1085), .A2(n1089), .ZN(n1086) );
  AND2_X1 U1046 ( .A1(n1090), .A2(n1091), .ZN(n1085) );
  OR2_X1 U1047 ( .A1(n1092), .A2(b_5_), .ZN(n1091) );
  OR2_X1 U1048 ( .A1(n1093), .A2(n1094), .ZN(Result_36_) );
  AND2_X1 U1049 ( .A1(n1095), .A2(Result_9_), .ZN(n1094) );
  OR2_X1 U1050 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
  INV_X1 U1051 ( .A(n1098), .ZN(n1097) );
  OR2_X1 U1052 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
  AND2_X1 U1053 ( .A1(n1100), .A2(n1099), .ZN(n1096) );
  AND3_X1 U1054 ( .A1(n1101), .A2(n1102), .A3(n713), .ZN(n1093) );
  INV_X1 U1055 ( .A(n1103), .ZN(n1102) );
  AND2_X1 U1056 ( .A1(n1104), .A2(n1100), .ZN(n1103) );
  OR2_X1 U1057 ( .A1(n1100), .A2(n1104), .ZN(n1101) );
  AND2_X1 U1058 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
  OR2_X1 U1059 ( .A1(n1107), .A2(b_4_), .ZN(n1106) );
  OR2_X1 U1060 ( .A1(n1108), .A2(n1109), .ZN(Result_35_) );
  AND2_X1 U1061 ( .A1(n1110), .A2(Result_9_), .ZN(n1109) );
  OR2_X1 U1062 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
  INV_X1 U1063 ( .A(n1113), .ZN(n1112) );
  OR2_X1 U1064 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
  AND2_X1 U1065 ( .A1(n1115), .A2(n1114), .ZN(n1111) );
  AND3_X1 U1066 ( .A1(n1116), .A2(n1117), .A3(n713), .ZN(n1108) );
  INV_X1 U1067 ( .A(n1118), .ZN(n1117) );
  AND2_X1 U1068 ( .A1(n1119), .A2(n1115), .ZN(n1118) );
  OR2_X1 U1069 ( .A1(n1115), .A2(n1119), .ZN(n1116) );
  AND2_X1 U1070 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
  OR2_X1 U1071 ( .A1(n1122), .A2(b_3_), .ZN(n1121) );
  OR2_X1 U1072 ( .A1(n1123), .A2(n1124), .ZN(Result_34_) );
  AND2_X1 U1073 ( .A1(n1125), .A2(Result_9_), .ZN(n1124) );
  OR2_X1 U1074 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
  INV_X1 U1075 ( .A(n1128), .ZN(n1127) );
  OR2_X1 U1076 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
  AND2_X1 U1077 ( .A1(n1130), .A2(n1129), .ZN(n1126) );
  AND3_X1 U1078 ( .A1(n1131), .A2(n1132), .A3(n713), .ZN(n1123) );
  INV_X1 U1079 ( .A(n1133), .ZN(n1132) );
  AND2_X1 U1080 ( .A1(n1134), .A2(n1130), .ZN(n1133) );
  OR2_X1 U1081 ( .A1(n1130), .A2(n1134), .ZN(n1131) );
  AND2_X1 U1082 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
  OR2_X1 U1083 ( .A1(n1137), .A2(b_2_), .ZN(n1136) );
  OR2_X1 U1084 ( .A1(n1138), .A2(n1139), .ZN(Result_33_) );
  AND2_X1 U1085 ( .A1(n1140), .A2(Result_9_), .ZN(n1139) );
  OR2_X1 U1086 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
  INV_X1 U1087 ( .A(n1143), .ZN(n1142) );
  OR2_X1 U1088 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
  AND2_X1 U1089 ( .A1(n1145), .A2(n1144), .ZN(n1141) );
  AND3_X1 U1090 ( .A1(n1146), .A2(n1147), .A3(n713), .ZN(n1138) );
  INV_X1 U1091 ( .A(n1148), .ZN(n1147) );
  AND2_X1 U1092 ( .A1(n1149), .A2(n1145), .ZN(n1148) );
  OR2_X1 U1093 ( .A1(n1145), .A2(n1149), .ZN(n1146) );
  AND2_X1 U1094 ( .A1(n1150), .A2(n1151), .ZN(n1145) );
  INV_X1 U1095 ( .A(n1152), .ZN(n1151) );
  OR2_X1 U1096 ( .A1(n1153), .A2(n1154), .ZN(Result_32_) );
  AND2_X1 U1097 ( .A1(n1155), .A2(Result_9_), .ZN(n1154) );
  OR2_X1 U1098 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
  INV_X1 U1099 ( .A(n1158), .ZN(n1156) );
  OR2_X1 U1100 ( .A1(n1159), .A2(n1152), .ZN(n1158) );
  AND2_X1 U1101 ( .A1(n1144), .A2(n1150), .ZN(n1159) );
  OR2_X1 U1102 ( .A1(n1160), .A2(n1161), .ZN(n1144) );
  AND2_X1 U1103 ( .A1(n1129), .A2(n1135), .ZN(n1160) );
  OR2_X1 U1104 ( .A1(n1162), .A2(n1163), .ZN(n1129) );
  AND2_X1 U1105 ( .A1(n1114), .A2(n1120), .ZN(n1162) );
  OR2_X1 U1106 ( .A1(n1164), .A2(n1165), .ZN(n1114) );
  AND2_X1 U1107 ( .A1(n1099), .A2(n1105), .ZN(n1164) );
  OR2_X1 U1108 ( .A1(n1166), .A2(n1167), .ZN(n1099) );
  AND2_X1 U1109 ( .A1(n1084), .A2(n1090), .ZN(n1166) );
  OR2_X1 U1110 ( .A1(n1168), .A2(n1169), .ZN(n1084) );
  AND2_X1 U1111 ( .A1(n1069), .A2(n1075), .ZN(n1168) );
  OR2_X1 U1112 ( .A1(n1170), .A2(n1171), .ZN(n1069) );
  AND2_X1 U1113 ( .A1(n1054), .A2(n1060), .ZN(n1170) );
  OR2_X1 U1114 ( .A1(n1172), .A2(n1173), .ZN(n1054) );
  AND2_X1 U1115 ( .A1(n1039), .A2(n1045), .ZN(n1172) );
  OR2_X1 U1116 ( .A1(n1174), .A2(n1175), .ZN(n1039) );
  AND2_X1 U1117 ( .A1(n1024), .A2(n1030), .ZN(n1174) );
  OR2_X1 U1118 ( .A1(n1176), .A2(n1177), .ZN(n1024) );
  AND2_X1 U1119 ( .A1(n1009), .A2(n1015), .ZN(n1176) );
  OR2_X1 U1120 ( .A1(n1178), .A2(n1179), .ZN(n1009) );
  AND2_X1 U1121 ( .A1(n994), .A2(n1000), .ZN(n1178) );
  OR2_X1 U1122 ( .A1(n1180), .A2(n1181), .ZN(n994) );
  AND2_X1 U1123 ( .A1(n979), .A2(n985), .ZN(n1180) );
  OR2_X1 U1124 ( .A1(n1182), .A2(n1183), .ZN(n979) );
  AND2_X1 U1125 ( .A1(n964), .A2(n970), .ZN(n1182) );
  OR2_X1 U1126 ( .A1(n1184), .A2(n1185), .ZN(n964) );
  AND2_X1 U1127 ( .A1(n949), .A2(n955), .ZN(n1184) );
  OR2_X1 U1128 ( .A1(n1186), .A2(n1187), .ZN(n949) );
  AND2_X1 U1129 ( .A1(n934), .A2(n940), .ZN(n1186) );
  OR2_X1 U1130 ( .A1(n1188), .A2(n1189), .ZN(n934) );
  AND2_X1 U1131 ( .A1(n919), .A2(n925), .ZN(n1188) );
  OR2_X1 U1132 ( .A1(n1190), .A2(n1191), .ZN(n919) );
  AND2_X1 U1133 ( .A1(n904), .A2(n910), .ZN(n1190) );
  OR2_X1 U1134 ( .A1(n1192), .A2(n1193), .ZN(n904) );
  AND2_X1 U1135 ( .A1(n889), .A2(n895), .ZN(n1192) );
  OR2_X1 U1136 ( .A1(n1194), .A2(n1195), .ZN(n889) );
  AND2_X1 U1137 ( .A1(n874), .A2(n880), .ZN(n1194) );
  OR2_X1 U1138 ( .A1(n1196), .A2(n1197), .ZN(n874) );
  AND2_X1 U1139 ( .A1(n859), .A2(n865), .ZN(n1196) );
  OR2_X1 U1140 ( .A1(n1198), .A2(n1199), .ZN(n859) );
  AND2_X1 U1141 ( .A1(n844), .A2(n850), .ZN(n1198) );
  OR2_X1 U1142 ( .A1(n1200), .A2(n1201), .ZN(n844) );
  AND2_X1 U1143 ( .A1(n829), .A2(n835), .ZN(n1200) );
  OR2_X1 U1144 ( .A1(n1202), .A2(n1203), .ZN(n829) );
  AND2_X1 U1145 ( .A1(n814), .A2(n820), .ZN(n1202) );
  OR2_X1 U1146 ( .A1(n1204), .A2(n1205), .ZN(n814) );
  AND2_X1 U1147 ( .A1(n799), .A2(n805), .ZN(n1204) );
  OR2_X1 U1148 ( .A1(n1206), .A2(n1207), .ZN(n799) );
  AND2_X1 U1149 ( .A1(n784), .A2(n790), .ZN(n1206) );
  OR2_X1 U1150 ( .A1(n1208), .A2(n1209), .ZN(n784) );
  AND2_X1 U1151 ( .A1(n769), .A2(n775), .ZN(n1208) );
  OR2_X1 U1152 ( .A1(n1210), .A2(n1211), .ZN(n769) );
  AND2_X1 U1153 ( .A1(n754), .A2(n760), .ZN(n1210) );
  OR2_X1 U1154 ( .A1(n1212), .A2(n1213), .ZN(n754) );
  AND2_X1 U1155 ( .A1(n739), .A2(n745), .ZN(n1212) );
  AND3_X1 U1156 ( .A1(n1214), .A2(n1215), .A3(n713), .ZN(n1153) );
  INV_X1 U1157 ( .A(n707), .ZN(n713) );
  OR2_X1 U1158 ( .A1(Result_9_), .A2(n1216), .ZN(n707) );
  AND2_X1 U1159 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
  AND4_X1 U1160 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218)
         );
  AND4_X1 U1161 ( .A1(n1120), .A2(n1135), .A3(n1150), .A4(n1223), .ZN(n1222)
         );
  AND4_X1 U1162 ( .A1(n1060), .A2(n1075), .A3(n1090), .A4(n1105), .ZN(n1221)
         );
  AND4_X1 U1163 ( .A1(n1000), .A2(n1015), .A3(n1030), .A4(n1045), .ZN(n1220)
         );
  AND4_X1 U1164 ( .A1(n940), .A2(n955), .A3(n970), .A4(n985), .ZN(n1219) );
  AND4_X1 U1165 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1217)
         );
  AND4_X1 U1166 ( .A1(n880), .A2(n895), .A3(n910), .A4(n925), .ZN(n1227) );
  AND4_X1 U1167 ( .A1(n820), .A2(n835), .A3(n850), .A4(n865), .ZN(n1226) );
  AND4_X1 U1168 ( .A1(n760), .A2(n775), .A3(n790), .A4(n805), .ZN(n1225) );
  AND4_X1 U1169 ( .A1(n698), .A2(n730), .A3(n715), .A4(n745), .ZN(n1224) );
  OR2_X1 U1170 ( .A1(a_31_), .A2(n1228), .ZN(n698) );
  AND2_X1 U1171 ( .A1(n1231), .A2(n1223), .ZN(n1229) );
  OR2_X1 U1172 ( .A1(n1232), .A2(n1152), .ZN(n1231) );
  AND2_X1 U1173 ( .A1(n1233), .A2(a_1_), .ZN(n1152) );
  AND2_X1 U1174 ( .A1(n1234), .A2(n1150), .ZN(n1232) );
  OR2_X1 U1175 ( .A1(a_1_), .A2(n1233), .ZN(n1150) );
  OR2_X1 U1176 ( .A1(n1235), .A2(n1161), .ZN(n1234) );
  AND2_X1 U1177 ( .A1(a_2_), .A2(n1236), .ZN(n1161) );
  AND2_X1 U1178 ( .A1(n1237), .A2(n1135), .ZN(n1235) );
  OR2_X1 U1179 ( .A1(a_2_), .A2(n1236), .ZN(n1135) );
  OR2_X1 U1180 ( .A1(n1238), .A2(n1163), .ZN(n1237) );
  AND2_X1 U1181 ( .A1(a_3_), .A2(n1239), .ZN(n1163) );
  AND3_X1 U1182 ( .A1(n1105), .A2(n1120), .A3(n1240), .ZN(n1238) );
  OR3_X1 U1183 ( .A1(n1241), .A2(n1165), .A3(n1167), .ZN(n1240) );
  AND2_X1 U1184 ( .A1(a_5_), .A2(n1242), .ZN(n1167) );
  AND2_X1 U1185 ( .A1(a_4_), .A2(n1243), .ZN(n1165) );
  AND3_X1 U1186 ( .A1(n1075), .A2(n1090), .A3(n1244), .ZN(n1241) );
  OR3_X1 U1187 ( .A1(n1245), .A2(n1169), .A3(n1171), .ZN(n1244) );
  AND2_X1 U1188 ( .A1(a_7_), .A2(n1246), .ZN(n1171) );
  AND2_X1 U1189 ( .A1(a_6_), .A2(n1247), .ZN(n1169) );
  AND3_X1 U1190 ( .A1(n1045), .A2(n1060), .A3(n1248), .ZN(n1245) );
  OR3_X1 U1191 ( .A1(n1249), .A2(n1173), .A3(n1175), .ZN(n1248) );
  AND2_X1 U1192 ( .A1(a_9_), .A2(n1250), .ZN(n1175) );
  AND2_X1 U1193 ( .A1(a_8_), .A2(n1251), .ZN(n1173) );
  AND3_X1 U1194 ( .A1(n1015), .A2(n1030), .A3(n1252), .ZN(n1249) );
  OR3_X1 U1195 ( .A1(n1253), .A2(n1177), .A3(n1179), .ZN(n1252) );
  AND2_X1 U1196 ( .A1(a_11_), .A2(n1254), .ZN(n1179) );
  AND2_X1 U1197 ( .A1(a_10_), .A2(n1255), .ZN(n1177) );
  AND3_X1 U1198 ( .A1(n985), .A2(n1000), .A3(n1256), .ZN(n1253) );
  OR3_X1 U1199 ( .A1(n1257), .A2(n1181), .A3(n1183), .ZN(n1256) );
  AND2_X1 U1200 ( .A1(a_13_), .A2(n1258), .ZN(n1183) );
  AND2_X1 U1201 ( .A1(a_12_), .A2(n1259), .ZN(n1181) );
  AND3_X1 U1202 ( .A1(n955), .A2(n970), .A3(n1260), .ZN(n1257) );
  OR3_X1 U1203 ( .A1(n1261), .A2(n1185), .A3(n1187), .ZN(n1260) );
  AND2_X1 U1204 ( .A1(a_15_), .A2(n1262), .ZN(n1187) );
  AND2_X1 U1205 ( .A1(a_14_), .A2(n1263), .ZN(n1185) );
  AND3_X1 U1206 ( .A1(n925), .A2(n940), .A3(n1264), .ZN(n1261) );
  OR3_X1 U1207 ( .A1(n1265), .A2(n1189), .A3(n1191), .ZN(n1264) );
  AND2_X1 U1208 ( .A1(a_17_), .A2(n1266), .ZN(n1191) );
  AND2_X1 U1209 ( .A1(a_16_), .A2(n1267), .ZN(n1189) );
  AND3_X1 U1210 ( .A1(n895), .A2(n910), .A3(n1268), .ZN(n1265) );
  OR3_X1 U1211 ( .A1(n1269), .A2(n1193), .A3(n1195), .ZN(n1268) );
  AND2_X1 U1212 ( .A1(a_19_), .A2(n1270), .ZN(n1195) );
  AND2_X1 U1213 ( .A1(a_18_), .A2(n1271), .ZN(n1193) );
  AND3_X1 U1214 ( .A1(n865), .A2(n880), .A3(n1272), .ZN(n1269) );
  OR3_X1 U1215 ( .A1(n1273), .A2(n1197), .A3(n1199), .ZN(n1272) );
  AND2_X1 U1216 ( .A1(a_21_), .A2(n1274), .ZN(n1199) );
  AND2_X1 U1217 ( .A1(a_20_), .A2(n1275), .ZN(n1197) );
  AND3_X1 U1218 ( .A1(n835), .A2(n850), .A3(n1276), .ZN(n1273) );
  OR3_X1 U1219 ( .A1(n1277), .A2(n1201), .A3(n1203), .ZN(n1276) );
  AND2_X1 U1220 ( .A1(a_23_), .A2(n1278), .ZN(n1203) );
  AND2_X1 U1221 ( .A1(a_22_), .A2(n1279), .ZN(n1201) );
  AND3_X1 U1222 ( .A1(n805), .A2(n820), .A3(n1280), .ZN(n1277) );
  OR3_X1 U1223 ( .A1(n1281), .A2(n1205), .A3(n1207), .ZN(n1280) );
  AND2_X1 U1224 ( .A1(a_25_), .A2(n1282), .ZN(n1207) );
  AND2_X1 U1225 ( .A1(a_24_), .A2(n1283), .ZN(n1205) );
  AND3_X1 U1226 ( .A1(n775), .A2(n790), .A3(n1284), .ZN(n1281) );
  OR3_X1 U1227 ( .A1(n1285), .A2(n1209), .A3(n1211), .ZN(n1284) );
  AND2_X1 U1228 ( .A1(a_27_), .A2(n1286), .ZN(n1211) );
  AND2_X1 U1229 ( .A1(a_26_), .A2(n1287), .ZN(n1209) );
  AND3_X1 U1230 ( .A1(n745), .A2(n760), .A3(n1288), .ZN(n1285) );
  OR2_X1 U1231 ( .A1(n1213), .A2(n739), .ZN(n1288) );
  OR2_X1 U1232 ( .A1(n1289), .A2(n1290), .ZN(n739) );
  AND2_X1 U1233 ( .A1(a_29_), .A2(n1291), .ZN(n1290) );
  AND2_X1 U1234 ( .A1(n730), .A2(n723), .ZN(n1289) );
  OR2_X1 U1235 ( .A1(n1292), .A2(n716), .ZN(n723) );
  AND2_X1 U1236 ( .A1(n1293), .A2(a_30_), .ZN(n716) );
  AND2_X1 U1237 ( .A1(n705), .A2(n715), .ZN(n1292) );
  OR2_X1 U1238 ( .A1(a_30_), .A2(n1293), .ZN(n715) );
  INV_X1 U1239 ( .A(b_30_), .ZN(n1293) );
  AND2_X1 U1240 ( .A1(n1228), .A2(a_31_), .ZN(n705) );
  INV_X1 U1241 ( .A(b_31_), .ZN(n1228) );
  OR2_X1 U1242 ( .A1(a_29_), .A2(n1291), .ZN(n730) );
  AND2_X1 U1243 ( .A1(a_28_), .A2(n1294), .ZN(n1213) );
  OR2_X1 U1244 ( .A1(a_27_), .A2(n1286), .ZN(n760) );
  OR2_X1 U1245 ( .A1(a_28_), .A2(n1294), .ZN(n745) );
  OR2_X1 U1246 ( .A1(a_25_), .A2(n1282), .ZN(n790) );
  OR2_X1 U1247 ( .A1(a_26_), .A2(n1287), .ZN(n775) );
  OR2_X1 U1248 ( .A1(a_23_), .A2(n1278), .ZN(n820) );
  OR2_X1 U1249 ( .A1(a_24_), .A2(n1283), .ZN(n805) );
  OR2_X1 U1250 ( .A1(a_21_), .A2(n1274), .ZN(n850) );
  OR2_X1 U1251 ( .A1(a_22_), .A2(n1279), .ZN(n835) );
  OR2_X1 U1252 ( .A1(a_19_), .A2(n1270), .ZN(n880) );
  OR2_X1 U1253 ( .A1(a_20_), .A2(n1275), .ZN(n865) );
  OR2_X1 U1254 ( .A1(a_17_), .A2(n1266), .ZN(n910) );
  OR2_X1 U1255 ( .A1(a_18_), .A2(n1271), .ZN(n895) );
  OR2_X1 U1256 ( .A1(a_15_), .A2(n1262), .ZN(n940) );
  OR2_X1 U1257 ( .A1(a_16_), .A2(n1267), .ZN(n925) );
  OR2_X1 U1258 ( .A1(a_13_), .A2(n1258), .ZN(n970) );
  OR2_X1 U1259 ( .A1(a_14_), .A2(n1263), .ZN(n955) );
  OR2_X1 U1260 ( .A1(a_11_), .A2(n1254), .ZN(n1000) );
  OR2_X1 U1261 ( .A1(a_12_), .A2(n1259), .ZN(n985) );
  OR2_X1 U1262 ( .A1(a_9_), .A2(n1250), .ZN(n1030) );
  OR2_X1 U1263 ( .A1(a_10_), .A2(n1255), .ZN(n1015) );
  OR2_X1 U1264 ( .A1(a_7_), .A2(n1246), .ZN(n1060) );
  OR2_X1 U1265 ( .A1(a_8_), .A2(n1251), .ZN(n1045) );
  OR2_X1 U1266 ( .A1(a_5_), .A2(n1242), .ZN(n1090) );
  OR2_X1 U1267 ( .A1(a_6_), .A2(n1247), .ZN(n1075) );
  OR2_X1 U1268 ( .A1(a_3_), .A2(n1239), .ZN(n1120) );
  OR2_X1 U1269 ( .A1(a_4_), .A2(n1243), .ZN(n1105) );
  INV_X1 U1270 ( .A(n1295), .ZN(n1215) );
  AND2_X1 U1271 ( .A1(n1296), .A2(n1157), .ZN(n1295) );
  OR2_X1 U1272 ( .A1(n1157), .A2(n1296), .ZN(n1214) );
  OR2_X1 U1273 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
  AND2_X1 U1274 ( .A1(n1149), .A2(n1299), .ZN(n1298) );
  AND2_X1 U1275 ( .A1(n1300), .A2(n1233), .ZN(n1297) );
  INV_X1 U1276 ( .A(b_1_), .ZN(n1233) );
  OR2_X1 U1277 ( .A1(n1299), .A2(n1149), .ZN(n1300) );
  OR2_X1 U1278 ( .A1(n1301), .A2(n1302), .ZN(n1149) );
  AND2_X1 U1279 ( .A1(n1134), .A2(n1137), .ZN(n1302) );
  AND2_X1 U1280 ( .A1(n1303), .A2(n1236), .ZN(n1301) );
  INV_X1 U1281 ( .A(b_2_), .ZN(n1236) );
  OR2_X1 U1282 ( .A1(n1137), .A2(n1134), .ZN(n1303) );
  OR2_X1 U1283 ( .A1(n1304), .A2(n1305), .ZN(n1134) );
  AND2_X1 U1284 ( .A1(n1119), .A2(n1122), .ZN(n1305) );
  AND2_X1 U1285 ( .A1(n1306), .A2(n1239), .ZN(n1304) );
  INV_X1 U1286 ( .A(b_3_), .ZN(n1239) );
  OR2_X1 U1287 ( .A1(n1122), .A2(n1119), .ZN(n1306) );
  OR2_X1 U1288 ( .A1(n1307), .A2(n1308), .ZN(n1119) );
  AND2_X1 U1289 ( .A1(n1104), .A2(n1107), .ZN(n1308) );
  AND2_X1 U1290 ( .A1(n1309), .A2(n1243), .ZN(n1307) );
  INV_X1 U1291 ( .A(b_4_), .ZN(n1243) );
  OR2_X1 U1292 ( .A1(n1107), .A2(n1104), .ZN(n1309) );
  OR2_X1 U1293 ( .A1(n1310), .A2(n1311), .ZN(n1104) );
  AND2_X1 U1294 ( .A1(n1089), .A2(n1092), .ZN(n1311) );
  AND2_X1 U1295 ( .A1(n1312), .A2(n1242), .ZN(n1310) );
  INV_X1 U1296 ( .A(b_5_), .ZN(n1242) );
  OR2_X1 U1297 ( .A1(n1092), .A2(n1089), .ZN(n1312) );
  OR2_X1 U1298 ( .A1(n1313), .A2(n1314), .ZN(n1089) );
  AND2_X1 U1299 ( .A1(n1074), .A2(n1077), .ZN(n1314) );
  AND2_X1 U1300 ( .A1(n1315), .A2(n1247), .ZN(n1313) );
  INV_X1 U1301 ( .A(b_6_), .ZN(n1247) );
  OR2_X1 U1302 ( .A1(n1077), .A2(n1074), .ZN(n1315) );
  OR2_X1 U1303 ( .A1(n1316), .A2(n1317), .ZN(n1074) );
  AND2_X1 U1304 ( .A1(n1059), .A2(n1062), .ZN(n1317) );
  AND2_X1 U1305 ( .A1(n1318), .A2(n1246), .ZN(n1316) );
  INV_X1 U1306 ( .A(b_7_), .ZN(n1246) );
  OR2_X1 U1307 ( .A1(n1062), .A2(n1059), .ZN(n1318) );
  OR2_X1 U1308 ( .A1(n1319), .A2(n1320), .ZN(n1059) );
  AND2_X1 U1309 ( .A1(n1044), .A2(n1047), .ZN(n1320) );
  AND2_X1 U1310 ( .A1(n1321), .A2(n1251), .ZN(n1319) );
  INV_X1 U1311 ( .A(b_8_), .ZN(n1251) );
  OR2_X1 U1312 ( .A1(n1047), .A2(n1044), .ZN(n1321) );
  OR2_X1 U1313 ( .A1(n1322), .A2(n1323), .ZN(n1044) );
  AND2_X1 U1314 ( .A1(n1029), .A2(n1032), .ZN(n1323) );
  AND2_X1 U1315 ( .A1(n1324), .A2(n1250), .ZN(n1322) );
  INV_X1 U1316 ( .A(b_9_), .ZN(n1250) );
  OR2_X1 U1317 ( .A1(n1032), .A2(n1029), .ZN(n1324) );
  OR2_X1 U1318 ( .A1(n1325), .A2(n1326), .ZN(n1029) );
  AND2_X1 U1319 ( .A1(n1014), .A2(n1017), .ZN(n1326) );
  AND2_X1 U1320 ( .A1(n1327), .A2(n1255), .ZN(n1325) );
  INV_X1 U1321 ( .A(b_10_), .ZN(n1255) );
  OR2_X1 U1322 ( .A1(n1017), .A2(n1014), .ZN(n1327) );
  OR2_X1 U1323 ( .A1(n1328), .A2(n1329), .ZN(n1014) );
  AND2_X1 U1324 ( .A1(n999), .A2(n1002), .ZN(n1329) );
  AND2_X1 U1325 ( .A1(n1330), .A2(n1254), .ZN(n1328) );
  INV_X1 U1326 ( .A(b_11_), .ZN(n1254) );
  OR2_X1 U1327 ( .A1(n1002), .A2(n999), .ZN(n1330) );
  OR2_X1 U1328 ( .A1(n1331), .A2(n1332), .ZN(n999) );
  AND2_X1 U1329 ( .A1(n984), .A2(n987), .ZN(n1332) );
  AND2_X1 U1330 ( .A1(n1333), .A2(n1259), .ZN(n1331) );
  INV_X1 U1331 ( .A(b_12_), .ZN(n1259) );
  OR2_X1 U1332 ( .A1(n987), .A2(n984), .ZN(n1333) );
  OR2_X1 U1333 ( .A1(n1334), .A2(n1335), .ZN(n984) );
  AND2_X1 U1334 ( .A1(n969), .A2(n972), .ZN(n1335) );
  AND2_X1 U1335 ( .A1(n1336), .A2(n1258), .ZN(n1334) );
  INV_X1 U1336 ( .A(b_13_), .ZN(n1258) );
  OR2_X1 U1337 ( .A1(n972), .A2(n969), .ZN(n1336) );
  OR2_X1 U1338 ( .A1(n1337), .A2(n1338), .ZN(n969) );
  AND2_X1 U1339 ( .A1(n954), .A2(n957), .ZN(n1338) );
  AND2_X1 U1340 ( .A1(n1339), .A2(n1263), .ZN(n1337) );
  INV_X1 U1341 ( .A(b_14_), .ZN(n1263) );
  OR2_X1 U1342 ( .A1(n957), .A2(n954), .ZN(n1339) );
  OR2_X1 U1343 ( .A1(n1340), .A2(n1341), .ZN(n954) );
  AND2_X1 U1344 ( .A1(n939), .A2(n942), .ZN(n1341) );
  AND2_X1 U1345 ( .A1(n1342), .A2(n1262), .ZN(n1340) );
  INV_X1 U1346 ( .A(b_15_), .ZN(n1262) );
  OR2_X1 U1347 ( .A1(n942), .A2(n939), .ZN(n1342) );
  OR2_X1 U1348 ( .A1(n1343), .A2(n1344), .ZN(n939) );
  AND2_X1 U1349 ( .A1(n924), .A2(n927), .ZN(n1344) );
  AND2_X1 U1350 ( .A1(n1345), .A2(n1267), .ZN(n1343) );
  INV_X1 U1351 ( .A(b_16_), .ZN(n1267) );
  OR2_X1 U1352 ( .A1(n927), .A2(n924), .ZN(n1345) );
  OR2_X1 U1353 ( .A1(n1346), .A2(n1347), .ZN(n924) );
  AND2_X1 U1354 ( .A1(n909), .A2(n912), .ZN(n1347) );
  AND2_X1 U1355 ( .A1(n1348), .A2(n1266), .ZN(n1346) );
  INV_X1 U1356 ( .A(b_17_), .ZN(n1266) );
  OR2_X1 U1357 ( .A1(n912), .A2(n909), .ZN(n1348) );
  OR2_X1 U1358 ( .A1(n1349), .A2(n1350), .ZN(n909) );
  AND2_X1 U1359 ( .A1(n894), .A2(n897), .ZN(n1350) );
  AND2_X1 U1360 ( .A1(n1351), .A2(n1271), .ZN(n1349) );
  INV_X1 U1361 ( .A(b_18_), .ZN(n1271) );
  OR2_X1 U1362 ( .A1(n897), .A2(n894), .ZN(n1351) );
  OR2_X1 U1363 ( .A1(n1352), .A2(n1353), .ZN(n894) );
  AND2_X1 U1364 ( .A1(n879), .A2(n882), .ZN(n1353) );
  AND2_X1 U1365 ( .A1(n1354), .A2(n1270), .ZN(n1352) );
  INV_X1 U1366 ( .A(b_19_), .ZN(n1270) );
  OR2_X1 U1367 ( .A1(n882), .A2(n879), .ZN(n1354) );
  OR2_X1 U1368 ( .A1(n1355), .A2(n1356), .ZN(n879) );
  AND2_X1 U1369 ( .A1(n864), .A2(n867), .ZN(n1356) );
  AND2_X1 U1370 ( .A1(n1357), .A2(n1275), .ZN(n1355) );
  INV_X1 U1371 ( .A(b_20_), .ZN(n1275) );
  OR2_X1 U1372 ( .A1(n867), .A2(n864), .ZN(n1357) );
  OR2_X1 U1373 ( .A1(n1358), .A2(n1359), .ZN(n864) );
  AND2_X1 U1374 ( .A1(n849), .A2(n852), .ZN(n1359) );
  AND2_X1 U1375 ( .A1(n1360), .A2(n1274), .ZN(n1358) );
  INV_X1 U1376 ( .A(b_21_), .ZN(n1274) );
  OR2_X1 U1377 ( .A1(n852), .A2(n849), .ZN(n1360) );
  OR2_X1 U1378 ( .A1(n1361), .A2(n1362), .ZN(n849) );
  AND2_X1 U1379 ( .A1(n834), .A2(n837), .ZN(n1362) );
  AND2_X1 U1380 ( .A1(n1363), .A2(n1279), .ZN(n1361) );
  INV_X1 U1381 ( .A(b_22_), .ZN(n1279) );
  OR2_X1 U1382 ( .A1(n837), .A2(n834), .ZN(n1363) );
  OR2_X1 U1383 ( .A1(n1364), .A2(n1365), .ZN(n834) );
  AND2_X1 U1384 ( .A1(n819), .A2(n822), .ZN(n1365) );
  AND2_X1 U1385 ( .A1(n1366), .A2(n1278), .ZN(n1364) );
  INV_X1 U1386 ( .A(b_23_), .ZN(n1278) );
  OR2_X1 U1387 ( .A1(n822), .A2(n819), .ZN(n1366) );
  OR2_X1 U1388 ( .A1(n1367), .A2(n1368), .ZN(n819) );
  AND2_X1 U1389 ( .A1(n804), .A2(n807), .ZN(n1368) );
  AND2_X1 U1390 ( .A1(n1369), .A2(n1283), .ZN(n1367) );
  INV_X1 U1391 ( .A(b_24_), .ZN(n1283) );
  OR2_X1 U1392 ( .A1(n807), .A2(n804), .ZN(n1369) );
  OR2_X1 U1393 ( .A1(n1370), .A2(n1371), .ZN(n804) );
  AND2_X1 U1394 ( .A1(n789), .A2(n792), .ZN(n1371) );
  AND2_X1 U1395 ( .A1(n1372), .A2(n1282), .ZN(n1370) );
  INV_X1 U1396 ( .A(b_25_), .ZN(n1282) );
  OR2_X1 U1397 ( .A1(n792), .A2(n789), .ZN(n1372) );
  OR2_X1 U1398 ( .A1(n1373), .A2(n1374), .ZN(n789) );
  AND2_X1 U1399 ( .A1(n774), .A2(n777), .ZN(n1374) );
  AND2_X1 U1400 ( .A1(n1375), .A2(n1287), .ZN(n1373) );
  INV_X1 U1401 ( .A(b_26_), .ZN(n1287) );
  OR2_X1 U1402 ( .A1(n777), .A2(n774), .ZN(n1375) );
  OR2_X1 U1403 ( .A1(n1376), .A2(n1377), .ZN(n774) );
  AND2_X1 U1404 ( .A1(n759), .A2(n762), .ZN(n1377) );
  AND2_X1 U1405 ( .A1(n1378), .A2(n1286), .ZN(n1376) );
  INV_X1 U1406 ( .A(b_27_), .ZN(n1286) );
  OR2_X1 U1407 ( .A1(n762), .A2(n759), .ZN(n1378) );
  OR2_X1 U1408 ( .A1(n1379), .A2(n1380), .ZN(n759) );
  AND2_X1 U1409 ( .A1(n744), .A2(n747), .ZN(n1380) );
  AND2_X1 U1410 ( .A1(n1381), .A2(n1294), .ZN(n1379) );
  INV_X1 U1411 ( .A(b_28_), .ZN(n1294) );
  OR2_X1 U1412 ( .A1(n747), .A2(n744), .ZN(n1381) );
  OR2_X1 U1413 ( .A1(n1382), .A2(n1383), .ZN(n744) );
  AND2_X1 U1414 ( .A1(n1384), .A2(n732), .ZN(n1383) );
  AND2_X1 U1415 ( .A1(n1385), .A2(n1291), .ZN(n1382) );
  INV_X1 U1416 ( .A(b_29_), .ZN(n1291) );
  OR2_X1 U1417 ( .A1(n1384), .A2(n732), .ZN(n1385) );
  INV_X1 U1418 ( .A(a_29_), .ZN(n732) );
  INV_X1 U1419 ( .A(n729), .ZN(n1384) );
  OR2_X1 U1420 ( .A1(n1386), .A2(n1387), .ZN(n729) );
  AND2_X1 U1421 ( .A1(a_30_), .A2(b_30_), .ZN(n1387) );
  AND3_X1 U1422 ( .A1(a_31_), .A2(n1388), .A3(b_31_), .ZN(n1386) );
  OR2_X1 U1423 ( .A1(a_30_), .A2(b_30_), .ZN(n1388) );
  INV_X1 U1424 ( .A(a_28_), .ZN(n747) );
  INV_X1 U1425 ( .A(a_27_), .ZN(n762) );
  INV_X1 U1426 ( .A(a_26_), .ZN(n777) );
  INV_X1 U1427 ( .A(a_25_), .ZN(n792) );
  INV_X1 U1428 ( .A(a_24_), .ZN(n807) );
  INV_X1 U1429 ( .A(a_23_), .ZN(n822) );
  INV_X1 U1430 ( .A(a_22_), .ZN(n837) );
  INV_X1 U1431 ( .A(a_21_), .ZN(n852) );
  INV_X1 U1432 ( .A(a_20_), .ZN(n867) );
  INV_X1 U1433 ( .A(a_19_), .ZN(n882) );
  INV_X1 U1434 ( .A(a_18_), .ZN(n897) );
  INV_X1 U1435 ( .A(a_17_), .ZN(n912) );
  INV_X1 U1436 ( .A(a_16_), .ZN(n927) );
  INV_X1 U1437 ( .A(a_15_), .ZN(n942) );
  INV_X1 U1438 ( .A(a_14_), .ZN(n957) );
  INV_X1 U1439 ( .A(a_13_), .ZN(n972) );
  INV_X1 U1440 ( .A(a_12_), .ZN(n987) );
  INV_X1 U1441 ( .A(a_11_), .ZN(n1002) );
  INV_X1 U1442 ( .A(a_10_), .ZN(n1017) );
  INV_X1 U1443 ( .A(a_9_), .ZN(n1032) );
  INV_X1 U1444 ( .A(a_8_), .ZN(n1047) );
  INV_X1 U1445 ( .A(a_7_), .ZN(n1062) );
  INV_X1 U1446 ( .A(a_6_), .ZN(n1077) );
  INV_X1 U1447 ( .A(a_5_), .ZN(n1092) );
  INV_X1 U1448 ( .A(a_4_), .ZN(n1107) );
  INV_X1 U1449 ( .A(a_3_), .ZN(n1122) );
  INV_X1 U1450 ( .A(a_2_), .ZN(n1137) );
  INV_X1 U1451 ( .A(a_1_), .ZN(n1299) );
  AND2_X1 U1452 ( .A1(n1223), .A2(n1389), .ZN(n1157) );
  INV_X1 U1453 ( .A(n1230), .ZN(n1389) );
  AND2_X1 U1454 ( .A1(a_0_), .A2(n1390), .ZN(n1230) );
  OR2_X1 U1455 ( .A1(a_0_), .A2(n1390), .ZN(n1223) );
  INV_X1 U1456 ( .A(b_0_), .ZN(n1390) );
endmodule

