module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n220_, new_n624_, new_n534_, new_n214_, new_n451_, new_n424_, new_n602_, new_n240_, new_n413_, new_n526_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n257_, new_n212_, new_n364_, new_n449_, new_n580_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n326_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n385_, new_n478_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n498_, new_n205_, new_n492_, new_n496_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n483_, new_n394_, new_n299_, new_n314_, new_n363_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n438_, new_n208_, new_n632_, new_n528_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n295_, new_n359_, new_n628_, new_n409_, new_n457_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n570_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n407_, new_n480_, new_n625_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n522_, new_n588_, new_n428_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n417_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n440_, new_n531_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n217_, new_n269_, new_n512_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n490_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n226_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n204_, new_n573_, new_n405_;

xor g000 ( new_n202_, N33, N49 );
xnor g001 ( new_n203_, new_n202_, keyIn_0_16 );
xor g002 ( new_n204_, N1, N17 );
xnor g003 ( new_n205_, new_n203_, new_n204_ );
and g004 ( new_n206_, N129, N137 );
xor g005 ( new_n207_, new_n206_, keyIn_0_9 );
xor g006 ( new_n208_, N73, N77 );
xnor g007 ( new_n209_, N65, N69 );
xnor g008 ( new_n210_, new_n208_, new_n209_ );
not g009 ( new_n211_, new_n210_ );
not g010 ( new_n212_, keyIn_0_6 );
xnor g011 ( new_n213_, N89, N93 );
xnor g012 ( new_n214_, new_n213_, new_n212_ );
xnor g013 ( new_n215_, N81, N85 );
xnor g014 ( new_n216_, new_n215_, keyIn_0_5 );
xnor g015 ( new_n217_, new_n214_, new_n216_ );
xnor g016 ( new_n218_, new_n217_, keyIn_0_28 );
xnor g017 ( new_n219_, new_n218_, new_n211_ );
xnor g018 ( new_n220_, new_n219_, keyIn_0_34 );
xnor g019 ( new_n221_, new_n220_, new_n207_ );
xnor g020 ( new_n222_, new_n221_, keyIn_0_36 );
xnor g021 ( new_n223_, new_n222_, new_n205_ );
xor g022 ( new_n224_, new_n223_, keyIn_0_40 );
not g023 ( new_n225_, keyIn_0_78 );
xnor g024 ( new_n226_, new_n224_, keyIn_0_49 );
xnor g025 ( new_n227_, N105, N109 );
xnor g026 ( new_n228_, new_n227_, keyIn_0_7 );
xnor g027 ( new_n229_, N97, N101 );
xnor g028 ( new_n230_, new_n228_, new_n229_ );
xnor g029 ( new_n231_, new_n230_, new_n210_ );
and g030 ( new_n232_, N131, N137 );
xnor g031 ( new_n233_, new_n232_, keyIn_0_11 );
xnor g032 ( new_n234_, new_n231_, new_n233_ );
xor g033 ( new_n235_, N41, N57 );
xnor g034 ( new_n236_, new_n235_, keyIn_0_19 );
xor g035 ( new_n237_, N9, N25 );
xnor g036 ( new_n238_, new_n236_, new_n237_ );
xnor g037 ( new_n239_, new_n238_, keyIn_0_29 );
xor g038 ( new_n240_, new_n234_, new_n239_ );
not g039 ( new_n241_, keyIn_0_41 );
xor g040 ( new_n242_, N13, N29 );
xnor g041 ( new_n243_, new_n242_, keyIn_0_20 );
xor g042 ( new_n244_, N45, N61 );
xnor g043 ( new_n245_, new_n243_, new_n244_ );
xor g044 ( new_n246_, new_n245_, keyIn_0_30 );
not g045 ( new_n247_, keyIn_0_37 );
and g046 ( new_n248_, N132, N137 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_12 );
xnor g048 ( new_n250_, N121, N125 );
xnor g049 ( new_n251_, new_n250_, keyIn_0_8 );
xnor g050 ( new_n252_, N113, N117 );
xnor g051 ( new_n253_, new_n251_, new_n252_ );
xnor g052 ( new_n254_, new_n218_, new_n253_ );
xnor g053 ( new_n255_, new_n254_, new_n249_ );
xnor g054 ( new_n256_, new_n255_, new_n247_ );
xnor g055 ( new_n257_, new_n256_, new_n246_ );
or g056 ( new_n258_, new_n257_, new_n241_ );
not g057 ( new_n259_, new_n256_ );
and g058 ( new_n260_, new_n259_, new_n246_ );
not g059 ( new_n261_, new_n246_ );
and g060 ( new_n262_, new_n256_, new_n261_ );
or g061 ( new_n263_, new_n262_, keyIn_0_41 );
or g062 ( new_n264_, new_n263_, new_n260_ );
and g063 ( new_n265_, new_n264_, new_n258_ );
and g064 ( new_n266_, new_n265_, new_n240_ );
xnor g065 ( new_n267_, new_n230_, new_n253_ );
xnor g066 ( new_n268_, new_n267_, keyIn_0_35 );
and g067 ( new_n269_, N130, N137 );
xor g068 ( new_n270_, new_n269_, keyIn_0_10 );
xnor g069 ( new_n271_, new_n268_, new_n270_ );
xor g070 ( new_n272_, N37, N53 );
xnor g071 ( new_n273_, new_n272_, keyIn_0_18 );
xor g072 ( new_n274_, N5, N21 );
xnor g073 ( new_n275_, new_n274_, keyIn_0_17 );
xnor g074 ( new_n276_, new_n273_, new_n275_ );
xor g075 ( new_n277_, new_n271_, new_n276_ );
xor g076 ( new_n278_, new_n277_, keyIn_0_50 );
and g077 ( new_n279_, new_n266_, new_n278_ );
and g078 ( new_n280_, new_n226_, new_n279_ );
xnor g079 ( new_n281_, new_n280_, keyIn_0_73 );
xnor g080 ( new_n282_, new_n224_, keyIn_0_46 );
not g081 ( new_n283_, new_n265_ );
xor g082 ( new_n284_, new_n277_, keyIn_0_47 );
xor g083 ( new_n285_, new_n240_, keyIn_0_48 );
and g084 ( new_n286_, new_n284_, new_n285_ );
and g085 ( new_n287_, new_n283_, new_n286_ );
and g086 ( new_n288_, new_n282_, new_n287_ );
xnor g087 ( new_n289_, new_n288_, keyIn_0_72 );
not g088 ( new_n290_, new_n224_ );
not g089 ( new_n291_, keyIn_0_52 );
xnor g090 ( new_n292_, new_n257_, new_n241_ );
and g091 ( new_n293_, new_n292_, new_n291_ );
xnor g092 ( new_n294_, new_n257_, keyIn_0_41 );
and g093 ( new_n295_, new_n294_, keyIn_0_52 );
xor g094 ( new_n296_, new_n240_, keyIn_0_51 );
and g095 ( new_n297_, new_n296_, new_n277_ );
not g096 ( new_n298_, new_n297_ );
or g097 ( new_n299_, new_n295_, new_n298_ );
or g098 ( new_n300_, new_n299_, new_n293_ );
or g099 ( new_n301_, new_n300_, new_n290_ );
or g100 ( new_n302_, new_n301_, keyIn_0_74 );
not g101 ( new_n303_, keyIn_0_74 );
and g102 ( new_n304_, new_n224_, new_n277_ );
or g103 ( new_n305_, new_n265_, keyIn_0_52 );
or g104 ( new_n306_, new_n292_, new_n291_ );
and g105 ( new_n307_, new_n306_, new_n296_ );
and g106 ( new_n308_, new_n307_, new_n305_ );
and g107 ( new_n309_, new_n308_, new_n304_ );
or g108 ( new_n310_, new_n309_, new_n303_ );
and g109 ( new_n311_, new_n302_, new_n310_ );
not g110 ( new_n312_, new_n240_ );
not g111 ( new_n313_, new_n277_ );
and g112 ( new_n314_, new_n313_, new_n312_ );
and g113 ( new_n315_, new_n294_, new_n314_ );
and g114 ( new_n316_, new_n290_, new_n315_ );
xnor g115 ( new_n317_, new_n316_, keyIn_0_75 );
not g116 ( new_n318_, new_n317_ );
and g117 ( new_n319_, new_n311_, new_n318_ );
and g118 ( new_n320_, new_n319_, new_n289_ );
and g119 ( new_n321_, new_n320_, new_n281_ );
or g120 ( new_n322_, new_n321_, new_n225_ );
not g121 ( new_n323_, new_n281_ );
not g122 ( new_n324_, new_n289_ );
not g123 ( new_n325_, new_n302_ );
or g124 ( new_n326_, new_n325_, keyIn_0_78 );
and g125 ( new_n327_, new_n301_, keyIn_0_74 );
or g126 ( new_n328_, new_n327_, new_n317_ );
or g127 ( new_n329_, new_n326_, new_n328_ );
or g128 ( new_n330_, new_n329_, new_n324_ );
or g129 ( new_n331_, new_n330_, new_n323_ );
and g130 ( new_n332_, new_n322_, new_n331_ );
not g131 ( new_n333_, keyIn_0_53 );
xnor g132 ( new_n334_, N49, N53 );
xnor g133 ( new_n335_, new_n334_, keyIn_0_3 );
xnor g134 ( new_n336_, N57, N61 );
xnor g135 ( new_n337_, new_n336_, keyIn_0_4 );
xnor g136 ( new_n338_, new_n335_, new_n337_ );
xnor g137 ( new_n339_, new_n338_, keyIn_0_27 );
xnor g138 ( new_n340_, N33, N37 );
xnor g139 ( new_n341_, new_n340_, keyIn_0_1 );
xor g140 ( new_n342_, N41, N45 );
xnor g141 ( new_n343_, new_n342_, keyIn_0_2 );
xnor g142 ( new_n344_, new_n343_, new_n341_ );
xor g143 ( new_n345_, new_n344_, keyIn_0_26 );
xnor g144 ( new_n346_, new_n345_, new_n339_ );
xnor g145 ( new_n347_, new_n346_, keyIn_0_33 );
and g146 ( new_n348_, N134, N137 );
xnor g147 ( new_n349_, new_n348_, keyIn_0_14 );
xnor g148 ( new_n350_, new_n347_, new_n349_ );
xnor g149 ( new_n351_, new_n350_, keyIn_0_39 );
xnor g150 ( new_n352_, N69, N85 );
xnor g151 ( new_n353_, new_n352_, keyIn_0_23 );
xnor g152 ( new_n354_, N101, N117 );
xnor g153 ( new_n355_, new_n354_, keyIn_0_24 );
xnor g154 ( new_n356_, new_n353_, new_n355_ );
xnor g155 ( new_n357_, new_n351_, new_n356_ );
xnor g156 ( new_n358_, new_n357_, keyIn_0_43 );
not g157 ( new_n359_, new_n358_ );
and g158 ( new_n360_, new_n359_, new_n333_ );
and g159 ( new_n361_, new_n358_, keyIn_0_53 );
xnor g160 ( new_n362_, N17, N21 );
xnor g161 ( new_n363_, new_n362_, keyIn_0_0 );
xnor g162 ( new_n364_, N25, N29 );
xnor g163 ( new_n365_, new_n363_, new_n364_ );
xnor g164 ( new_n366_, new_n365_, keyIn_0_25 );
xor g165 ( new_n367_, N9, N13 );
xnor g166 ( new_n368_, N1, N5 );
xnor g167 ( new_n369_, new_n367_, new_n368_ );
xnor g168 ( new_n370_, new_n366_, new_n369_ );
and g169 ( new_n371_, N133, N137 );
xnor g170 ( new_n372_, new_n371_, keyIn_0_13 );
xnor g171 ( new_n373_, new_n370_, new_n372_ );
xnor g172 ( new_n374_, new_n373_, keyIn_0_38 );
xnor g173 ( new_n375_, N97, N113 );
xor g174 ( new_n376_, new_n375_, keyIn_0_22 );
xor g175 ( new_n377_, N65, N81 );
xnor g176 ( new_n378_, new_n377_, keyIn_0_21 );
xnor g177 ( new_n379_, new_n376_, new_n378_ );
xnor g178 ( new_n380_, new_n374_, new_n379_ );
xor g179 ( new_n381_, new_n380_, keyIn_0_42 );
not g180 ( new_n382_, new_n381_ );
not g181 ( new_n383_, keyIn_0_54 );
xnor g182 ( new_n384_, new_n339_, new_n366_ );
and g183 ( new_n385_, N136, N137 );
xnor g184 ( new_n386_, new_n385_, keyIn_0_15 );
xnor g185 ( new_n387_, new_n384_, new_n386_ );
xnor g186 ( new_n388_, N109, N125 );
xnor g187 ( new_n389_, N77, N93 );
xnor g188 ( new_n390_, new_n388_, new_n389_ );
xnor g189 ( new_n391_, new_n390_, keyIn_0_32 );
xnor g190 ( new_n392_, new_n387_, new_n391_ );
xor g191 ( new_n393_, new_n392_, keyIn_0_45 );
and g192 ( new_n394_, new_n393_, new_n383_ );
not g193 ( new_n395_, new_n393_ );
and g194 ( new_n396_, new_n395_, keyIn_0_54 );
xnor g195 ( new_n397_, new_n345_, new_n369_ );
and g196 ( new_n398_, N135, N137 );
xnor g197 ( new_n399_, new_n397_, new_n398_ );
xnor g198 ( new_n400_, N105, N121 );
xnor g199 ( new_n401_, N73, N89 );
xnor g200 ( new_n402_, new_n400_, new_n401_ );
xnor g201 ( new_n403_, new_n402_, keyIn_0_31 );
xnor g202 ( new_n404_, new_n399_, new_n403_ );
xnor g203 ( new_n405_, new_n404_, keyIn_0_44 );
not g204 ( new_n406_, new_n405_ );
or g205 ( new_n407_, new_n396_, new_n406_ );
or g206 ( new_n408_, new_n407_, new_n394_ );
or g207 ( new_n409_, new_n408_, new_n382_ );
or g208 ( new_n410_, new_n409_, new_n361_ );
or g209 ( new_n411_, new_n410_, new_n360_ );
or g210 ( new_n412_, new_n332_, new_n411_ );
or g211 ( new_n413_, new_n412_, new_n224_ );
xor g212 ( new_n414_, new_n413_, N1 );
xnor g213 ( N724, new_n414_, keyIn_0_107 );
or g214 ( new_n416_, new_n412_, new_n313_ );
xnor g215 ( new_n417_, new_n416_, keyIn_0_86 );
xnor g216 ( new_n418_, new_n417_, N5 );
xnor g217 ( N725, new_n418_, keyIn_0_108 );
or g218 ( new_n420_, new_n412_, new_n312_ );
xnor g219 ( new_n421_, new_n420_, keyIn_0_87 );
xnor g220 ( new_n422_, new_n421_, N9 );
xor g221 ( N726, new_n422_, keyIn_0_109 );
or g222 ( new_n424_, new_n412_, new_n294_ );
xor g223 ( new_n425_, new_n424_, keyIn_0_88 );
xnor g224 ( new_n426_, new_n425_, N13 );
xnor g225 ( N727, new_n426_, keyIn_0_110 );
xor g226 ( new_n428_, new_n358_, keyIn_0_55 );
or g227 ( new_n429_, new_n395_, new_n405_ );
or g228 ( new_n430_, new_n382_, new_n429_ );
or g229 ( new_n431_, new_n428_, new_n430_ );
or g230 ( new_n432_, new_n332_, new_n431_ );
xnor g231 ( new_n433_, new_n432_, keyIn_0_80 );
and g232 ( new_n434_, new_n433_, new_n290_ );
xor g233 ( N728, new_n434_, N17 );
and g234 ( new_n436_, new_n433_, new_n277_ );
xor g235 ( N729, new_n436_, N21 );
and g236 ( new_n438_, new_n433_, new_n240_ );
xor g237 ( N730, new_n438_, N25 );
and g238 ( new_n440_, new_n433_, new_n292_ );
xnor g239 ( new_n441_, new_n440_, N29 );
xor g240 ( N731, new_n441_, keyIn_0_111 );
and g241 ( new_n443_, new_n381_, keyIn_0_56 );
not g242 ( new_n444_, keyIn_0_56 );
and g243 ( new_n445_, new_n382_, new_n444_ );
or g244 ( new_n446_, new_n406_, new_n393_ );
or g245 ( new_n447_, new_n445_, new_n446_ );
or g246 ( new_n448_, new_n447_, new_n443_ );
or g247 ( new_n449_, new_n448_, new_n358_ );
or g248 ( new_n450_, new_n332_, new_n449_ );
or g249 ( new_n451_, new_n450_, new_n224_ );
xnor g250 ( new_n452_, new_n451_, keyIn_0_89 );
xnor g251 ( new_n453_, new_n452_, N33 );
xnor g252 ( N732, new_n453_, keyIn_0_112 );
or g253 ( new_n455_, new_n450_, new_n313_ );
xnor g254 ( new_n456_, new_n455_, keyIn_0_90 );
xnor g255 ( new_n457_, new_n456_, N37 );
xor g256 ( N733, new_n457_, keyIn_0_113 );
or g257 ( new_n459_, new_n450_, new_n312_ );
xnor g258 ( new_n460_, new_n459_, keyIn_0_91 );
xnor g259 ( N734, new_n460_, N41 );
or g260 ( new_n462_, new_n450_, new_n265_ );
xnor g261 ( new_n463_, new_n462_, N45 );
xor g262 ( N735, new_n463_, keyIn_0_114 );
not g263 ( new_n465_, keyIn_0_81 );
not g264 ( new_n466_, keyIn_0_57 );
and g265 ( new_n467_, new_n382_, new_n466_ );
and g266 ( new_n468_, new_n381_, keyIn_0_57 );
and g267 ( new_n469_, new_n406_, keyIn_0_58 );
not g268 ( new_n470_, keyIn_0_58 );
and g269 ( new_n471_, new_n405_, new_n470_ );
or g270 ( new_n472_, new_n471_, new_n395_ );
or g271 ( new_n473_, new_n472_, new_n469_ );
or g272 ( new_n474_, new_n473_, new_n468_ );
or g273 ( new_n475_, new_n474_, new_n467_ );
or g274 ( new_n476_, new_n475_, new_n358_ );
or g275 ( new_n477_, new_n332_, new_n476_ );
xnor g276 ( new_n478_, new_n477_, new_n465_ );
and g277 ( new_n479_, new_n478_, new_n290_ );
xnor g278 ( new_n480_, new_n479_, keyIn_0_92 );
xor g279 ( N736, new_n480_, N49 );
and g280 ( new_n482_, new_n478_, new_n277_ );
xnor g281 ( new_n483_, new_n482_, keyIn_0_93 );
xor g282 ( N737, new_n483_, N53 );
not g283 ( new_n485_, keyIn_0_115 );
and g284 ( new_n486_, new_n478_, new_n240_ );
xnor g285 ( new_n487_, new_n486_, keyIn_0_94 );
xnor g286 ( new_n488_, new_n487_, N57 );
xnor g287 ( N738, new_n488_, new_n485_ );
and g288 ( new_n490_, new_n478_, new_n292_ );
xnor g289 ( new_n491_, new_n490_, keyIn_0_95 );
xnor g290 ( new_n492_, new_n491_, N61 );
xnor g291 ( N739, new_n492_, keyIn_0_116 );
not g292 ( new_n494_, keyIn_0_79 );
not g293 ( new_n495_, keyIn_0_59 );
and g294 ( new_n496_, new_n359_, new_n495_ );
and g295 ( new_n497_, new_n358_, keyIn_0_59 );
and g296 ( new_n498_, new_n406_, keyIn_0_60 );
not g297 ( new_n499_, keyIn_0_60 );
and g298 ( new_n500_, new_n405_, new_n499_ );
or g299 ( new_n501_, new_n500_, new_n395_ );
or g300 ( new_n502_, new_n501_, new_n498_ );
or g301 ( new_n503_, new_n502_, new_n381_ );
or g302 ( new_n504_, new_n503_, new_n497_ );
or g303 ( new_n505_, new_n504_, new_n496_ );
xnor g304 ( new_n506_, new_n505_, keyIn_0_76 );
not g305 ( new_n507_, keyIn_0_62 );
or g306 ( new_n508_, new_n382_, new_n507_ );
or g307 ( new_n509_, new_n381_, keyIn_0_62 );
xor g308 ( new_n510_, new_n405_, keyIn_0_63 );
xor g309 ( new_n511_, new_n393_, keyIn_0_64 );
and g310 ( new_n512_, new_n510_, new_n511_ );
and g311 ( new_n513_, new_n512_, new_n509_ );
and g312 ( new_n514_, new_n513_, new_n508_ );
and g313 ( new_n515_, new_n514_, new_n359_ );
not g314 ( new_n516_, new_n515_ );
not g315 ( new_n517_, keyIn_0_61 );
and g316 ( new_n518_, new_n395_, new_n517_ );
and g317 ( new_n519_, new_n393_, keyIn_0_61 );
or g318 ( new_n520_, new_n519_, new_n406_ );
or g319 ( new_n521_, new_n520_, new_n518_ );
or g320 ( new_n522_, new_n521_, new_n381_ );
or g321 ( new_n523_, new_n522_, new_n359_ );
and g322 ( new_n524_, new_n516_, new_n523_ );
xnor g323 ( new_n525_, new_n405_, keyIn_0_65 );
xnor g324 ( new_n526_, new_n393_, keyIn_0_66 );
and g325 ( new_n527_, new_n526_, new_n381_ );
and g326 ( new_n528_, new_n527_, new_n525_ );
and g327 ( new_n529_, new_n528_, new_n358_ );
xor g328 ( new_n530_, new_n529_, keyIn_0_77 );
and g329 ( new_n531_, new_n524_, new_n530_ );
and g330 ( new_n532_, new_n531_, new_n506_ );
xnor g331 ( new_n533_, new_n532_, new_n494_ );
not g332 ( new_n534_, keyIn_0_68 );
or g333 ( new_n535_, new_n294_, new_n534_ );
or g334 ( new_n536_, new_n292_, keyIn_0_68 );
or g335 ( new_n537_, new_n313_, keyIn_0_67 );
not g336 ( new_n538_, keyIn_0_67 );
or g337 ( new_n539_, new_n277_, new_n538_ );
and g338 ( new_n540_, new_n539_, new_n240_ );
and g339 ( new_n541_, new_n540_, new_n537_ );
and g340 ( new_n542_, new_n536_, new_n541_ );
and g341 ( new_n543_, new_n542_, new_n535_ );
and g342 ( new_n544_, new_n543_, new_n290_ );
and g343 ( new_n545_, new_n533_, new_n544_ );
xnor g344 ( new_n546_, new_n545_, keyIn_0_82 );
and g345 ( new_n547_, new_n546_, new_n381_ );
xor g346 ( new_n548_, new_n547_, keyIn_0_96 );
xnor g347 ( new_n549_, new_n548_, N65 );
xor g348 ( N740, new_n549_, keyIn_0_117 );
and g349 ( new_n551_, new_n546_, new_n359_ );
xnor g350 ( new_n552_, new_n551_, keyIn_0_97 );
xnor g351 ( new_n553_, new_n552_, N69 );
xor g352 ( N741, new_n553_, keyIn_0_118 );
and g353 ( new_n555_, new_n546_, new_n405_ );
xnor g354 ( new_n556_, new_n555_, keyIn_0_98 );
xnor g355 ( N742, new_n556_, N73 );
and g356 ( new_n558_, new_n546_, new_n393_ );
xnor g357 ( new_n559_, new_n558_, N77 );
xnor g358 ( N743, new_n559_, keyIn_0_119 );
xnor g359 ( new_n561_, new_n277_, keyIn_0_69 );
xnor g360 ( new_n562_, new_n240_, keyIn_0_70 );
and g361 ( new_n563_, new_n561_, new_n562_ );
and g362 ( new_n564_, new_n283_, new_n563_ );
and g363 ( new_n565_, new_n290_, new_n564_ );
and g364 ( new_n566_, new_n533_, new_n565_ );
xnor g365 ( new_n567_, new_n566_, keyIn_0_83 );
not g366 ( new_n568_, keyIn_0_83 );
or g367 ( new_n569_, new_n564_, new_n568_ );
and g368 ( new_n570_, new_n567_, new_n569_ );
or g369 ( new_n571_, new_n382_, keyIn_0_99 );
or g370 ( new_n572_, new_n570_, new_n571_ );
not g371 ( new_n573_, keyIn_0_99 );
not g372 ( new_n574_, new_n567_ );
and g373 ( new_n575_, new_n574_, new_n381_ );
or g374 ( new_n576_, new_n575_, new_n573_ );
and g375 ( new_n577_, new_n576_, new_n572_ );
xnor g376 ( new_n578_, new_n577_, N81 );
xnor g377 ( N744, new_n578_, keyIn_0_120 );
and g378 ( new_n580_, new_n574_, new_n359_ );
xnor g379 ( new_n581_, new_n580_, N85 );
xor g380 ( N745, new_n581_, keyIn_0_121 );
or g381 ( new_n583_, new_n406_, keyIn_0_100 );
or g382 ( new_n584_, new_n570_, new_n583_ );
not g383 ( new_n585_, keyIn_0_100 );
and g384 ( new_n586_, new_n574_, new_n405_ );
or g385 ( new_n587_, new_n586_, new_n585_ );
and g386 ( new_n588_, new_n587_, new_n584_ );
xnor g387 ( new_n589_, new_n588_, N89 );
xnor g388 ( N746, new_n589_, keyIn_0_122 );
and g389 ( new_n591_, new_n574_, new_n393_ );
xnor g390 ( new_n592_, new_n591_, keyIn_0_101 );
xnor g391 ( N747, new_n592_, N93 );
and g392 ( new_n594_, new_n304_, new_n266_ );
and g393 ( new_n595_, new_n533_, new_n594_ );
xnor g394 ( new_n596_, new_n595_, keyIn_0_84 );
and g395 ( new_n597_, new_n596_, new_n381_ );
xnor g396 ( new_n598_, new_n597_, keyIn_0_102 );
xnor g397 ( N748, new_n598_, N97 );
not g398 ( new_n600_, keyIn_0_84 );
or g399 ( new_n601_, new_n266_, new_n600_ );
and g400 ( new_n602_, new_n596_, new_n601_ );
and g401 ( new_n603_, new_n602_, new_n359_ );
xnor g402 ( new_n604_, new_n603_, keyIn_0_103 );
xnor g403 ( N749, new_n604_, N101 );
not g404 ( new_n606_, keyIn_0_123 );
not g405 ( new_n607_, new_n596_ );
not g406 ( new_n608_, keyIn_0_104 );
or g407 ( new_n609_, new_n406_, new_n608_ );
or g408 ( new_n610_, new_n607_, new_n609_ );
and g409 ( new_n611_, new_n602_, new_n405_ );
or g410 ( new_n612_, new_n611_, keyIn_0_104 );
and g411 ( new_n613_, new_n612_, new_n610_ );
xnor g412 ( new_n614_, new_n613_, N105 );
xnor g413 ( N750, new_n614_, new_n606_ );
and g414 ( new_n616_, new_n602_, new_n393_ );
xor g415 ( N751, new_n616_, N109 );
xor g416 ( new_n618_, new_n240_, keyIn_0_71 );
and g417 ( new_n619_, new_n292_, new_n618_ );
and g418 ( new_n620_, new_n304_, new_n619_ );
and g419 ( new_n621_, new_n533_, new_n620_ );
xor g420 ( new_n622_, new_n621_, keyIn_0_85 );
and g421 ( new_n623_, new_n622_, new_n381_ );
xnor g422 ( new_n624_, new_n623_, keyIn_0_105 );
xnor g423 ( new_n625_, new_n624_, N113 );
xor g424 ( N752, new_n625_, keyIn_0_124 );
and g425 ( new_n627_, new_n622_, new_n359_ );
xnor g426 ( new_n628_, new_n627_, keyIn_0_106 );
xnor g427 ( new_n629_, new_n628_, N117 );
xor g428 ( N753, new_n629_, keyIn_0_125 );
and g429 ( new_n631_, new_n622_, new_n405_ );
xnor g430 ( new_n632_, new_n631_, N121 );
xnor g431 ( N754, new_n632_, keyIn_0_126 );
and g432 ( new_n634_, new_n622_, new_n393_ );
xnor g433 ( new_n635_, new_n634_, N125 );
xnor g434 ( N755, new_n635_, keyIn_0_127 );
endmodule