module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n108_, keyIn_0_14 );
or g001 ( new_n109_, keyIn_0_6, N89 );
not g002 ( new_n110_, N95 );
and g003 ( new_n111_, keyIn_0_6, N89 );
or g004 ( new_n112_, new_n111_, new_n110_ );
not g005 ( new_n113_, new_n112_ );
and g006 ( new_n114_, new_n113_, new_n109_ );
and g007 ( new_n115_, new_n114_, keyIn_0_12 );
not g008 ( new_n116_, new_n115_ );
or g009 ( new_n117_, new_n114_, keyIn_0_12 );
and g010 ( new_n118_, new_n116_, new_n117_ );
not g011 ( new_n119_, new_n118_ );
not g012 ( new_n120_, N30 );
not g013 ( new_n121_, keyIn_0_1 );
or g014 ( new_n122_, new_n121_, N24 );
not g015 ( new_n123_, N24 );
or g016 ( new_n124_, new_n123_, keyIn_0_1 );
and g017 ( new_n125_, new_n122_, new_n124_ );
or g018 ( new_n126_, new_n125_, new_n120_ );
and g019 ( new_n127_, new_n126_, keyIn_0_8 );
not g020 ( new_n128_, keyIn_0_8 );
and g021 ( new_n129_, new_n123_, keyIn_0_1 );
and g022 ( new_n130_, new_n121_, N24 );
or g023 ( new_n131_, new_n129_, new_n130_ );
and g024 ( new_n132_, new_n131_, N30 );
and g025 ( new_n133_, new_n132_, new_n128_ );
or g026 ( new_n134_, new_n127_, new_n133_ );
not g027 ( new_n135_, keyIn_0_10 );
not g028 ( new_n136_, N56 );
and g029 ( new_n137_, keyIn_0_4, N50 );
not g030 ( new_n138_, new_n137_ );
or g031 ( new_n139_, keyIn_0_4, N50 );
and g032 ( new_n140_, new_n138_, new_n139_ );
or g033 ( new_n141_, new_n140_, new_n136_ );
and g034 ( new_n142_, new_n141_, new_n135_ );
not g035 ( new_n143_, keyIn_0_4 );
not g036 ( new_n144_, N50 );
and g037 ( new_n145_, new_n143_, new_n144_ );
or g038 ( new_n146_, new_n145_, new_n137_ );
and g039 ( new_n147_, new_n146_, N56 );
and g040 ( new_n148_, new_n147_, keyIn_0_10 );
or g041 ( new_n149_, new_n142_, new_n148_ );
and g042 ( new_n150_, new_n134_, new_n149_ );
and g043 ( new_n151_, new_n150_, new_n119_ );
not g044 ( new_n152_, N43 );
not g045 ( new_n153_, keyIn_0_2 );
or g046 ( new_n154_, new_n153_, N37 );
not g047 ( new_n155_, N37 );
or g048 ( new_n156_, new_n155_, keyIn_0_2 );
and g049 ( new_n157_, new_n154_, new_n156_ );
or g050 ( new_n158_, new_n157_, new_n152_ );
and g051 ( new_n159_, new_n158_, keyIn_0_9 );
not g052 ( new_n160_, keyIn_0_9 );
and g053 ( new_n161_, new_n155_, keyIn_0_2 );
and g054 ( new_n162_, new_n153_, N37 );
or g055 ( new_n163_, new_n161_, new_n162_ );
and g056 ( new_n164_, new_n163_, N43 );
and g057 ( new_n165_, new_n164_, new_n160_ );
or g058 ( new_n166_, new_n159_, new_n165_ );
not g059 ( new_n167_, keyIn_0_0 );
and g060 ( new_n168_, new_n167_, N1 );
not g061 ( new_n169_, new_n168_ );
or g062 ( new_n170_, new_n167_, N1 );
and g063 ( new_n171_, new_n170_, N4 );
and g064 ( new_n172_, new_n171_, new_n169_ );
not g065 ( new_n173_, N11 );
and g066 ( new_n174_, new_n173_, N17 );
not g067 ( new_n175_, N63 );
and g068 ( new_n176_, new_n175_, N69 );
or g069 ( new_n177_, new_n174_, new_n176_ );
or g070 ( new_n178_, new_n172_, new_n177_ );
not g071 ( new_n179_, new_n178_ );
and g072 ( new_n180_, new_n166_, new_n179_ );
not g073 ( new_n181_, keyIn_0_7 );
and g074 ( new_n182_, new_n181_, N102 );
not g075 ( new_n183_, N108 );
not g076 ( new_n184_, N102 );
and g077 ( new_n185_, new_n184_, keyIn_0_7 );
or g078 ( new_n186_, new_n185_, new_n183_ );
or g079 ( new_n187_, new_n186_, new_n182_ );
and g080 ( new_n188_, new_n187_, keyIn_0_13 );
not g081 ( new_n189_, keyIn_0_13 );
not g082 ( new_n190_, new_n182_ );
or g083 ( new_n191_, new_n181_, N102 );
and g084 ( new_n192_, new_n191_, N108 );
and g085 ( new_n193_, new_n192_, new_n190_ );
and g086 ( new_n194_, new_n193_, new_n189_ );
or g087 ( new_n195_, new_n188_, new_n194_ );
not g088 ( new_n196_, N76 );
and g089 ( new_n197_, new_n196_, keyIn_0_5 );
not g090 ( new_n198_, keyIn_0_5 );
and g091 ( new_n199_, new_n198_, N76 );
or g092 ( new_n200_, new_n197_, new_n199_ );
and g093 ( new_n201_, new_n200_, N82 );
and g094 ( new_n202_, new_n201_, keyIn_0_11 );
not g095 ( new_n203_, keyIn_0_11 );
not g096 ( new_n204_, N82 );
or g097 ( new_n205_, new_n198_, N76 );
or g098 ( new_n206_, new_n196_, keyIn_0_5 );
and g099 ( new_n207_, new_n205_, new_n206_ );
or g100 ( new_n208_, new_n207_, new_n204_ );
and g101 ( new_n209_, new_n208_, new_n203_ );
or g102 ( new_n210_, new_n209_, new_n202_ );
and g103 ( new_n211_, new_n210_, new_n195_ );
and g104 ( new_n212_, new_n180_, new_n211_ );
and g105 ( new_n213_, new_n212_, new_n151_ );
and g106 ( new_n214_, new_n213_, new_n108_ );
not g107 ( new_n215_, new_n214_ );
or g108 ( new_n216_, new_n213_, new_n108_ );
and g109 ( N223, new_n215_, new_n216_ );
not g110 ( new_n218_, keyIn_0_28 );
not g111 ( new_n219_, keyIn_0_26 );
not g112 ( new_n220_, keyIn_0_20 );
or g113 ( new_n221_, new_n132_, new_n128_ );
or g114 ( new_n222_, new_n126_, keyIn_0_8 );
and g115 ( new_n223_, new_n222_, new_n221_ );
or g116 ( new_n224_, new_n147_, keyIn_0_10 );
or g117 ( new_n225_, new_n141_, new_n135_ );
and g118 ( new_n226_, new_n224_, new_n225_ );
or g119 ( new_n227_, new_n223_, new_n226_ );
or g120 ( new_n228_, new_n227_, new_n118_ );
or g121 ( new_n229_, new_n164_, new_n160_ );
or g122 ( new_n230_, new_n158_, keyIn_0_9 );
and g123 ( new_n231_, new_n230_, new_n229_ );
or g124 ( new_n232_, new_n231_, new_n178_ );
or g125 ( new_n233_, new_n193_, new_n189_ );
or g126 ( new_n234_, new_n187_, keyIn_0_13 );
and g127 ( new_n235_, new_n234_, new_n233_ );
or g128 ( new_n236_, new_n208_, new_n203_ );
or g129 ( new_n237_, new_n201_, keyIn_0_11 );
and g130 ( new_n238_, new_n236_, new_n237_ );
or g131 ( new_n239_, new_n238_, new_n235_ );
or g132 ( new_n240_, new_n239_, new_n232_ );
or g133 ( new_n241_, new_n240_, new_n228_ );
and g134 ( new_n242_, new_n241_, keyIn_0_14 );
or g135 ( new_n243_, new_n242_, new_n214_ );
and g136 ( new_n244_, new_n243_, keyIn_0_15 );
not g137 ( new_n245_, keyIn_0_15 );
and g138 ( new_n246_, N223, new_n245_ );
or g139 ( new_n247_, new_n244_, new_n246_ );
and g140 ( new_n248_, new_n247_, new_n176_ );
not g141 ( new_n249_, new_n248_ );
or g142 ( new_n250_, new_n247_, new_n176_ );
and g143 ( new_n251_, new_n249_, new_n250_ );
and g144 ( new_n252_, new_n251_, new_n220_ );
not g145 ( new_n253_, new_n252_ );
or g146 ( new_n254_, new_n251_, new_n220_ );
and g147 ( new_n255_, new_n253_, new_n254_ );
not g148 ( new_n256_, N73 );
and g149 ( new_n257_, new_n256_, N69 );
and g150 ( new_n258_, new_n255_, new_n257_ );
and g151 ( new_n259_, new_n258_, new_n219_ );
not g152 ( new_n260_, new_n259_ );
or g153 ( new_n261_, new_n258_, new_n219_ );
and g154 ( new_n262_, new_n260_, new_n261_ );
and g155 ( new_n263_, new_n247_, new_n172_ );
not g156 ( new_n264_, new_n172_ );
or g157 ( new_n265_, N223, new_n245_ );
or g158 ( new_n266_, new_n243_, keyIn_0_15 );
and g159 ( new_n267_, new_n266_, new_n265_ );
and g160 ( new_n268_, new_n267_, new_n264_ );
or g161 ( new_n269_, new_n263_, new_n268_ );
and g162 ( new_n270_, new_n269_, keyIn_0_16 );
not g163 ( new_n271_, keyIn_0_16 );
or g164 ( new_n272_, new_n267_, new_n264_ );
or g165 ( new_n273_, new_n247_, new_n172_ );
and g166 ( new_n274_, new_n273_, new_n272_ );
and g167 ( new_n275_, new_n274_, new_n271_ );
or g168 ( new_n276_, new_n270_, new_n275_ );
not g169 ( new_n277_, N8 );
and g170 ( new_n278_, new_n277_, N4 );
not g171 ( new_n279_, new_n278_ );
or g172 ( new_n280_, new_n276_, new_n279_ );
or g173 ( new_n281_, new_n280_, keyIn_0_22 );
not g174 ( new_n282_, keyIn_0_22 );
or g175 ( new_n283_, new_n274_, new_n271_ );
or g176 ( new_n284_, new_n269_, keyIn_0_16 );
and g177 ( new_n285_, new_n284_, new_n283_ );
and g178 ( new_n286_, new_n285_, new_n278_ );
or g179 ( new_n287_, new_n286_, new_n282_ );
and g180 ( new_n288_, new_n281_, new_n287_ );
not g181 ( new_n289_, keyIn_0_25 );
not g182 ( new_n290_, keyIn_0_19 );
and g183 ( new_n291_, new_n247_, new_n226_ );
and g184 ( new_n292_, new_n267_, new_n149_ );
or g185 ( new_n293_, new_n291_, new_n292_ );
or g186 ( new_n294_, new_n293_, new_n290_ );
or g187 ( new_n295_, new_n267_, new_n149_ );
or g188 ( new_n296_, new_n247_, new_n226_ );
and g189 ( new_n297_, new_n296_, new_n295_ );
or g190 ( new_n298_, new_n297_, keyIn_0_19 );
and g191 ( new_n299_, new_n294_, new_n298_ );
not g192 ( new_n300_, N60 );
and g193 ( new_n301_, new_n300_, N56 );
not g194 ( new_n302_, new_n301_ );
or g195 ( new_n303_, new_n299_, new_n302_ );
or g196 ( new_n304_, new_n303_, new_n289_ );
and g197 ( new_n305_, new_n297_, keyIn_0_19 );
and g198 ( new_n306_, new_n293_, new_n290_ );
or g199 ( new_n307_, new_n306_, new_n305_ );
and g200 ( new_n308_, new_n307_, new_n301_ );
or g201 ( new_n309_, new_n308_, keyIn_0_25 );
and g202 ( new_n310_, new_n304_, new_n309_ );
or g203 ( new_n311_, new_n288_, new_n310_ );
or g204 ( new_n312_, new_n311_, new_n262_ );
and g205 ( new_n313_, new_n247_, new_n235_ );
and g206 ( new_n314_, new_n267_, new_n195_ );
or g207 ( new_n315_, new_n313_, new_n314_ );
and g208 ( new_n316_, new_n315_, keyIn_0_21 );
not g209 ( new_n317_, keyIn_0_21 );
or g210 ( new_n318_, new_n267_, new_n195_ );
or g211 ( new_n319_, new_n247_, new_n235_ );
and g212 ( new_n320_, new_n319_, new_n318_ );
and g213 ( new_n321_, new_n320_, new_n317_ );
or g214 ( new_n322_, new_n316_, new_n321_ );
not g215 ( new_n323_, N112 );
and g216 ( new_n324_, new_n323_, N108 );
not g217 ( new_n325_, new_n324_ );
or g218 ( new_n326_, new_n322_, new_n325_ );
or g219 ( new_n327_, new_n326_, keyIn_0_27 );
not g220 ( new_n328_, keyIn_0_27 );
or g221 ( new_n329_, new_n320_, new_n317_ );
or g222 ( new_n330_, new_n315_, keyIn_0_21 );
and g223 ( new_n331_, new_n330_, new_n329_ );
and g224 ( new_n332_, new_n331_, new_n324_ );
or g225 ( new_n333_, new_n332_, new_n328_ );
and g226 ( new_n334_, new_n327_, new_n333_ );
not g227 ( new_n335_, N86 );
and g228 ( new_n336_, new_n247_, new_n238_ );
and g229 ( new_n337_, new_n267_, new_n210_ );
or g230 ( new_n338_, new_n336_, new_n337_ );
and g231 ( new_n339_, new_n338_, N82 );
and g232 ( new_n340_, new_n339_, new_n335_ );
not g233 ( new_n341_, new_n340_ );
not g234 ( new_n342_, N34 );
and g235 ( new_n343_, new_n247_, new_n223_ );
and g236 ( new_n344_, new_n267_, new_n134_ );
or g237 ( new_n345_, new_n343_, new_n344_ );
and g238 ( new_n346_, new_n345_, N30 );
and g239 ( new_n347_, new_n346_, new_n342_ );
not g240 ( new_n348_, new_n347_ );
not g241 ( new_n349_, N99 );
and g242 ( new_n350_, new_n247_, new_n118_ );
and g243 ( new_n351_, new_n267_, new_n119_ );
or g244 ( new_n352_, new_n350_, new_n351_ );
and g245 ( new_n353_, new_n352_, N95 );
and g246 ( new_n354_, new_n353_, new_n349_ );
not g247 ( new_n355_, new_n354_ );
and g248 ( new_n356_, new_n348_, new_n355_ );
and g249 ( new_n357_, new_n356_, new_n341_ );
not g250 ( new_n358_, new_n357_ );
or g251 ( new_n359_, new_n334_, new_n358_ );
and g252 ( new_n360_, new_n247_, new_n231_ );
and g253 ( new_n361_, new_n267_, new_n166_ );
or g254 ( new_n362_, new_n360_, new_n361_ );
or g255 ( new_n363_, new_n362_, keyIn_0_18 );
not g256 ( new_n364_, keyIn_0_18 );
or g257 ( new_n365_, new_n267_, new_n166_ );
or g258 ( new_n366_, new_n247_, new_n231_ );
and g259 ( new_n367_, new_n366_, new_n365_ );
or g260 ( new_n368_, new_n367_, new_n364_ );
and g261 ( new_n369_, new_n363_, new_n368_ );
not g262 ( new_n370_, N47 );
and g263 ( new_n371_, keyIn_0_3, N43 );
not g264 ( new_n372_, new_n371_ );
or g265 ( new_n373_, keyIn_0_3, N43 );
and g266 ( new_n374_, new_n372_, new_n373_ );
not g267 ( new_n375_, new_n374_ );
and g268 ( new_n376_, new_n375_, new_n370_ );
not g269 ( new_n377_, new_n376_ );
or g270 ( new_n378_, new_n369_, new_n377_ );
or g271 ( new_n379_, new_n378_, keyIn_0_24 );
not g272 ( new_n380_, keyIn_0_24 );
and g273 ( new_n381_, new_n367_, new_n364_ );
and g274 ( new_n382_, new_n362_, keyIn_0_18 );
or g275 ( new_n383_, new_n382_, new_n381_ );
and g276 ( new_n384_, new_n383_, new_n376_ );
or g277 ( new_n385_, new_n384_, new_n380_ );
and g278 ( new_n386_, new_n379_, new_n385_ );
not g279 ( new_n387_, keyIn_0_23 );
not g280 ( new_n388_, keyIn_0_17 );
and g281 ( new_n389_, new_n247_, new_n174_ );
not g282 ( new_n390_, new_n174_ );
and g283 ( new_n391_, new_n267_, new_n390_ );
or g284 ( new_n392_, new_n389_, new_n391_ );
or g285 ( new_n393_, new_n392_, new_n388_ );
or g286 ( new_n394_, new_n267_, new_n390_ );
or g287 ( new_n395_, new_n247_, new_n174_ );
and g288 ( new_n396_, new_n395_, new_n394_ );
or g289 ( new_n397_, new_n396_, keyIn_0_17 );
and g290 ( new_n398_, new_n393_, new_n397_ );
not g291 ( new_n399_, N21 );
and g292 ( new_n400_, new_n399_, N17 );
not g293 ( new_n401_, new_n400_ );
or g294 ( new_n402_, new_n398_, new_n401_ );
and g295 ( new_n403_, new_n402_, new_n387_ );
and g296 ( new_n404_, new_n396_, keyIn_0_17 );
and g297 ( new_n405_, new_n392_, new_n388_ );
or g298 ( new_n406_, new_n405_, new_n404_ );
and g299 ( new_n407_, new_n406_, new_n400_ );
and g300 ( new_n408_, new_n407_, keyIn_0_23 );
or g301 ( new_n409_, new_n403_, new_n408_ );
or g302 ( new_n410_, new_n409_, new_n386_ );
or g303 ( new_n411_, new_n410_, new_n359_ );
or g304 ( new_n412_, new_n411_, new_n312_ );
and g305 ( new_n413_, new_n412_, new_n218_ );
not g306 ( new_n414_, new_n258_ );
and g307 ( new_n415_, new_n414_, keyIn_0_26 );
or g308 ( new_n416_, new_n415_, new_n259_ );
and g309 ( new_n417_, new_n286_, new_n282_ );
and g310 ( new_n418_, new_n280_, keyIn_0_22 );
or g311 ( new_n419_, new_n418_, new_n417_ );
and g312 ( new_n420_, new_n308_, keyIn_0_25 );
and g313 ( new_n421_, new_n303_, new_n289_ );
or g314 ( new_n422_, new_n421_, new_n420_ );
and g315 ( new_n423_, new_n422_, new_n419_ );
and g316 ( new_n424_, new_n423_, new_n416_ );
and g317 ( new_n425_, new_n332_, new_n328_ );
and g318 ( new_n426_, new_n326_, keyIn_0_27 );
or g319 ( new_n427_, new_n426_, new_n425_ );
and g320 ( new_n428_, new_n427_, new_n357_ );
and g321 ( new_n429_, new_n384_, new_n380_ );
and g322 ( new_n430_, new_n378_, keyIn_0_24 );
or g323 ( new_n431_, new_n430_, new_n429_ );
or g324 ( new_n432_, new_n407_, keyIn_0_23 );
or g325 ( new_n433_, new_n402_, new_n387_ );
and g326 ( new_n434_, new_n433_, new_n432_ );
and g327 ( new_n435_, new_n431_, new_n434_ );
and g328 ( new_n436_, new_n435_, new_n428_ );
and g329 ( new_n437_, new_n424_, new_n436_ );
and g330 ( new_n438_, new_n437_, keyIn_0_28 );
or g331 ( N329, new_n413_, new_n438_ );
not g332 ( new_n440_, keyIn_0_43 );
not g333 ( new_n441_, keyIn_0_31 );
and g334 ( new_n442_, N329, new_n441_ );
or g335 ( new_n443_, new_n437_, keyIn_0_28 );
not g336 ( new_n444_, new_n438_ );
and g337 ( new_n445_, new_n444_, new_n443_ );
and g338 ( new_n446_, new_n445_, keyIn_0_31 );
or g339 ( new_n447_, new_n442_, new_n446_ );
and g340 ( new_n448_, new_n447_, new_n427_ );
or g341 ( new_n449_, new_n445_, keyIn_0_31 );
or g342 ( new_n450_, N329, new_n441_ );
and g343 ( new_n451_, new_n450_, new_n449_ );
and g344 ( new_n452_, new_n451_, new_n334_ );
or g345 ( new_n453_, new_n448_, new_n452_ );
not g346 ( new_n454_, new_n453_ );
and g347 ( new_n455_, new_n454_, keyIn_0_37 );
not g348 ( new_n456_, new_n455_ );
or g349 ( new_n457_, new_n454_, keyIn_0_37 );
not g350 ( new_n458_, N115 );
and g351 ( new_n459_, new_n458_, N108 );
and g352 ( new_n460_, new_n331_, new_n459_ );
not g353 ( new_n461_, new_n460_ );
and g354 ( new_n462_, new_n461_, keyIn_0_30 );
not g355 ( new_n463_, new_n462_ );
or g356 ( new_n464_, new_n461_, keyIn_0_30 );
and g357 ( new_n465_, new_n463_, new_n464_ );
not g358 ( new_n466_, new_n465_ );
and g359 ( new_n467_, new_n457_, new_n466_ );
and g360 ( new_n468_, new_n467_, new_n456_ );
and g361 ( new_n469_, new_n468_, new_n440_ );
not g362 ( new_n470_, new_n469_ );
or g363 ( new_n471_, new_n468_, new_n440_ );
and g364 ( new_n472_, new_n470_, new_n471_ );
not g365 ( new_n473_, keyIn_0_38 );
not g366 ( new_n474_, keyIn_0_32 );
or g367 ( new_n475_, new_n451_, new_n409_ );
or g368 ( new_n476_, new_n447_, new_n434_ );
and g369 ( new_n477_, new_n476_, new_n475_ );
and g370 ( new_n478_, new_n477_, new_n474_ );
not g371 ( new_n479_, new_n478_ );
or g372 ( new_n480_, new_n477_, new_n474_ );
not g373 ( new_n481_, N27 );
and g374 ( new_n482_, new_n481_, N17 );
and g375 ( new_n483_, new_n406_, new_n482_ );
and g376 ( new_n484_, new_n480_, new_n483_ );
and g377 ( new_n485_, new_n484_, new_n479_ );
and g378 ( new_n486_, new_n485_, new_n473_ );
not g379 ( new_n487_, new_n486_ );
or g380 ( new_n488_, new_n485_, new_n473_ );
and g381 ( new_n489_, new_n487_, new_n488_ );
not g382 ( new_n490_, keyIn_0_41 );
not g383 ( new_n491_, keyIn_0_35 );
or g384 ( new_n492_, new_n451_, new_n262_ );
or g385 ( new_n493_, new_n447_, new_n416_ );
and g386 ( new_n494_, new_n493_, new_n492_ );
and g387 ( new_n495_, new_n494_, new_n491_ );
and g388 ( new_n496_, new_n447_, new_n416_ );
and g389 ( new_n497_, new_n451_, new_n262_ );
or g390 ( new_n498_, new_n496_, new_n497_ );
and g391 ( new_n499_, new_n498_, keyIn_0_35 );
not g392 ( new_n500_, keyIn_0_29 );
not g393 ( new_n501_, N79 );
and g394 ( new_n502_, new_n501_, N69 );
and g395 ( new_n503_, new_n255_, new_n502_ );
not g396 ( new_n504_, new_n503_ );
and g397 ( new_n505_, new_n504_, new_n500_ );
and g398 ( new_n506_, new_n503_, keyIn_0_29 );
or g399 ( new_n507_, new_n505_, new_n506_ );
not g400 ( new_n508_, new_n507_ );
or g401 ( new_n509_, new_n499_, new_n508_ );
or g402 ( new_n510_, new_n509_, new_n495_ );
or g403 ( new_n511_, new_n510_, new_n490_ );
not g404 ( new_n512_, new_n495_ );
or g405 ( new_n513_, new_n494_, new_n491_ );
and g406 ( new_n514_, new_n513_, new_n507_ );
and g407 ( new_n515_, new_n514_, new_n512_ );
or g408 ( new_n516_, new_n515_, keyIn_0_41 );
and g409 ( new_n517_, new_n511_, new_n516_ );
or g410 ( new_n518_, new_n489_, new_n517_ );
or g411 ( new_n519_, new_n518_, new_n472_ );
not g412 ( new_n520_, keyIn_0_42 );
or g413 ( new_n521_, new_n451_, new_n354_ );
or g414 ( new_n522_, new_n447_, new_n355_ );
and g415 ( new_n523_, new_n522_, new_n521_ );
and g416 ( new_n524_, new_n523_, keyIn_0_36 );
not g417 ( new_n525_, new_n524_ );
or g418 ( new_n526_, new_n523_, keyIn_0_36 );
not g419 ( new_n527_, N105 );
and g420 ( new_n528_, new_n353_, new_n527_ );
and g421 ( new_n529_, new_n526_, new_n528_ );
and g422 ( new_n530_, new_n529_, new_n525_ );
and g423 ( new_n531_, new_n530_, new_n520_ );
not g424 ( new_n532_, keyIn_0_36 );
and g425 ( new_n533_, new_n447_, new_n355_ );
and g426 ( new_n534_, new_n451_, new_n354_ );
or g427 ( new_n535_, new_n533_, new_n534_ );
and g428 ( new_n536_, new_n535_, new_n532_ );
not g429 ( new_n537_, new_n528_ );
or g430 ( new_n538_, new_n536_, new_n537_ );
or g431 ( new_n539_, new_n538_, new_n524_ );
and g432 ( new_n540_, new_n539_, keyIn_0_42 );
not g433 ( new_n541_, keyIn_0_33 );
or g434 ( new_n542_, new_n451_, new_n347_ );
or g435 ( new_n543_, new_n447_, new_n348_ );
and g436 ( new_n544_, new_n543_, new_n542_ );
and g437 ( new_n545_, new_n544_, new_n541_ );
not g438 ( new_n546_, new_n545_ );
or g439 ( new_n547_, new_n544_, new_n541_ );
not g440 ( new_n548_, N40 );
and g441 ( new_n549_, new_n346_, new_n548_ );
and g442 ( new_n550_, new_n547_, new_n549_ );
and g443 ( new_n551_, new_n550_, new_n546_ );
and g444 ( new_n552_, new_n551_, keyIn_0_39 );
or g445 ( new_n553_, new_n540_, new_n552_ );
or g446 ( new_n554_, new_n553_, new_n531_ );
not g447 ( new_n555_, keyIn_0_39 );
and g448 ( new_n556_, new_n447_, new_n348_ );
and g449 ( new_n557_, new_n451_, new_n347_ );
or g450 ( new_n558_, new_n556_, new_n557_ );
and g451 ( new_n559_, new_n558_, keyIn_0_33 );
not g452 ( new_n560_, new_n549_ );
or g453 ( new_n561_, new_n559_, new_n560_ );
or g454 ( new_n562_, new_n561_, new_n545_ );
and g455 ( new_n563_, new_n562_, new_n555_ );
and g456 ( new_n564_, new_n447_, new_n419_ );
and g457 ( new_n565_, new_n451_, new_n288_ );
or g458 ( new_n566_, new_n564_, new_n565_ );
not g459 ( new_n567_, N14 );
and g460 ( new_n568_, new_n567_, N4 );
and g461 ( new_n569_, new_n285_, new_n568_ );
and g462 ( new_n570_, new_n566_, new_n569_ );
and g463 ( new_n571_, new_n447_, new_n431_ );
and g464 ( new_n572_, new_n451_, new_n386_ );
or g465 ( new_n573_, new_n571_, new_n572_ );
not g466 ( new_n574_, N53 );
and g467 ( new_n575_, new_n375_, new_n574_ );
and g468 ( new_n576_, new_n383_, new_n575_ );
and g469 ( new_n577_, new_n573_, new_n576_ );
and g470 ( new_n578_, new_n447_, new_n341_ );
and g471 ( new_n579_, new_n451_, new_n340_ );
or g472 ( new_n580_, new_n578_, new_n579_ );
not g473 ( new_n581_, N92 );
and g474 ( new_n582_, new_n339_, new_n581_ );
and g475 ( new_n583_, new_n580_, new_n582_ );
or g476 ( new_n584_, new_n577_, new_n583_ );
or g477 ( new_n585_, new_n584_, new_n570_ );
or g478 ( new_n586_, new_n563_, new_n585_ );
not g479 ( new_n587_, keyIn_0_34 );
or g480 ( new_n588_, new_n451_, new_n310_ );
or g481 ( new_n589_, new_n447_, new_n422_ );
and g482 ( new_n590_, new_n589_, new_n588_ );
and g483 ( new_n591_, new_n590_, new_n587_ );
and g484 ( new_n592_, new_n447_, new_n422_ );
and g485 ( new_n593_, new_n451_, new_n310_ );
or g486 ( new_n594_, new_n592_, new_n593_ );
and g487 ( new_n595_, new_n594_, keyIn_0_34 );
not g488 ( new_n596_, N66 );
and g489 ( new_n597_, new_n596_, N56 );
and g490 ( new_n598_, new_n307_, new_n597_ );
not g491 ( new_n599_, new_n598_ );
or g492 ( new_n600_, new_n595_, new_n599_ );
or g493 ( new_n601_, new_n600_, new_n591_ );
and g494 ( new_n602_, new_n601_, keyIn_0_40 );
not g495 ( new_n603_, keyIn_0_40 );
not g496 ( new_n604_, new_n591_ );
or g497 ( new_n605_, new_n590_, new_n587_ );
and g498 ( new_n606_, new_n605_, new_n598_ );
and g499 ( new_n607_, new_n606_, new_n604_ );
and g500 ( new_n608_, new_n607_, new_n603_ );
or g501 ( new_n609_, new_n602_, new_n608_ );
or g502 ( new_n610_, new_n586_, new_n609_ );
or g503 ( new_n611_, new_n610_, new_n554_ );
or g504 ( new_n612_, new_n519_, new_n611_ );
and g505 ( new_n613_, new_n612_, keyIn_0_44 );
not g506 ( new_n614_, keyIn_0_44 );
not g507 ( new_n615_, new_n471_ );
or g508 ( new_n616_, new_n615_, new_n469_ );
and g509 ( new_n617_, new_n447_, new_n434_ );
and g510 ( new_n618_, new_n451_, new_n409_ );
or g511 ( new_n619_, new_n617_, new_n618_ );
and g512 ( new_n620_, new_n619_, keyIn_0_32 );
not g513 ( new_n621_, new_n483_ );
or g514 ( new_n622_, new_n620_, new_n621_ );
or g515 ( new_n623_, new_n622_, new_n478_ );
and g516 ( new_n624_, new_n623_, keyIn_0_38 );
or g517 ( new_n625_, new_n624_, new_n486_ );
and g518 ( new_n626_, new_n515_, keyIn_0_41 );
and g519 ( new_n627_, new_n510_, new_n490_ );
or g520 ( new_n628_, new_n627_, new_n626_ );
and g521 ( new_n629_, new_n625_, new_n628_ );
and g522 ( new_n630_, new_n629_, new_n616_ );
not g523 ( new_n631_, new_n531_ );
or g524 ( new_n632_, new_n530_, new_n520_ );
or g525 ( new_n633_, new_n562_, new_n555_ );
and g526 ( new_n634_, new_n633_, new_n632_ );
and g527 ( new_n635_, new_n634_, new_n631_ );
or g528 ( new_n636_, new_n551_, keyIn_0_39 );
not g529 ( new_n637_, new_n585_ );
and g530 ( new_n638_, new_n636_, new_n637_ );
or g531 ( new_n639_, new_n607_, new_n603_ );
or g532 ( new_n640_, new_n601_, keyIn_0_40 );
and g533 ( new_n641_, new_n640_, new_n639_ );
and g534 ( new_n642_, new_n641_, new_n638_ );
and g535 ( new_n643_, new_n635_, new_n642_ );
and g536 ( new_n644_, new_n630_, new_n643_ );
and g537 ( new_n645_, new_n644_, new_n614_ );
or g538 ( N370, new_n613_, new_n645_ );
not g539 ( new_n647_, keyIn_0_58 );
not g540 ( new_n648_, keyIn_0_49 );
not g541 ( new_n649_, keyIn_0_45 );
or g542 ( new_n650_, new_n644_, new_n614_ );
not g543 ( new_n651_, new_n645_ );
and g544 ( new_n652_, new_n651_, new_n650_ );
and g545 ( new_n653_, new_n652_, new_n649_ );
and g546 ( new_n654_, N370, keyIn_0_45 );
or g547 ( new_n655_, new_n654_, new_n653_ );
and g548 ( new_n656_, new_n655_, N66 );
and g549 ( new_n657_, new_n656_, new_n648_ );
or g550 ( new_n658_, N370, keyIn_0_45 );
or g551 ( new_n659_, new_n652_, new_n649_ );
and g552 ( new_n660_, new_n658_, new_n659_ );
or g553 ( new_n661_, new_n660_, new_n596_ );
and g554 ( new_n662_, new_n661_, keyIn_0_49 );
or g555 ( new_n663_, new_n662_, new_n657_ );
and g556 ( new_n664_, N329, N60 );
and g557 ( new_n665_, N223, N50 );
or g558 ( new_n666_, new_n665_, new_n136_ );
or g559 ( new_n667_, new_n664_, new_n666_ );
not g560 ( new_n668_, new_n667_ );
and g561 ( new_n669_, new_n663_, new_n668_ );
and g562 ( new_n670_, new_n669_, keyIn_0_54 );
not g563 ( new_n671_, keyIn_0_54 );
or g564 ( new_n672_, new_n661_, keyIn_0_49 );
or g565 ( new_n673_, new_n656_, new_n648_ );
and g566 ( new_n674_, new_n672_, new_n673_ );
or g567 ( new_n675_, new_n674_, new_n667_ );
and g568 ( new_n676_, new_n675_, new_n671_ );
or g569 ( new_n677_, new_n676_, new_n670_ );
not g570 ( new_n678_, keyIn_0_48 );
and g571 ( new_n679_, new_n655_, N53 );
and g572 ( new_n680_, new_n679_, new_n678_ );
or g573 ( new_n681_, new_n660_, new_n574_ );
and g574 ( new_n682_, new_n681_, keyIn_0_48 );
or g575 ( new_n683_, new_n682_, new_n680_ );
and g576 ( new_n684_, N329, N47 );
and g577 ( new_n685_, N223, N37 );
or g578 ( new_n686_, new_n685_, new_n152_ );
or g579 ( new_n687_, new_n684_, new_n686_ );
not g580 ( new_n688_, new_n687_ );
and g581 ( new_n689_, new_n683_, new_n688_ );
or g582 ( new_n690_, new_n689_, keyIn_0_53 );
and g583 ( new_n691_, new_n689_, keyIn_0_53 );
not g584 ( new_n692_, new_n691_ );
and g585 ( new_n693_, new_n692_, new_n690_ );
and g586 ( new_n694_, new_n693_, new_n677_ );
and g587 ( new_n695_, new_n655_, N40 );
and g588 ( new_n696_, new_n695_, keyIn_0_47 );
not g589 ( new_n697_, keyIn_0_47 );
or g590 ( new_n698_, new_n660_, new_n548_ );
and g591 ( new_n699_, new_n698_, new_n697_ );
or g592 ( new_n700_, new_n699_, new_n696_ );
and g593 ( new_n701_, N329, N34 );
and g594 ( new_n702_, N223, N24 );
or g595 ( new_n703_, new_n702_, new_n120_ );
or g596 ( new_n704_, new_n701_, new_n703_ );
not g597 ( new_n705_, new_n704_ );
and g598 ( new_n706_, new_n700_, new_n705_ );
or g599 ( new_n707_, new_n706_, keyIn_0_52 );
not g600 ( new_n708_, keyIn_0_52 );
or g601 ( new_n709_, new_n698_, new_n697_ );
or g602 ( new_n710_, new_n695_, keyIn_0_47 );
and g603 ( new_n711_, new_n709_, new_n710_ );
or g604 ( new_n712_, new_n711_, new_n704_ );
or g605 ( new_n713_, new_n712_, new_n708_ );
and g606 ( new_n714_, new_n713_, new_n707_ );
not g607 ( new_n715_, keyIn_0_46 );
and g608 ( new_n716_, new_n655_, N27 );
and g609 ( new_n717_, new_n716_, new_n715_ );
or g610 ( new_n718_, new_n660_, new_n481_ );
and g611 ( new_n719_, new_n718_, keyIn_0_46 );
or g612 ( new_n720_, new_n719_, new_n717_ );
and g613 ( new_n721_, N329, N21 );
not g614 ( new_n722_, new_n721_ );
and g615 ( new_n723_, N223, N11 );
not g616 ( new_n724_, new_n723_ );
and g617 ( new_n725_, new_n724_, N17 );
and g618 ( new_n726_, new_n722_, new_n725_ );
and g619 ( new_n727_, new_n720_, new_n726_ );
or g620 ( new_n728_, new_n727_, keyIn_0_51 );
not g621 ( new_n729_, keyIn_0_51 );
or g622 ( new_n730_, new_n718_, keyIn_0_46 );
or g623 ( new_n731_, new_n716_, new_n715_ );
and g624 ( new_n732_, new_n730_, new_n731_ );
not g625 ( new_n733_, new_n726_ );
or g626 ( new_n734_, new_n732_, new_n733_ );
or g627 ( new_n735_, new_n734_, new_n729_ );
and g628 ( new_n736_, new_n735_, new_n728_ );
and g629 ( new_n737_, new_n714_, new_n736_ );
not g630 ( new_n738_, keyIn_0_55 );
not g631 ( new_n739_, keyIn_0_50 );
and g632 ( new_n740_, new_n655_, N79 );
and g633 ( new_n741_, new_n740_, new_n739_ );
or g634 ( new_n742_, new_n660_, new_n501_ );
and g635 ( new_n743_, new_n742_, keyIn_0_50 );
or g636 ( new_n744_, new_n743_, new_n741_ );
and g637 ( new_n745_, N329, N73 );
not g638 ( new_n746_, new_n745_ );
and g639 ( new_n747_, N223, N63 );
not g640 ( new_n748_, new_n747_ );
and g641 ( new_n749_, new_n748_, N69 );
and g642 ( new_n750_, new_n746_, new_n749_ );
and g643 ( new_n751_, new_n744_, new_n750_ );
and g644 ( new_n752_, new_n751_, new_n738_ );
or g645 ( new_n753_, new_n742_, keyIn_0_50 );
or g646 ( new_n754_, new_n740_, new_n739_ );
and g647 ( new_n755_, new_n753_, new_n754_ );
not g648 ( new_n756_, new_n750_ );
or g649 ( new_n757_, new_n755_, new_n756_ );
and g650 ( new_n758_, new_n757_, keyIn_0_55 );
or g651 ( new_n759_, new_n758_, new_n752_ );
and g652 ( new_n760_, new_n655_, N115 );
and g653 ( new_n761_, N329, N112 );
and g654 ( new_n762_, N223, N102 );
or g655 ( new_n763_, new_n762_, new_n183_ );
or g656 ( new_n764_, new_n761_, new_n763_ );
or g657 ( new_n765_, new_n760_, new_n764_ );
and g658 ( new_n766_, new_n655_, N92 );
and g659 ( new_n767_, N329, N86 );
and g660 ( new_n768_, N223, N76 );
or g661 ( new_n769_, new_n768_, new_n204_ );
or g662 ( new_n770_, new_n767_, new_n769_ );
or g663 ( new_n771_, new_n766_, new_n770_ );
and g664 ( new_n772_, new_n655_, N105 );
and g665 ( new_n773_, N329, N99 );
and g666 ( new_n774_, N223, N89 );
or g667 ( new_n775_, new_n774_, new_n110_ );
or g668 ( new_n776_, new_n773_, new_n775_ );
or g669 ( new_n777_, new_n772_, new_n776_ );
and g670 ( new_n778_, new_n771_, new_n777_ );
and g671 ( new_n779_, new_n778_, new_n765_ );
and g672 ( new_n780_, new_n759_, new_n779_ );
and g673 ( new_n781_, new_n737_, new_n780_ );
and g674 ( new_n782_, new_n781_, new_n694_ );
not g675 ( new_n783_, new_n782_ );
and g676 ( new_n784_, new_n783_, keyIn_0_56 );
not g677 ( new_n785_, keyIn_0_56 );
and g678 ( new_n786_, new_n782_, new_n785_ );
or g679 ( new_n787_, new_n784_, new_n786_ );
and g680 ( new_n788_, new_n655_, N14 );
and g681 ( new_n789_, N329, N8 );
not g682 ( new_n790_, N4 );
and g683 ( new_n791_, N223, N1 );
or g684 ( new_n792_, new_n791_, new_n790_ );
or g685 ( new_n793_, new_n789_, new_n792_ );
or g686 ( new_n794_, new_n788_, new_n793_ );
and g687 ( new_n795_, new_n787_, new_n794_ );
and g688 ( new_n796_, new_n795_, new_n647_ );
or g689 ( new_n797_, new_n782_, new_n785_ );
not g690 ( new_n798_, new_n786_ );
and g691 ( new_n799_, new_n798_, new_n797_ );
not g692 ( new_n800_, new_n794_ );
or g693 ( new_n801_, new_n799_, new_n800_ );
and g694 ( new_n802_, new_n801_, keyIn_0_58 );
or g695 ( N421, new_n802_, new_n796_ );
not g696 ( new_n804_, keyIn_0_61 );
and g697 ( new_n805_, new_n693_, keyIn_0_57 );
not g698 ( new_n806_, new_n805_ );
or g699 ( new_n807_, new_n693_, keyIn_0_57 );
and g700 ( new_n808_, new_n807_, new_n714_ );
and g701 ( new_n809_, new_n808_, new_n806_ );
or g702 ( new_n810_, new_n809_, keyIn_0_59 );
not g703 ( new_n811_, keyIn_0_59 );
and g704 ( new_n812_, new_n712_, new_n708_ );
and g705 ( new_n813_, new_n706_, keyIn_0_52 );
or g706 ( new_n814_, new_n812_, new_n813_ );
not g707 ( new_n815_, keyIn_0_57 );
not g708 ( new_n816_, keyIn_0_53 );
or g709 ( new_n817_, new_n681_, keyIn_0_48 );
or g710 ( new_n818_, new_n679_, new_n678_ );
and g711 ( new_n819_, new_n817_, new_n818_ );
or g712 ( new_n820_, new_n819_, new_n687_ );
and g713 ( new_n821_, new_n820_, new_n816_ );
or g714 ( new_n822_, new_n821_, new_n691_ );
and g715 ( new_n823_, new_n822_, new_n815_ );
or g716 ( new_n824_, new_n823_, new_n814_ );
or g717 ( new_n825_, new_n824_, new_n805_ );
or g718 ( new_n826_, new_n825_, new_n811_ );
and g719 ( new_n827_, new_n810_, new_n826_ );
and g720 ( new_n828_, new_n737_, new_n677_ );
not g721 ( new_n829_, new_n828_ );
or g722 ( new_n830_, new_n827_, new_n829_ );
and g723 ( new_n831_, new_n830_, new_n804_ );
and g724 ( new_n832_, new_n825_, new_n811_ );
and g725 ( new_n833_, new_n809_, keyIn_0_59 );
or g726 ( new_n834_, new_n833_, new_n832_ );
and g727 ( new_n835_, new_n834_, new_n828_ );
and g728 ( new_n836_, new_n835_, keyIn_0_61 );
or g729 ( N430, new_n831_, new_n836_ );
or g730 ( new_n838_, new_n675_, new_n671_ );
or g731 ( new_n839_, new_n669_, keyIn_0_54 );
and g732 ( new_n840_, new_n838_, new_n839_ );
or g733 ( new_n841_, new_n822_, new_n840_ );
or g734 ( new_n842_, new_n814_, new_n759_ );
or g735 ( new_n843_, new_n842_, new_n841_ );
or g736 ( new_n844_, new_n843_, keyIn_0_60 );
not g737 ( new_n845_, keyIn_0_60 );
or g738 ( new_n846_, new_n757_, keyIn_0_55 );
or g739 ( new_n847_, new_n751_, new_n738_ );
and g740 ( new_n848_, new_n846_, new_n847_ );
and g741 ( new_n849_, new_n714_, new_n848_ );
and g742 ( new_n850_, new_n694_, new_n849_ );
or g743 ( new_n851_, new_n850_, new_n845_ );
and g744 ( new_n852_, new_n844_, new_n851_ );
and g745 ( new_n853_, new_n734_, new_n729_ );
and g746 ( new_n854_, new_n727_, keyIn_0_51 );
or g747 ( new_n855_, new_n853_, new_n854_ );
or g748 ( new_n856_, new_n814_, new_n855_ );
not g749 ( new_n857_, new_n771_ );
and g750 ( new_n858_, new_n694_, new_n857_ );
or g751 ( new_n859_, new_n858_, new_n856_ );
or g752 ( new_n860_, new_n852_, new_n859_ );
not g753 ( new_n861_, new_n860_ );
and g754 ( new_n862_, new_n861_, keyIn_0_62 );
not g755 ( new_n863_, keyIn_0_62 );
and g756 ( new_n864_, new_n860_, new_n863_ );
or g757 ( N431, new_n862_, new_n864_ );
not g758 ( new_n866_, keyIn_0_63 );
or g759 ( new_n867_, new_n857_, new_n777_ );
or g760 ( new_n868_, new_n814_, new_n867_ );
or g761 ( new_n869_, new_n868_, new_n822_ );
and g762 ( new_n870_, new_n869_, new_n736_ );
not g763 ( new_n871_, new_n870_ );
or g764 ( new_n872_, new_n852_, new_n871_ );
or g765 ( new_n873_, new_n872_, new_n827_ );
and g766 ( new_n874_, new_n873_, new_n866_ );
and g767 ( new_n875_, new_n850_, new_n845_ );
and g768 ( new_n876_, new_n843_, keyIn_0_60 );
or g769 ( new_n877_, new_n876_, new_n875_ );
and g770 ( new_n878_, new_n877_, new_n870_ );
and g771 ( new_n879_, new_n878_, new_n834_ );
and g772 ( new_n880_, new_n879_, keyIn_0_63 );
or g773 ( N432, new_n874_, new_n880_ );
endmodule