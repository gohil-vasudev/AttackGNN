module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945;

  AND2_X2 U7925 ( .A1(n8726), .A2(n8727), .ZN(n7900) );
  AND2_X2 U7926 ( .A1(n8726), .A2(operation_0_), .ZN(n7899) );
  AND2_X2 U7927 ( .A1(n8727), .A2(operation_1_), .ZN(n7898) );
  AND2_X2 U7928 ( .A1(operation_0_), .A2(operation_1_), .ZN(n7864) );
  INV_X2 U7929 ( .A(b_1_), .ZN(n8731) );
  INV_X2 U7930 ( .A(b_26_), .ZN(n8830) );
  INV_X2 U7931 ( .A(b_3_), .ZN(n8739) );
  INV_X2 U7932 ( .A(b_4_), .ZN(n8743) );
  INV_X2 U7933 ( .A(b_5_), .ZN(n8747) );
  INV_X2 U7934 ( .A(b_8_), .ZN(n8759) );
  INV_X2 U7935 ( .A(b_23_), .ZN(n8818) );
  INV_X2 U7936 ( .A(b_24_), .ZN(n8822) );
  INV_X2 U7937 ( .A(b_25_), .ZN(n8826) );
  INV_X2 U7938 ( .A(b_6_), .ZN(n8751) );
  INV_X2 U7939 ( .A(b_7_), .ZN(n8755) );
  INV_X2 U7940 ( .A(b_2_), .ZN(n8735) );
  INV_X2 U7941 ( .A(b_11_), .ZN(n8771) );
  INV_X2 U7942 ( .A(b_12_), .ZN(n8775) );
  INV_X2 U7943 ( .A(b_13_), .ZN(n8779) );
  INV_X2 U7944 ( .A(b_14_), .ZN(n8783) );
  INV_X2 U7945 ( .A(b_16_), .ZN(n8791) );
  INV_X2 U7946 ( .A(b_17_), .ZN(n8795) );
  INV_X2 U7947 ( .A(b_18_), .ZN(n8799) );
  INV_X2 U7948 ( .A(b_19_), .ZN(n8803) );
  INV_X2 U7949 ( .A(b_20_), .ZN(n8807) );
  INV_X2 U7950 ( .A(b_21_), .ZN(n8811) );
  INV_X2 U7951 ( .A(b_27_), .ZN(n8834) );
  INV_X2 U7952 ( .A(b_9_), .ZN(n8763) );
  INV_X2 U7953 ( .A(b_22_), .ZN(n8814) );
  INV_X2 U7954 ( .A(b_29_), .ZN(n8842) );
  INV_X2 U7955 ( .A(b_15_), .ZN(n8787) );
  INV_X2 U7956 ( .A(b_28_), .ZN(n8838) );
  INV_X2 U7957 ( .A(b_10_), .ZN(n8767) );
  INV_X2 U7958 ( .A(b_0_), .ZN(n9126) );
  INV_X2 U7959 ( .A(a_29_), .ZN(n7954) );
  INV_X2 U7960 ( .A(a_22_), .ZN(n8140) );
  INV_X2 U7961 ( .A(a_23_), .ZN(n8115) );
  INV_X2 U7962 ( .A(a_24_), .ZN(n8090) );
  INV_X2 U7963 ( .A(a_25_), .ZN(n8065) );
  INV_X2 U7964 ( .A(a_26_), .ZN(n8040) );
  INV_X2 U7965 ( .A(a_27_), .ZN(n8015) );
  INV_X2 U7966 ( .A(a_28_), .ZN(n7979) );
  INV_X2 U7967 ( .A(b_30_), .ZN(n7908) );
  OR2_X1 U7968 ( .A1(n7861), .A2(n7862), .ZN(Result_9_) );
  AND2_X1 U7969 ( .A1(n7863), .A2(n7864), .ZN(n7861) );
  XOR2_X1 U7970 ( .A(n7865), .B(n7866), .Z(n7863) );
  AND2_X1 U7971 ( .A1(n7867), .A2(n7868), .ZN(n7866) );
  OR2_X1 U7972 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
  AND2_X1 U7973 ( .A1(n7871), .A2(n7872), .ZN(n7870) );
  INV_X1 U7974 ( .A(n7873), .ZN(n7867) );
  OR2_X1 U7975 ( .A1(n7874), .A2(n7862), .ZN(Result_8_) );
  AND2_X1 U7976 ( .A1(n7875), .A2(n7864), .ZN(n7874) );
  XOR2_X1 U7977 ( .A(n7876), .B(n7877), .Z(n7875) );
  OR2_X1 U7978 ( .A1(n7878), .A2(n7862), .ZN(Result_7_) );
  AND2_X1 U7979 ( .A1(n7864), .A2(n7879), .ZN(n7878) );
  XOR2_X1 U7980 ( .A(n7880), .B(n7881), .Z(n7879) );
  AND2_X1 U7981 ( .A1(n7882), .A2(n7883), .ZN(n7881) );
  OR2_X1 U7982 ( .A1(n7884), .A2(n7885), .ZN(n7883) );
  AND2_X1 U7983 ( .A1(n7886), .A2(n7887), .ZN(n7885) );
  INV_X1 U7984 ( .A(n7888), .ZN(n7882) );
  OR2_X1 U7985 ( .A1(n7889), .A2(n7862), .ZN(Result_6_) );
  AND2_X1 U7986 ( .A1(n7890), .A2(n7864), .ZN(n7889) );
  XOR2_X1 U7987 ( .A(n7891), .B(n7892), .Z(n7890) );
  OR2_X1 U7988 ( .A1(n7893), .A2(n7894), .ZN(Result_63_) );
  AND2_X1 U7989 ( .A1(n7895), .A2(n7864), .ZN(n7894) );
  AND2_X1 U7990 ( .A1(n7896), .A2(n7897), .ZN(n7893) );
  OR3_X1 U7991 ( .A1(n7898), .A2(n7899), .A3(n7900), .ZN(n7897) );
  OR2_X1 U7992 ( .A1(n7901), .A2(n7902), .ZN(n7896) );
  OR3_X1 U7993 ( .A1(n7903), .A2(n7904), .A3(n7905), .ZN(Result_62_) );
  AND3_X1 U7994 ( .A1(a_30_), .A2(n7906), .A3(n7864), .ZN(n7905) );
  OR2_X1 U7995 ( .A1(n7907), .A2(n7902), .ZN(n7906) );
  AND2_X1 U7996 ( .A1(b_31_), .A2(n7908), .ZN(n7907) );
  AND2_X1 U7997 ( .A1(n7909), .A2(n7908), .ZN(n7904) );
  OR2_X1 U7998 ( .A1(n7910), .A2(n7911), .ZN(n7909) );
  AND2_X1 U7999 ( .A1(a_30_), .A2(n7912), .ZN(n7911) );
  AND2_X1 U8000 ( .A1(n7913), .A2(n7914), .ZN(n7910) );
  AND2_X1 U8001 ( .A1(b_30_), .A2(n7915), .ZN(n7903) );
  OR3_X1 U8002 ( .A1(n7916), .A2(n7917), .A3(n7918), .ZN(n7915) );
  AND2_X1 U8003 ( .A1(n7864), .A2(n7919), .ZN(n7918) );
  OR2_X1 U8004 ( .A1(n7901), .A2(n7920), .ZN(n7919) );
  AND2_X1 U8005 ( .A1(n7912), .A2(n7914), .ZN(n7917) );
  OR3_X1 U8006 ( .A1(n7921), .A2(n7922), .A3(n7923), .ZN(n7912) );
  AND2_X1 U8007 ( .A1(n7898), .A2(n7924), .ZN(n7923) );
  AND2_X1 U8008 ( .A1(n7899), .A2(n7925), .ZN(n7922) );
  AND2_X1 U8009 ( .A1(n7900), .A2(n7926), .ZN(n7921) );
  AND2_X1 U8010 ( .A1(a_30_), .A2(n7913), .ZN(n7916) );
  OR3_X1 U8011 ( .A1(n7927), .A2(n7928), .A3(n7929), .ZN(n7913) );
  AND2_X1 U8012 ( .A1(n7898), .A2(n7902), .ZN(n7929) );
  AND2_X1 U8013 ( .A1(n7899), .A2(n7901), .ZN(n7928) );
  AND2_X1 U8014 ( .A1(n7900), .A2(n7895), .ZN(n7927) );
  INV_X1 U8015 ( .A(n7926), .ZN(n7895) );
  OR3_X1 U8016 ( .A1(n7930), .A2(n7931), .A3(n7932), .ZN(Result_61_) );
  AND2_X1 U8017 ( .A1(n7933), .A2(n7864), .ZN(n7932) );
  XOR2_X1 U8018 ( .A(n7934), .B(n7935), .Z(n7933) );
  XOR2_X1 U8019 ( .A(n7936), .B(n7937), .Z(n7935) );
  AND2_X1 U8020 ( .A1(n7938), .A2(n7939), .ZN(n7931) );
  OR3_X1 U8021 ( .A1(n7940), .A2(n7941), .A3(n7942), .ZN(n7939) );
  AND2_X1 U8022 ( .A1(n7898), .A2(n7943), .ZN(n7942) );
  AND2_X1 U8023 ( .A1(n7899), .A2(n7944), .ZN(n7941) );
  AND2_X1 U8024 ( .A1(n7900), .A2(n7945), .ZN(n7940) );
  INV_X1 U8025 ( .A(n7946), .ZN(n7945) );
  INV_X1 U8026 ( .A(n7947), .ZN(n7938) );
  AND2_X1 U8027 ( .A1(n7947), .A2(n7948), .ZN(n7930) );
  OR3_X1 U8028 ( .A1(n7949), .A2(n7950), .A3(n7951), .ZN(n7948) );
  AND2_X1 U8029 ( .A1(n7898), .A2(n7952), .ZN(n7951) );
  INV_X1 U8030 ( .A(n7943), .ZN(n7952) );
  AND2_X1 U8031 ( .A1(n7899), .A2(n7953), .ZN(n7950) );
  INV_X1 U8032 ( .A(n7944), .ZN(n7953) );
  AND2_X1 U8033 ( .A1(n7946), .A2(n7900), .ZN(n7949) );
  XNOR2_X1 U8034 ( .A(n7954), .B(b_29_), .ZN(n7947) );
  OR3_X1 U8035 ( .A1(n7955), .A2(n7956), .A3(n7957), .ZN(Result_60_) );
  AND2_X1 U8036 ( .A1(n7958), .A2(n7864), .ZN(n7957) );
  XNOR2_X1 U8037 ( .A(n7959), .B(n7960), .ZN(n7958) );
  XOR2_X1 U8038 ( .A(n7961), .B(n7962), .Z(n7960) );
  AND2_X1 U8039 ( .A1(n7963), .A2(n7964), .ZN(n7956) );
  OR3_X1 U8040 ( .A1(n7965), .A2(n7966), .A3(n7967), .ZN(n7964) );
  AND2_X1 U8041 ( .A1(n7898), .A2(n7968), .ZN(n7967) );
  AND2_X1 U8042 ( .A1(n7899), .A2(n7969), .ZN(n7966) );
  AND2_X1 U8043 ( .A1(n7970), .A2(n7900), .ZN(n7965) );
  INV_X1 U8044 ( .A(n7971), .ZN(n7970) );
  INV_X1 U8045 ( .A(n7972), .ZN(n7963) );
  AND2_X1 U8046 ( .A1(n7972), .A2(n7973), .ZN(n7955) );
  OR3_X1 U8047 ( .A1(n7974), .A2(n7975), .A3(n7976), .ZN(n7973) );
  AND2_X1 U8048 ( .A1(n7898), .A2(n7977), .ZN(n7976) );
  INV_X1 U8049 ( .A(n7968), .ZN(n7977) );
  AND2_X1 U8050 ( .A1(n7899), .A2(n7978), .ZN(n7975) );
  INV_X1 U8051 ( .A(n7969), .ZN(n7978) );
  AND2_X1 U8052 ( .A1(n7900), .A2(n7971), .ZN(n7974) );
  XNOR2_X1 U8053 ( .A(n7979), .B(b_28_), .ZN(n7972) );
  OR2_X1 U8054 ( .A1(n7980), .A2(n7862), .ZN(Result_5_) );
  AND2_X1 U8055 ( .A1(n7864), .A2(n7981), .ZN(n7980) );
  XOR2_X1 U8056 ( .A(n7982), .B(n7983), .Z(n7981) );
  AND2_X1 U8057 ( .A1(n7984), .A2(n7985), .ZN(n7983) );
  OR2_X1 U8058 ( .A1(n7986), .A2(n7987), .ZN(n7985) );
  AND2_X1 U8059 ( .A1(n7988), .A2(n7989), .ZN(n7987) );
  INV_X1 U8060 ( .A(n7990), .ZN(n7984) );
  OR3_X1 U8061 ( .A1(n7991), .A2(n7992), .A3(n7993), .ZN(Result_59_) );
  AND2_X1 U8062 ( .A1(n7994), .A2(n7864), .ZN(n7993) );
  XNOR2_X1 U8063 ( .A(n7995), .B(n7996), .ZN(n7994) );
  XOR2_X1 U8064 ( .A(n7997), .B(n7998), .Z(n7996) );
  AND2_X1 U8065 ( .A1(n7999), .A2(n8000), .ZN(n7992) );
  OR3_X1 U8066 ( .A1(n8001), .A2(n8002), .A3(n8003), .ZN(n8000) );
  AND2_X1 U8067 ( .A1(n7898), .A2(n8004), .ZN(n8003) );
  AND2_X1 U8068 ( .A1(n7899), .A2(n8005), .ZN(n8002) );
  AND2_X1 U8069 ( .A1(n8006), .A2(n7900), .ZN(n8001) );
  INV_X1 U8070 ( .A(n8007), .ZN(n8006) );
  INV_X1 U8071 ( .A(n8008), .ZN(n7999) );
  AND2_X1 U8072 ( .A1(n8008), .A2(n8009), .ZN(n7991) );
  OR3_X1 U8073 ( .A1(n8010), .A2(n8011), .A3(n8012), .ZN(n8009) );
  AND2_X1 U8074 ( .A1(n7898), .A2(n8013), .ZN(n8012) );
  INV_X1 U8075 ( .A(n8004), .ZN(n8013) );
  AND2_X1 U8076 ( .A1(n7899), .A2(n8014), .ZN(n8011) );
  INV_X1 U8077 ( .A(n8005), .ZN(n8014) );
  AND2_X1 U8078 ( .A1(n7900), .A2(n8007), .ZN(n8010) );
  XNOR2_X1 U8079 ( .A(n8015), .B(b_27_), .ZN(n8008) );
  OR3_X1 U8080 ( .A1(n8016), .A2(n8017), .A3(n8018), .ZN(Result_58_) );
  AND2_X1 U8081 ( .A1(n8019), .A2(n7864), .ZN(n8018) );
  XNOR2_X1 U8082 ( .A(n8020), .B(n8021), .ZN(n8019) );
  XOR2_X1 U8083 ( .A(n8022), .B(n8023), .Z(n8021) );
  AND2_X1 U8084 ( .A1(n8024), .A2(n8025), .ZN(n8017) );
  OR3_X1 U8085 ( .A1(n8026), .A2(n8027), .A3(n8028), .ZN(n8025) );
  AND2_X1 U8086 ( .A1(n7898), .A2(n8029), .ZN(n8028) );
  AND2_X1 U8087 ( .A1(n7899), .A2(n8030), .ZN(n8027) );
  AND2_X1 U8088 ( .A1(n8031), .A2(n7900), .ZN(n8026) );
  INV_X1 U8089 ( .A(n8032), .ZN(n8031) );
  INV_X1 U8090 ( .A(n8033), .ZN(n8024) );
  AND2_X1 U8091 ( .A1(n8033), .A2(n8034), .ZN(n8016) );
  OR3_X1 U8092 ( .A1(n8035), .A2(n8036), .A3(n8037), .ZN(n8034) );
  AND2_X1 U8093 ( .A1(n7898), .A2(n8038), .ZN(n8037) );
  INV_X1 U8094 ( .A(n8029), .ZN(n8038) );
  AND2_X1 U8095 ( .A1(n7899), .A2(n8039), .ZN(n8036) );
  INV_X1 U8096 ( .A(n8030), .ZN(n8039) );
  AND2_X1 U8097 ( .A1(n7900), .A2(n8032), .ZN(n8035) );
  XNOR2_X1 U8098 ( .A(n8040), .B(b_26_), .ZN(n8033) );
  OR3_X1 U8099 ( .A1(n8041), .A2(n8042), .A3(n8043), .ZN(Result_57_) );
  AND2_X1 U8100 ( .A1(n8044), .A2(n7864), .ZN(n8043) );
  XNOR2_X1 U8101 ( .A(n8045), .B(n8046), .ZN(n8044) );
  XOR2_X1 U8102 ( .A(n8047), .B(n8048), .Z(n8046) );
  AND2_X1 U8103 ( .A1(n8049), .A2(n8050), .ZN(n8042) );
  OR3_X1 U8104 ( .A1(n8051), .A2(n8052), .A3(n8053), .ZN(n8050) );
  AND2_X1 U8105 ( .A1(n7898), .A2(n8054), .ZN(n8053) );
  AND2_X1 U8106 ( .A1(n7899), .A2(n8055), .ZN(n8052) );
  AND2_X1 U8107 ( .A1(n8056), .A2(n7900), .ZN(n8051) );
  INV_X1 U8108 ( .A(n8057), .ZN(n8056) );
  INV_X1 U8109 ( .A(n8058), .ZN(n8049) );
  AND2_X1 U8110 ( .A1(n8058), .A2(n8059), .ZN(n8041) );
  OR3_X1 U8111 ( .A1(n8060), .A2(n8061), .A3(n8062), .ZN(n8059) );
  AND2_X1 U8112 ( .A1(n7898), .A2(n8063), .ZN(n8062) );
  INV_X1 U8113 ( .A(n8054), .ZN(n8063) );
  AND2_X1 U8114 ( .A1(n7899), .A2(n8064), .ZN(n8061) );
  INV_X1 U8115 ( .A(n8055), .ZN(n8064) );
  AND2_X1 U8116 ( .A1(n7900), .A2(n8057), .ZN(n8060) );
  XNOR2_X1 U8117 ( .A(n8065), .B(b_25_), .ZN(n8058) );
  OR3_X1 U8118 ( .A1(n8066), .A2(n8067), .A3(n8068), .ZN(Result_56_) );
  AND2_X1 U8119 ( .A1(n8069), .A2(n7864), .ZN(n8068) );
  XNOR2_X1 U8120 ( .A(n8070), .B(n8071), .ZN(n8069) );
  XOR2_X1 U8121 ( .A(n8072), .B(n8073), .Z(n8071) );
  AND2_X1 U8122 ( .A1(n8074), .A2(n8075), .ZN(n8067) );
  OR3_X1 U8123 ( .A1(n8076), .A2(n8077), .A3(n8078), .ZN(n8075) );
  AND2_X1 U8124 ( .A1(n7898), .A2(n8079), .ZN(n8078) );
  AND2_X1 U8125 ( .A1(n7899), .A2(n8080), .ZN(n8077) );
  AND2_X1 U8126 ( .A1(n8081), .A2(n7900), .ZN(n8076) );
  INV_X1 U8127 ( .A(n8082), .ZN(n8081) );
  INV_X1 U8128 ( .A(n8083), .ZN(n8074) );
  AND2_X1 U8129 ( .A1(n8083), .A2(n8084), .ZN(n8066) );
  OR3_X1 U8130 ( .A1(n8085), .A2(n8086), .A3(n8087), .ZN(n8084) );
  AND2_X1 U8131 ( .A1(n7898), .A2(n8088), .ZN(n8087) );
  INV_X1 U8132 ( .A(n8079), .ZN(n8088) );
  AND2_X1 U8133 ( .A1(n7899), .A2(n8089), .ZN(n8086) );
  INV_X1 U8134 ( .A(n8080), .ZN(n8089) );
  AND2_X1 U8135 ( .A1(n7900), .A2(n8082), .ZN(n8085) );
  XNOR2_X1 U8136 ( .A(n8090), .B(b_24_), .ZN(n8083) );
  OR3_X1 U8137 ( .A1(n8091), .A2(n8092), .A3(n8093), .ZN(Result_55_) );
  AND2_X1 U8138 ( .A1(n8094), .A2(n7864), .ZN(n8093) );
  XNOR2_X1 U8139 ( .A(n8095), .B(n8096), .ZN(n8094) );
  XOR2_X1 U8140 ( .A(n8097), .B(n8098), .Z(n8096) );
  AND2_X1 U8141 ( .A1(n8099), .A2(n8100), .ZN(n8092) );
  OR3_X1 U8142 ( .A1(n8101), .A2(n8102), .A3(n8103), .ZN(n8100) );
  AND2_X1 U8143 ( .A1(n7898), .A2(n8104), .ZN(n8103) );
  AND2_X1 U8144 ( .A1(n7899), .A2(n8105), .ZN(n8102) );
  AND2_X1 U8145 ( .A1(n8106), .A2(n7900), .ZN(n8101) );
  INV_X1 U8146 ( .A(n8107), .ZN(n8106) );
  INV_X1 U8147 ( .A(n8108), .ZN(n8099) );
  AND2_X1 U8148 ( .A1(n8108), .A2(n8109), .ZN(n8091) );
  OR3_X1 U8149 ( .A1(n8110), .A2(n8111), .A3(n8112), .ZN(n8109) );
  AND2_X1 U8150 ( .A1(n7898), .A2(n8113), .ZN(n8112) );
  INV_X1 U8151 ( .A(n8104), .ZN(n8113) );
  AND2_X1 U8152 ( .A1(n7899), .A2(n8114), .ZN(n8111) );
  INV_X1 U8153 ( .A(n8105), .ZN(n8114) );
  AND2_X1 U8154 ( .A1(n7900), .A2(n8107), .ZN(n8110) );
  XNOR2_X1 U8155 ( .A(n8115), .B(b_23_), .ZN(n8108) );
  OR3_X1 U8156 ( .A1(n8116), .A2(n8117), .A3(n8118), .ZN(Result_54_) );
  AND2_X1 U8157 ( .A1(n8119), .A2(n7864), .ZN(n8118) );
  XNOR2_X1 U8158 ( .A(n8120), .B(n8121), .ZN(n8119) );
  XOR2_X1 U8159 ( .A(n8122), .B(n8123), .Z(n8121) );
  AND2_X1 U8160 ( .A1(n8124), .A2(n8125), .ZN(n8117) );
  OR3_X1 U8161 ( .A1(n8126), .A2(n8127), .A3(n8128), .ZN(n8125) );
  AND2_X1 U8162 ( .A1(n7898), .A2(n8129), .ZN(n8128) );
  AND2_X1 U8163 ( .A1(n7899), .A2(n8130), .ZN(n8127) );
  AND2_X1 U8164 ( .A1(n8131), .A2(n7900), .ZN(n8126) );
  INV_X1 U8165 ( .A(n8132), .ZN(n8131) );
  INV_X1 U8166 ( .A(n8133), .ZN(n8124) );
  AND2_X1 U8167 ( .A1(n8133), .A2(n8134), .ZN(n8116) );
  OR3_X1 U8168 ( .A1(n8135), .A2(n8136), .A3(n8137), .ZN(n8134) );
  AND2_X1 U8169 ( .A1(n7898), .A2(n8138), .ZN(n8137) );
  INV_X1 U8170 ( .A(n8129), .ZN(n8138) );
  AND2_X1 U8171 ( .A1(n7899), .A2(n8139), .ZN(n8136) );
  INV_X1 U8172 ( .A(n8130), .ZN(n8139) );
  AND2_X1 U8173 ( .A1(n7900), .A2(n8132), .ZN(n8135) );
  XNOR2_X1 U8174 ( .A(n8140), .B(b_22_), .ZN(n8133) );
  OR3_X1 U8175 ( .A1(n8141), .A2(n8142), .A3(n8143), .ZN(Result_53_) );
  AND2_X1 U8176 ( .A1(n8144), .A2(n7864), .ZN(n8143) );
  XNOR2_X1 U8177 ( .A(n8145), .B(n8146), .ZN(n8144) );
  XOR2_X1 U8178 ( .A(n8147), .B(n8148), .Z(n8146) );
  AND2_X1 U8179 ( .A1(n8149), .A2(n8150), .ZN(n8142) );
  OR3_X1 U8180 ( .A1(n8151), .A2(n8152), .A3(n8153), .ZN(n8150) );
  AND2_X1 U8181 ( .A1(n7898), .A2(n8154), .ZN(n8153) );
  INV_X1 U8182 ( .A(n8155), .ZN(n8154) );
  AND2_X1 U8183 ( .A1(n7899), .A2(n8156), .ZN(n8152) );
  INV_X1 U8184 ( .A(n8157), .ZN(n8156) );
  AND2_X1 U8185 ( .A1(n7900), .A2(n8158), .ZN(n8151) );
  AND2_X1 U8186 ( .A1(n8159), .A2(n8160), .ZN(n8141) );
  INV_X1 U8187 ( .A(n8149), .ZN(n8160) );
  AND2_X1 U8188 ( .A1(n8161), .A2(n8162), .ZN(n8149) );
  OR2_X1 U8189 ( .A1(a_21_), .A2(b_21_), .ZN(n8161) );
  OR3_X1 U8190 ( .A1(n8163), .A2(n8164), .A3(n8165), .ZN(n8159) );
  AND2_X1 U8191 ( .A1(n7898), .A2(n8155), .ZN(n8165) );
  AND2_X1 U8192 ( .A1(n7899), .A2(n8157), .ZN(n8164) );
  AND2_X1 U8193 ( .A1(n8166), .A2(n7900), .ZN(n8163) );
  INV_X1 U8194 ( .A(n8158), .ZN(n8166) );
  OR3_X1 U8195 ( .A1(n8167), .A2(n8168), .A3(n8169), .ZN(Result_52_) );
  AND2_X1 U8196 ( .A1(n8170), .A2(n7864), .ZN(n8169) );
  XNOR2_X1 U8197 ( .A(n8171), .B(n8172), .ZN(n8170) );
  XOR2_X1 U8198 ( .A(n8173), .B(n8174), .Z(n8172) );
  AND2_X1 U8199 ( .A1(n8175), .A2(n8176), .ZN(n8168) );
  OR3_X1 U8200 ( .A1(n8177), .A2(n8178), .A3(n8179), .ZN(n8176) );
  AND2_X1 U8201 ( .A1(n7898), .A2(n8180), .ZN(n8179) );
  INV_X1 U8202 ( .A(n8181), .ZN(n8180) );
  AND2_X1 U8203 ( .A1(n7899), .A2(n8182), .ZN(n8178) );
  INV_X1 U8204 ( .A(n8183), .ZN(n8182) );
  AND2_X1 U8205 ( .A1(n7900), .A2(n8184), .ZN(n8177) );
  AND2_X1 U8206 ( .A1(n8185), .A2(n8186), .ZN(n8167) );
  INV_X1 U8207 ( .A(n8175), .ZN(n8186) );
  AND2_X1 U8208 ( .A1(n8187), .A2(n8188), .ZN(n8175) );
  OR2_X1 U8209 ( .A1(a_20_), .A2(b_20_), .ZN(n8187) );
  OR3_X1 U8210 ( .A1(n8189), .A2(n8190), .A3(n8191), .ZN(n8185) );
  AND2_X1 U8211 ( .A1(n7898), .A2(n8181), .ZN(n8191) );
  AND2_X1 U8212 ( .A1(n7899), .A2(n8183), .ZN(n8190) );
  AND2_X1 U8213 ( .A1(n8192), .A2(n7900), .ZN(n8189) );
  INV_X1 U8214 ( .A(n8184), .ZN(n8192) );
  OR3_X1 U8215 ( .A1(n8193), .A2(n8194), .A3(n8195), .ZN(Result_51_) );
  AND2_X1 U8216 ( .A1(n8196), .A2(n7864), .ZN(n8195) );
  XNOR2_X1 U8217 ( .A(n8197), .B(n8198), .ZN(n8196) );
  XOR2_X1 U8218 ( .A(n8199), .B(n8200), .Z(n8198) );
  AND2_X1 U8219 ( .A1(n8201), .A2(n8202), .ZN(n8194) );
  OR3_X1 U8220 ( .A1(n8203), .A2(n8204), .A3(n8205), .ZN(n8202) );
  AND2_X1 U8221 ( .A1(n7898), .A2(n8206), .ZN(n8205) );
  INV_X1 U8222 ( .A(n8207), .ZN(n8206) );
  AND2_X1 U8223 ( .A1(n7899), .A2(n8208), .ZN(n8204) );
  INV_X1 U8224 ( .A(n8209), .ZN(n8208) );
  AND2_X1 U8225 ( .A1(n7900), .A2(n8210), .ZN(n8203) );
  AND2_X1 U8226 ( .A1(n8211), .A2(n8212), .ZN(n8193) );
  INV_X1 U8227 ( .A(n8201), .ZN(n8212) );
  AND2_X1 U8228 ( .A1(n8213), .A2(n8214), .ZN(n8201) );
  OR2_X1 U8229 ( .A1(a_19_), .A2(b_19_), .ZN(n8213) );
  OR3_X1 U8230 ( .A1(n8215), .A2(n8216), .A3(n8217), .ZN(n8211) );
  AND2_X1 U8231 ( .A1(n7898), .A2(n8207), .ZN(n8217) );
  AND2_X1 U8232 ( .A1(n7899), .A2(n8209), .ZN(n8216) );
  AND2_X1 U8233 ( .A1(n8218), .A2(n7900), .ZN(n8215) );
  INV_X1 U8234 ( .A(n8210), .ZN(n8218) );
  OR3_X1 U8235 ( .A1(n8219), .A2(n8220), .A3(n8221), .ZN(Result_50_) );
  AND2_X1 U8236 ( .A1(n8222), .A2(n7864), .ZN(n8221) );
  XNOR2_X1 U8237 ( .A(n8223), .B(n8224), .ZN(n8222) );
  XOR2_X1 U8238 ( .A(n8225), .B(n8226), .Z(n8224) );
  AND2_X1 U8239 ( .A1(n8227), .A2(n8228), .ZN(n8220) );
  OR3_X1 U8240 ( .A1(n8229), .A2(n8230), .A3(n8231), .ZN(n8228) );
  AND2_X1 U8241 ( .A1(n7898), .A2(n8232), .ZN(n8231) );
  INV_X1 U8242 ( .A(n8233), .ZN(n8232) );
  AND2_X1 U8243 ( .A1(n7899), .A2(n8234), .ZN(n8230) );
  INV_X1 U8244 ( .A(n8235), .ZN(n8234) );
  AND2_X1 U8245 ( .A1(n7900), .A2(n8236), .ZN(n8229) );
  AND2_X1 U8246 ( .A1(n8237), .A2(n8238), .ZN(n8219) );
  INV_X1 U8247 ( .A(n8227), .ZN(n8238) );
  AND2_X1 U8248 ( .A1(n8239), .A2(n8240), .ZN(n8227) );
  OR2_X1 U8249 ( .A1(a_18_), .A2(b_18_), .ZN(n8239) );
  OR3_X1 U8250 ( .A1(n8241), .A2(n8242), .A3(n8243), .ZN(n8237) );
  AND2_X1 U8251 ( .A1(n7898), .A2(n8233), .ZN(n8243) );
  AND2_X1 U8252 ( .A1(n7899), .A2(n8235), .ZN(n8242) );
  AND2_X1 U8253 ( .A1(n8244), .A2(n7900), .ZN(n8241) );
  INV_X1 U8254 ( .A(n8236), .ZN(n8244) );
  OR2_X1 U8255 ( .A1(n8245), .A2(n7862), .ZN(Result_4_) );
  AND2_X1 U8256 ( .A1(n8246), .A2(n7864), .ZN(n8245) );
  XOR2_X1 U8257 ( .A(n8247), .B(n8248), .Z(n8246) );
  OR3_X1 U8258 ( .A1(n8249), .A2(n8250), .A3(n8251), .ZN(Result_49_) );
  AND2_X1 U8259 ( .A1(n8252), .A2(n7864), .ZN(n8251) );
  XNOR2_X1 U8260 ( .A(n8253), .B(n8254), .ZN(n8252) );
  XOR2_X1 U8261 ( .A(n8255), .B(n8256), .Z(n8254) );
  AND2_X1 U8262 ( .A1(n8257), .A2(n8258), .ZN(n8250) );
  OR3_X1 U8263 ( .A1(n8259), .A2(n8260), .A3(n8261), .ZN(n8258) );
  AND2_X1 U8264 ( .A1(n7898), .A2(n8262), .ZN(n8261) );
  INV_X1 U8265 ( .A(n8263), .ZN(n8262) );
  AND2_X1 U8266 ( .A1(n7899), .A2(n8264), .ZN(n8260) );
  INV_X1 U8267 ( .A(n8265), .ZN(n8264) );
  AND2_X1 U8268 ( .A1(n7900), .A2(n8266), .ZN(n8259) );
  AND2_X1 U8269 ( .A1(n8267), .A2(n8268), .ZN(n8249) );
  INV_X1 U8270 ( .A(n8257), .ZN(n8268) );
  AND2_X1 U8271 ( .A1(n8269), .A2(n8270), .ZN(n8257) );
  OR2_X1 U8272 ( .A1(a_17_), .A2(b_17_), .ZN(n8269) );
  OR3_X1 U8273 ( .A1(n8271), .A2(n8272), .A3(n8273), .ZN(n8267) );
  AND2_X1 U8274 ( .A1(n7898), .A2(n8263), .ZN(n8273) );
  AND2_X1 U8275 ( .A1(n7899), .A2(n8265), .ZN(n8272) );
  AND2_X1 U8276 ( .A1(n8274), .A2(n7900), .ZN(n8271) );
  INV_X1 U8277 ( .A(n8266), .ZN(n8274) );
  OR3_X1 U8278 ( .A1(n8275), .A2(n8276), .A3(n8277), .ZN(Result_48_) );
  AND2_X1 U8279 ( .A1(n8278), .A2(n7864), .ZN(n8277) );
  XNOR2_X1 U8280 ( .A(n8279), .B(n8280), .ZN(n8278) );
  XOR2_X1 U8281 ( .A(n8281), .B(n8282), .Z(n8280) );
  AND2_X1 U8282 ( .A1(n8283), .A2(n8284), .ZN(n8276) );
  OR3_X1 U8283 ( .A1(n8285), .A2(n8286), .A3(n8287), .ZN(n8284) );
  AND2_X1 U8284 ( .A1(n7898), .A2(n8288), .ZN(n8287) );
  INV_X1 U8285 ( .A(n8289), .ZN(n8288) );
  AND2_X1 U8286 ( .A1(n7899), .A2(n8290), .ZN(n8286) );
  INV_X1 U8287 ( .A(n8291), .ZN(n8290) );
  AND2_X1 U8288 ( .A1(n7900), .A2(n8292), .ZN(n8285) );
  AND2_X1 U8289 ( .A1(n8293), .A2(n8294), .ZN(n8275) );
  INV_X1 U8290 ( .A(n8283), .ZN(n8294) );
  AND2_X1 U8291 ( .A1(n8295), .A2(n8296), .ZN(n8283) );
  OR2_X1 U8292 ( .A1(a_16_), .A2(b_16_), .ZN(n8295) );
  OR3_X1 U8293 ( .A1(n8297), .A2(n8298), .A3(n8299), .ZN(n8293) );
  AND2_X1 U8294 ( .A1(n7898), .A2(n8289), .ZN(n8299) );
  AND2_X1 U8295 ( .A1(n7899), .A2(n8291), .ZN(n8298) );
  AND2_X1 U8296 ( .A1(n8300), .A2(n7900), .ZN(n8297) );
  INV_X1 U8297 ( .A(n8292), .ZN(n8300) );
  OR3_X1 U8298 ( .A1(n8301), .A2(n8302), .A3(n8303), .ZN(Result_47_) );
  AND2_X1 U8299 ( .A1(n8304), .A2(n7864), .ZN(n8303) );
  XNOR2_X1 U8300 ( .A(n8305), .B(n8306), .ZN(n8304) );
  XOR2_X1 U8301 ( .A(n8307), .B(n8308), .Z(n8306) );
  AND2_X1 U8302 ( .A1(n8309), .A2(n8310), .ZN(n8302) );
  OR3_X1 U8303 ( .A1(n8311), .A2(n8312), .A3(n8313), .ZN(n8310) );
  AND2_X1 U8304 ( .A1(n7898), .A2(n8314), .ZN(n8313) );
  INV_X1 U8305 ( .A(n8315), .ZN(n8314) );
  AND2_X1 U8306 ( .A1(n7899), .A2(n8316), .ZN(n8312) );
  INV_X1 U8307 ( .A(n8317), .ZN(n8316) );
  AND2_X1 U8308 ( .A1(n7900), .A2(n8318), .ZN(n8311) );
  AND2_X1 U8309 ( .A1(n8319), .A2(n8320), .ZN(n8301) );
  INV_X1 U8310 ( .A(n8309), .ZN(n8320) );
  AND2_X1 U8311 ( .A1(n8321), .A2(n8322), .ZN(n8309) );
  OR2_X1 U8312 ( .A1(a_15_), .A2(b_15_), .ZN(n8321) );
  OR3_X1 U8313 ( .A1(n8323), .A2(n8324), .A3(n8325), .ZN(n8319) );
  AND2_X1 U8314 ( .A1(n7898), .A2(n8315), .ZN(n8325) );
  AND2_X1 U8315 ( .A1(n7899), .A2(n8317), .ZN(n8324) );
  AND2_X1 U8316 ( .A1(n8326), .A2(n7900), .ZN(n8323) );
  INV_X1 U8317 ( .A(n8318), .ZN(n8326) );
  OR3_X1 U8318 ( .A1(n8327), .A2(n8328), .A3(n8329), .ZN(Result_46_) );
  AND2_X1 U8319 ( .A1(n8330), .A2(n7864), .ZN(n8329) );
  XNOR2_X1 U8320 ( .A(n8331), .B(n8332), .ZN(n8330) );
  XOR2_X1 U8321 ( .A(n8333), .B(n8334), .Z(n8332) );
  AND2_X1 U8322 ( .A1(n8335), .A2(n8336), .ZN(n8328) );
  OR3_X1 U8323 ( .A1(n8337), .A2(n8338), .A3(n8339), .ZN(n8336) );
  AND2_X1 U8324 ( .A1(n7898), .A2(n8340), .ZN(n8339) );
  INV_X1 U8325 ( .A(n8341), .ZN(n8340) );
  AND2_X1 U8326 ( .A1(n7899), .A2(n8342), .ZN(n8338) );
  INV_X1 U8327 ( .A(n8343), .ZN(n8342) );
  AND2_X1 U8328 ( .A1(n7900), .A2(n8344), .ZN(n8337) );
  AND2_X1 U8329 ( .A1(n8345), .A2(n8346), .ZN(n8327) );
  INV_X1 U8330 ( .A(n8335), .ZN(n8346) );
  AND2_X1 U8331 ( .A1(n8347), .A2(n8348), .ZN(n8335) );
  OR2_X1 U8332 ( .A1(a_14_), .A2(b_14_), .ZN(n8347) );
  OR3_X1 U8333 ( .A1(n8349), .A2(n8350), .A3(n8351), .ZN(n8345) );
  AND2_X1 U8334 ( .A1(n7898), .A2(n8341), .ZN(n8351) );
  AND2_X1 U8335 ( .A1(n7899), .A2(n8343), .ZN(n8350) );
  AND2_X1 U8336 ( .A1(n8352), .A2(n7900), .ZN(n8349) );
  INV_X1 U8337 ( .A(n8344), .ZN(n8352) );
  OR3_X1 U8338 ( .A1(n8353), .A2(n8354), .A3(n8355), .ZN(Result_45_) );
  AND2_X1 U8339 ( .A1(n8356), .A2(n7864), .ZN(n8355) );
  XNOR2_X1 U8340 ( .A(n8357), .B(n8358), .ZN(n8356) );
  XOR2_X1 U8341 ( .A(n8359), .B(n8360), .Z(n8358) );
  AND2_X1 U8342 ( .A1(n8361), .A2(n8362), .ZN(n8354) );
  OR3_X1 U8343 ( .A1(n8363), .A2(n8364), .A3(n8365), .ZN(n8362) );
  AND2_X1 U8344 ( .A1(n7898), .A2(n8366), .ZN(n8365) );
  INV_X1 U8345 ( .A(n8367), .ZN(n8366) );
  AND2_X1 U8346 ( .A1(n7899), .A2(n8368), .ZN(n8364) );
  INV_X1 U8347 ( .A(n8369), .ZN(n8368) );
  AND2_X1 U8348 ( .A1(n7900), .A2(n8370), .ZN(n8363) );
  AND2_X1 U8349 ( .A1(n8371), .A2(n8372), .ZN(n8353) );
  INV_X1 U8350 ( .A(n8361), .ZN(n8372) );
  AND2_X1 U8351 ( .A1(n8373), .A2(n8374), .ZN(n8361) );
  OR2_X1 U8352 ( .A1(a_13_), .A2(b_13_), .ZN(n8373) );
  OR3_X1 U8353 ( .A1(n8375), .A2(n8376), .A3(n8377), .ZN(n8371) );
  AND2_X1 U8354 ( .A1(n7898), .A2(n8367), .ZN(n8377) );
  AND2_X1 U8355 ( .A1(n7899), .A2(n8369), .ZN(n8376) );
  AND2_X1 U8356 ( .A1(n8378), .A2(n7900), .ZN(n8375) );
  INV_X1 U8357 ( .A(n8370), .ZN(n8378) );
  OR3_X1 U8358 ( .A1(n8379), .A2(n8380), .A3(n8381), .ZN(Result_44_) );
  AND2_X1 U8359 ( .A1(n8382), .A2(n7864), .ZN(n8381) );
  XNOR2_X1 U8360 ( .A(n8383), .B(n8384), .ZN(n8382) );
  XOR2_X1 U8361 ( .A(n8385), .B(n8386), .Z(n8384) );
  AND2_X1 U8362 ( .A1(n8387), .A2(n8388), .ZN(n8380) );
  OR3_X1 U8363 ( .A1(n8389), .A2(n8390), .A3(n8391), .ZN(n8388) );
  AND2_X1 U8364 ( .A1(n7898), .A2(n8392), .ZN(n8391) );
  INV_X1 U8365 ( .A(n8393), .ZN(n8392) );
  AND2_X1 U8366 ( .A1(n7899), .A2(n8394), .ZN(n8390) );
  INV_X1 U8367 ( .A(n8395), .ZN(n8394) );
  AND2_X1 U8368 ( .A1(n7900), .A2(n8396), .ZN(n8389) );
  AND2_X1 U8369 ( .A1(n8397), .A2(n8398), .ZN(n8379) );
  INV_X1 U8370 ( .A(n8387), .ZN(n8398) );
  AND2_X1 U8371 ( .A1(n8399), .A2(n8400), .ZN(n8387) );
  OR2_X1 U8372 ( .A1(a_12_), .A2(b_12_), .ZN(n8399) );
  OR3_X1 U8373 ( .A1(n8401), .A2(n8402), .A3(n8403), .ZN(n8397) );
  AND2_X1 U8374 ( .A1(n7898), .A2(n8393), .ZN(n8403) );
  AND2_X1 U8375 ( .A1(n7899), .A2(n8395), .ZN(n8402) );
  AND2_X1 U8376 ( .A1(n8404), .A2(n7900), .ZN(n8401) );
  INV_X1 U8377 ( .A(n8396), .ZN(n8404) );
  OR3_X1 U8378 ( .A1(n8405), .A2(n8406), .A3(n8407), .ZN(Result_43_) );
  AND2_X1 U8379 ( .A1(n8408), .A2(n7864), .ZN(n8407) );
  XNOR2_X1 U8380 ( .A(n8409), .B(n8410), .ZN(n8408) );
  XOR2_X1 U8381 ( .A(n8411), .B(n8412), .Z(n8410) );
  AND2_X1 U8382 ( .A1(n8413), .A2(n8414), .ZN(n8406) );
  OR3_X1 U8383 ( .A1(n8415), .A2(n8416), .A3(n8417), .ZN(n8414) );
  AND2_X1 U8384 ( .A1(n7898), .A2(n8418), .ZN(n8417) );
  INV_X1 U8385 ( .A(n8419), .ZN(n8418) );
  AND2_X1 U8386 ( .A1(n7899), .A2(n8420), .ZN(n8416) );
  INV_X1 U8387 ( .A(n8421), .ZN(n8420) );
  AND2_X1 U8388 ( .A1(n7900), .A2(n8422), .ZN(n8415) );
  AND2_X1 U8389 ( .A1(n8423), .A2(n8424), .ZN(n8405) );
  INV_X1 U8390 ( .A(n8413), .ZN(n8424) );
  AND2_X1 U8391 ( .A1(n8425), .A2(n8426), .ZN(n8413) );
  OR2_X1 U8392 ( .A1(a_11_), .A2(b_11_), .ZN(n8425) );
  OR3_X1 U8393 ( .A1(n8427), .A2(n8428), .A3(n8429), .ZN(n8423) );
  AND2_X1 U8394 ( .A1(n7898), .A2(n8419), .ZN(n8429) );
  AND2_X1 U8395 ( .A1(n7899), .A2(n8421), .ZN(n8428) );
  AND2_X1 U8396 ( .A1(n8430), .A2(n7900), .ZN(n8427) );
  INV_X1 U8397 ( .A(n8422), .ZN(n8430) );
  OR3_X1 U8398 ( .A1(n8431), .A2(n8432), .A3(n8433), .ZN(Result_42_) );
  AND2_X1 U8399 ( .A1(n8434), .A2(n7864), .ZN(n8433) );
  XNOR2_X1 U8400 ( .A(n8435), .B(n8436), .ZN(n8434) );
  XOR2_X1 U8401 ( .A(n8437), .B(n8438), .Z(n8436) );
  AND2_X1 U8402 ( .A1(n8439), .A2(n8440), .ZN(n8432) );
  OR3_X1 U8403 ( .A1(n8441), .A2(n8442), .A3(n8443), .ZN(n8440) );
  AND2_X1 U8404 ( .A1(n7898), .A2(n8444), .ZN(n8443) );
  INV_X1 U8405 ( .A(n8445), .ZN(n8444) );
  AND2_X1 U8406 ( .A1(n7899), .A2(n8446), .ZN(n8442) );
  INV_X1 U8407 ( .A(n8447), .ZN(n8446) );
  AND2_X1 U8408 ( .A1(n7900), .A2(n8448), .ZN(n8441) );
  AND2_X1 U8409 ( .A1(n8449), .A2(n8450), .ZN(n8431) );
  INV_X1 U8410 ( .A(n8439), .ZN(n8450) );
  AND2_X1 U8411 ( .A1(n8451), .A2(n8452), .ZN(n8439) );
  OR2_X1 U8412 ( .A1(a_10_), .A2(b_10_), .ZN(n8451) );
  OR3_X1 U8413 ( .A1(n8453), .A2(n8454), .A3(n8455), .ZN(n8449) );
  AND2_X1 U8414 ( .A1(n7898), .A2(n8445), .ZN(n8455) );
  AND2_X1 U8415 ( .A1(n7899), .A2(n8447), .ZN(n8454) );
  AND2_X1 U8416 ( .A1(n8456), .A2(n7900), .ZN(n8453) );
  INV_X1 U8417 ( .A(n8448), .ZN(n8456) );
  OR3_X1 U8418 ( .A1(n8457), .A2(n8458), .A3(n8459), .ZN(Result_41_) );
  AND2_X1 U8419 ( .A1(n8460), .A2(n7864), .ZN(n8459) );
  XNOR2_X1 U8420 ( .A(n8461), .B(n8462), .ZN(n8460) );
  XOR2_X1 U8421 ( .A(n8463), .B(n8464), .Z(n8462) );
  AND2_X1 U8422 ( .A1(n8465), .A2(n8466), .ZN(n8458) );
  OR3_X1 U8423 ( .A1(n8467), .A2(n8468), .A3(n8469), .ZN(n8466) );
  AND2_X1 U8424 ( .A1(n7898), .A2(n8470), .ZN(n8469) );
  INV_X1 U8425 ( .A(n8471), .ZN(n8470) );
  AND2_X1 U8426 ( .A1(n7899), .A2(n8472), .ZN(n8468) );
  INV_X1 U8427 ( .A(n8473), .ZN(n8472) );
  AND2_X1 U8428 ( .A1(n7900), .A2(n8474), .ZN(n8467) );
  AND2_X1 U8429 ( .A1(n8475), .A2(n8476), .ZN(n8457) );
  INV_X1 U8430 ( .A(n8465), .ZN(n8476) );
  AND2_X1 U8431 ( .A1(n8477), .A2(n8478), .ZN(n8465) );
  OR2_X1 U8432 ( .A1(a_9_), .A2(b_9_), .ZN(n8477) );
  OR3_X1 U8433 ( .A1(n8479), .A2(n8480), .A3(n8481), .ZN(n8475) );
  AND2_X1 U8434 ( .A1(n7898), .A2(n8471), .ZN(n8481) );
  AND2_X1 U8435 ( .A1(n7899), .A2(n8473), .ZN(n8480) );
  AND2_X1 U8436 ( .A1(n8482), .A2(n7900), .ZN(n8479) );
  INV_X1 U8437 ( .A(n8474), .ZN(n8482) );
  OR3_X1 U8438 ( .A1(n8483), .A2(n8484), .A3(n8485), .ZN(Result_40_) );
  AND2_X1 U8439 ( .A1(n8486), .A2(n7864), .ZN(n8485) );
  XNOR2_X1 U8440 ( .A(n8487), .B(n8488), .ZN(n8486) );
  XOR2_X1 U8441 ( .A(n8489), .B(n8490), .Z(n8488) );
  AND2_X1 U8442 ( .A1(n8491), .A2(n8492), .ZN(n8484) );
  OR3_X1 U8443 ( .A1(n8493), .A2(n8494), .A3(n8495), .ZN(n8492) );
  AND2_X1 U8444 ( .A1(n7898), .A2(n8496), .ZN(n8495) );
  INV_X1 U8445 ( .A(n8497), .ZN(n8496) );
  AND2_X1 U8446 ( .A1(n7899), .A2(n8498), .ZN(n8494) );
  INV_X1 U8447 ( .A(n8499), .ZN(n8498) );
  AND2_X1 U8448 ( .A1(n7900), .A2(n8500), .ZN(n8493) );
  AND2_X1 U8449 ( .A1(n8501), .A2(n8502), .ZN(n8483) );
  INV_X1 U8450 ( .A(n8491), .ZN(n8502) );
  AND2_X1 U8451 ( .A1(n8503), .A2(n8504), .ZN(n8491) );
  OR2_X1 U8452 ( .A1(a_8_), .A2(b_8_), .ZN(n8503) );
  OR3_X1 U8453 ( .A1(n8505), .A2(n8506), .A3(n8507), .ZN(n8501) );
  AND2_X1 U8454 ( .A1(n7898), .A2(n8497), .ZN(n8507) );
  AND2_X1 U8455 ( .A1(n7899), .A2(n8499), .ZN(n8506) );
  AND2_X1 U8456 ( .A1(n8508), .A2(n7900), .ZN(n8505) );
  INV_X1 U8457 ( .A(n8500), .ZN(n8508) );
  OR2_X1 U8458 ( .A1(n8509), .A2(n7862), .ZN(Result_3_) );
  AND2_X1 U8459 ( .A1(n7864), .A2(n8510), .ZN(n8509) );
  XOR2_X1 U8460 ( .A(n8511), .B(n8512), .Z(n8510) );
  AND2_X1 U8461 ( .A1(n8513), .A2(n8514), .ZN(n8512) );
  OR2_X1 U8462 ( .A1(n8515), .A2(n8516), .ZN(n8514) );
  AND2_X1 U8463 ( .A1(n8517), .A2(n8518), .ZN(n8516) );
  INV_X1 U8464 ( .A(n8519), .ZN(n8513) );
  OR3_X1 U8465 ( .A1(n8520), .A2(n8521), .A3(n8522), .ZN(Result_39_) );
  AND2_X1 U8466 ( .A1(n8523), .A2(n7864), .ZN(n8522) );
  XNOR2_X1 U8467 ( .A(n8524), .B(n8525), .ZN(n8523) );
  XOR2_X1 U8468 ( .A(n8526), .B(n8527), .Z(n8525) );
  AND2_X1 U8469 ( .A1(n8528), .A2(n8529), .ZN(n8521) );
  OR3_X1 U8470 ( .A1(n8530), .A2(n8531), .A3(n8532), .ZN(n8529) );
  AND2_X1 U8471 ( .A1(n7898), .A2(n8533), .ZN(n8532) );
  INV_X1 U8472 ( .A(n8534), .ZN(n8533) );
  AND2_X1 U8473 ( .A1(n7899), .A2(n8535), .ZN(n8531) );
  INV_X1 U8474 ( .A(n8536), .ZN(n8535) );
  AND2_X1 U8475 ( .A1(n7900), .A2(n8537), .ZN(n8530) );
  AND2_X1 U8476 ( .A1(n8538), .A2(n8539), .ZN(n8520) );
  INV_X1 U8477 ( .A(n8528), .ZN(n8539) );
  AND2_X1 U8478 ( .A1(n8540), .A2(n8541), .ZN(n8528) );
  OR2_X1 U8479 ( .A1(a_7_), .A2(b_7_), .ZN(n8540) );
  OR3_X1 U8480 ( .A1(n8542), .A2(n8543), .A3(n8544), .ZN(n8538) );
  AND2_X1 U8481 ( .A1(n7898), .A2(n8534), .ZN(n8544) );
  AND2_X1 U8482 ( .A1(n7899), .A2(n8536), .ZN(n8543) );
  AND2_X1 U8483 ( .A1(n8545), .A2(n7900), .ZN(n8542) );
  INV_X1 U8484 ( .A(n8537), .ZN(n8545) );
  OR3_X1 U8485 ( .A1(n8546), .A2(n8547), .A3(n8548), .ZN(Result_38_) );
  AND2_X1 U8486 ( .A1(n8549), .A2(n7864), .ZN(n8548) );
  XNOR2_X1 U8487 ( .A(n8550), .B(n8551), .ZN(n8549) );
  XOR2_X1 U8488 ( .A(n8552), .B(n8553), .Z(n8551) );
  AND2_X1 U8489 ( .A1(n8554), .A2(n8555), .ZN(n8547) );
  OR3_X1 U8490 ( .A1(n8556), .A2(n8557), .A3(n8558), .ZN(n8555) );
  AND2_X1 U8491 ( .A1(n7898), .A2(n8559), .ZN(n8558) );
  INV_X1 U8492 ( .A(n8560), .ZN(n8559) );
  AND2_X1 U8493 ( .A1(n7899), .A2(n8561), .ZN(n8557) );
  INV_X1 U8494 ( .A(n8562), .ZN(n8561) );
  AND2_X1 U8495 ( .A1(n7900), .A2(n8563), .ZN(n8556) );
  AND2_X1 U8496 ( .A1(n8564), .A2(n8565), .ZN(n8546) );
  INV_X1 U8497 ( .A(n8554), .ZN(n8565) );
  AND2_X1 U8498 ( .A1(n8566), .A2(n8567), .ZN(n8554) );
  OR2_X1 U8499 ( .A1(a_6_), .A2(b_6_), .ZN(n8566) );
  OR3_X1 U8500 ( .A1(n8568), .A2(n8569), .A3(n8570), .ZN(n8564) );
  AND2_X1 U8501 ( .A1(n7898), .A2(n8560), .ZN(n8570) );
  AND2_X1 U8502 ( .A1(n7899), .A2(n8562), .ZN(n8569) );
  AND2_X1 U8503 ( .A1(n8571), .A2(n7900), .ZN(n8568) );
  INV_X1 U8504 ( .A(n8563), .ZN(n8571) );
  OR3_X1 U8505 ( .A1(n8572), .A2(n8573), .A3(n8574), .ZN(Result_37_) );
  AND2_X1 U8506 ( .A1(n8575), .A2(n7864), .ZN(n8574) );
  XNOR2_X1 U8507 ( .A(n8576), .B(n8577), .ZN(n8575) );
  XOR2_X1 U8508 ( .A(n8578), .B(n8579), .Z(n8577) );
  AND2_X1 U8509 ( .A1(n8580), .A2(n8581), .ZN(n8573) );
  OR3_X1 U8510 ( .A1(n8582), .A2(n8583), .A3(n8584), .ZN(n8581) );
  AND2_X1 U8511 ( .A1(n7898), .A2(n8585), .ZN(n8584) );
  INV_X1 U8512 ( .A(n8586), .ZN(n8585) );
  AND2_X1 U8513 ( .A1(n7899), .A2(n8587), .ZN(n8583) );
  INV_X1 U8514 ( .A(n8588), .ZN(n8587) );
  AND2_X1 U8515 ( .A1(n7900), .A2(n8589), .ZN(n8582) );
  AND2_X1 U8516 ( .A1(n8590), .A2(n8591), .ZN(n8572) );
  INV_X1 U8517 ( .A(n8580), .ZN(n8591) );
  AND2_X1 U8518 ( .A1(n8592), .A2(n8593), .ZN(n8580) );
  OR2_X1 U8519 ( .A1(a_5_), .A2(b_5_), .ZN(n8592) );
  OR3_X1 U8520 ( .A1(n8594), .A2(n8595), .A3(n8596), .ZN(n8590) );
  AND2_X1 U8521 ( .A1(n7898), .A2(n8586), .ZN(n8596) );
  AND2_X1 U8522 ( .A1(n7899), .A2(n8588), .ZN(n8595) );
  AND2_X1 U8523 ( .A1(n8597), .A2(n7900), .ZN(n8594) );
  INV_X1 U8524 ( .A(n8589), .ZN(n8597) );
  OR3_X1 U8525 ( .A1(n8598), .A2(n8599), .A3(n8600), .ZN(Result_36_) );
  AND2_X1 U8526 ( .A1(n8601), .A2(n7864), .ZN(n8600) );
  XNOR2_X1 U8527 ( .A(n8602), .B(n8603), .ZN(n8601) );
  XOR2_X1 U8528 ( .A(n8604), .B(n8605), .Z(n8603) );
  AND2_X1 U8529 ( .A1(n8606), .A2(n8607), .ZN(n8599) );
  OR3_X1 U8530 ( .A1(n8608), .A2(n8609), .A3(n8610), .ZN(n8607) );
  AND2_X1 U8531 ( .A1(n7898), .A2(n8611), .ZN(n8610) );
  INV_X1 U8532 ( .A(n8612), .ZN(n8611) );
  AND2_X1 U8533 ( .A1(n7899), .A2(n8613), .ZN(n8609) );
  INV_X1 U8534 ( .A(n8614), .ZN(n8613) );
  AND2_X1 U8535 ( .A1(n7900), .A2(n8615), .ZN(n8608) );
  AND2_X1 U8536 ( .A1(n8616), .A2(n8617), .ZN(n8598) );
  INV_X1 U8537 ( .A(n8606), .ZN(n8617) );
  AND2_X1 U8538 ( .A1(n8618), .A2(n8619), .ZN(n8606) );
  OR2_X1 U8539 ( .A1(a_4_), .A2(b_4_), .ZN(n8618) );
  OR3_X1 U8540 ( .A1(n8620), .A2(n8621), .A3(n8622), .ZN(n8616) );
  AND2_X1 U8541 ( .A1(n7898), .A2(n8612), .ZN(n8622) );
  AND2_X1 U8542 ( .A1(n7899), .A2(n8614), .ZN(n8621) );
  AND2_X1 U8543 ( .A1(n8623), .A2(n7900), .ZN(n8620) );
  INV_X1 U8544 ( .A(n8615), .ZN(n8623) );
  OR3_X1 U8545 ( .A1(n8624), .A2(n8625), .A3(n8626), .ZN(Result_35_) );
  AND2_X1 U8546 ( .A1(n8627), .A2(n7864), .ZN(n8626) );
  XNOR2_X1 U8547 ( .A(n8628), .B(n8629), .ZN(n8627) );
  XOR2_X1 U8548 ( .A(n8630), .B(n8631), .Z(n8629) );
  AND2_X1 U8549 ( .A1(n8632), .A2(n8633), .ZN(n8625) );
  OR3_X1 U8550 ( .A1(n8634), .A2(n8635), .A3(n8636), .ZN(n8633) );
  AND2_X1 U8551 ( .A1(n7898), .A2(n8637), .ZN(n8636) );
  INV_X1 U8552 ( .A(n8638), .ZN(n8637) );
  AND2_X1 U8553 ( .A1(n7899), .A2(n8639), .ZN(n8635) );
  INV_X1 U8554 ( .A(n8640), .ZN(n8639) );
  AND2_X1 U8555 ( .A1(n7900), .A2(n8641), .ZN(n8634) );
  AND2_X1 U8556 ( .A1(n8642), .A2(n8643), .ZN(n8624) );
  INV_X1 U8557 ( .A(n8632), .ZN(n8643) );
  AND2_X1 U8558 ( .A1(n8644), .A2(n8645), .ZN(n8632) );
  OR2_X1 U8559 ( .A1(a_3_), .A2(b_3_), .ZN(n8644) );
  OR3_X1 U8560 ( .A1(n8646), .A2(n8647), .A3(n8648), .ZN(n8642) );
  AND2_X1 U8561 ( .A1(n7898), .A2(n8638), .ZN(n8648) );
  AND2_X1 U8562 ( .A1(n7899), .A2(n8640), .ZN(n8647) );
  AND2_X1 U8563 ( .A1(n8649), .A2(n7900), .ZN(n8646) );
  INV_X1 U8564 ( .A(n8641), .ZN(n8649) );
  OR3_X1 U8565 ( .A1(n8650), .A2(n8651), .A3(n8652), .ZN(Result_34_) );
  AND2_X1 U8566 ( .A1(n8653), .A2(n7864), .ZN(n8652) );
  XNOR2_X1 U8567 ( .A(n8654), .B(n8655), .ZN(n8653) );
  XOR2_X1 U8568 ( .A(n8656), .B(n8657), .Z(n8655) );
  AND2_X1 U8569 ( .A1(n8658), .A2(n8659), .ZN(n8651) );
  OR3_X1 U8570 ( .A1(n8660), .A2(n8661), .A3(n8662), .ZN(n8659) );
  AND2_X1 U8571 ( .A1(n7898), .A2(n8663), .ZN(n8662) );
  INV_X1 U8572 ( .A(n8664), .ZN(n8663) );
  AND2_X1 U8573 ( .A1(n7899), .A2(n8665), .ZN(n8661) );
  INV_X1 U8574 ( .A(n8666), .ZN(n8665) );
  AND2_X1 U8575 ( .A1(n7900), .A2(n8667), .ZN(n8660) );
  AND2_X1 U8576 ( .A1(n8668), .A2(n8669), .ZN(n8650) );
  INV_X1 U8577 ( .A(n8658), .ZN(n8669) );
  AND2_X1 U8578 ( .A1(n8670), .A2(n8671), .ZN(n8658) );
  OR2_X1 U8579 ( .A1(a_2_), .A2(b_2_), .ZN(n8670) );
  OR3_X1 U8580 ( .A1(n8672), .A2(n8673), .A3(n8674), .ZN(n8668) );
  AND2_X1 U8581 ( .A1(n7898), .A2(n8664), .ZN(n8674) );
  AND2_X1 U8582 ( .A1(n7899), .A2(n8666), .ZN(n8673) );
  AND2_X1 U8583 ( .A1(n8675), .A2(n7900), .ZN(n8672) );
  INV_X1 U8584 ( .A(n8667), .ZN(n8675) );
  OR3_X1 U8585 ( .A1(n8676), .A2(n8677), .A3(n8678), .ZN(Result_33_) );
  AND2_X1 U8586 ( .A1(n8679), .A2(n7864), .ZN(n8678) );
  XNOR2_X1 U8587 ( .A(n8680), .B(n8681), .ZN(n8679) );
  XOR2_X1 U8588 ( .A(n8682), .B(n8683), .Z(n8681) );
  AND2_X1 U8589 ( .A1(n8684), .A2(n8685), .ZN(n8677) );
  OR3_X1 U8590 ( .A1(n8686), .A2(n8687), .A3(n8688), .ZN(n8685) );
  AND2_X1 U8591 ( .A1(n7898), .A2(n8689), .ZN(n8688) );
  INV_X1 U8592 ( .A(n8690), .ZN(n8689) );
  AND2_X1 U8593 ( .A1(n7899), .A2(n8691), .ZN(n8687) );
  INV_X1 U8594 ( .A(n8692), .ZN(n8691) );
  AND2_X1 U8595 ( .A1(n7900), .A2(n8693), .ZN(n8686) );
  AND2_X1 U8596 ( .A1(n8694), .A2(n8695), .ZN(n8676) );
  INV_X1 U8597 ( .A(n8684), .ZN(n8695) );
  AND2_X1 U8598 ( .A1(n8696), .A2(n8697), .ZN(n8684) );
  OR2_X1 U8599 ( .A1(a_1_), .A2(b_1_), .ZN(n8696) );
  OR3_X1 U8600 ( .A1(n8698), .A2(n8699), .A3(n8700), .ZN(n8694) );
  AND2_X1 U8601 ( .A1(n7898), .A2(n8690), .ZN(n8700) );
  AND2_X1 U8602 ( .A1(n7899), .A2(n8692), .ZN(n8699) );
  AND2_X1 U8603 ( .A1(n8701), .A2(n7900), .ZN(n8698) );
  INV_X1 U8604 ( .A(n8693), .ZN(n8701) );
  OR3_X1 U8605 ( .A1(n8702), .A2(n8703), .A3(n8704), .ZN(Result_32_) );
  AND2_X1 U8606 ( .A1(n8705), .A2(n7864), .ZN(n8704) );
  XNOR2_X1 U8607 ( .A(n8706), .B(n8707), .ZN(n8705) );
  XOR2_X1 U8608 ( .A(n8708), .B(n8709), .Z(n8707) );
  AND2_X1 U8609 ( .A1(n8710), .A2(n8711), .ZN(n8703) );
  OR3_X1 U8610 ( .A1(n8712), .A2(n8713), .A3(n8714), .ZN(n8710) );
  AND2_X1 U8611 ( .A1(n8715), .A2(n7898), .ZN(n8714) );
  AND2_X1 U8612 ( .A1(n7899), .A2(n8716), .ZN(n8713) );
  INV_X1 U8613 ( .A(n8717), .ZN(n8716) );
  AND2_X1 U8614 ( .A1(n7900), .A2(n8718), .ZN(n8712) );
  AND2_X1 U8615 ( .A1(n8719), .A2(n8720), .ZN(n8702) );
  OR3_X1 U8616 ( .A1(n8721), .A2(n8722), .A3(n8723), .ZN(n8720) );
  AND2_X1 U8617 ( .A1(n7898), .A2(n8724), .ZN(n8723) );
  AND2_X1 U8618 ( .A1(n7899), .A2(n8717), .ZN(n8722) );
  AND2_X1 U8619 ( .A1(n8725), .A2(n7900), .ZN(n8721) );
  INV_X1 U8620 ( .A(n8718), .ZN(n8725) );
  OR2_X1 U8621 ( .A1(n8728), .A2(n8729), .ZN(n8718) );
  AND2_X1 U8622 ( .A1(n8730), .A2(n8731), .ZN(n8729) );
  AND2_X1 U8623 ( .A1(n8693), .A2(n8697), .ZN(n8728) );
  OR2_X1 U8624 ( .A1(n8732), .A2(n8733), .ZN(n8693) );
  AND2_X1 U8625 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  AND2_X1 U8626 ( .A1(n8667), .A2(n8671), .ZN(n8732) );
  OR2_X1 U8627 ( .A1(n8736), .A2(n8737), .ZN(n8667) );
  AND2_X1 U8628 ( .A1(n8738), .A2(n8739), .ZN(n8737) );
  AND2_X1 U8629 ( .A1(n8641), .A2(n8645), .ZN(n8736) );
  OR2_X1 U8630 ( .A1(n8740), .A2(n8741), .ZN(n8641) );
  AND2_X1 U8631 ( .A1(n8742), .A2(n8743), .ZN(n8741) );
  AND2_X1 U8632 ( .A1(n8615), .A2(n8619), .ZN(n8740) );
  OR2_X1 U8633 ( .A1(n8744), .A2(n8745), .ZN(n8615) );
  AND2_X1 U8634 ( .A1(n8746), .A2(n8747), .ZN(n8745) );
  AND2_X1 U8635 ( .A1(n8589), .A2(n8593), .ZN(n8744) );
  OR2_X1 U8636 ( .A1(n8748), .A2(n8749), .ZN(n8589) );
  AND2_X1 U8637 ( .A1(n8750), .A2(n8751), .ZN(n8749) );
  AND2_X1 U8638 ( .A1(n8563), .A2(n8567), .ZN(n8748) );
  OR2_X1 U8639 ( .A1(n8752), .A2(n8753), .ZN(n8563) );
  AND2_X1 U8640 ( .A1(n8754), .A2(n8755), .ZN(n8753) );
  AND2_X1 U8641 ( .A1(n8537), .A2(n8541), .ZN(n8752) );
  OR2_X1 U8642 ( .A1(n8756), .A2(n8757), .ZN(n8537) );
  AND2_X1 U8643 ( .A1(n8758), .A2(n8759), .ZN(n8757) );
  AND2_X1 U8644 ( .A1(n8500), .A2(n8504), .ZN(n8756) );
  OR2_X1 U8645 ( .A1(n8760), .A2(n8761), .ZN(n8500) );
  AND2_X1 U8646 ( .A1(n8762), .A2(n8763), .ZN(n8761) );
  AND2_X1 U8647 ( .A1(n8474), .A2(n8478), .ZN(n8760) );
  OR2_X1 U8648 ( .A1(n8764), .A2(n8765), .ZN(n8474) );
  AND2_X1 U8649 ( .A1(n8766), .A2(n8767), .ZN(n8765) );
  AND2_X1 U8650 ( .A1(n8448), .A2(n8452), .ZN(n8764) );
  OR2_X1 U8651 ( .A1(n8768), .A2(n8769), .ZN(n8448) );
  AND2_X1 U8652 ( .A1(n8770), .A2(n8771), .ZN(n8769) );
  AND2_X1 U8653 ( .A1(n8422), .A2(n8426), .ZN(n8768) );
  OR2_X1 U8654 ( .A1(n8772), .A2(n8773), .ZN(n8422) );
  AND2_X1 U8655 ( .A1(n8774), .A2(n8775), .ZN(n8773) );
  AND2_X1 U8656 ( .A1(n8396), .A2(n8400), .ZN(n8772) );
  OR2_X1 U8657 ( .A1(n8776), .A2(n8777), .ZN(n8396) );
  AND2_X1 U8658 ( .A1(n8778), .A2(n8779), .ZN(n8777) );
  AND2_X1 U8659 ( .A1(n8370), .A2(n8374), .ZN(n8776) );
  OR2_X1 U8660 ( .A1(n8780), .A2(n8781), .ZN(n8370) );
  AND2_X1 U8661 ( .A1(n8782), .A2(n8783), .ZN(n8781) );
  AND2_X1 U8662 ( .A1(n8344), .A2(n8348), .ZN(n8780) );
  OR2_X1 U8663 ( .A1(n8784), .A2(n8785), .ZN(n8344) );
  AND2_X1 U8664 ( .A1(n8786), .A2(n8787), .ZN(n8785) );
  AND2_X1 U8665 ( .A1(n8318), .A2(n8322), .ZN(n8784) );
  OR2_X1 U8666 ( .A1(n8788), .A2(n8789), .ZN(n8318) );
  AND2_X1 U8667 ( .A1(n8790), .A2(n8791), .ZN(n8789) );
  AND2_X1 U8668 ( .A1(n8292), .A2(n8296), .ZN(n8788) );
  OR2_X1 U8669 ( .A1(n8792), .A2(n8793), .ZN(n8292) );
  AND2_X1 U8670 ( .A1(n8794), .A2(n8795), .ZN(n8793) );
  AND2_X1 U8671 ( .A1(n8266), .A2(n8270), .ZN(n8792) );
  OR2_X1 U8672 ( .A1(n8796), .A2(n8797), .ZN(n8266) );
  AND2_X1 U8673 ( .A1(n8798), .A2(n8799), .ZN(n8797) );
  AND2_X1 U8674 ( .A1(n8236), .A2(n8240), .ZN(n8796) );
  OR2_X1 U8675 ( .A1(n8800), .A2(n8801), .ZN(n8236) );
  AND2_X1 U8676 ( .A1(n8802), .A2(n8803), .ZN(n8801) );
  AND2_X1 U8677 ( .A1(n8210), .A2(n8214), .ZN(n8800) );
  OR2_X1 U8678 ( .A1(n8804), .A2(n8805), .ZN(n8210) );
  AND2_X1 U8679 ( .A1(n8806), .A2(n8807), .ZN(n8805) );
  AND2_X1 U8680 ( .A1(n8184), .A2(n8188), .ZN(n8804) );
  OR2_X1 U8681 ( .A1(n8808), .A2(n8809), .ZN(n8184) );
  AND2_X1 U8682 ( .A1(n8810), .A2(n8811), .ZN(n8809) );
  AND2_X1 U8683 ( .A1(n8158), .A2(n8162), .ZN(n8808) );
  OR2_X1 U8684 ( .A1(n8812), .A2(n8813), .ZN(n8158) );
  AND2_X1 U8685 ( .A1(n8140), .A2(n8814), .ZN(n8813) );
  AND2_X1 U8686 ( .A1(n8132), .A2(n8815), .ZN(n8812) );
  OR2_X1 U8687 ( .A1(n8816), .A2(n8817), .ZN(n8132) );
  AND2_X1 U8688 ( .A1(n8115), .A2(n8818), .ZN(n8817) );
  AND2_X1 U8689 ( .A1(n8107), .A2(n8819), .ZN(n8816) );
  OR2_X1 U8690 ( .A1(n8820), .A2(n8821), .ZN(n8107) );
  AND2_X1 U8691 ( .A1(n8090), .A2(n8822), .ZN(n8821) );
  AND2_X1 U8692 ( .A1(n8082), .A2(n8823), .ZN(n8820) );
  OR2_X1 U8693 ( .A1(n8824), .A2(n8825), .ZN(n8082) );
  AND2_X1 U8694 ( .A1(n8065), .A2(n8826), .ZN(n8825) );
  AND2_X1 U8695 ( .A1(n8057), .A2(n8827), .ZN(n8824) );
  OR2_X1 U8696 ( .A1(n8828), .A2(n8829), .ZN(n8057) );
  AND2_X1 U8697 ( .A1(n8040), .A2(n8830), .ZN(n8829) );
  AND2_X1 U8698 ( .A1(n8032), .A2(n8831), .ZN(n8828) );
  OR2_X1 U8699 ( .A1(n8832), .A2(n8833), .ZN(n8032) );
  AND2_X1 U8700 ( .A1(n8015), .A2(n8834), .ZN(n8833) );
  AND2_X1 U8701 ( .A1(n8007), .A2(n8835), .ZN(n8832) );
  OR2_X1 U8702 ( .A1(n8836), .A2(n8837), .ZN(n8007) );
  AND2_X1 U8703 ( .A1(n7979), .A2(n8838), .ZN(n8837) );
  AND2_X1 U8704 ( .A1(n7971), .A2(n8839), .ZN(n8836) );
  OR2_X1 U8705 ( .A1(n8840), .A2(n8841), .ZN(n7971) );
  AND2_X1 U8706 ( .A1(n7954), .A2(n8842), .ZN(n8841) );
  AND2_X1 U8707 ( .A1(n7946), .A2(n8843), .ZN(n8840) );
  AND2_X1 U8708 ( .A1(n8844), .A2(n8845), .ZN(n7946) );
  OR2_X1 U8709 ( .A1(n7908), .A2(n8846), .ZN(n8845) );
  AND2_X1 U8710 ( .A1(n7914), .A2(n7926), .ZN(n8846) );
  OR2_X1 U8711 ( .A1(n8847), .A2(n8848), .ZN(n7926) );
  INV_X1 U8712 ( .A(n8711), .ZN(n8719) );
  OR2_X1 U8713 ( .A1(n8849), .A2(n8850), .ZN(n8711) );
  INV_X1 U8714 ( .A(n8851), .ZN(n8849) );
  OR2_X1 U8715 ( .A1(n8852), .A2(n7862), .ZN(Result_31_) );
  AND2_X1 U8716 ( .A1(n7864), .A2(n8853), .ZN(n8852) );
  XOR2_X1 U8717 ( .A(n8854), .B(n8855), .Z(n8853) );
  OR2_X1 U8718 ( .A1(n8856), .A2(n7862), .ZN(Result_30_) );
  AND2_X1 U8719 ( .A1(n8857), .A2(n8858), .ZN(n8856) );
  OR2_X1 U8720 ( .A1(n8859), .A2(n8860), .ZN(n8858) );
  AND2_X1 U8721 ( .A1(n8854), .A2(n8855), .ZN(n8859) );
  OR2_X1 U8722 ( .A1(n8861), .A2(n7862), .ZN(Result_2_) );
  AND2_X1 U8723 ( .A1(n8862), .A2(n7864), .ZN(n8861) );
  XOR2_X1 U8724 ( .A(n8863), .B(n8864), .Z(n8862) );
  OR3_X1 U8725 ( .A1(n8865), .A2(n8866), .A3(n7862), .ZN(Result_29_) );
  AND2_X1 U8726 ( .A1(n8867), .A2(n8857), .ZN(n8866) );
  AND2_X1 U8727 ( .A1(n8868), .A2(n7864), .ZN(n8857) );
  AND3_X1 U8728 ( .A1(n7864), .A2(n8869), .A3(n8870), .ZN(n8865) );
  INV_X1 U8729 ( .A(n8867), .ZN(n8870) );
  AND2_X1 U8730 ( .A1(n8871), .A2(n8872), .ZN(n8867) );
  INV_X1 U8731 ( .A(n8873), .ZN(n8872) );
  OR2_X1 U8732 ( .A1(n8874), .A2(n7862), .ZN(Result_28_) );
  AND2_X1 U8733 ( .A1(n8875), .A2(n7864), .ZN(n8874) );
  XNOR2_X1 U8734 ( .A(n8876), .B(n8877), .ZN(n8875) );
  AND2_X1 U8735 ( .A1(n8878), .A2(n8879), .ZN(n8877) );
  INV_X1 U8736 ( .A(n8880), .ZN(n8879) );
  OR2_X1 U8737 ( .A1(n8881), .A2(n7862), .ZN(Result_27_) );
  AND2_X1 U8738 ( .A1(n8882), .A2(n7864), .ZN(n8881) );
  XOR2_X1 U8739 ( .A(n8883), .B(n8884), .Z(n8882) );
  AND2_X1 U8740 ( .A1(n8885), .A2(n8886), .ZN(n8884) );
  INV_X1 U8741 ( .A(n8887), .ZN(n8886) );
  OR2_X1 U8742 ( .A1(n8888), .A2(n7862), .ZN(Result_26_) );
  AND2_X1 U8743 ( .A1(n8889), .A2(n7864), .ZN(n8888) );
  XOR2_X1 U8744 ( .A(n8890), .B(n8891), .Z(n8889) );
  AND2_X1 U8745 ( .A1(n8892), .A2(n8893), .ZN(n8891) );
  INV_X1 U8746 ( .A(n8894), .ZN(n8893) );
  OR2_X1 U8747 ( .A1(n8895), .A2(n7862), .ZN(Result_25_) );
  AND2_X1 U8748 ( .A1(n8896), .A2(n7864), .ZN(n8895) );
  XOR2_X1 U8749 ( .A(n8897), .B(n8898), .Z(n8896) );
  AND2_X1 U8750 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  INV_X1 U8751 ( .A(n8901), .ZN(n8899) );
  OR2_X1 U8752 ( .A1(n8902), .A2(n7862), .ZN(Result_24_) );
  AND2_X1 U8753 ( .A1(n8903), .A2(n7864), .ZN(n8902) );
  XOR2_X1 U8754 ( .A(n8904), .B(n8905), .Z(n8903) );
  AND2_X1 U8755 ( .A1(n8906), .A2(n8907), .ZN(n8905) );
  OR2_X1 U8756 ( .A1(n8908), .A2(n7862), .ZN(Result_23_) );
  AND2_X1 U8757 ( .A1(n8909), .A2(n7864), .ZN(n8908) );
  XOR2_X1 U8758 ( .A(n8910), .B(n8911), .Z(n8909) );
  AND2_X1 U8759 ( .A1(n8912), .A2(n8913), .ZN(n8911) );
  OR2_X1 U8760 ( .A1(n8914), .A2(n7862), .ZN(Result_22_) );
  AND2_X1 U8761 ( .A1(n8915), .A2(n7864), .ZN(n8914) );
  XOR2_X1 U8762 ( .A(n8916), .B(n8917), .Z(n8915) );
  AND2_X1 U8763 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  OR2_X1 U8764 ( .A1(n8920), .A2(n7862), .ZN(Result_21_) );
  AND2_X1 U8765 ( .A1(n8921), .A2(n7864), .ZN(n8920) );
  XOR2_X1 U8766 ( .A(n8922), .B(n8923), .Z(n8921) );
  AND2_X1 U8767 ( .A1(n8924), .A2(n8925), .ZN(n8923) );
  INV_X1 U8768 ( .A(n8926), .ZN(n8924) );
  OR2_X1 U8769 ( .A1(n8927), .A2(n7862), .ZN(Result_20_) );
  AND2_X1 U8770 ( .A1(n8928), .A2(n7864), .ZN(n8927) );
  XOR2_X1 U8771 ( .A(n8929), .B(n8930), .Z(n8928) );
  AND2_X1 U8772 ( .A1(n8931), .A2(n8932), .ZN(n8930) );
  OR2_X1 U8773 ( .A1(n8933), .A2(n7862), .ZN(Result_1_) );
  AND2_X1 U8774 ( .A1(n7864), .A2(n8934), .ZN(n8933) );
  XOR2_X1 U8775 ( .A(n8935), .B(n8936), .Z(n8934) );
  AND2_X1 U8776 ( .A1(n8937), .A2(n8938), .ZN(n8936) );
  OR2_X1 U8777 ( .A1(n8939), .A2(n8940), .ZN(n8938) );
  AND2_X1 U8778 ( .A1(n8941), .A2(n8942), .ZN(n8939) );
  INV_X1 U8779 ( .A(n8943), .ZN(n8937) );
  OR2_X1 U8780 ( .A1(n8944), .A2(n7862), .ZN(Result_19_) );
  AND2_X1 U8781 ( .A1(n8945), .A2(n7864), .ZN(n8944) );
  XOR2_X1 U8782 ( .A(n8946), .B(n8947), .Z(n8945) );
  AND2_X1 U8783 ( .A1(n8948), .A2(n8949), .ZN(n8947) );
  OR2_X1 U8784 ( .A1(n8950), .A2(n7862), .ZN(Result_18_) );
  AND2_X1 U8785 ( .A1(n8951), .A2(n7864), .ZN(n8950) );
  XOR2_X1 U8786 ( .A(n8952), .B(n8953), .Z(n8951) );
  AND2_X1 U8787 ( .A1(n8954), .A2(n8955), .ZN(n8953) );
  OR2_X1 U8788 ( .A1(n8956), .A2(n7862), .ZN(Result_17_) );
  AND2_X1 U8789 ( .A1(n8957), .A2(n7864), .ZN(n8956) );
  XOR2_X1 U8790 ( .A(n8958), .B(n8959), .Z(n8957) );
  AND2_X1 U8791 ( .A1(n8960), .A2(n8961), .ZN(n8959) );
  OR2_X1 U8792 ( .A1(n8962), .A2(n7862), .ZN(Result_16_) );
  AND2_X1 U8793 ( .A1(n8963), .A2(n7864), .ZN(n8962) );
  XOR2_X1 U8794 ( .A(n8964), .B(n8965), .Z(n8963) );
  AND2_X1 U8795 ( .A1(n8966), .A2(n8967), .ZN(n8965) );
  OR2_X1 U8796 ( .A1(n8968), .A2(n7862), .ZN(Result_15_) );
  AND2_X1 U8797 ( .A1(n8969), .A2(n7864), .ZN(n8968) );
  XOR2_X1 U8798 ( .A(n8970), .B(n8971), .Z(n8969) );
  AND2_X1 U8799 ( .A1(n8972), .A2(n8973), .ZN(n8971) );
  OR2_X1 U8800 ( .A1(n8974), .A2(n7862), .ZN(Result_14_) );
  AND2_X1 U8801 ( .A1(n8975), .A2(n7864), .ZN(n8974) );
  XOR2_X1 U8802 ( .A(n8976), .B(n8977), .Z(n8975) );
  AND2_X1 U8803 ( .A1(n8978), .A2(n8979), .ZN(n8977) );
  INV_X1 U8804 ( .A(n8980), .ZN(n8979) );
  OR2_X1 U8805 ( .A1(n8981), .A2(n8982), .ZN(n8978) );
  AND2_X1 U8806 ( .A1(n8983), .A2(n8984), .ZN(n8981) );
  OR2_X1 U8807 ( .A1(n8985), .A2(n7862), .ZN(Result_13_) );
  AND2_X1 U8808 ( .A1(n8986), .A2(n7864), .ZN(n8985) );
  XOR2_X1 U8809 ( .A(n8987), .B(n8988), .Z(n8986) );
  AND2_X1 U8810 ( .A1(n8989), .A2(n8990), .ZN(n8988) );
  INV_X1 U8811 ( .A(n8991), .ZN(n8990) );
  OR2_X1 U8812 ( .A1(n8992), .A2(n8993), .ZN(n8989) );
  AND2_X1 U8813 ( .A1(n8994), .A2(n8995), .ZN(n8992) );
  OR2_X1 U8814 ( .A1(n8996), .A2(n7862), .ZN(Result_12_) );
  AND2_X1 U8815 ( .A1(n8997), .A2(n7864), .ZN(n8996) );
  XOR2_X1 U8816 ( .A(n8998), .B(n8999), .Z(n8997) );
  AND2_X1 U8817 ( .A1(n9000), .A2(n9001), .ZN(n8999) );
  INV_X1 U8818 ( .A(n9002), .ZN(n9001) );
  OR2_X1 U8819 ( .A1(n9003), .A2(n9004), .ZN(n9000) );
  AND2_X1 U8820 ( .A1(n9005), .A2(n9006), .ZN(n9003) );
  OR2_X1 U8821 ( .A1(n9007), .A2(n7862), .ZN(Result_11_) );
  AND2_X1 U8822 ( .A1(n9008), .A2(n7864), .ZN(n9007) );
  XOR2_X1 U8823 ( .A(n9009), .B(n9010), .Z(n9008) );
  AND2_X1 U8824 ( .A1(n9011), .A2(n9012), .ZN(n9010) );
  INV_X1 U8825 ( .A(n9013), .ZN(n9012) );
  OR2_X1 U8826 ( .A1(n9014), .A2(n9015), .ZN(n9011) );
  AND2_X1 U8827 ( .A1(n9016), .A2(n9017), .ZN(n9014) );
  OR2_X1 U8828 ( .A1(n9018), .A2(n7862), .ZN(Result_10_) );
  AND2_X1 U8829 ( .A1(n9019), .A2(n7864), .ZN(n9018) );
  XOR2_X1 U8830 ( .A(n9020), .B(n9021), .Z(n9019) );
  AND2_X1 U8831 ( .A1(n9022), .A2(n9023), .ZN(n9021) );
  INV_X1 U8832 ( .A(n9024), .ZN(n9023) );
  OR2_X1 U8833 ( .A1(n9025), .A2(n9026), .ZN(n9022) );
  AND2_X1 U8834 ( .A1(n9027), .A2(n9028), .ZN(n9025) );
  OR2_X1 U8835 ( .A1(n9029), .A2(n7862), .ZN(Result_0_) );
  OR2_X1 U8836 ( .A1(n9030), .A2(n9031), .ZN(n7862) );
  AND2_X1 U8837 ( .A1(n7898), .A2(n9032), .ZN(n9031) );
  INV_X1 U8838 ( .A(n9033), .ZN(n9032) );
  AND2_X1 U8839 ( .A1(n9034), .A2(n8851), .ZN(n9033) );
  OR2_X1 U8840 ( .A1(n8715), .A2(n8850), .ZN(n9034) );
  INV_X1 U8841 ( .A(n8724), .ZN(n8715) );
  OR2_X1 U8842 ( .A1(n9035), .A2(n9036), .ZN(n8724) );
  AND2_X1 U8843 ( .A1(n8690), .A2(n8730), .ZN(n9036) );
  AND2_X1 U8844 ( .A1(b_1_), .A2(n9037), .ZN(n9035) );
  OR2_X1 U8845 ( .A1(n8730), .A2(n8690), .ZN(n9037) );
  OR2_X1 U8846 ( .A1(n9038), .A2(n9039), .ZN(n8690) );
  AND2_X1 U8847 ( .A1(n8664), .A2(n8734), .ZN(n9039) );
  AND2_X1 U8848 ( .A1(b_2_), .A2(n9040), .ZN(n9038) );
  OR2_X1 U8849 ( .A1(n8734), .A2(n8664), .ZN(n9040) );
  OR2_X1 U8850 ( .A1(n9041), .A2(n9042), .ZN(n8664) );
  AND2_X1 U8851 ( .A1(n8638), .A2(n8738), .ZN(n9042) );
  AND2_X1 U8852 ( .A1(b_3_), .A2(n9043), .ZN(n9041) );
  OR2_X1 U8853 ( .A1(n8738), .A2(n8638), .ZN(n9043) );
  OR2_X1 U8854 ( .A1(n9044), .A2(n9045), .ZN(n8638) );
  AND2_X1 U8855 ( .A1(n8612), .A2(n8742), .ZN(n9045) );
  AND2_X1 U8856 ( .A1(b_4_), .A2(n9046), .ZN(n9044) );
  OR2_X1 U8857 ( .A1(n8742), .A2(n8612), .ZN(n9046) );
  OR2_X1 U8858 ( .A1(n9047), .A2(n9048), .ZN(n8612) );
  AND2_X1 U8859 ( .A1(n8586), .A2(n8746), .ZN(n9048) );
  AND2_X1 U8860 ( .A1(b_5_), .A2(n9049), .ZN(n9047) );
  OR2_X1 U8861 ( .A1(n8746), .A2(n8586), .ZN(n9049) );
  OR2_X1 U8862 ( .A1(n9050), .A2(n9051), .ZN(n8586) );
  AND2_X1 U8863 ( .A1(n8560), .A2(n8750), .ZN(n9051) );
  AND2_X1 U8864 ( .A1(b_6_), .A2(n9052), .ZN(n9050) );
  OR2_X1 U8865 ( .A1(n8750), .A2(n8560), .ZN(n9052) );
  OR2_X1 U8866 ( .A1(n9053), .A2(n9054), .ZN(n8560) );
  AND2_X1 U8867 ( .A1(n8534), .A2(n8754), .ZN(n9054) );
  AND2_X1 U8868 ( .A1(b_7_), .A2(n9055), .ZN(n9053) );
  OR2_X1 U8869 ( .A1(n8754), .A2(n8534), .ZN(n9055) );
  OR2_X1 U8870 ( .A1(n9056), .A2(n9057), .ZN(n8534) );
  AND2_X1 U8871 ( .A1(n8497), .A2(n8758), .ZN(n9057) );
  AND2_X1 U8872 ( .A1(b_8_), .A2(n9058), .ZN(n9056) );
  OR2_X1 U8873 ( .A1(n8758), .A2(n8497), .ZN(n9058) );
  OR2_X1 U8874 ( .A1(n9059), .A2(n9060), .ZN(n8497) );
  AND2_X1 U8875 ( .A1(n8471), .A2(n8762), .ZN(n9060) );
  AND2_X1 U8876 ( .A1(b_9_), .A2(n9061), .ZN(n9059) );
  OR2_X1 U8877 ( .A1(n8762), .A2(n8471), .ZN(n9061) );
  OR2_X1 U8878 ( .A1(n9062), .A2(n9063), .ZN(n8471) );
  AND2_X1 U8879 ( .A1(n8445), .A2(n8766), .ZN(n9063) );
  AND2_X1 U8880 ( .A1(b_10_), .A2(n9064), .ZN(n9062) );
  OR2_X1 U8881 ( .A1(n8766), .A2(n8445), .ZN(n9064) );
  OR2_X1 U8882 ( .A1(n9065), .A2(n9066), .ZN(n8445) );
  AND2_X1 U8883 ( .A1(n8419), .A2(n8770), .ZN(n9066) );
  AND2_X1 U8884 ( .A1(b_11_), .A2(n9067), .ZN(n9065) );
  OR2_X1 U8885 ( .A1(n8770), .A2(n8419), .ZN(n9067) );
  OR2_X1 U8886 ( .A1(n9068), .A2(n9069), .ZN(n8419) );
  AND2_X1 U8887 ( .A1(n8393), .A2(n8774), .ZN(n9069) );
  AND2_X1 U8888 ( .A1(b_12_), .A2(n9070), .ZN(n9068) );
  OR2_X1 U8889 ( .A1(n8774), .A2(n8393), .ZN(n9070) );
  OR2_X1 U8890 ( .A1(n9071), .A2(n9072), .ZN(n8393) );
  AND2_X1 U8891 ( .A1(n8367), .A2(n8778), .ZN(n9072) );
  AND2_X1 U8892 ( .A1(b_13_), .A2(n9073), .ZN(n9071) );
  OR2_X1 U8893 ( .A1(n8778), .A2(n8367), .ZN(n9073) );
  OR2_X1 U8894 ( .A1(n9074), .A2(n9075), .ZN(n8367) );
  AND2_X1 U8895 ( .A1(n8341), .A2(n8782), .ZN(n9075) );
  AND2_X1 U8896 ( .A1(b_14_), .A2(n9076), .ZN(n9074) );
  OR2_X1 U8897 ( .A1(n8782), .A2(n8341), .ZN(n9076) );
  OR2_X1 U8898 ( .A1(n9077), .A2(n9078), .ZN(n8341) );
  AND2_X1 U8899 ( .A1(n8315), .A2(n8786), .ZN(n9078) );
  AND2_X1 U8900 ( .A1(b_15_), .A2(n9079), .ZN(n9077) );
  OR2_X1 U8901 ( .A1(n8786), .A2(n8315), .ZN(n9079) );
  OR2_X1 U8902 ( .A1(n9080), .A2(n9081), .ZN(n8315) );
  AND2_X1 U8903 ( .A1(n8289), .A2(n8790), .ZN(n9081) );
  AND2_X1 U8904 ( .A1(b_16_), .A2(n9082), .ZN(n9080) );
  OR2_X1 U8905 ( .A1(n8790), .A2(n8289), .ZN(n9082) );
  OR2_X1 U8906 ( .A1(n9083), .A2(n9084), .ZN(n8289) );
  AND2_X1 U8907 ( .A1(n8263), .A2(n8794), .ZN(n9084) );
  AND2_X1 U8908 ( .A1(b_17_), .A2(n9085), .ZN(n9083) );
  OR2_X1 U8909 ( .A1(n8794), .A2(n8263), .ZN(n9085) );
  OR2_X1 U8910 ( .A1(n9086), .A2(n9087), .ZN(n8263) );
  AND2_X1 U8911 ( .A1(n8233), .A2(n8798), .ZN(n9087) );
  AND2_X1 U8912 ( .A1(b_18_), .A2(n9088), .ZN(n9086) );
  OR2_X1 U8913 ( .A1(n8798), .A2(n8233), .ZN(n9088) );
  OR2_X1 U8914 ( .A1(n9089), .A2(n9090), .ZN(n8233) );
  AND2_X1 U8915 ( .A1(n8207), .A2(n8802), .ZN(n9090) );
  AND2_X1 U8916 ( .A1(b_19_), .A2(n9091), .ZN(n9089) );
  OR2_X1 U8917 ( .A1(n8802), .A2(n8207), .ZN(n9091) );
  OR2_X1 U8918 ( .A1(n9092), .A2(n9093), .ZN(n8207) );
  AND2_X1 U8919 ( .A1(n8181), .A2(n8806), .ZN(n9093) );
  AND2_X1 U8920 ( .A1(b_20_), .A2(n9094), .ZN(n9092) );
  OR2_X1 U8921 ( .A1(n8806), .A2(n8181), .ZN(n9094) );
  OR2_X1 U8922 ( .A1(n9095), .A2(n9096), .ZN(n8181) );
  AND2_X1 U8923 ( .A1(n8155), .A2(n8810), .ZN(n9096) );
  AND2_X1 U8924 ( .A1(b_21_), .A2(n9097), .ZN(n9095) );
  OR2_X1 U8925 ( .A1(n8810), .A2(n8155), .ZN(n9097) );
  OR2_X1 U8926 ( .A1(n9098), .A2(n9099), .ZN(n8155) );
  AND2_X1 U8927 ( .A1(n8129), .A2(n8140), .ZN(n9099) );
  AND2_X1 U8928 ( .A1(b_22_), .A2(n9100), .ZN(n9098) );
  OR2_X1 U8929 ( .A1(n8140), .A2(n8129), .ZN(n9100) );
  OR2_X1 U8930 ( .A1(n9101), .A2(n9102), .ZN(n8129) );
  AND2_X1 U8931 ( .A1(n8104), .A2(n8115), .ZN(n9102) );
  AND2_X1 U8932 ( .A1(b_23_), .A2(n9103), .ZN(n9101) );
  OR2_X1 U8933 ( .A1(n8115), .A2(n8104), .ZN(n9103) );
  OR2_X1 U8934 ( .A1(n9104), .A2(n9105), .ZN(n8104) );
  AND2_X1 U8935 ( .A1(n8079), .A2(n8090), .ZN(n9105) );
  AND2_X1 U8936 ( .A1(b_24_), .A2(n9106), .ZN(n9104) );
  OR2_X1 U8937 ( .A1(n8090), .A2(n8079), .ZN(n9106) );
  OR2_X1 U8938 ( .A1(n9107), .A2(n9108), .ZN(n8079) );
  AND2_X1 U8939 ( .A1(n8054), .A2(n8065), .ZN(n9108) );
  AND2_X1 U8940 ( .A1(b_25_), .A2(n9109), .ZN(n9107) );
  OR2_X1 U8941 ( .A1(n8065), .A2(n8054), .ZN(n9109) );
  OR2_X1 U8942 ( .A1(n9110), .A2(n9111), .ZN(n8054) );
  AND2_X1 U8943 ( .A1(n8029), .A2(n8040), .ZN(n9111) );
  AND2_X1 U8944 ( .A1(b_26_), .A2(n9112), .ZN(n9110) );
  OR2_X1 U8945 ( .A1(n8040), .A2(n8029), .ZN(n9112) );
  OR2_X1 U8946 ( .A1(n9113), .A2(n9114), .ZN(n8029) );
  AND2_X1 U8947 ( .A1(n8004), .A2(n8015), .ZN(n9114) );
  AND2_X1 U8948 ( .A1(b_27_), .A2(n9115), .ZN(n9113) );
  OR2_X1 U8949 ( .A1(n8015), .A2(n8004), .ZN(n9115) );
  OR2_X1 U8950 ( .A1(n9116), .A2(n9117), .ZN(n8004) );
  AND2_X1 U8951 ( .A1(n7968), .A2(n7979), .ZN(n9117) );
  AND2_X1 U8952 ( .A1(b_28_), .A2(n9118), .ZN(n9116) );
  OR2_X1 U8953 ( .A1(n7979), .A2(n7968), .ZN(n9118) );
  OR2_X1 U8954 ( .A1(n9119), .A2(n9120), .ZN(n7968) );
  AND2_X1 U8955 ( .A1(n7943), .A2(n7954), .ZN(n9120) );
  AND2_X1 U8956 ( .A1(b_29_), .A2(n9121), .ZN(n9119) );
  OR2_X1 U8957 ( .A1(n7954), .A2(n7943), .ZN(n9121) );
  OR2_X1 U8958 ( .A1(n9122), .A2(n9123), .ZN(n7943) );
  AND2_X1 U8959 ( .A1(n7902), .A2(n7914), .ZN(n9123) );
  AND2_X1 U8960 ( .A1(b_30_), .A2(n9124), .ZN(n9122) );
  OR2_X1 U8961 ( .A1(n7902), .A2(n7914), .ZN(n9124) );
  INV_X1 U8962 ( .A(n7924), .ZN(n7902) );
  OR2_X1 U8963 ( .A1(a_31_), .A2(n8848), .ZN(n7924) );
  INV_X1 U8964 ( .A(operation_0_), .ZN(n8727) );
  AND3_X1 U8965 ( .A1(n9125), .A2(n8851), .A3(n7899), .ZN(n9030) );
  INV_X1 U8966 ( .A(operation_1_), .ZN(n8726) );
  OR2_X1 U8967 ( .A1(a_0_), .A2(n9126), .ZN(n8851) );
  OR2_X1 U8968 ( .A1(n8850), .A2(n8717), .ZN(n9125) );
  OR2_X1 U8969 ( .A1(n9127), .A2(n9128), .ZN(n8717) );
  AND2_X1 U8970 ( .A1(a_1_), .A2(n8692), .ZN(n9128) );
  AND2_X1 U8971 ( .A1(n9129), .A2(n8731), .ZN(n9127) );
  OR2_X1 U8972 ( .A1(a_1_), .A2(n8692), .ZN(n9129) );
  OR2_X1 U8973 ( .A1(n9130), .A2(n9131), .ZN(n8692) );
  AND2_X1 U8974 ( .A1(a_2_), .A2(n8666), .ZN(n9131) );
  AND2_X1 U8975 ( .A1(n9132), .A2(n8735), .ZN(n9130) );
  OR2_X1 U8976 ( .A1(a_2_), .A2(n8666), .ZN(n9132) );
  OR2_X1 U8977 ( .A1(n9133), .A2(n9134), .ZN(n8666) );
  AND2_X1 U8978 ( .A1(a_3_), .A2(n8640), .ZN(n9134) );
  AND2_X1 U8979 ( .A1(n9135), .A2(n8739), .ZN(n9133) );
  OR2_X1 U8980 ( .A1(a_3_), .A2(n8640), .ZN(n9135) );
  OR2_X1 U8981 ( .A1(n9136), .A2(n9137), .ZN(n8640) );
  AND2_X1 U8982 ( .A1(a_4_), .A2(n8614), .ZN(n9137) );
  AND2_X1 U8983 ( .A1(n9138), .A2(n8743), .ZN(n9136) );
  OR2_X1 U8984 ( .A1(a_4_), .A2(n8614), .ZN(n9138) );
  OR2_X1 U8985 ( .A1(n9139), .A2(n9140), .ZN(n8614) );
  AND2_X1 U8986 ( .A1(a_5_), .A2(n8588), .ZN(n9140) );
  AND2_X1 U8987 ( .A1(n9141), .A2(n8747), .ZN(n9139) );
  OR2_X1 U8988 ( .A1(a_5_), .A2(n8588), .ZN(n9141) );
  OR2_X1 U8989 ( .A1(n9142), .A2(n9143), .ZN(n8588) );
  AND2_X1 U8990 ( .A1(a_6_), .A2(n8562), .ZN(n9143) );
  AND2_X1 U8991 ( .A1(n9144), .A2(n8751), .ZN(n9142) );
  OR2_X1 U8992 ( .A1(a_6_), .A2(n8562), .ZN(n9144) );
  OR2_X1 U8993 ( .A1(n9145), .A2(n9146), .ZN(n8562) );
  AND2_X1 U8994 ( .A1(a_7_), .A2(n8536), .ZN(n9146) );
  AND2_X1 U8995 ( .A1(n9147), .A2(n8755), .ZN(n9145) );
  OR2_X1 U8996 ( .A1(a_7_), .A2(n8536), .ZN(n9147) );
  OR2_X1 U8997 ( .A1(n9148), .A2(n9149), .ZN(n8536) );
  AND2_X1 U8998 ( .A1(a_8_), .A2(n8499), .ZN(n9149) );
  AND2_X1 U8999 ( .A1(n9150), .A2(n8759), .ZN(n9148) );
  OR2_X1 U9000 ( .A1(a_8_), .A2(n8499), .ZN(n9150) );
  OR2_X1 U9001 ( .A1(n9151), .A2(n9152), .ZN(n8499) );
  AND2_X1 U9002 ( .A1(a_9_), .A2(n8473), .ZN(n9152) );
  AND2_X1 U9003 ( .A1(n9153), .A2(n8763), .ZN(n9151) );
  OR2_X1 U9004 ( .A1(a_9_), .A2(n8473), .ZN(n9153) );
  OR2_X1 U9005 ( .A1(n9154), .A2(n9155), .ZN(n8473) );
  AND2_X1 U9006 ( .A1(a_10_), .A2(n8447), .ZN(n9155) );
  AND2_X1 U9007 ( .A1(n9156), .A2(n8767), .ZN(n9154) );
  OR2_X1 U9008 ( .A1(a_10_), .A2(n8447), .ZN(n9156) );
  OR2_X1 U9009 ( .A1(n9157), .A2(n9158), .ZN(n8447) );
  AND2_X1 U9010 ( .A1(a_11_), .A2(n8421), .ZN(n9158) );
  AND2_X1 U9011 ( .A1(n9159), .A2(n8771), .ZN(n9157) );
  OR2_X1 U9012 ( .A1(a_11_), .A2(n8421), .ZN(n9159) );
  OR2_X1 U9013 ( .A1(n9160), .A2(n9161), .ZN(n8421) );
  AND2_X1 U9014 ( .A1(a_12_), .A2(n8395), .ZN(n9161) );
  AND2_X1 U9015 ( .A1(n9162), .A2(n8775), .ZN(n9160) );
  OR2_X1 U9016 ( .A1(a_12_), .A2(n8395), .ZN(n9162) );
  OR2_X1 U9017 ( .A1(n9163), .A2(n9164), .ZN(n8395) );
  AND2_X1 U9018 ( .A1(a_13_), .A2(n8369), .ZN(n9164) );
  AND2_X1 U9019 ( .A1(n9165), .A2(n8779), .ZN(n9163) );
  OR2_X1 U9020 ( .A1(a_13_), .A2(n8369), .ZN(n9165) );
  OR2_X1 U9021 ( .A1(n9166), .A2(n9167), .ZN(n8369) );
  AND2_X1 U9022 ( .A1(a_14_), .A2(n8343), .ZN(n9167) );
  AND2_X1 U9023 ( .A1(n9168), .A2(n8783), .ZN(n9166) );
  OR2_X1 U9024 ( .A1(a_14_), .A2(n8343), .ZN(n9168) );
  OR2_X1 U9025 ( .A1(n9169), .A2(n9170), .ZN(n8343) );
  AND2_X1 U9026 ( .A1(a_15_), .A2(n8317), .ZN(n9170) );
  AND2_X1 U9027 ( .A1(n9171), .A2(n8787), .ZN(n9169) );
  OR2_X1 U9028 ( .A1(a_15_), .A2(n8317), .ZN(n9171) );
  OR2_X1 U9029 ( .A1(n9172), .A2(n9173), .ZN(n8317) );
  AND2_X1 U9030 ( .A1(a_16_), .A2(n8291), .ZN(n9173) );
  AND2_X1 U9031 ( .A1(n9174), .A2(n8791), .ZN(n9172) );
  OR2_X1 U9032 ( .A1(a_16_), .A2(n8291), .ZN(n9174) );
  OR2_X1 U9033 ( .A1(n9175), .A2(n9176), .ZN(n8291) );
  AND2_X1 U9034 ( .A1(a_17_), .A2(n8265), .ZN(n9176) );
  AND2_X1 U9035 ( .A1(n9177), .A2(n8795), .ZN(n9175) );
  OR2_X1 U9036 ( .A1(a_17_), .A2(n8265), .ZN(n9177) );
  OR2_X1 U9037 ( .A1(n9178), .A2(n9179), .ZN(n8265) );
  AND2_X1 U9038 ( .A1(a_18_), .A2(n8235), .ZN(n9179) );
  AND2_X1 U9039 ( .A1(n9180), .A2(n8799), .ZN(n9178) );
  OR2_X1 U9040 ( .A1(a_18_), .A2(n8235), .ZN(n9180) );
  OR2_X1 U9041 ( .A1(n9181), .A2(n9182), .ZN(n8235) );
  AND2_X1 U9042 ( .A1(a_19_), .A2(n8209), .ZN(n9182) );
  AND2_X1 U9043 ( .A1(n9183), .A2(n8803), .ZN(n9181) );
  OR2_X1 U9044 ( .A1(a_19_), .A2(n8209), .ZN(n9183) );
  OR2_X1 U9045 ( .A1(n9184), .A2(n9185), .ZN(n8209) );
  AND2_X1 U9046 ( .A1(a_20_), .A2(n8183), .ZN(n9185) );
  AND2_X1 U9047 ( .A1(n9186), .A2(n8807), .ZN(n9184) );
  OR2_X1 U9048 ( .A1(a_20_), .A2(n8183), .ZN(n9186) );
  OR2_X1 U9049 ( .A1(n9187), .A2(n9188), .ZN(n8183) );
  AND2_X1 U9050 ( .A1(a_21_), .A2(n8157), .ZN(n9188) );
  AND2_X1 U9051 ( .A1(n9189), .A2(n8811), .ZN(n9187) );
  OR2_X1 U9052 ( .A1(a_21_), .A2(n8157), .ZN(n9189) );
  OR2_X1 U9053 ( .A1(n9190), .A2(n9191), .ZN(n8157) );
  AND2_X1 U9054 ( .A1(a_22_), .A2(n8130), .ZN(n9191) );
  AND2_X1 U9055 ( .A1(n9192), .A2(n8814), .ZN(n9190) );
  OR2_X1 U9056 ( .A1(a_22_), .A2(n8130), .ZN(n9192) );
  OR2_X1 U9057 ( .A1(n9193), .A2(n9194), .ZN(n8130) );
  AND2_X1 U9058 ( .A1(a_23_), .A2(n8105), .ZN(n9194) );
  AND2_X1 U9059 ( .A1(n9195), .A2(n8818), .ZN(n9193) );
  OR2_X1 U9060 ( .A1(a_23_), .A2(n8105), .ZN(n9195) );
  OR2_X1 U9061 ( .A1(n9196), .A2(n9197), .ZN(n8105) );
  AND2_X1 U9062 ( .A1(a_24_), .A2(n8080), .ZN(n9197) );
  AND2_X1 U9063 ( .A1(n9198), .A2(n8822), .ZN(n9196) );
  OR2_X1 U9064 ( .A1(a_24_), .A2(n8080), .ZN(n9198) );
  OR2_X1 U9065 ( .A1(n9199), .A2(n9200), .ZN(n8080) );
  AND2_X1 U9066 ( .A1(a_25_), .A2(n8055), .ZN(n9200) );
  AND2_X1 U9067 ( .A1(n9201), .A2(n8826), .ZN(n9199) );
  OR2_X1 U9068 ( .A1(a_25_), .A2(n8055), .ZN(n9201) );
  OR2_X1 U9069 ( .A1(n9202), .A2(n9203), .ZN(n8055) );
  AND2_X1 U9070 ( .A1(a_26_), .A2(n8030), .ZN(n9203) );
  AND2_X1 U9071 ( .A1(n9204), .A2(n8830), .ZN(n9202) );
  OR2_X1 U9072 ( .A1(a_26_), .A2(n8030), .ZN(n9204) );
  OR2_X1 U9073 ( .A1(n9205), .A2(n9206), .ZN(n8030) );
  AND2_X1 U9074 ( .A1(a_27_), .A2(n8005), .ZN(n9206) );
  AND2_X1 U9075 ( .A1(n9207), .A2(n8834), .ZN(n9205) );
  OR2_X1 U9076 ( .A1(a_27_), .A2(n8005), .ZN(n9207) );
  OR2_X1 U9077 ( .A1(n9208), .A2(n9209), .ZN(n8005) );
  AND2_X1 U9078 ( .A1(a_28_), .A2(n7969), .ZN(n9209) );
  AND2_X1 U9079 ( .A1(n9210), .A2(n8838), .ZN(n9208) );
  OR2_X1 U9080 ( .A1(a_28_), .A2(n7969), .ZN(n9210) );
  OR2_X1 U9081 ( .A1(n9211), .A2(n9212), .ZN(n7969) );
  AND2_X1 U9082 ( .A1(a_29_), .A2(n7944), .ZN(n9212) );
  AND2_X1 U9083 ( .A1(n9213), .A2(n8842), .ZN(n9211) );
  OR2_X1 U9084 ( .A1(a_29_), .A2(n7944), .ZN(n9213) );
  OR2_X1 U9085 ( .A1(n9214), .A2(n9215), .ZN(n7944) );
  AND2_X1 U9086 ( .A1(a_30_), .A2(n7901), .ZN(n9215) );
  AND2_X1 U9087 ( .A1(n9216), .A2(n7908), .ZN(n9214) );
  OR2_X1 U9088 ( .A1(n7901), .A2(a_30_), .ZN(n9216) );
  INV_X1 U9089 ( .A(n7925), .ZN(n7901) );
  OR2_X1 U9090 ( .A1(b_31_), .A2(n8847), .ZN(n7925) );
  AND2_X1 U9091 ( .A1(n9126), .A2(a_0_), .ZN(n8850) );
  AND2_X1 U9092 ( .A1(n7864), .A2(n9217), .ZN(n9029) );
  OR3_X1 U9093 ( .A1(n8943), .A2(n9218), .A3(n9219), .ZN(n9217) );
  AND2_X1 U9094 ( .A1(n9220), .A2(a_0_), .ZN(n9219) );
  INV_X1 U9095 ( .A(n9221), .ZN(n9220) );
  AND2_X1 U9096 ( .A1(n8935), .A2(n8940), .ZN(n9218) );
  AND2_X1 U9097 ( .A1(n8863), .A2(n8864), .ZN(n8935) );
  XOR2_X1 U9098 ( .A(n8942), .B(n8941), .Z(n8864) );
  OR2_X1 U9099 ( .A1(n9222), .A2(n9223), .ZN(n8863) );
  INV_X1 U9100 ( .A(n9224), .ZN(n9223) );
  OR2_X1 U9101 ( .A1(n9225), .A2(n8519), .ZN(n9222) );
  AND3_X1 U9102 ( .A1(n8518), .A2(n8517), .A3(n8515), .ZN(n8519) );
  AND2_X1 U9103 ( .A1(n8511), .A2(n8515), .ZN(n9225) );
  AND2_X1 U9104 ( .A1(n9226), .A2(n9224), .ZN(n8515) );
  OR2_X1 U9105 ( .A1(n9227), .A2(n9228), .ZN(n9224) );
  INV_X1 U9106 ( .A(n9229), .ZN(n9226) );
  AND2_X1 U9107 ( .A1(n9227), .A2(n9228), .ZN(n9229) );
  OR2_X1 U9108 ( .A1(n9230), .A2(n9231), .ZN(n9228) );
  AND2_X1 U9109 ( .A1(n9232), .A2(n9233), .ZN(n9231) );
  AND2_X1 U9110 ( .A1(n9234), .A2(n9235), .ZN(n9230) );
  OR2_X1 U9111 ( .A1(n9233), .A2(n9232), .ZN(n9235) );
  XOR2_X1 U9112 ( .A(n9236), .B(n9237), .Z(n9227) );
  XOR2_X1 U9113 ( .A(n9238), .B(n9239), .Z(n9237) );
  AND2_X1 U9114 ( .A1(n8247), .A2(n8248), .ZN(n8511) );
  XOR2_X1 U9115 ( .A(n8518), .B(n8517), .Z(n8248) );
  INV_X1 U9116 ( .A(n9240), .ZN(n8517) );
  OR2_X1 U9117 ( .A1(n9241), .A2(n9242), .ZN(n9240) );
  AND2_X1 U9118 ( .A1(n9243), .A2(n9244), .ZN(n9242) );
  AND2_X1 U9119 ( .A1(n9245), .A2(n9246), .ZN(n9241) );
  OR2_X1 U9120 ( .A1(n9244), .A2(n9243), .ZN(n9246) );
  XNOR2_X1 U9121 ( .A(n9234), .B(n9247), .ZN(n8518) );
  XOR2_X1 U9122 ( .A(n9233), .B(n9232), .Z(n9247) );
  OR2_X1 U9123 ( .A1(n9248), .A2(n8739), .ZN(n9232) );
  OR2_X1 U9124 ( .A1(n9249), .A2(n9250), .ZN(n9233) );
  AND2_X1 U9125 ( .A1(n9251), .A2(n9252), .ZN(n9250) );
  AND2_X1 U9126 ( .A1(n9253), .A2(n9254), .ZN(n9249) );
  OR2_X1 U9127 ( .A1(n9252), .A2(n9251), .ZN(n9254) );
  XOR2_X1 U9128 ( .A(n9255), .B(n9256), .Z(n9234) );
  XOR2_X1 U9129 ( .A(n9257), .B(n9258), .Z(n9256) );
  OR2_X1 U9130 ( .A1(n9259), .A2(n9260), .ZN(n8247) );
  INV_X1 U9131 ( .A(n9261), .ZN(n9260) );
  OR2_X1 U9132 ( .A1(n9262), .A2(n7990), .ZN(n9259) );
  AND3_X1 U9133 ( .A1(n7989), .A2(n7988), .A3(n7986), .ZN(n7990) );
  AND2_X1 U9134 ( .A1(n7982), .A2(n7986), .ZN(n9262) );
  AND2_X1 U9135 ( .A1(n9263), .A2(n9261), .ZN(n7986) );
  OR2_X1 U9136 ( .A1(n9264), .A2(n9265), .ZN(n9261) );
  INV_X1 U9137 ( .A(n9266), .ZN(n9263) );
  AND2_X1 U9138 ( .A1(n9264), .A2(n9265), .ZN(n9266) );
  OR2_X1 U9139 ( .A1(n9267), .A2(n9268), .ZN(n9265) );
  AND2_X1 U9140 ( .A1(n9269), .A2(n9270), .ZN(n9268) );
  AND2_X1 U9141 ( .A1(n9271), .A2(n9272), .ZN(n9267) );
  OR2_X1 U9142 ( .A1(n9270), .A2(n9269), .ZN(n9272) );
  XOR2_X1 U9143 ( .A(n9245), .B(n9273), .Z(n9264) );
  XOR2_X1 U9144 ( .A(n9244), .B(n9243), .Z(n9273) );
  OR2_X1 U9145 ( .A1(n9248), .A2(n8743), .ZN(n9243) );
  OR2_X1 U9146 ( .A1(n9274), .A2(n9275), .ZN(n9244) );
  AND2_X1 U9147 ( .A1(n9276), .A2(n9277), .ZN(n9275) );
  AND2_X1 U9148 ( .A1(n9278), .A2(n9279), .ZN(n9274) );
  OR2_X1 U9149 ( .A1(n9277), .A2(n9276), .ZN(n9279) );
  XOR2_X1 U9150 ( .A(n9253), .B(n9280), .Z(n9245) );
  XOR2_X1 U9151 ( .A(n9252), .B(n9251), .Z(n9280) );
  OR2_X1 U9152 ( .A1(n8730), .A2(n8739), .ZN(n9251) );
  OR2_X1 U9153 ( .A1(n9281), .A2(n9282), .ZN(n9252) );
  AND2_X1 U9154 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  AND2_X1 U9155 ( .A1(n9285), .A2(n9286), .ZN(n9281) );
  OR2_X1 U9156 ( .A1(n9284), .A2(n9283), .ZN(n9286) );
  XOR2_X1 U9157 ( .A(n9287), .B(n9288), .Z(n9253) );
  XOR2_X1 U9158 ( .A(n9289), .B(n8671), .Z(n9288) );
  AND2_X1 U9159 ( .A1(n7891), .A2(n7892), .ZN(n7982) );
  XOR2_X1 U9160 ( .A(n7989), .B(n7988), .Z(n7892) );
  INV_X1 U9161 ( .A(n9290), .ZN(n7988) );
  OR2_X1 U9162 ( .A1(n9291), .A2(n9292), .ZN(n9290) );
  AND2_X1 U9163 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  AND2_X1 U9164 ( .A1(n9295), .A2(n9296), .ZN(n9291) );
  OR2_X1 U9165 ( .A1(n9294), .A2(n9293), .ZN(n9296) );
  XNOR2_X1 U9166 ( .A(n9271), .B(n9297), .ZN(n7989) );
  XOR2_X1 U9167 ( .A(n9270), .B(n9269), .Z(n9297) );
  OR2_X1 U9168 ( .A1(n9248), .A2(n8747), .ZN(n9269) );
  OR2_X1 U9169 ( .A1(n9298), .A2(n9299), .ZN(n9270) );
  AND2_X1 U9170 ( .A1(n9300), .A2(n9301), .ZN(n9299) );
  AND2_X1 U9171 ( .A1(n9302), .A2(n9303), .ZN(n9298) );
  OR2_X1 U9172 ( .A1(n9301), .A2(n9300), .ZN(n9303) );
  XOR2_X1 U9173 ( .A(n9278), .B(n9304), .Z(n9271) );
  XOR2_X1 U9174 ( .A(n9277), .B(n9276), .Z(n9304) );
  OR2_X1 U9175 ( .A1(n8730), .A2(n8743), .ZN(n9276) );
  OR2_X1 U9176 ( .A1(n9305), .A2(n9306), .ZN(n9277) );
  AND2_X1 U9177 ( .A1(n9307), .A2(n9308), .ZN(n9306) );
  AND2_X1 U9178 ( .A1(n9309), .A2(n9310), .ZN(n9305) );
  OR2_X1 U9179 ( .A1(n9308), .A2(n9307), .ZN(n9310) );
  XOR2_X1 U9180 ( .A(n9285), .B(n9311), .Z(n9278) );
  XOR2_X1 U9181 ( .A(n9284), .B(n9283), .Z(n9311) );
  OR2_X1 U9182 ( .A1(n8734), .A2(n8739), .ZN(n9283) );
  OR2_X1 U9183 ( .A1(n9312), .A2(n9313), .ZN(n9284) );
  AND2_X1 U9184 ( .A1(n8645), .A2(n9314), .ZN(n9313) );
  AND2_X1 U9185 ( .A1(n9315), .A2(n9316), .ZN(n9312) );
  OR2_X1 U9186 ( .A1(n9314), .A2(n8645), .ZN(n9316) );
  XOR2_X1 U9187 ( .A(n9317), .B(n9318), .Z(n9285) );
  XOR2_X1 U9188 ( .A(n9319), .B(n9320), .Z(n9318) );
  OR2_X1 U9189 ( .A1(n9321), .A2(n9322), .ZN(n7891) );
  INV_X1 U9190 ( .A(n9323), .ZN(n9322) );
  OR2_X1 U9191 ( .A1(n9324), .A2(n7888), .ZN(n9321) );
  AND3_X1 U9192 ( .A1(n7887), .A2(n7886), .A3(n7884), .ZN(n7888) );
  AND2_X1 U9193 ( .A1(n7880), .A2(n7884), .ZN(n9324) );
  AND2_X1 U9194 ( .A1(n9325), .A2(n9323), .ZN(n7884) );
  OR2_X1 U9195 ( .A1(n9326), .A2(n9327), .ZN(n9323) );
  INV_X1 U9196 ( .A(n9328), .ZN(n9325) );
  AND2_X1 U9197 ( .A1(n9326), .A2(n9327), .ZN(n9328) );
  OR2_X1 U9198 ( .A1(n9329), .A2(n9330), .ZN(n9327) );
  AND2_X1 U9199 ( .A1(n9331), .A2(n9332), .ZN(n9330) );
  AND2_X1 U9200 ( .A1(n9333), .A2(n9334), .ZN(n9329) );
  OR2_X1 U9201 ( .A1(n9332), .A2(n9331), .ZN(n9334) );
  XOR2_X1 U9202 ( .A(n9295), .B(n9335), .Z(n9326) );
  XOR2_X1 U9203 ( .A(n9294), .B(n9293), .Z(n9335) );
  OR2_X1 U9204 ( .A1(n9248), .A2(n8751), .ZN(n9293) );
  OR2_X1 U9205 ( .A1(n9336), .A2(n9337), .ZN(n9294) );
  AND2_X1 U9206 ( .A1(n9338), .A2(n9339), .ZN(n9337) );
  AND2_X1 U9207 ( .A1(n9340), .A2(n9341), .ZN(n9336) );
  OR2_X1 U9208 ( .A1(n9339), .A2(n9338), .ZN(n9341) );
  XOR2_X1 U9209 ( .A(n9302), .B(n9342), .Z(n9295) );
  XOR2_X1 U9210 ( .A(n9301), .B(n9300), .Z(n9342) );
  OR2_X1 U9211 ( .A1(n8730), .A2(n8747), .ZN(n9300) );
  OR2_X1 U9212 ( .A1(n9343), .A2(n9344), .ZN(n9301) );
  AND2_X1 U9213 ( .A1(n9345), .A2(n9346), .ZN(n9344) );
  AND2_X1 U9214 ( .A1(n9347), .A2(n9348), .ZN(n9343) );
  OR2_X1 U9215 ( .A1(n9346), .A2(n9345), .ZN(n9348) );
  XOR2_X1 U9216 ( .A(n9309), .B(n9349), .Z(n9302) );
  XOR2_X1 U9217 ( .A(n9308), .B(n9307), .Z(n9349) );
  OR2_X1 U9218 ( .A1(n8734), .A2(n8743), .ZN(n9307) );
  OR2_X1 U9219 ( .A1(n9350), .A2(n9351), .ZN(n9308) );
  AND2_X1 U9220 ( .A1(n9352), .A2(n9353), .ZN(n9351) );
  AND2_X1 U9221 ( .A1(n9354), .A2(n9355), .ZN(n9350) );
  OR2_X1 U9222 ( .A1(n9353), .A2(n9352), .ZN(n9355) );
  XOR2_X1 U9223 ( .A(n9315), .B(n9356), .Z(n9309) );
  XOR2_X1 U9224 ( .A(n9314), .B(n8645), .Z(n9356) );
  OR2_X1 U9225 ( .A1(n8738), .A2(n8739), .ZN(n8645) );
  OR2_X1 U9226 ( .A1(n9357), .A2(n9358), .ZN(n9314) );
  AND2_X1 U9227 ( .A1(n9359), .A2(n9360), .ZN(n9358) );
  AND2_X1 U9228 ( .A1(n9361), .A2(n9362), .ZN(n9357) );
  OR2_X1 U9229 ( .A1(n9360), .A2(n9359), .ZN(n9362) );
  XOR2_X1 U9230 ( .A(n9363), .B(n9364), .Z(n9315) );
  XOR2_X1 U9231 ( .A(n9365), .B(n9366), .Z(n9364) );
  AND2_X1 U9232 ( .A1(n7876), .A2(n7877), .ZN(n7880) );
  XOR2_X1 U9233 ( .A(n7887), .B(n7886), .Z(n7877) );
  INV_X1 U9234 ( .A(n9367), .ZN(n7886) );
  OR2_X1 U9235 ( .A1(n9368), .A2(n9369), .ZN(n9367) );
  AND2_X1 U9236 ( .A1(n9370), .A2(n9371), .ZN(n9369) );
  AND2_X1 U9237 ( .A1(n9372), .A2(n9373), .ZN(n9368) );
  OR2_X1 U9238 ( .A1(n9371), .A2(n9370), .ZN(n9373) );
  XNOR2_X1 U9239 ( .A(n9333), .B(n9374), .ZN(n7887) );
  XOR2_X1 U9240 ( .A(n9332), .B(n9331), .Z(n9374) );
  OR2_X1 U9241 ( .A1(n9248), .A2(n8755), .ZN(n9331) );
  OR2_X1 U9242 ( .A1(n9375), .A2(n9376), .ZN(n9332) );
  AND2_X1 U9243 ( .A1(n9377), .A2(n9378), .ZN(n9376) );
  AND2_X1 U9244 ( .A1(n9379), .A2(n9380), .ZN(n9375) );
  OR2_X1 U9245 ( .A1(n9378), .A2(n9377), .ZN(n9380) );
  XOR2_X1 U9246 ( .A(n9340), .B(n9381), .Z(n9333) );
  XOR2_X1 U9247 ( .A(n9339), .B(n9338), .Z(n9381) );
  OR2_X1 U9248 ( .A1(n8730), .A2(n8751), .ZN(n9338) );
  OR2_X1 U9249 ( .A1(n9382), .A2(n9383), .ZN(n9339) );
  AND2_X1 U9250 ( .A1(n9384), .A2(n9385), .ZN(n9383) );
  AND2_X1 U9251 ( .A1(n9386), .A2(n9387), .ZN(n9382) );
  OR2_X1 U9252 ( .A1(n9385), .A2(n9384), .ZN(n9387) );
  XOR2_X1 U9253 ( .A(n9347), .B(n9388), .Z(n9340) );
  XOR2_X1 U9254 ( .A(n9346), .B(n9345), .Z(n9388) );
  OR2_X1 U9255 ( .A1(n8734), .A2(n8747), .ZN(n9345) );
  OR2_X1 U9256 ( .A1(n9389), .A2(n9390), .ZN(n9346) );
  AND2_X1 U9257 ( .A1(n9391), .A2(n9392), .ZN(n9390) );
  AND2_X1 U9258 ( .A1(n9393), .A2(n9394), .ZN(n9389) );
  OR2_X1 U9259 ( .A1(n9392), .A2(n9391), .ZN(n9394) );
  XOR2_X1 U9260 ( .A(n9354), .B(n9395), .Z(n9347) );
  XOR2_X1 U9261 ( .A(n9353), .B(n9352), .Z(n9395) );
  OR2_X1 U9262 ( .A1(n8738), .A2(n8743), .ZN(n9352) );
  OR2_X1 U9263 ( .A1(n9396), .A2(n9397), .ZN(n9353) );
  AND2_X1 U9264 ( .A1(n8619), .A2(n9398), .ZN(n9397) );
  AND2_X1 U9265 ( .A1(n9399), .A2(n9400), .ZN(n9396) );
  OR2_X1 U9266 ( .A1(n9398), .A2(n8619), .ZN(n9400) );
  XOR2_X1 U9267 ( .A(n9361), .B(n9401), .Z(n9354) );
  XOR2_X1 U9268 ( .A(n9360), .B(n9359), .Z(n9401) );
  OR2_X1 U9269 ( .A1(n8742), .A2(n8739), .ZN(n9359) );
  OR2_X1 U9270 ( .A1(n9402), .A2(n9403), .ZN(n9360) );
  AND2_X1 U9271 ( .A1(n9404), .A2(n9405), .ZN(n9403) );
  AND2_X1 U9272 ( .A1(n9406), .A2(n9407), .ZN(n9402) );
  OR2_X1 U9273 ( .A1(n9405), .A2(n9404), .ZN(n9407) );
  XOR2_X1 U9274 ( .A(n9408), .B(n9409), .Z(n9361) );
  XOR2_X1 U9275 ( .A(n9410), .B(n9411), .Z(n9409) );
  OR2_X1 U9276 ( .A1(n9412), .A2(n9413), .ZN(n7876) );
  INV_X1 U9277 ( .A(n9414), .ZN(n9413) );
  OR2_X1 U9278 ( .A1(n9415), .A2(n7873), .ZN(n9412) );
  AND3_X1 U9279 ( .A1(n7872), .A2(n7871), .A3(n7869), .ZN(n7873) );
  AND2_X1 U9280 ( .A1(n7869), .A2(n7865), .ZN(n9415) );
  OR2_X1 U9281 ( .A1(n9416), .A2(n9024), .ZN(n7865) );
  AND3_X1 U9282 ( .A1(n9028), .A2(n9026), .A3(n9027), .ZN(n9024) );
  AND2_X1 U9283 ( .A1(n9026), .A2(n9020), .ZN(n9416) );
  OR2_X1 U9284 ( .A1(n9417), .A2(n9013), .ZN(n9020) );
  AND3_X1 U9285 ( .A1(n9017), .A2(n9015), .A3(n9016), .ZN(n9013) );
  AND2_X1 U9286 ( .A1(n9015), .A2(n9009), .ZN(n9417) );
  OR2_X1 U9287 ( .A1(n9418), .A2(n9002), .ZN(n9009) );
  AND3_X1 U9288 ( .A1(n9006), .A2(n9004), .A3(n9005), .ZN(n9002) );
  AND2_X1 U9289 ( .A1(n9004), .A2(n8998), .ZN(n9418) );
  OR2_X1 U9290 ( .A1(n9419), .A2(n8991), .ZN(n8998) );
  AND3_X1 U9291 ( .A1(n8995), .A2(n8993), .A3(n8994), .ZN(n8991) );
  AND2_X1 U9292 ( .A1(n8993), .A2(n8987), .ZN(n9419) );
  OR2_X1 U9293 ( .A1(n9420), .A2(n8980), .ZN(n8987) );
  AND3_X1 U9294 ( .A1(n8984), .A2(n8982), .A3(n8983), .ZN(n8980) );
  INV_X1 U9295 ( .A(n9421), .ZN(n8983) );
  AND2_X1 U9296 ( .A1(n8982), .A2(n8976), .ZN(n9420) );
  OR2_X1 U9297 ( .A1(n9422), .A2(n9423), .ZN(n8976) );
  INV_X1 U9298 ( .A(n8973), .ZN(n9423) );
  OR3_X1 U9299 ( .A1(n9424), .A2(n9425), .A3(n9426), .ZN(n8973) );
  AND2_X1 U9300 ( .A1(n8970), .A2(n8972), .ZN(n9422) );
  INV_X1 U9301 ( .A(n9427), .ZN(n8972) );
  AND2_X1 U9302 ( .A1(n9428), .A2(n9425), .ZN(n9427) );
  XOR2_X1 U9303 ( .A(n8984), .B(n9421), .Z(n9425) );
  OR2_X1 U9304 ( .A1(n9429), .A2(n9430), .ZN(n9421) );
  AND2_X1 U9305 ( .A1(n9431), .A2(n9432), .ZN(n9430) );
  AND2_X1 U9306 ( .A1(n9433), .A2(n9434), .ZN(n9429) );
  OR2_X1 U9307 ( .A1(n9432), .A2(n9431), .ZN(n9434) );
  XNOR2_X1 U9308 ( .A(n9435), .B(n9436), .ZN(n8984) );
  XOR2_X1 U9309 ( .A(n9437), .B(n9438), .Z(n9436) );
  OR2_X1 U9310 ( .A1(n9426), .A2(n9424), .ZN(n9428) );
  OR2_X1 U9311 ( .A1(n9439), .A2(n9440), .ZN(n8970) );
  INV_X1 U9312 ( .A(n8966), .ZN(n9440) );
  OR3_X1 U9313 ( .A1(n9441), .A2(n9442), .A3(n9443), .ZN(n8966) );
  AND2_X1 U9314 ( .A1(n8964), .A2(n8967), .ZN(n9439) );
  INV_X1 U9315 ( .A(n9444), .ZN(n8967) );
  AND2_X1 U9316 ( .A1(n9445), .A2(n9442), .ZN(n9444) );
  XNOR2_X1 U9317 ( .A(n9424), .B(n9426), .ZN(n9442) );
  OR2_X1 U9318 ( .A1(n9446), .A2(n9447), .ZN(n9426) );
  AND2_X1 U9319 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
  AND2_X1 U9320 ( .A1(n9450), .A2(n9451), .ZN(n9446) );
  OR2_X1 U9321 ( .A1(n9448), .A2(n9449), .ZN(n9451) );
  XOR2_X1 U9322 ( .A(n9433), .B(n9452), .Z(n9424) );
  XOR2_X1 U9323 ( .A(n9432), .B(n9431), .Z(n9452) );
  OR2_X1 U9324 ( .A1(n9248), .A2(n8787), .ZN(n9431) );
  OR2_X1 U9325 ( .A1(n9453), .A2(n9454), .ZN(n9432) );
  AND2_X1 U9326 ( .A1(n9455), .A2(n9456), .ZN(n9454) );
  AND2_X1 U9327 ( .A1(n9457), .A2(n9458), .ZN(n9453) );
  OR2_X1 U9328 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  XOR2_X1 U9329 ( .A(n9459), .B(n9460), .Z(n9433) );
  XOR2_X1 U9330 ( .A(n9461), .B(n9462), .Z(n9460) );
  OR2_X1 U9331 ( .A1(n9443), .A2(n9441), .ZN(n9445) );
  OR2_X1 U9332 ( .A1(n9463), .A2(n9464), .ZN(n8964) );
  INV_X1 U9333 ( .A(n8960), .ZN(n9464) );
  OR3_X1 U9334 ( .A1(n9465), .A2(n9466), .A3(n9467), .ZN(n8960) );
  AND2_X1 U9335 ( .A1(n8958), .A2(n8961), .ZN(n9463) );
  INV_X1 U9336 ( .A(n9468), .ZN(n8961) );
  AND2_X1 U9337 ( .A1(n9469), .A2(n9466), .ZN(n9468) );
  XNOR2_X1 U9338 ( .A(n9441), .B(n9443), .ZN(n9466) );
  OR2_X1 U9339 ( .A1(n9470), .A2(n9471), .ZN(n9443) );
  AND2_X1 U9340 ( .A1(n9472), .A2(n9473), .ZN(n9471) );
  AND2_X1 U9341 ( .A1(n9474), .A2(n9475), .ZN(n9470) );
  OR2_X1 U9342 ( .A1(n9472), .A2(n9473), .ZN(n9475) );
  XOR2_X1 U9343 ( .A(n9450), .B(n9476), .Z(n9441) );
  XOR2_X1 U9344 ( .A(n9449), .B(n9448), .Z(n9476) );
  OR2_X1 U9345 ( .A1(n9248), .A2(n8791), .ZN(n9448) );
  OR2_X1 U9346 ( .A1(n9477), .A2(n9478), .ZN(n9449) );
  AND2_X1 U9347 ( .A1(n9479), .A2(n9480), .ZN(n9478) );
  AND2_X1 U9348 ( .A1(n9481), .A2(n9482), .ZN(n9477) );
  OR2_X1 U9349 ( .A1(n9479), .A2(n9480), .ZN(n9482) );
  XOR2_X1 U9350 ( .A(n9457), .B(n9483), .Z(n9450) );
  XOR2_X1 U9351 ( .A(n9456), .B(n9455), .Z(n9483) );
  OR2_X1 U9352 ( .A1(n8730), .A2(n8787), .ZN(n9455) );
  OR2_X1 U9353 ( .A1(n9484), .A2(n9485), .ZN(n9456) );
  AND2_X1 U9354 ( .A1(n9486), .A2(n9487), .ZN(n9485) );
  AND2_X1 U9355 ( .A1(n9488), .A2(n9489), .ZN(n9484) );
  OR2_X1 U9356 ( .A1(n9487), .A2(n9486), .ZN(n9489) );
  XOR2_X1 U9357 ( .A(n9490), .B(n9491), .Z(n9457) );
  XOR2_X1 U9358 ( .A(n9492), .B(n9493), .Z(n9491) );
  OR2_X1 U9359 ( .A1(n9467), .A2(n9465), .ZN(n9469) );
  OR2_X1 U9360 ( .A1(n9494), .A2(n9495), .ZN(n8958) );
  INV_X1 U9361 ( .A(n8955), .ZN(n9495) );
  OR3_X1 U9362 ( .A1(n9496), .A2(n9497), .A3(n9498), .ZN(n8955) );
  AND2_X1 U9363 ( .A1(n8952), .A2(n8954), .ZN(n9494) );
  INV_X1 U9364 ( .A(n9499), .ZN(n8954) );
  AND2_X1 U9365 ( .A1(n9500), .A2(n9497), .ZN(n9499) );
  XNOR2_X1 U9366 ( .A(n9465), .B(n9467), .ZN(n9497) );
  OR2_X1 U9367 ( .A1(n9501), .A2(n9502), .ZN(n9467) );
  AND2_X1 U9368 ( .A1(n9503), .A2(n9504), .ZN(n9502) );
  AND2_X1 U9369 ( .A1(n9505), .A2(n9506), .ZN(n9501) );
  OR2_X1 U9370 ( .A1(n9503), .A2(n9504), .ZN(n9506) );
  XOR2_X1 U9371 ( .A(n9474), .B(n9507), .Z(n9465) );
  XOR2_X1 U9372 ( .A(n9473), .B(n9472), .Z(n9507) );
  OR2_X1 U9373 ( .A1(n9248), .A2(n8795), .ZN(n9472) );
  OR2_X1 U9374 ( .A1(n9508), .A2(n9509), .ZN(n9473) );
  AND2_X1 U9375 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  AND2_X1 U9376 ( .A1(n9512), .A2(n9513), .ZN(n9508) );
  OR2_X1 U9377 ( .A1(n9510), .A2(n9511), .ZN(n9513) );
  XOR2_X1 U9378 ( .A(n9481), .B(n9514), .Z(n9474) );
  XOR2_X1 U9379 ( .A(n9480), .B(n9479), .Z(n9514) );
  OR2_X1 U9380 ( .A1(n8730), .A2(n8791), .ZN(n9479) );
  OR2_X1 U9381 ( .A1(n9515), .A2(n9516), .ZN(n9480) );
  AND2_X1 U9382 ( .A1(n9517), .A2(n9518), .ZN(n9516) );
  AND2_X1 U9383 ( .A1(n9519), .A2(n9520), .ZN(n9515) );
  OR2_X1 U9384 ( .A1(n9517), .A2(n9518), .ZN(n9520) );
  XOR2_X1 U9385 ( .A(n9488), .B(n9521), .Z(n9481) );
  XOR2_X1 U9386 ( .A(n9487), .B(n9486), .Z(n9521) );
  OR2_X1 U9387 ( .A1(n8734), .A2(n8787), .ZN(n9486) );
  OR2_X1 U9388 ( .A1(n9522), .A2(n9523), .ZN(n9487) );
  AND2_X1 U9389 ( .A1(n9524), .A2(n9525), .ZN(n9523) );
  AND2_X1 U9390 ( .A1(n9526), .A2(n9527), .ZN(n9522) );
  OR2_X1 U9391 ( .A1(n9525), .A2(n9524), .ZN(n9527) );
  XOR2_X1 U9392 ( .A(n9528), .B(n9529), .Z(n9488) );
  XOR2_X1 U9393 ( .A(n9530), .B(n9531), .Z(n9529) );
  OR2_X1 U9394 ( .A1(n9498), .A2(n9496), .ZN(n9500) );
  OR2_X1 U9395 ( .A1(n9532), .A2(n9533), .ZN(n8952) );
  INV_X1 U9396 ( .A(n8948), .ZN(n9533) );
  OR3_X1 U9397 ( .A1(n9534), .A2(n9535), .A3(n9536), .ZN(n8948) );
  AND2_X1 U9398 ( .A1(n8946), .A2(n8949), .ZN(n9532) );
  INV_X1 U9399 ( .A(n9537), .ZN(n8949) );
  AND2_X1 U9400 ( .A1(n9538), .A2(n9535), .ZN(n9537) );
  XNOR2_X1 U9401 ( .A(n9496), .B(n9498), .ZN(n9535) );
  OR2_X1 U9402 ( .A1(n9539), .A2(n9540), .ZN(n9498) );
  AND2_X1 U9403 ( .A1(n9541), .A2(n9542), .ZN(n9540) );
  AND2_X1 U9404 ( .A1(n9543), .A2(n9544), .ZN(n9539) );
  OR2_X1 U9405 ( .A1(n9541), .A2(n9542), .ZN(n9544) );
  XOR2_X1 U9406 ( .A(n9505), .B(n9545), .Z(n9496) );
  XOR2_X1 U9407 ( .A(n9504), .B(n9503), .Z(n9545) );
  OR2_X1 U9408 ( .A1(n9248), .A2(n8799), .ZN(n9503) );
  OR2_X1 U9409 ( .A1(n9546), .A2(n9547), .ZN(n9504) );
  AND2_X1 U9410 ( .A1(n9548), .A2(n9549), .ZN(n9547) );
  AND2_X1 U9411 ( .A1(n9550), .A2(n9551), .ZN(n9546) );
  OR2_X1 U9412 ( .A1(n9548), .A2(n9549), .ZN(n9551) );
  XOR2_X1 U9413 ( .A(n9512), .B(n9552), .Z(n9505) );
  XOR2_X1 U9414 ( .A(n9511), .B(n9510), .Z(n9552) );
  OR2_X1 U9415 ( .A1(n8730), .A2(n8795), .ZN(n9510) );
  OR2_X1 U9416 ( .A1(n9553), .A2(n9554), .ZN(n9511) );
  AND2_X1 U9417 ( .A1(n9555), .A2(n9556), .ZN(n9554) );
  AND2_X1 U9418 ( .A1(n9557), .A2(n9558), .ZN(n9553) );
  OR2_X1 U9419 ( .A1(n9555), .A2(n9556), .ZN(n9558) );
  XOR2_X1 U9420 ( .A(n9519), .B(n9559), .Z(n9512) );
  XOR2_X1 U9421 ( .A(n9518), .B(n9517), .Z(n9559) );
  OR2_X1 U9422 ( .A1(n8734), .A2(n8791), .ZN(n9517) );
  OR2_X1 U9423 ( .A1(n9560), .A2(n9561), .ZN(n9518) );
  AND2_X1 U9424 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  AND2_X1 U9425 ( .A1(n9564), .A2(n9565), .ZN(n9560) );
  OR2_X1 U9426 ( .A1(n9562), .A2(n9563), .ZN(n9565) );
  XOR2_X1 U9427 ( .A(n9526), .B(n9566), .Z(n9519) );
  XOR2_X1 U9428 ( .A(n9525), .B(n9524), .Z(n9566) );
  OR2_X1 U9429 ( .A1(n8738), .A2(n8787), .ZN(n9524) );
  OR2_X1 U9430 ( .A1(n9567), .A2(n9568), .ZN(n9525) );
  AND2_X1 U9431 ( .A1(n9569), .A2(n9570), .ZN(n9568) );
  AND2_X1 U9432 ( .A1(n9571), .A2(n9572), .ZN(n9567) );
  OR2_X1 U9433 ( .A1(n9570), .A2(n9569), .ZN(n9572) );
  XOR2_X1 U9434 ( .A(n9573), .B(n9574), .Z(n9526) );
  XOR2_X1 U9435 ( .A(n9575), .B(n9576), .Z(n9574) );
  OR2_X1 U9436 ( .A1(n9536), .A2(n9534), .ZN(n9538) );
  OR2_X1 U9437 ( .A1(n9577), .A2(n9578), .ZN(n8946) );
  INV_X1 U9438 ( .A(n8931), .ZN(n9578) );
  OR3_X1 U9439 ( .A1(n9579), .A2(n9580), .A3(n9581), .ZN(n8931) );
  AND2_X1 U9440 ( .A1(n8929), .A2(n8932), .ZN(n9577) );
  INV_X1 U9441 ( .A(n9582), .ZN(n8932) );
  AND2_X1 U9442 ( .A1(n9583), .A2(n9580), .ZN(n9582) );
  XNOR2_X1 U9443 ( .A(n9534), .B(n9536), .ZN(n9580) );
  OR2_X1 U9444 ( .A1(n9584), .A2(n9585), .ZN(n9536) );
  AND2_X1 U9445 ( .A1(n9586), .A2(n9587), .ZN(n9585) );
  AND2_X1 U9446 ( .A1(n9588), .A2(n9589), .ZN(n9584) );
  OR2_X1 U9447 ( .A1(n9586), .A2(n9587), .ZN(n9589) );
  XOR2_X1 U9448 ( .A(n9543), .B(n9590), .Z(n9534) );
  XOR2_X1 U9449 ( .A(n9542), .B(n9541), .Z(n9590) );
  OR2_X1 U9450 ( .A1(n9248), .A2(n8803), .ZN(n9541) );
  OR2_X1 U9451 ( .A1(n9591), .A2(n9592), .ZN(n9542) );
  AND2_X1 U9452 ( .A1(n9593), .A2(n9594), .ZN(n9592) );
  AND2_X1 U9453 ( .A1(n9595), .A2(n9596), .ZN(n9591) );
  OR2_X1 U9454 ( .A1(n9593), .A2(n9594), .ZN(n9596) );
  XOR2_X1 U9455 ( .A(n9550), .B(n9597), .Z(n9543) );
  XOR2_X1 U9456 ( .A(n9549), .B(n9548), .Z(n9597) );
  OR2_X1 U9457 ( .A1(n8730), .A2(n8799), .ZN(n9548) );
  OR2_X1 U9458 ( .A1(n9598), .A2(n9599), .ZN(n9549) );
  AND2_X1 U9459 ( .A1(n9600), .A2(n9601), .ZN(n9599) );
  AND2_X1 U9460 ( .A1(n9602), .A2(n9603), .ZN(n9598) );
  OR2_X1 U9461 ( .A1(n9600), .A2(n9601), .ZN(n9603) );
  XOR2_X1 U9462 ( .A(n9557), .B(n9604), .Z(n9550) );
  XOR2_X1 U9463 ( .A(n9556), .B(n9555), .Z(n9604) );
  OR2_X1 U9464 ( .A1(n8734), .A2(n8795), .ZN(n9555) );
  OR2_X1 U9465 ( .A1(n9605), .A2(n9606), .ZN(n9556) );
  AND2_X1 U9466 ( .A1(n9607), .A2(n9608), .ZN(n9606) );
  AND2_X1 U9467 ( .A1(n9609), .A2(n9610), .ZN(n9605) );
  OR2_X1 U9468 ( .A1(n9607), .A2(n9608), .ZN(n9610) );
  XOR2_X1 U9469 ( .A(n9564), .B(n9611), .Z(n9557) );
  XOR2_X1 U9470 ( .A(n9563), .B(n9562), .Z(n9611) );
  OR2_X1 U9471 ( .A1(n8738), .A2(n8791), .ZN(n9562) );
  OR2_X1 U9472 ( .A1(n9612), .A2(n9613), .ZN(n9563) );
  AND2_X1 U9473 ( .A1(n9614), .A2(n9615), .ZN(n9613) );
  AND2_X1 U9474 ( .A1(n9616), .A2(n9617), .ZN(n9612) );
  OR2_X1 U9475 ( .A1(n9614), .A2(n9615), .ZN(n9617) );
  XOR2_X1 U9476 ( .A(n9571), .B(n9618), .Z(n9564) );
  XOR2_X1 U9477 ( .A(n9570), .B(n9569), .Z(n9618) );
  OR2_X1 U9478 ( .A1(n8742), .A2(n8787), .ZN(n9569) );
  OR2_X1 U9479 ( .A1(n9619), .A2(n9620), .ZN(n9570) );
  AND2_X1 U9480 ( .A1(n9621), .A2(n9622), .ZN(n9620) );
  AND2_X1 U9481 ( .A1(n9623), .A2(n9624), .ZN(n9619) );
  OR2_X1 U9482 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  XOR2_X1 U9483 ( .A(n9625), .B(n9626), .Z(n9571) );
  XOR2_X1 U9484 ( .A(n9627), .B(n9628), .Z(n9626) );
  OR2_X1 U9485 ( .A1(n9581), .A2(n9579), .ZN(n9583) );
  OR2_X1 U9486 ( .A1(n9629), .A2(n8926), .ZN(n8929) );
  AND3_X1 U9487 ( .A1(n9630), .A2(n9631), .A3(n9632), .ZN(n8926) );
  AND2_X1 U9488 ( .A1(n8925), .A2(n8922), .ZN(n9629) );
  OR2_X1 U9489 ( .A1(n9633), .A2(n9634), .ZN(n8922) );
  INV_X1 U9490 ( .A(n8919), .ZN(n9634) );
  OR3_X1 U9491 ( .A1(n9635), .A2(n9636), .A3(n9637), .ZN(n8919) );
  AND2_X1 U9492 ( .A1(n8916), .A2(n8918), .ZN(n9633) );
  INV_X1 U9493 ( .A(n9638), .ZN(n8918) );
  AND2_X1 U9494 ( .A1(n9639), .A2(n9636), .ZN(n9638) );
  XOR2_X1 U9495 ( .A(n9630), .B(n9640), .Z(n9636) );
  OR2_X1 U9496 ( .A1(n9637), .A2(n9635), .ZN(n9639) );
  OR2_X1 U9497 ( .A1(n9641), .A2(n9642), .ZN(n8916) );
  INV_X1 U9498 ( .A(n8912), .ZN(n9642) );
  OR3_X1 U9499 ( .A1(n9643), .A2(n9644), .A3(n9645), .ZN(n8912) );
  AND2_X1 U9500 ( .A1(n8910), .A2(n8913), .ZN(n9641) );
  INV_X1 U9501 ( .A(n9646), .ZN(n8913) );
  AND2_X1 U9502 ( .A1(n9647), .A2(n9644), .ZN(n9646) );
  XNOR2_X1 U9503 ( .A(n9635), .B(n9637), .ZN(n9644) );
  OR2_X1 U9504 ( .A1(n9648), .A2(n9649), .ZN(n9637) );
  AND2_X1 U9505 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  AND2_X1 U9506 ( .A1(n9652), .A2(n9653), .ZN(n9648) );
  OR2_X1 U9507 ( .A1(n9650), .A2(n9651), .ZN(n9653) );
  XOR2_X1 U9508 ( .A(n9654), .B(n9655), .Z(n9635) );
  XOR2_X1 U9509 ( .A(n9656), .B(n9657), .Z(n9655) );
  OR2_X1 U9510 ( .A1(n9645), .A2(n9643), .ZN(n9647) );
  OR2_X1 U9511 ( .A1(n9658), .A2(n9659), .ZN(n8910) );
  INV_X1 U9512 ( .A(n8906), .ZN(n9659) );
  OR3_X1 U9513 ( .A1(n9660), .A2(n9661), .A3(n9662), .ZN(n8906) );
  AND2_X1 U9514 ( .A1(n8904), .A2(n8907), .ZN(n9658) );
  INV_X1 U9515 ( .A(n9663), .ZN(n8907) );
  AND2_X1 U9516 ( .A1(n9664), .A2(n9661), .ZN(n9663) );
  XNOR2_X1 U9517 ( .A(n9643), .B(n9645), .ZN(n9661) );
  OR2_X1 U9518 ( .A1(n9665), .A2(n9666), .ZN(n9645) );
  AND2_X1 U9519 ( .A1(n9667), .A2(n9668), .ZN(n9666) );
  AND2_X1 U9520 ( .A1(n9669), .A2(n9670), .ZN(n9665) );
  OR2_X1 U9521 ( .A1(n9667), .A2(n9668), .ZN(n9670) );
  XOR2_X1 U9522 ( .A(n9652), .B(n9671), .Z(n9643) );
  XOR2_X1 U9523 ( .A(n9651), .B(n9650), .Z(n9671) );
  OR2_X1 U9524 ( .A1(n9248), .A2(n8818), .ZN(n9650) );
  OR2_X1 U9525 ( .A1(n9672), .A2(n9673), .ZN(n9651) );
  AND2_X1 U9526 ( .A1(n9674), .A2(n9675), .ZN(n9673) );
  AND2_X1 U9527 ( .A1(n9676), .A2(n9677), .ZN(n9672) );
  OR2_X1 U9528 ( .A1(n9674), .A2(n9675), .ZN(n9677) );
  XOR2_X1 U9529 ( .A(n9678), .B(n9679), .Z(n9652) );
  XOR2_X1 U9530 ( .A(n9680), .B(n9681), .Z(n9679) );
  OR2_X1 U9531 ( .A1(n9662), .A2(n9660), .ZN(n9664) );
  OR2_X1 U9532 ( .A1(n9682), .A2(n8901), .ZN(n8904) );
  AND3_X1 U9533 ( .A1(n9683), .A2(n9684), .A3(n9685), .ZN(n8901) );
  AND2_X1 U9534 ( .A1(n8900), .A2(n8897), .ZN(n9682) );
  OR2_X1 U9535 ( .A1(n9686), .A2(n8894), .ZN(n8897) );
  AND2_X1 U9536 ( .A1(n9687), .A2(n9688), .ZN(n8894) );
  AND2_X1 U9537 ( .A1(n8892), .A2(n8890), .ZN(n9686) );
  OR2_X1 U9538 ( .A1(n9689), .A2(n8887), .ZN(n8890) );
  AND3_X1 U9539 ( .A1(n9690), .A2(n9691), .A3(n9692), .ZN(n8887) );
  AND2_X1 U9540 ( .A1(n8885), .A2(n8883), .ZN(n9689) );
  OR2_X1 U9541 ( .A1(n9693), .A2(n8880), .ZN(n8883) );
  AND3_X1 U9542 ( .A1(n9694), .A2(n9695), .A3(n9696), .ZN(n8880) );
  AND2_X1 U9543 ( .A1(n8878), .A2(n9697), .ZN(n9693) );
  INV_X1 U9544 ( .A(n8876), .ZN(n9697) );
  AND2_X1 U9545 ( .A1(n9698), .A2(n8871), .ZN(n8876) );
  OR3_X1 U9546 ( .A1(n9699), .A2(n9700), .A3(n9701), .ZN(n8871) );
  OR2_X1 U9547 ( .A1(n8868), .A2(n8873), .ZN(n9698) );
  AND2_X1 U9548 ( .A1(n9702), .A2(n9699), .ZN(n8873) );
  XOR2_X1 U9549 ( .A(n9694), .B(n9703), .Z(n9699) );
  OR2_X1 U9550 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  INV_X1 U9551 ( .A(n8869), .ZN(n8868) );
  AND3_X1 U9552 ( .A1(n8855), .A2(n8860), .A3(n8854), .ZN(n8869) );
  INV_X1 U9553 ( .A(n9704), .ZN(n8854) );
  OR2_X1 U9554 ( .A1(n9705), .A2(n9706), .ZN(n9704) );
  AND2_X1 U9555 ( .A1(n8709), .A2(n8708), .ZN(n9706) );
  AND2_X1 U9556 ( .A1(n8706), .A2(n9707), .ZN(n9705) );
  OR2_X1 U9557 ( .A1(n8709), .A2(n8708), .ZN(n9707) );
  OR2_X1 U9558 ( .A1(n9708), .A2(n9709), .ZN(n8708) );
  AND2_X1 U9559 ( .A1(n8683), .A2(n8682), .ZN(n9709) );
  AND2_X1 U9560 ( .A1(n8680), .A2(n9710), .ZN(n9708) );
  OR2_X1 U9561 ( .A1(n8683), .A2(n8682), .ZN(n9710) );
  OR2_X1 U9562 ( .A1(n9711), .A2(n9712), .ZN(n8682) );
  AND2_X1 U9563 ( .A1(n8657), .A2(n8656), .ZN(n9712) );
  AND2_X1 U9564 ( .A1(n8654), .A2(n9713), .ZN(n9711) );
  OR2_X1 U9565 ( .A1(n8657), .A2(n8656), .ZN(n9713) );
  OR2_X1 U9566 ( .A1(n9714), .A2(n9715), .ZN(n8656) );
  AND2_X1 U9567 ( .A1(n8631), .A2(n8630), .ZN(n9715) );
  AND2_X1 U9568 ( .A1(n8628), .A2(n9716), .ZN(n9714) );
  OR2_X1 U9569 ( .A1(n8631), .A2(n8630), .ZN(n9716) );
  OR2_X1 U9570 ( .A1(n9717), .A2(n9718), .ZN(n8630) );
  AND2_X1 U9571 ( .A1(n8605), .A2(n8604), .ZN(n9718) );
  AND2_X1 U9572 ( .A1(n8602), .A2(n9719), .ZN(n9717) );
  OR2_X1 U9573 ( .A1(n8605), .A2(n8604), .ZN(n9719) );
  OR2_X1 U9574 ( .A1(n9720), .A2(n9721), .ZN(n8604) );
  AND2_X1 U9575 ( .A1(n8579), .A2(n8578), .ZN(n9721) );
  AND2_X1 U9576 ( .A1(n8576), .A2(n9722), .ZN(n9720) );
  OR2_X1 U9577 ( .A1(n8579), .A2(n8578), .ZN(n9722) );
  OR2_X1 U9578 ( .A1(n9723), .A2(n9724), .ZN(n8578) );
  AND2_X1 U9579 ( .A1(n8553), .A2(n8552), .ZN(n9724) );
  AND2_X1 U9580 ( .A1(n8550), .A2(n9725), .ZN(n9723) );
  OR2_X1 U9581 ( .A1(n8553), .A2(n8552), .ZN(n9725) );
  OR2_X1 U9582 ( .A1(n9726), .A2(n9727), .ZN(n8552) );
  AND2_X1 U9583 ( .A1(n8527), .A2(n8526), .ZN(n9727) );
  AND2_X1 U9584 ( .A1(n8524), .A2(n9728), .ZN(n9726) );
  OR2_X1 U9585 ( .A1(n8527), .A2(n8526), .ZN(n9728) );
  OR2_X1 U9586 ( .A1(n9729), .A2(n9730), .ZN(n8526) );
  AND2_X1 U9587 ( .A1(n8490), .A2(n8489), .ZN(n9730) );
  AND2_X1 U9588 ( .A1(n8487), .A2(n9731), .ZN(n9729) );
  OR2_X1 U9589 ( .A1(n8490), .A2(n8489), .ZN(n9731) );
  OR2_X1 U9590 ( .A1(n9732), .A2(n9733), .ZN(n8489) );
  AND2_X1 U9591 ( .A1(n8464), .A2(n8463), .ZN(n9733) );
  AND2_X1 U9592 ( .A1(n8461), .A2(n9734), .ZN(n9732) );
  OR2_X1 U9593 ( .A1(n8464), .A2(n8463), .ZN(n9734) );
  OR2_X1 U9594 ( .A1(n9735), .A2(n9736), .ZN(n8463) );
  AND2_X1 U9595 ( .A1(n8438), .A2(n8437), .ZN(n9736) );
  AND2_X1 U9596 ( .A1(n8435), .A2(n9737), .ZN(n9735) );
  OR2_X1 U9597 ( .A1(n8438), .A2(n8437), .ZN(n9737) );
  OR2_X1 U9598 ( .A1(n9738), .A2(n9739), .ZN(n8437) );
  AND2_X1 U9599 ( .A1(n8412), .A2(n8411), .ZN(n9739) );
  AND2_X1 U9600 ( .A1(n8409), .A2(n9740), .ZN(n9738) );
  OR2_X1 U9601 ( .A1(n8412), .A2(n8411), .ZN(n9740) );
  OR2_X1 U9602 ( .A1(n9741), .A2(n9742), .ZN(n8411) );
  AND2_X1 U9603 ( .A1(n8386), .A2(n8385), .ZN(n9742) );
  AND2_X1 U9604 ( .A1(n8383), .A2(n9743), .ZN(n9741) );
  OR2_X1 U9605 ( .A1(n8386), .A2(n8385), .ZN(n9743) );
  OR2_X1 U9606 ( .A1(n9744), .A2(n9745), .ZN(n8385) );
  AND2_X1 U9607 ( .A1(n8360), .A2(n8359), .ZN(n9745) );
  AND2_X1 U9608 ( .A1(n8357), .A2(n9746), .ZN(n9744) );
  OR2_X1 U9609 ( .A1(n8360), .A2(n8359), .ZN(n9746) );
  OR2_X1 U9610 ( .A1(n9747), .A2(n9748), .ZN(n8359) );
  AND2_X1 U9611 ( .A1(n8334), .A2(n8333), .ZN(n9748) );
  AND2_X1 U9612 ( .A1(n8331), .A2(n9749), .ZN(n9747) );
  OR2_X1 U9613 ( .A1(n8334), .A2(n8333), .ZN(n9749) );
  OR2_X1 U9614 ( .A1(n9750), .A2(n9751), .ZN(n8333) );
  AND2_X1 U9615 ( .A1(n8308), .A2(n8307), .ZN(n9751) );
  AND2_X1 U9616 ( .A1(n8305), .A2(n9752), .ZN(n9750) );
  OR2_X1 U9617 ( .A1(n8308), .A2(n8307), .ZN(n9752) );
  OR2_X1 U9618 ( .A1(n9753), .A2(n9754), .ZN(n8307) );
  AND2_X1 U9619 ( .A1(n8282), .A2(n8281), .ZN(n9754) );
  AND2_X1 U9620 ( .A1(n8279), .A2(n9755), .ZN(n9753) );
  OR2_X1 U9621 ( .A1(n8282), .A2(n8281), .ZN(n9755) );
  OR2_X1 U9622 ( .A1(n9756), .A2(n9757), .ZN(n8281) );
  AND2_X1 U9623 ( .A1(n8256), .A2(n8255), .ZN(n9757) );
  AND2_X1 U9624 ( .A1(n8253), .A2(n9758), .ZN(n9756) );
  OR2_X1 U9625 ( .A1(n8256), .A2(n8255), .ZN(n9758) );
  OR2_X1 U9626 ( .A1(n9759), .A2(n9760), .ZN(n8255) );
  AND2_X1 U9627 ( .A1(n8226), .A2(n8225), .ZN(n9760) );
  AND2_X1 U9628 ( .A1(n8223), .A2(n9761), .ZN(n9759) );
  OR2_X1 U9629 ( .A1(n8226), .A2(n8225), .ZN(n9761) );
  OR2_X1 U9630 ( .A1(n9762), .A2(n9763), .ZN(n8225) );
  AND2_X1 U9631 ( .A1(n8200), .A2(n8199), .ZN(n9763) );
  AND2_X1 U9632 ( .A1(n8197), .A2(n9764), .ZN(n9762) );
  OR2_X1 U9633 ( .A1(n8200), .A2(n8199), .ZN(n9764) );
  OR2_X1 U9634 ( .A1(n9765), .A2(n9766), .ZN(n8199) );
  AND2_X1 U9635 ( .A1(n8174), .A2(n8173), .ZN(n9766) );
  AND2_X1 U9636 ( .A1(n8171), .A2(n9767), .ZN(n9765) );
  OR2_X1 U9637 ( .A1(n8174), .A2(n8173), .ZN(n9767) );
  OR2_X1 U9638 ( .A1(n9768), .A2(n9769), .ZN(n8173) );
  AND2_X1 U9639 ( .A1(n8148), .A2(n8147), .ZN(n9769) );
  AND2_X1 U9640 ( .A1(n8145), .A2(n9770), .ZN(n9768) );
  OR2_X1 U9641 ( .A1(n8148), .A2(n8147), .ZN(n9770) );
  OR2_X1 U9642 ( .A1(n9771), .A2(n9772), .ZN(n8147) );
  AND2_X1 U9643 ( .A1(n8123), .A2(n8122), .ZN(n9772) );
  AND2_X1 U9644 ( .A1(n8120), .A2(n9773), .ZN(n9771) );
  OR2_X1 U9645 ( .A1(n8123), .A2(n8122), .ZN(n9773) );
  OR2_X1 U9646 ( .A1(n9774), .A2(n9775), .ZN(n8122) );
  AND2_X1 U9647 ( .A1(n8098), .A2(n8097), .ZN(n9775) );
  AND2_X1 U9648 ( .A1(n8095), .A2(n9776), .ZN(n9774) );
  OR2_X1 U9649 ( .A1(n8098), .A2(n8097), .ZN(n9776) );
  OR2_X1 U9650 ( .A1(n9777), .A2(n9778), .ZN(n8097) );
  AND2_X1 U9651 ( .A1(n8073), .A2(n8072), .ZN(n9778) );
  AND2_X1 U9652 ( .A1(n8070), .A2(n9779), .ZN(n9777) );
  OR2_X1 U9653 ( .A1(n8073), .A2(n8072), .ZN(n9779) );
  OR2_X1 U9654 ( .A1(n9780), .A2(n9781), .ZN(n8072) );
  AND2_X1 U9655 ( .A1(n8048), .A2(n8047), .ZN(n9781) );
  AND2_X1 U9656 ( .A1(n8045), .A2(n9782), .ZN(n9780) );
  OR2_X1 U9657 ( .A1(n8048), .A2(n8047), .ZN(n9782) );
  OR2_X1 U9658 ( .A1(n9783), .A2(n9784), .ZN(n8047) );
  AND2_X1 U9659 ( .A1(n8023), .A2(n8022), .ZN(n9784) );
  AND2_X1 U9660 ( .A1(n8020), .A2(n9785), .ZN(n9783) );
  OR2_X1 U9661 ( .A1(n8023), .A2(n8022), .ZN(n9785) );
  OR2_X1 U9662 ( .A1(n9786), .A2(n9787), .ZN(n8022) );
  AND2_X1 U9663 ( .A1(n7998), .A2(n7997), .ZN(n9787) );
  AND2_X1 U9664 ( .A1(n7995), .A2(n9788), .ZN(n9786) );
  OR2_X1 U9665 ( .A1(n7998), .A2(n7997), .ZN(n9788) );
  OR2_X1 U9666 ( .A1(n9789), .A2(n9790), .ZN(n7997) );
  AND2_X1 U9667 ( .A1(n7962), .A2(n7961), .ZN(n9790) );
  AND2_X1 U9668 ( .A1(n7959), .A2(n9791), .ZN(n9789) );
  OR2_X1 U9669 ( .A1(n7962), .A2(n7961), .ZN(n9791) );
  OR2_X1 U9670 ( .A1(n9792), .A2(n9793), .ZN(n7961) );
  AND2_X1 U9671 ( .A1(n7934), .A2(n7937), .ZN(n9793) );
  AND2_X1 U9672 ( .A1(n9794), .A2(n9795), .ZN(n9792) );
  OR2_X1 U9673 ( .A1(n7934), .A2(n7937), .ZN(n9795) );
  OR2_X1 U9674 ( .A1(n7954), .A2(n8848), .ZN(n7937) );
  OR2_X1 U9675 ( .A1(n7908), .A2(n8844), .ZN(n7934) );
  OR2_X1 U9676 ( .A1(n8848), .A2(n9796), .ZN(n8844) );
  INV_X1 U9677 ( .A(n7936), .ZN(n9794) );
  OR2_X1 U9678 ( .A1(n9797), .A2(n9798), .ZN(n7936) );
  AND2_X1 U9679 ( .A1(b_30_), .A2(n9799), .ZN(n9798) );
  OR2_X1 U9680 ( .A1(n9800), .A2(n9801), .ZN(n9799) );
  AND2_X1 U9681 ( .A1(a_30_), .A2(n8842), .ZN(n9800) );
  AND2_X1 U9682 ( .A1(b_29_), .A2(n9802), .ZN(n9797) );
  OR2_X1 U9683 ( .A1(n9803), .A2(n7920), .ZN(n9802) );
  AND2_X1 U9684 ( .A1(a_31_), .A2(n7908), .ZN(n9803) );
  OR2_X1 U9685 ( .A1(n7979), .A2(n8848), .ZN(n7962) );
  XNOR2_X1 U9686 ( .A(n9804), .B(n9805), .ZN(n7959) );
  XOR2_X1 U9687 ( .A(n9806), .B(n9807), .Z(n9805) );
  OR2_X1 U9688 ( .A1(n8015), .A2(n8848), .ZN(n7998) );
  XOR2_X1 U9689 ( .A(n9808), .B(n9809), .Z(n7995) );
  XOR2_X1 U9690 ( .A(n9810), .B(n9811), .Z(n9809) );
  OR2_X1 U9691 ( .A1(n8040), .A2(n8848), .ZN(n8023) );
  XOR2_X1 U9692 ( .A(n9812), .B(n9813), .Z(n8020) );
  XOR2_X1 U9693 ( .A(n9814), .B(n9815), .Z(n9813) );
  OR2_X1 U9694 ( .A1(n8065), .A2(n8848), .ZN(n8048) );
  XOR2_X1 U9695 ( .A(n9816), .B(n9817), .Z(n8045) );
  XOR2_X1 U9696 ( .A(n9818), .B(n9819), .Z(n9817) );
  OR2_X1 U9697 ( .A1(n8090), .A2(n8848), .ZN(n8073) );
  XOR2_X1 U9698 ( .A(n9820), .B(n9821), .Z(n8070) );
  XOR2_X1 U9699 ( .A(n9822), .B(n9823), .Z(n9821) );
  OR2_X1 U9700 ( .A1(n8115), .A2(n8848), .ZN(n8098) );
  XOR2_X1 U9701 ( .A(n9824), .B(n9825), .Z(n8095) );
  XOR2_X1 U9702 ( .A(n9826), .B(n9827), .Z(n9825) );
  OR2_X1 U9703 ( .A1(n8140), .A2(n8848), .ZN(n8123) );
  XOR2_X1 U9704 ( .A(n9828), .B(n9829), .Z(n8120) );
  XOR2_X1 U9705 ( .A(n9830), .B(n9831), .Z(n9829) );
  OR2_X1 U9706 ( .A1(n8810), .A2(n8848), .ZN(n8148) );
  XOR2_X1 U9707 ( .A(n9832), .B(n9833), .Z(n8145) );
  XOR2_X1 U9708 ( .A(n9834), .B(n9835), .Z(n9833) );
  OR2_X1 U9709 ( .A1(n8806), .A2(n8848), .ZN(n8174) );
  XOR2_X1 U9710 ( .A(n9836), .B(n9837), .Z(n8171) );
  XOR2_X1 U9711 ( .A(n9838), .B(n9839), .Z(n9837) );
  OR2_X1 U9712 ( .A1(n8802), .A2(n8848), .ZN(n8200) );
  XOR2_X1 U9713 ( .A(n9840), .B(n9841), .Z(n8197) );
  XOR2_X1 U9714 ( .A(n9842), .B(n9843), .Z(n9841) );
  OR2_X1 U9715 ( .A1(n8798), .A2(n8848), .ZN(n8226) );
  XOR2_X1 U9716 ( .A(n9844), .B(n9845), .Z(n8223) );
  XOR2_X1 U9717 ( .A(n9846), .B(n9847), .Z(n9845) );
  OR2_X1 U9718 ( .A1(n8794), .A2(n8848), .ZN(n8256) );
  XOR2_X1 U9719 ( .A(n9848), .B(n9849), .Z(n8253) );
  XOR2_X1 U9720 ( .A(n9850), .B(n9851), .Z(n9849) );
  OR2_X1 U9721 ( .A1(n8790), .A2(n8848), .ZN(n8282) );
  XOR2_X1 U9722 ( .A(n9852), .B(n9853), .Z(n8279) );
  XOR2_X1 U9723 ( .A(n9854), .B(n9855), .Z(n9853) );
  OR2_X1 U9724 ( .A1(n8786), .A2(n8848), .ZN(n8308) );
  XOR2_X1 U9725 ( .A(n9856), .B(n9857), .Z(n8305) );
  XOR2_X1 U9726 ( .A(n9858), .B(n9859), .Z(n9857) );
  OR2_X1 U9727 ( .A1(n8782), .A2(n8848), .ZN(n8334) );
  XOR2_X1 U9728 ( .A(n9860), .B(n9861), .Z(n8331) );
  XOR2_X1 U9729 ( .A(n9862), .B(n9863), .Z(n9861) );
  OR2_X1 U9730 ( .A1(n8778), .A2(n8848), .ZN(n8360) );
  XOR2_X1 U9731 ( .A(n9864), .B(n9865), .Z(n8357) );
  XOR2_X1 U9732 ( .A(n9866), .B(n9867), .Z(n9865) );
  OR2_X1 U9733 ( .A1(n8774), .A2(n8848), .ZN(n8386) );
  XOR2_X1 U9734 ( .A(n9868), .B(n9869), .Z(n8383) );
  XOR2_X1 U9735 ( .A(n9870), .B(n9871), .Z(n9869) );
  OR2_X1 U9736 ( .A1(n8770), .A2(n8848), .ZN(n8412) );
  XOR2_X1 U9737 ( .A(n9872), .B(n9873), .Z(n8409) );
  XOR2_X1 U9738 ( .A(n9874), .B(n9875), .Z(n9873) );
  OR2_X1 U9739 ( .A1(n8766), .A2(n8848), .ZN(n8438) );
  XOR2_X1 U9740 ( .A(n9876), .B(n9877), .Z(n8435) );
  XOR2_X1 U9741 ( .A(n9878), .B(n9879), .Z(n9877) );
  OR2_X1 U9742 ( .A1(n8762), .A2(n8848), .ZN(n8464) );
  XOR2_X1 U9743 ( .A(n9880), .B(n9881), .Z(n8461) );
  XOR2_X1 U9744 ( .A(n9882), .B(n9883), .Z(n9881) );
  OR2_X1 U9745 ( .A1(n8758), .A2(n8848), .ZN(n8490) );
  XOR2_X1 U9746 ( .A(n9884), .B(n9885), .Z(n8487) );
  XOR2_X1 U9747 ( .A(n9886), .B(n9887), .Z(n9885) );
  OR2_X1 U9748 ( .A1(n8754), .A2(n8848), .ZN(n8527) );
  XOR2_X1 U9749 ( .A(n9888), .B(n9889), .Z(n8524) );
  XOR2_X1 U9750 ( .A(n9890), .B(n9891), .Z(n9889) );
  OR2_X1 U9751 ( .A1(n8750), .A2(n8848), .ZN(n8553) );
  XOR2_X1 U9752 ( .A(n9892), .B(n9893), .Z(n8550) );
  XOR2_X1 U9753 ( .A(n9894), .B(n9895), .Z(n9893) );
  OR2_X1 U9754 ( .A1(n8746), .A2(n8848), .ZN(n8579) );
  XOR2_X1 U9755 ( .A(n9896), .B(n9897), .Z(n8576) );
  XOR2_X1 U9756 ( .A(n9898), .B(n9899), .Z(n9897) );
  OR2_X1 U9757 ( .A1(n8742), .A2(n8848), .ZN(n8605) );
  XOR2_X1 U9758 ( .A(n9900), .B(n9901), .Z(n8602) );
  XOR2_X1 U9759 ( .A(n9902), .B(n9903), .Z(n9901) );
  OR2_X1 U9760 ( .A1(n8738), .A2(n8848), .ZN(n8631) );
  XOR2_X1 U9761 ( .A(n9904), .B(n9905), .Z(n8628) );
  XOR2_X1 U9762 ( .A(n9906), .B(n9907), .Z(n9905) );
  OR2_X1 U9763 ( .A1(n8734), .A2(n8848), .ZN(n8657) );
  XOR2_X1 U9764 ( .A(n9908), .B(n9909), .Z(n8654) );
  XOR2_X1 U9765 ( .A(n9910), .B(n9911), .Z(n9909) );
  OR2_X1 U9766 ( .A1(n8730), .A2(n8848), .ZN(n8683) );
  XOR2_X1 U9767 ( .A(n9912), .B(n9913), .Z(n8680) );
  XOR2_X1 U9768 ( .A(n9914), .B(n9915), .Z(n9913) );
  OR2_X1 U9769 ( .A1(n9248), .A2(n8848), .ZN(n8709) );
  INV_X1 U9770 ( .A(b_31_), .ZN(n8848) );
  XOR2_X1 U9771 ( .A(n9916), .B(n9917), .Z(n8706) );
  XOR2_X1 U9772 ( .A(n9918), .B(n9919), .Z(n9917) );
  XOR2_X1 U9773 ( .A(n9700), .B(n9701), .Z(n8860) );
  OR2_X1 U9774 ( .A1(n9920), .A2(n9921), .ZN(n9701) );
  AND2_X1 U9775 ( .A1(n9922), .A2(n9923), .ZN(n9921) );
  AND2_X1 U9776 ( .A1(n9924), .A2(n9925), .ZN(n9920) );
  OR2_X1 U9777 ( .A1(n9922), .A2(n9923), .ZN(n9925) );
  XOR2_X1 U9778 ( .A(n9926), .B(n9927), .Z(n9700) );
  XOR2_X1 U9779 ( .A(n9928), .B(n9929), .Z(n9927) );
  XNOR2_X1 U9780 ( .A(n9924), .B(n9930), .ZN(n8855) );
  XOR2_X1 U9781 ( .A(n9923), .B(n9922), .Z(n9930) );
  OR2_X1 U9782 ( .A1(n9248), .A2(n7908), .ZN(n9922) );
  OR2_X1 U9783 ( .A1(n9931), .A2(n9932), .ZN(n9923) );
  AND2_X1 U9784 ( .A1(n9916), .A2(n9919), .ZN(n9932) );
  AND2_X1 U9785 ( .A1(n9933), .A2(n9918), .ZN(n9931) );
  OR2_X1 U9786 ( .A1(n9934), .A2(n9935), .ZN(n9918) );
  AND2_X1 U9787 ( .A1(n9912), .A2(n9915), .ZN(n9935) );
  AND2_X1 U9788 ( .A1(n9936), .A2(n9914), .ZN(n9934) );
  OR2_X1 U9789 ( .A1(n9937), .A2(n9938), .ZN(n9914) );
  AND2_X1 U9790 ( .A1(n9908), .A2(n9911), .ZN(n9938) );
  AND2_X1 U9791 ( .A1(n9939), .A2(n9910), .ZN(n9937) );
  OR2_X1 U9792 ( .A1(n9940), .A2(n9941), .ZN(n9910) );
  AND2_X1 U9793 ( .A1(n9904), .A2(n9907), .ZN(n9941) );
  AND2_X1 U9794 ( .A1(n9942), .A2(n9906), .ZN(n9940) );
  OR2_X1 U9795 ( .A1(n9943), .A2(n9944), .ZN(n9906) );
  AND2_X1 U9796 ( .A1(n9900), .A2(n9903), .ZN(n9944) );
  AND2_X1 U9797 ( .A1(n9945), .A2(n9902), .ZN(n9943) );
  OR2_X1 U9798 ( .A1(n9946), .A2(n9947), .ZN(n9902) );
  AND2_X1 U9799 ( .A1(n9896), .A2(n9899), .ZN(n9947) );
  AND2_X1 U9800 ( .A1(n9948), .A2(n9898), .ZN(n9946) );
  OR2_X1 U9801 ( .A1(n9949), .A2(n9950), .ZN(n9898) );
  AND2_X1 U9802 ( .A1(n9892), .A2(n9895), .ZN(n9950) );
  AND2_X1 U9803 ( .A1(n9951), .A2(n9894), .ZN(n9949) );
  OR2_X1 U9804 ( .A1(n9952), .A2(n9953), .ZN(n9894) );
  AND2_X1 U9805 ( .A1(n9888), .A2(n9891), .ZN(n9953) );
  AND2_X1 U9806 ( .A1(n9954), .A2(n9890), .ZN(n9952) );
  OR2_X1 U9807 ( .A1(n9955), .A2(n9956), .ZN(n9890) );
  AND2_X1 U9808 ( .A1(n9884), .A2(n9887), .ZN(n9956) );
  AND2_X1 U9809 ( .A1(n9957), .A2(n9886), .ZN(n9955) );
  OR2_X1 U9810 ( .A1(n9958), .A2(n9959), .ZN(n9886) );
  AND2_X1 U9811 ( .A1(n9880), .A2(n9883), .ZN(n9959) );
  AND2_X1 U9812 ( .A1(n9960), .A2(n9882), .ZN(n9958) );
  OR2_X1 U9813 ( .A1(n9961), .A2(n9962), .ZN(n9882) );
  AND2_X1 U9814 ( .A1(n9876), .A2(n9879), .ZN(n9962) );
  AND2_X1 U9815 ( .A1(n9963), .A2(n9878), .ZN(n9961) );
  OR2_X1 U9816 ( .A1(n9964), .A2(n9965), .ZN(n9878) );
  AND2_X1 U9817 ( .A1(n9872), .A2(n9875), .ZN(n9965) );
  AND2_X1 U9818 ( .A1(n9966), .A2(n9874), .ZN(n9964) );
  OR2_X1 U9819 ( .A1(n9967), .A2(n9968), .ZN(n9874) );
  AND2_X1 U9820 ( .A1(n9868), .A2(n9871), .ZN(n9968) );
  AND2_X1 U9821 ( .A1(n9969), .A2(n9870), .ZN(n9967) );
  OR2_X1 U9822 ( .A1(n9970), .A2(n9971), .ZN(n9870) );
  AND2_X1 U9823 ( .A1(n9864), .A2(n9867), .ZN(n9971) );
  AND2_X1 U9824 ( .A1(n9972), .A2(n9866), .ZN(n9970) );
  OR2_X1 U9825 ( .A1(n9973), .A2(n9974), .ZN(n9866) );
  AND2_X1 U9826 ( .A1(n9860), .A2(n9863), .ZN(n9974) );
  AND2_X1 U9827 ( .A1(n9975), .A2(n9862), .ZN(n9973) );
  OR2_X1 U9828 ( .A1(n9976), .A2(n9977), .ZN(n9862) );
  AND2_X1 U9829 ( .A1(n9856), .A2(n9859), .ZN(n9977) );
  AND2_X1 U9830 ( .A1(n9978), .A2(n9858), .ZN(n9976) );
  OR2_X1 U9831 ( .A1(n9979), .A2(n9980), .ZN(n9858) );
  AND2_X1 U9832 ( .A1(n9852), .A2(n9855), .ZN(n9980) );
  AND2_X1 U9833 ( .A1(n9981), .A2(n9854), .ZN(n9979) );
  OR2_X1 U9834 ( .A1(n9982), .A2(n9983), .ZN(n9854) );
  AND2_X1 U9835 ( .A1(n9848), .A2(n9851), .ZN(n9983) );
  AND2_X1 U9836 ( .A1(n9984), .A2(n9850), .ZN(n9982) );
  OR2_X1 U9837 ( .A1(n9985), .A2(n9986), .ZN(n9850) );
  AND2_X1 U9838 ( .A1(n9844), .A2(n9847), .ZN(n9986) );
  AND2_X1 U9839 ( .A1(n9987), .A2(n9846), .ZN(n9985) );
  OR2_X1 U9840 ( .A1(n9988), .A2(n9989), .ZN(n9846) );
  AND2_X1 U9841 ( .A1(n9840), .A2(n9843), .ZN(n9989) );
  AND2_X1 U9842 ( .A1(n9990), .A2(n9842), .ZN(n9988) );
  OR2_X1 U9843 ( .A1(n9991), .A2(n9992), .ZN(n9842) );
  AND2_X1 U9844 ( .A1(n9836), .A2(n9839), .ZN(n9992) );
  AND2_X1 U9845 ( .A1(n9993), .A2(n9838), .ZN(n9991) );
  OR2_X1 U9846 ( .A1(n9994), .A2(n9995), .ZN(n9838) );
  AND2_X1 U9847 ( .A1(n9832), .A2(n9835), .ZN(n9995) );
  AND2_X1 U9848 ( .A1(n9996), .A2(n9834), .ZN(n9994) );
  OR2_X1 U9849 ( .A1(n9997), .A2(n9998), .ZN(n9834) );
  AND2_X1 U9850 ( .A1(n9828), .A2(n9831), .ZN(n9998) );
  AND2_X1 U9851 ( .A1(n9999), .A2(n9830), .ZN(n9997) );
  OR2_X1 U9852 ( .A1(n10000), .A2(n10001), .ZN(n9830) );
  AND2_X1 U9853 ( .A1(n9824), .A2(n9827), .ZN(n10001) );
  AND2_X1 U9854 ( .A1(n10002), .A2(n9826), .ZN(n10000) );
  OR2_X1 U9855 ( .A1(n10003), .A2(n10004), .ZN(n9826) );
  AND2_X1 U9856 ( .A1(n9820), .A2(n9823), .ZN(n10004) );
  AND2_X1 U9857 ( .A1(n10005), .A2(n9822), .ZN(n10003) );
  OR2_X1 U9858 ( .A1(n10006), .A2(n10007), .ZN(n9822) );
  AND2_X1 U9859 ( .A1(n9816), .A2(n9819), .ZN(n10007) );
  AND2_X1 U9860 ( .A1(n10008), .A2(n9818), .ZN(n10006) );
  OR2_X1 U9861 ( .A1(n10009), .A2(n10010), .ZN(n9818) );
  AND2_X1 U9862 ( .A1(n9812), .A2(n9815), .ZN(n10010) );
  AND2_X1 U9863 ( .A1(n10011), .A2(n9814), .ZN(n10009) );
  OR2_X1 U9864 ( .A1(n10012), .A2(n10013), .ZN(n9814) );
  AND2_X1 U9865 ( .A1(n9808), .A2(n9811), .ZN(n10013) );
  AND2_X1 U9866 ( .A1(n10014), .A2(n9810), .ZN(n10012) );
  OR2_X1 U9867 ( .A1(n10015), .A2(n10016), .ZN(n9810) );
  AND2_X1 U9868 ( .A1(n9804), .A2(n9807), .ZN(n10016) );
  AND2_X1 U9869 ( .A1(n10017), .A2(n10018), .ZN(n10015) );
  OR2_X1 U9870 ( .A1(n9807), .A2(n9804), .ZN(n10018) );
  OR2_X1 U9871 ( .A1(n7954), .A2(n7908), .ZN(n9804) );
  OR3_X1 U9872 ( .A1(n7908), .A2(n8842), .A3(n9796), .ZN(n9807) );
  INV_X1 U9873 ( .A(n9806), .ZN(n10017) );
  OR2_X1 U9874 ( .A1(n10019), .A2(n10020), .ZN(n9806) );
  AND2_X1 U9875 ( .A1(b_29_), .A2(n10021), .ZN(n10020) );
  OR2_X1 U9876 ( .A1(n10022), .A2(n9801), .ZN(n10021) );
  AND2_X1 U9877 ( .A1(a_30_), .A2(n8838), .ZN(n10022) );
  AND2_X1 U9878 ( .A1(b_28_), .A2(n10023), .ZN(n10019) );
  OR2_X1 U9879 ( .A1(n10024), .A2(n7920), .ZN(n10023) );
  AND2_X1 U9880 ( .A1(a_31_), .A2(n8842), .ZN(n10024) );
  OR2_X1 U9881 ( .A1(n9811), .A2(n9808), .ZN(n10014) );
  XNOR2_X1 U9882 ( .A(n8843), .B(n10025), .ZN(n9808) );
  XOR2_X1 U9883 ( .A(n10026), .B(n10027), .Z(n10025) );
  OR2_X1 U9884 ( .A1(n7979), .A2(n7908), .ZN(n9811) );
  OR2_X1 U9885 ( .A1(n9815), .A2(n9812), .ZN(n10011) );
  XOR2_X1 U9886 ( .A(n10028), .B(n10029), .Z(n9812) );
  XOR2_X1 U9887 ( .A(n10030), .B(n10031), .Z(n10029) );
  OR2_X1 U9888 ( .A1(n8015), .A2(n7908), .ZN(n9815) );
  OR2_X1 U9889 ( .A1(n9819), .A2(n9816), .ZN(n10008) );
  XOR2_X1 U9890 ( .A(n10032), .B(n10033), .Z(n9816) );
  XOR2_X1 U9891 ( .A(n10034), .B(n10035), .Z(n10033) );
  OR2_X1 U9892 ( .A1(n8040), .A2(n7908), .ZN(n9819) );
  OR2_X1 U9893 ( .A1(n9823), .A2(n9820), .ZN(n10005) );
  XOR2_X1 U9894 ( .A(n10036), .B(n10037), .Z(n9820) );
  XOR2_X1 U9895 ( .A(n10038), .B(n10039), .Z(n10037) );
  OR2_X1 U9896 ( .A1(n8065), .A2(n7908), .ZN(n9823) );
  OR2_X1 U9897 ( .A1(n9827), .A2(n9824), .ZN(n10002) );
  XOR2_X1 U9898 ( .A(n10040), .B(n10041), .Z(n9824) );
  XOR2_X1 U9899 ( .A(n10042), .B(n10043), .Z(n10041) );
  OR2_X1 U9900 ( .A1(n8090), .A2(n7908), .ZN(n9827) );
  OR2_X1 U9901 ( .A1(n9831), .A2(n9828), .ZN(n9999) );
  XOR2_X1 U9902 ( .A(n10044), .B(n10045), .Z(n9828) );
  XOR2_X1 U9903 ( .A(n10046), .B(n10047), .Z(n10045) );
  OR2_X1 U9904 ( .A1(n8115), .A2(n7908), .ZN(n9831) );
  OR2_X1 U9905 ( .A1(n9835), .A2(n9832), .ZN(n9996) );
  XOR2_X1 U9906 ( .A(n10048), .B(n10049), .Z(n9832) );
  XOR2_X1 U9907 ( .A(n10050), .B(n10051), .Z(n10049) );
  OR2_X1 U9908 ( .A1(n8140), .A2(n7908), .ZN(n9835) );
  OR2_X1 U9909 ( .A1(n9839), .A2(n9836), .ZN(n9993) );
  XOR2_X1 U9910 ( .A(n10052), .B(n10053), .Z(n9836) );
  XOR2_X1 U9911 ( .A(n10054), .B(n10055), .Z(n10053) );
  OR2_X1 U9912 ( .A1(n8810), .A2(n7908), .ZN(n9839) );
  OR2_X1 U9913 ( .A1(n9843), .A2(n9840), .ZN(n9990) );
  XOR2_X1 U9914 ( .A(n10056), .B(n10057), .Z(n9840) );
  XOR2_X1 U9915 ( .A(n10058), .B(n10059), .Z(n10057) );
  OR2_X1 U9916 ( .A1(n8806), .A2(n7908), .ZN(n9843) );
  OR2_X1 U9917 ( .A1(n9847), .A2(n9844), .ZN(n9987) );
  XOR2_X1 U9918 ( .A(n10060), .B(n10061), .Z(n9844) );
  XOR2_X1 U9919 ( .A(n10062), .B(n10063), .Z(n10061) );
  OR2_X1 U9920 ( .A1(n8802), .A2(n7908), .ZN(n9847) );
  OR2_X1 U9921 ( .A1(n9851), .A2(n9848), .ZN(n9984) );
  XOR2_X1 U9922 ( .A(n10064), .B(n10065), .Z(n9848) );
  XOR2_X1 U9923 ( .A(n10066), .B(n10067), .Z(n10065) );
  OR2_X1 U9924 ( .A1(n8798), .A2(n7908), .ZN(n9851) );
  OR2_X1 U9925 ( .A1(n9855), .A2(n9852), .ZN(n9981) );
  XOR2_X1 U9926 ( .A(n10068), .B(n10069), .Z(n9852) );
  XOR2_X1 U9927 ( .A(n10070), .B(n10071), .Z(n10069) );
  OR2_X1 U9928 ( .A1(n8794), .A2(n7908), .ZN(n9855) );
  OR2_X1 U9929 ( .A1(n9859), .A2(n9856), .ZN(n9978) );
  XOR2_X1 U9930 ( .A(n10072), .B(n10073), .Z(n9856) );
  XOR2_X1 U9931 ( .A(n10074), .B(n10075), .Z(n10073) );
  OR2_X1 U9932 ( .A1(n8790), .A2(n7908), .ZN(n9859) );
  OR2_X1 U9933 ( .A1(n9863), .A2(n9860), .ZN(n9975) );
  XOR2_X1 U9934 ( .A(n10076), .B(n10077), .Z(n9860) );
  XOR2_X1 U9935 ( .A(n10078), .B(n10079), .Z(n10077) );
  OR2_X1 U9936 ( .A1(n8786), .A2(n7908), .ZN(n9863) );
  OR2_X1 U9937 ( .A1(n9867), .A2(n9864), .ZN(n9972) );
  XOR2_X1 U9938 ( .A(n10080), .B(n10081), .Z(n9864) );
  XOR2_X1 U9939 ( .A(n10082), .B(n10083), .Z(n10081) );
  OR2_X1 U9940 ( .A1(n8782), .A2(n7908), .ZN(n9867) );
  OR2_X1 U9941 ( .A1(n9871), .A2(n9868), .ZN(n9969) );
  XOR2_X1 U9942 ( .A(n10084), .B(n10085), .Z(n9868) );
  XOR2_X1 U9943 ( .A(n10086), .B(n10087), .Z(n10085) );
  OR2_X1 U9944 ( .A1(n8778), .A2(n7908), .ZN(n9871) );
  OR2_X1 U9945 ( .A1(n9875), .A2(n9872), .ZN(n9966) );
  XOR2_X1 U9946 ( .A(n10088), .B(n10089), .Z(n9872) );
  XOR2_X1 U9947 ( .A(n10090), .B(n10091), .Z(n10089) );
  OR2_X1 U9948 ( .A1(n8774), .A2(n7908), .ZN(n9875) );
  OR2_X1 U9949 ( .A1(n9879), .A2(n9876), .ZN(n9963) );
  XOR2_X1 U9950 ( .A(n10092), .B(n10093), .Z(n9876) );
  XOR2_X1 U9951 ( .A(n10094), .B(n10095), .Z(n10093) );
  OR2_X1 U9952 ( .A1(n8770), .A2(n7908), .ZN(n9879) );
  OR2_X1 U9953 ( .A1(n9883), .A2(n9880), .ZN(n9960) );
  XOR2_X1 U9954 ( .A(n10096), .B(n10097), .Z(n9880) );
  XOR2_X1 U9955 ( .A(n10098), .B(n10099), .Z(n10097) );
  OR2_X1 U9956 ( .A1(n8766), .A2(n7908), .ZN(n9883) );
  OR2_X1 U9957 ( .A1(n9887), .A2(n9884), .ZN(n9957) );
  XOR2_X1 U9958 ( .A(n10100), .B(n10101), .Z(n9884) );
  XOR2_X1 U9959 ( .A(n10102), .B(n10103), .Z(n10101) );
  OR2_X1 U9960 ( .A1(n8762), .A2(n7908), .ZN(n9887) );
  OR2_X1 U9961 ( .A1(n9891), .A2(n9888), .ZN(n9954) );
  XOR2_X1 U9962 ( .A(n10104), .B(n10105), .Z(n9888) );
  XOR2_X1 U9963 ( .A(n10106), .B(n10107), .Z(n10105) );
  OR2_X1 U9964 ( .A1(n8758), .A2(n7908), .ZN(n9891) );
  OR2_X1 U9965 ( .A1(n9895), .A2(n9892), .ZN(n9951) );
  XOR2_X1 U9966 ( .A(n10108), .B(n10109), .Z(n9892) );
  XOR2_X1 U9967 ( .A(n10110), .B(n10111), .Z(n10109) );
  OR2_X1 U9968 ( .A1(n8754), .A2(n7908), .ZN(n9895) );
  OR2_X1 U9969 ( .A1(n9899), .A2(n9896), .ZN(n9948) );
  XOR2_X1 U9970 ( .A(n10112), .B(n10113), .Z(n9896) );
  XOR2_X1 U9971 ( .A(n10114), .B(n10115), .Z(n10113) );
  OR2_X1 U9972 ( .A1(n8750), .A2(n7908), .ZN(n9899) );
  OR2_X1 U9973 ( .A1(n9903), .A2(n9900), .ZN(n9945) );
  XOR2_X1 U9974 ( .A(n10116), .B(n10117), .Z(n9900) );
  XOR2_X1 U9975 ( .A(n10118), .B(n10119), .Z(n10117) );
  OR2_X1 U9976 ( .A1(n8746), .A2(n7908), .ZN(n9903) );
  OR2_X1 U9977 ( .A1(n9907), .A2(n9904), .ZN(n9942) );
  XOR2_X1 U9978 ( .A(n10120), .B(n10121), .Z(n9904) );
  XOR2_X1 U9979 ( .A(n10122), .B(n10123), .Z(n10121) );
  OR2_X1 U9980 ( .A1(n8742), .A2(n7908), .ZN(n9907) );
  OR2_X1 U9981 ( .A1(n9911), .A2(n9908), .ZN(n9939) );
  XOR2_X1 U9982 ( .A(n10124), .B(n10125), .Z(n9908) );
  XOR2_X1 U9983 ( .A(n10126), .B(n10127), .Z(n10125) );
  OR2_X1 U9984 ( .A1(n8738), .A2(n7908), .ZN(n9911) );
  OR2_X1 U9985 ( .A1(n9915), .A2(n9912), .ZN(n9936) );
  XOR2_X1 U9986 ( .A(n10128), .B(n10129), .Z(n9912) );
  XOR2_X1 U9987 ( .A(n10130), .B(n10131), .Z(n10129) );
  OR2_X1 U9988 ( .A1(n8734), .A2(n7908), .ZN(n9915) );
  OR2_X1 U9989 ( .A1(n9919), .A2(n9916), .ZN(n9933) );
  XNOR2_X1 U9990 ( .A(n10132), .B(n10133), .ZN(n9916) );
  XNOR2_X1 U9991 ( .A(n10134), .B(n10135), .ZN(n10132) );
  OR2_X1 U9992 ( .A1(n8730), .A2(n7908), .ZN(n9919) );
  XOR2_X1 U9993 ( .A(n10136), .B(n10137), .Z(n9924) );
  XOR2_X1 U9994 ( .A(n10138), .B(n10139), .Z(n10137) );
  OR2_X1 U9995 ( .A1(n10140), .A2(n9695), .ZN(n8878) );
  XOR2_X1 U9996 ( .A(n9690), .B(n9691), .Z(n9695) );
  AND2_X1 U9997 ( .A1(n9696), .A2(n9694), .ZN(n10140) );
  XNOR2_X1 U9998 ( .A(n10141), .B(n10142), .ZN(n9694) );
  XOR2_X1 U9999 ( .A(n10143), .B(n10144), .Z(n10142) );
  INV_X1 U10000 ( .A(n9703), .ZN(n9696) );
  OR2_X1 U10001 ( .A1(n10145), .A2(n10146), .ZN(n9703) );
  AND2_X1 U10002 ( .A1(n9929), .A2(n9928), .ZN(n10146) );
  AND2_X1 U10003 ( .A1(n9926), .A2(n10147), .ZN(n10145) );
  OR2_X1 U10004 ( .A1(n9928), .A2(n9929), .ZN(n10147) );
  OR2_X1 U10005 ( .A1(n9248), .A2(n8842), .ZN(n9929) );
  OR2_X1 U10006 ( .A1(n10148), .A2(n10149), .ZN(n9928) );
  AND2_X1 U10007 ( .A1(n10139), .A2(n10138), .ZN(n10149) );
  AND2_X1 U10008 ( .A1(n10136), .A2(n10150), .ZN(n10148) );
  OR2_X1 U10009 ( .A1(n10138), .A2(n10139), .ZN(n10150) );
  OR2_X1 U10010 ( .A1(n8730), .A2(n8842), .ZN(n10139) );
  OR2_X1 U10011 ( .A1(n10151), .A2(n10152), .ZN(n10138) );
  AND2_X1 U10012 ( .A1(n10135), .A2(n10134), .ZN(n10152) );
  AND2_X1 U10013 ( .A1(n10133), .A2(n10153), .ZN(n10151) );
  OR2_X1 U10014 ( .A1(n10134), .A2(n10135), .ZN(n10153) );
  OR2_X1 U10015 ( .A1(n10154), .A2(n10155), .ZN(n10135) );
  AND2_X1 U10016 ( .A1(n10131), .A2(n10130), .ZN(n10155) );
  AND2_X1 U10017 ( .A1(n10128), .A2(n10156), .ZN(n10154) );
  OR2_X1 U10018 ( .A1(n10130), .A2(n10131), .ZN(n10156) );
  OR2_X1 U10019 ( .A1(n8738), .A2(n8842), .ZN(n10131) );
  OR2_X1 U10020 ( .A1(n10157), .A2(n10158), .ZN(n10130) );
  AND2_X1 U10021 ( .A1(n10127), .A2(n10126), .ZN(n10158) );
  AND2_X1 U10022 ( .A1(n10124), .A2(n10159), .ZN(n10157) );
  OR2_X1 U10023 ( .A1(n10126), .A2(n10127), .ZN(n10159) );
  OR2_X1 U10024 ( .A1(n8742), .A2(n8842), .ZN(n10127) );
  OR2_X1 U10025 ( .A1(n10160), .A2(n10161), .ZN(n10126) );
  AND2_X1 U10026 ( .A1(n10123), .A2(n10122), .ZN(n10161) );
  AND2_X1 U10027 ( .A1(n10120), .A2(n10162), .ZN(n10160) );
  OR2_X1 U10028 ( .A1(n10122), .A2(n10123), .ZN(n10162) );
  OR2_X1 U10029 ( .A1(n8746), .A2(n8842), .ZN(n10123) );
  OR2_X1 U10030 ( .A1(n10163), .A2(n10164), .ZN(n10122) );
  AND2_X1 U10031 ( .A1(n10119), .A2(n10118), .ZN(n10164) );
  AND2_X1 U10032 ( .A1(n10116), .A2(n10165), .ZN(n10163) );
  OR2_X1 U10033 ( .A1(n10118), .A2(n10119), .ZN(n10165) );
  OR2_X1 U10034 ( .A1(n8750), .A2(n8842), .ZN(n10119) );
  OR2_X1 U10035 ( .A1(n10166), .A2(n10167), .ZN(n10118) );
  AND2_X1 U10036 ( .A1(n10115), .A2(n10114), .ZN(n10167) );
  AND2_X1 U10037 ( .A1(n10112), .A2(n10168), .ZN(n10166) );
  OR2_X1 U10038 ( .A1(n10114), .A2(n10115), .ZN(n10168) );
  OR2_X1 U10039 ( .A1(n8754), .A2(n8842), .ZN(n10115) );
  OR2_X1 U10040 ( .A1(n10169), .A2(n10170), .ZN(n10114) );
  AND2_X1 U10041 ( .A1(n10111), .A2(n10110), .ZN(n10170) );
  AND2_X1 U10042 ( .A1(n10108), .A2(n10171), .ZN(n10169) );
  OR2_X1 U10043 ( .A1(n10110), .A2(n10111), .ZN(n10171) );
  OR2_X1 U10044 ( .A1(n8758), .A2(n8842), .ZN(n10111) );
  OR2_X1 U10045 ( .A1(n10172), .A2(n10173), .ZN(n10110) );
  AND2_X1 U10046 ( .A1(n10107), .A2(n10106), .ZN(n10173) );
  AND2_X1 U10047 ( .A1(n10104), .A2(n10174), .ZN(n10172) );
  OR2_X1 U10048 ( .A1(n10106), .A2(n10107), .ZN(n10174) );
  OR2_X1 U10049 ( .A1(n8762), .A2(n8842), .ZN(n10107) );
  OR2_X1 U10050 ( .A1(n10175), .A2(n10176), .ZN(n10106) );
  AND2_X1 U10051 ( .A1(n10103), .A2(n10102), .ZN(n10176) );
  AND2_X1 U10052 ( .A1(n10100), .A2(n10177), .ZN(n10175) );
  OR2_X1 U10053 ( .A1(n10102), .A2(n10103), .ZN(n10177) );
  OR2_X1 U10054 ( .A1(n8766), .A2(n8842), .ZN(n10103) );
  OR2_X1 U10055 ( .A1(n10178), .A2(n10179), .ZN(n10102) );
  AND2_X1 U10056 ( .A1(n10099), .A2(n10098), .ZN(n10179) );
  AND2_X1 U10057 ( .A1(n10096), .A2(n10180), .ZN(n10178) );
  OR2_X1 U10058 ( .A1(n10098), .A2(n10099), .ZN(n10180) );
  OR2_X1 U10059 ( .A1(n8770), .A2(n8842), .ZN(n10099) );
  OR2_X1 U10060 ( .A1(n10181), .A2(n10182), .ZN(n10098) );
  AND2_X1 U10061 ( .A1(n10095), .A2(n10094), .ZN(n10182) );
  AND2_X1 U10062 ( .A1(n10092), .A2(n10183), .ZN(n10181) );
  OR2_X1 U10063 ( .A1(n10094), .A2(n10095), .ZN(n10183) );
  OR2_X1 U10064 ( .A1(n8774), .A2(n8842), .ZN(n10095) );
  OR2_X1 U10065 ( .A1(n10184), .A2(n10185), .ZN(n10094) );
  AND2_X1 U10066 ( .A1(n10091), .A2(n10090), .ZN(n10185) );
  AND2_X1 U10067 ( .A1(n10088), .A2(n10186), .ZN(n10184) );
  OR2_X1 U10068 ( .A1(n10090), .A2(n10091), .ZN(n10186) );
  OR2_X1 U10069 ( .A1(n8778), .A2(n8842), .ZN(n10091) );
  OR2_X1 U10070 ( .A1(n10187), .A2(n10188), .ZN(n10090) );
  AND2_X1 U10071 ( .A1(n10087), .A2(n10086), .ZN(n10188) );
  AND2_X1 U10072 ( .A1(n10084), .A2(n10189), .ZN(n10187) );
  OR2_X1 U10073 ( .A1(n10086), .A2(n10087), .ZN(n10189) );
  OR2_X1 U10074 ( .A1(n8782), .A2(n8842), .ZN(n10087) );
  OR2_X1 U10075 ( .A1(n10190), .A2(n10191), .ZN(n10086) );
  AND2_X1 U10076 ( .A1(n10083), .A2(n10082), .ZN(n10191) );
  AND2_X1 U10077 ( .A1(n10080), .A2(n10192), .ZN(n10190) );
  OR2_X1 U10078 ( .A1(n10082), .A2(n10083), .ZN(n10192) );
  OR2_X1 U10079 ( .A1(n8786), .A2(n8842), .ZN(n10083) );
  OR2_X1 U10080 ( .A1(n10193), .A2(n10194), .ZN(n10082) );
  AND2_X1 U10081 ( .A1(n10079), .A2(n10078), .ZN(n10194) );
  AND2_X1 U10082 ( .A1(n10076), .A2(n10195), .ZN(n10193) );
  OR2_X1 U10083 ( .A1(n10078), .A2(n10079), .ZN(n10195) );
  OR2_X1 U10084 ( .A1(n8790), .A2(n8842), .ZN(n10079) );
  OR2_X1 U10085 ( .A1(n10196), .A2(n10197), .ZN(n10078) );
  AND2_X1 U10086 ( .A1(n10075), .A2(n10074), .ZN(n10197) );
  AND2_X1 U10087 ( .A1(n10072), .A2(n10198), .ZN(n10196) );
  OR2_X1 U10088 ( .A1(n10074), .A2(n10075), .ZN(n10198) );
  OR2_X1 U10089 ( .A1(n8794), .A2(n8842), .ZN(n10075) );
  OR2_X1 U10090 ( .A1(n10199), .A2(n10200), .ZN(n10074) );
  AND2_X1 U10091 ( .A1(n10071), .A2(n10070), .ZN(n10200) );
  AND2_X1 U10092 ( .A1(n10068), .A2(n10201), .ZN(n10199) );
  OR2_X1 U10093 ( .A1(n10070), .A2(n10071), .ZN(n10201) );
  OR2_X1 U10094 ( .A1(n8798), .A2(n8842), .ZN(n10071) );
  OR2_X1 U10095 ( .A1(n10202), .A2(n10203), .ZN(n10070) );
  AND2_X1 U10096 ( .A1(n10067), .A2(n10066), .ZN(n10203) );
  AND2_X1 U10097 ( .A1(n10064), .A2(n10204), .ZN(n10202) );
  OR2_X1 U10098 ( .A1(n10066), .A2(n10067), .ZN(n10204) );
  OR2_X1 U10099 ( .A1(n8802), .A2(n8842), .ZN(n10067) );
  OR2_X1 U10100 ( .A1(n10205), .A2(n10206), .ZN(n10066) );
  AND2_X1 U10101 ( .A1(n10063), .A2(n10062), .ZN(n10206) );
  AND2_X1 U10102 ( .A1(n10060), .A2(n10207), .ZN(n10205) );
  OR2_X1 U10103 ( .A1(n10062), .A2(n10063), .ZN(n10207) );
  OR2_X1 U10104 ( .A1(n8806), .A2(n8842), .ZN(n10063) );
  OR2_X1 U10105 ( .A1(n10208), .A2(n10209), .ZN(n10062) );
  AND2_X1 U10106 ( .A1(n10059), .A2(n10058), .ZN(n10209) );
  AND2_X1 U10107 ( .A1(n10056), .A2(n10210), .ZN(n10208) );
  OR2_X1 U10108 ( .A1(n10058), .A2(n10059), .ZN(n10210) );
  OR2_X1 U10109 ( .A1(n8810), .A2(n8842), .ZN(n10059) );
  OR2_X1 U10110 ( .A1(n10211), .A2(n10212), .ZN(n10058) );
  AND2_X1 U10111 ( .A1(n10055), .A2(n10054), .ZN(n10212) );
  AND2_X1 U10112 ( .A1(n10052), .A2(n10213), .ZN(n10211) );
  OR2_X1 U10113 ( .A1(n10054), .A2(n10055), .ZN(n10213) );
  OR2_X1 U10114 ( .A1(n8140), .A2(n8842), .ZN(n10055) );
  OR2_X1 U10115 ( .A1(n10214), .A2(n10215), .ZN(n10054) );
  AND2_X1 U10116 ( .A1(n10051), .A2(n10050), .ZN(n10215) );
  AND2_X1 U10117 ( .A1(n10048), .A2(n10216), .ZN(n10214) );
  OR2_X1 U10118 ( .A1(n10050), .A2(n10051), .ZN(n10216) );
  OR2_X1 U10119 ( .A1(n8115), .A2(n8842), .ZN(n10051) );
  OR2_X1 U10120 ( .A1(n10217), .A2(n10218), .ZN(n10050) );
  AND2_X1 U10121 ( .A1(n10047), .A2(n10046), .ZN(n10218) );
  AND2_X1 U10122 ( .A1(n10044), .A2(n10219), .ZN(n10217) );
  OR2_X1 U10123 ( .A1(n10046), .A2(n10047), .ZN(n10219) );
  OR2_X1 U10124 ( .A1(n8090), .A2(n8842), .ZN(n10047) );
  OR2_X1 U10125 ( .A1(n10220), .A2(n10221), .ZN(n10046) );
  AND2_X1 U10126 ( .A1(n10043), .A2(n10042), .ZN(n10221) );
  AND2_X1 U10127 ( .A1(n10040), .A2(n10222), .ZN(n10220) );
  OR2_X1 U10128 ( .A1(n10042), .A2(n10043), .ZN(n10222) );
  OR2_X1 U10129 ( .A1(n8065), .A2(n8842), .ZN(n10043) );
  OR2_X1 U10130 ( .A1(n10223), .A2(n10224), .ZN(n10042) );
  AND2_X1 U10131 ( .A1(n10039), .A2(n10038), .ZN(n10224) );
  AND2_X1 U10132 ( .A1(n10036), .A2(n10225), .ZN(n10223) );
  OR2_X1 U10133 ( .A1(n10038), .A2(n10039), .ZN(n10225) );
  OR2_X1 U10134 ( .A1(n8040), .A2(n8842), .ZN(n10039) );
  OR2_X1 U10135 ( .A1(n10226), .A2(n10227), .ZN(n10038) );
  AND2_X1 U10136 ( .A1(n10035), .A2(n10034), .ZN(n10227) );
  AND2_X1 U10137 ( .A1(n10032), .A2(n10228), .ZN(n10226) );
  OR2_X1 U10138 ( .A1(n10034), .A2(n10035), .ZN(n10228) );
  OR2_X1 U10139 ( .A1(n8015), .A2(n8842), .ZN(n10035) );
  OR2_X1 U10140 ( .A1(n10229), .A2(n10230), .ZN(n10034) );
  AND2_X1 U10141 ( .A1(n10031), .A2(n10030), .ZN(n10230) );
  AND2_X1 U10142 ( .A1(n10028), .A2(n10231), .ZN(n10229) );
  OR2_X1 U10143 ( .A1(n10030), .A2(n10031), .ZN(n10231) );
  OR2_X1 U10144 ( .A1(n7979), .A2(n8842), .ZN(n10031) );
  OR2_X1 U10145 ( .A1(n10232), .A2(n10233), .ZN(n10030) );
  AND2_X1 U10146 ( .A1(n8843), .A2(n10027), .ZN(n10233) );
  AND2_X1 U10147 ( .A1(n10234), .A2(n10235), .ZN(n10232) );
  OR2_X1 U10148 ( .A1(n10027), .A2(n8843), .ZN(n10235) );
  OR2_X1 U10149 ( .A1(n7954), .A2(n8842), .ZN(n8843) );
  OR3_X1 U10150 ( .A1(n8842), .A2(n8838), .A3(n9796), .ZN(n10027) );
  INV_X1 U10151 ( .A(n10026), .ZN(n10234) );
  OR2_X1 U10152 ( .A1(n10236), .A2(n10237), .ZN(n10026) );
  AND2_X1 U10153 ( .A1(b_28_), .A2(n10238), .ZN(n10237) );
  OR2_X1 U10154 ( .A1(n10239), .A2(n9801), .ZN(n10238) );
  AND2_X1 U10155 ( .A1(a_30_), .A2(n8834), .ZN(n10239) );
  AND2_X1 U10156 ( .A1(b_27_), .A2(n10240), .ZN(n10236) );
  OR2_X1 U10157 ( .A1(n10241), .A2(n7920), .ZN(n10240) );
  AND2_X1 U10158 ( .A1(a_31_), .A2(n8838), .ZN(n10241) );
  XNOR2_X1 U10159 ( .A(n10242), .B(n10243), .ZN(n10028) );
  XOR2_X1 U10160 ( .A(n10244), .B(n10245), .Z(n10243) );
  XOR2_X1 U10161 ( .A(n10246), .B(n10247), .Z(n10032) );
  XOR2_X1 U10162 ( .A(n10248), .B(n8839), .Z(n10247) );
  XOR2_X1 U10163 ( .A(n10249), .B(n10250), .Z(n10036) );
  XOR2_X1 U10164 ( .A(n10251), .B(n10252), .Z(n10250) );
  XOR2_X1 U10165 ( .A(n10253), .B(n10254), .Z(n10040) );
  XOR2_X1 U10166 ( .A(n10255), .B(n10256), .Z(n10254) );
  XOR2_X1 U10167 ( .A(n10257), .B(n10258), .Z(n10044) );
  XOR2_X1 U10168 ( .A(n10259), .B(n10260), .Z(n10258) );
  XOR2_X1 U10169 ( .A(n10261), .B(n10262), .Z(n10048) );
  XOR2_X1 U10170 ( .A(n10263), .B(n10264), .Z(n10262) );
  XOR2_X1 U10171 ( .A(n10265), .B(n10266), .Z(n10052) );
  XOR2_X1 U10172 ( .A(n10267), .B(n10268), .Z(n10266) );
  XOR2_X1 U10173 ( .A(n10269), .B(n10270), .Z(n10056) );
  XOR2_X1 U10174 ( .A(n10271), .B(n10272), .Z(n10270) );
  XOR2_X1 U10175 ( .A(n10273), .B(n10274), .Z(n10060) );
  XOR2_X1 U10176 ( .A(n10275), .B(n10276), .Z(n10274) );
  XOR2_X1 U10177 ( .A(n10277), .B(n10278), .Z(n10064) );
  XOR2_X1 U10178 ( .A(n10279), .B(n10280), .Z(n10278) );
  XOR2_X1 U10179 ( .A(n10281), .B(n10282), .Z(n10068) );
  XOR2_X1 U10180 ( .A(n10283), .B(n10284), .Z(n10282) );
  XOR2_X1 U10181 ( .A(n10285), .B(n10286), .Z(n10072) );
  XOR2_X1 U10182 ( .A(n10287), .B(n10288), .Z(n10286) );
  XOR2_X1 U10183 ( .A(n10289), .B(n10290), .Z(n10076) );
  XOR2_X1 U10184 ( .A(n10291), .B(n10292), .Z(n10290) );
  XOR2_X1 U10185 ( .A(n10293), .B(n10294), .Z(n10080) );
  XOR2_X1 U10186 ( .A(n10295), .B(n10296), .Z(n10294) );
  XOR2_X1 U10187 ( .A(n10297), .B(n10298), .Z(n10084) );
  XOR2_X1 U10188 ( .A(n10299), .B(n10300), .Z(n10298) );
  XOR2_X1 U10189 ( .A(n10301), .B(n10302), .Z(n10088) );
  XOR2_X1 U10190 ( .A(n10303), .B(n10304), .Z(n10302) );
  XOR2_X1 U10191 ( .A(n10305), .B(n10306), .Z(n10092) );
  XOR2_X1 U10192 ( .A(n10307), .B(n10308), .Z(n10306) );
  XOR2_X1 U10193 ( .A(n10309), .B(n10310), .Z(n10096) );
  XOR2_X1 U10194 ( .A(n10311), .B(n10312), .Z(n10310) );
  XOR2_X1 U10195 ( .A(n10313), .B(n10314), .Z(n10100) );
  XOR2_X1 U10196 ( .A(n10315), .B(n10316), .Z(n10314) );
  XOR2_X1 U10197 ( .A(n10317), .B(n10318), .Z(n10104) );
  XOR2_X1 U10198 ( .A(n10319), .B(n10320), .Z(n10318) );
  XOR2_X1 U10199 ( .A(n10321), .B(n10322), .Z(n10108) );
  XOR2_X1 U10200 ( .A(n10323), .B(n10324), .Z(n10322) );
  XOR2_X1 U10201 ( .A(n10325), .B(n10326), .Z(n10112) );
  XOR2_X1 U10202 ( .A(n10327), .B(n10328), .Z(n10326) );
  XOR2_X1 U10203 ( .A(n10329), .B(n10330), .Z(n10116) );
  XOR2_X1 U10204 ( .A(n10331), .B(n10332), .Z(n10330) );
  XOR2_X1 U10205 ( .A(n10333), .B(n10334), .Z(n10120) );
  XOR2_X1 U10206 ( .A(n10335), .B(n10336), .Z(n10334) );
  XOR2_X1 U10207 ( .A(n10337), .B(n10338), .Z(n10124) );
  XOR2_X1 U10208 ( .A(n10339), .B(n10340), .Z(n10338) );
  XOR2_X1 U10209 ( .A(n10341), .B(n10342), .Z(n10128) );
  XOR2_X1 U10210 ( .A(n10343), .B(n10344), .Z(n10342) );
  OR2_X1 U10211 ( .A1(n8734), .A2(n8842), .ZN(n10134) );
  XOR2_X1 U10212 ( .A(n10345), .B(n10346), .Z(n10133) );
  XOR2_X1 U10213 ( .A(n10347), .B(n10348), .Z(n10346) );
  XNOR2_X1 U10214 ( .A(n10349), .B(n10350), .ZN(n10136) );
  XNOR2_X1 U10215 ( .A(n10351), .B(n10352), .ZN(n10349) );
  XOR2_X1 U10216 ( .A(n10353), .B(n10354), .Z(n9926) );
  XOR2_X1 U10217 ( .A(n10355), .B(n10356), .Z(n10354) );
  OR2_X1 U10218 ( .A1(n10357), .A2(n9692), .ZN(n8885) );
  AND2_X1 U10219 ( .A1(n10358), .A2(n10359), .ZN(n9692) );
  INV_X1 U10220 ( .A(n10360), .ZN(n10358) );
  AND2_X1 U10221 ( .A1(n10361), .A2(n10362), .ZN(n10360) );
  AND2_X1 U10222 ( .A1(n9691), .A2(n9690), .ZN(n10357) );
  XNOR2_X1 U10223 ( .A(n10363), .B(n10364), .ZN(n9690) );
  XOR2_X1 U10224 ( .A(n10365), .B(n10366), .Z(n10364) );
  INV_X1 U10225 ( .A(n10367), .ZN(n9691) );
  OR2_X1 U10226 ( .A1(n10368), .A2(n10369), .ZN(n10367) );
  AND2_X1 U10227 ( .A1(n10144), .A2(n10143), .ZN(n10369) );
  AND2_X1 U10228 ( .A1(n10141), .A2(n10370), .ZN(n10368) );
  OR2_X1 U10229 ( .A1(n10143), .A2(n10144), .ZN(n10370) );
  OR2_X1 U10230 ( .A1(n9248), .A2(n8838), .ZN(n10144) );
  OR2_X1 U10231 ( .A1(n10371), .A2(n10372), .ZN(n10143) );
  AND2_X1 U10232 ( .A1(n10356), .A2(n10355), .ZN(n10372) );
  AND2_X1 U10233 ( .A1(n10353), .A2(n10373), .ZN(n10371) );
  OR2_X1 U10234 ( .A1(n10355), .A2(n10356), .ZN(n10373) );
  OR2_X1 U10235 ( .A1(n8730), .A2(n8838), .ZN(n10356) );
  OR2_X1 U10236 ( .A1(n10374), .A2(n10375), .ZN(n10355) );
  AND2_X1 U10237 ( .A1(n10352), .A2(n10351), .ZN(n10375) );
  AND2_X1 U10238 ( .A1(n10350), .A2(n10376), .ZN(n10374) );
  OR2_X1 U10239 ( .A1(n10351), .A2(n10352), .ZN(n10376) );
  OR2_X1 U10240 ( .A1(n10377), .A2(n10378), .ZN(n10352) );
  AND2_X1 U10241 ( .A1(n10348), .A2(n10347), .ZN(n10378) );
  AND2_X1 U10242 ( .A1(n10345), .A2(n10379), .ZN(n10377) );
  OR2_X1 U10243 ( .A1(n10347), .A2(n10348), .ZN(n10379) );
  OR2_X1 U10244 ( .A1(n8738), .A2(n8838), .ZN(n10348) );
  OR2_X1 U10245 ( .A1(n10380), .A2(n10381), .ZN(n10347) );
  AND2_X1 U10246 ( .A1(n10344), .A2(n10343), .ZN(n10381) );
  AND2_X1 U10247 ( .A1(n10341), .A2(n10382), .ZN(n10380) );
  OR2_X1 U10248 ( .A1(n10343), .A2(n10344), .ZN(n10382) );
  OR2_X1 U10249 ( .A1(n8742), .A2(n8838), .ZN(n10344) );
  OR2_X1 U10250 ( .A1(n10383), .A2(n10384), .ZN(n10343) );
  AND2_X1 U10251 ( .A1(n10340), .A2(n10339), .ZN(n10384) );
  AND2_X1 U10252 ( .A1(n10337), .A2(n10385), .ZN(n10383) );
  OR2_X1 U10253 ( .A1(n10339), .A2(n10340), .ZN(n10385) );
  OR2_X1 U10254 ( .A1(n8746), .A2(n8838), .ZN(n10340) );
  OR2_X1 U10255 ( .A1(n10386), .A2(n10387), .ZN(n10339) );
  AND2_X1 U10256 ( .A1(n10336), .A2(n10335), .ZN(n10387) );
  AND2_X1 U10257 ( .A1(n10333), .A2(n10388), .ZN(n10386) );
  OR2_X1 U10258 ( .A1(n10335), .A2(n10336), .ZN(n10388) );
  OR2_X1 U10259 ( .A1(n8750), .A2(n8838), .ZN(n10336) );
  OR2_X1 U10260 ( .A1(n10389), .A2(n10390), .ZN(n10335) );
  AND2_X1 U10261 ( .A1(n10332), .A2(n10331), .ZN(n10390) );
  AND2_X1 U10262 ( .A1(n10329), .A2(n10391), .ZN(n10389) );
  OR2_X1 U10263 ( .A1(n10331), .A2(n10332), .ZN(n10391) );
  OR2_X1 U10264 ( .A1(n8754), .A2(n8838), .ZN(n10332) );
  OR2_X1 U10265 ( .A1(n10392), .A2(n10393), .ZN(n10331) );
  AND2_X1 U10266 ( .A1(n10328), .A2(n10327), .ZN(n10393) );
  AND2_X1 U10267 ( .A1(n10325), .A2(n10394), .ZN(n10392) );
  OR2_X1 U10268 ( .A1(n10327), .A2(n10328), .ZN(n10394) );
  OR2_X1 U10269 ( .A1(n8758), .A2(n8838), .ZN(n10328) );
  OR2_X1 U10270 ( .A1(n10395), .A2(n10396), .ZN(n10327) );
  AND2_X1 U10271 ( .A1(n10324), .A2(n10323), .ZN(n10396) );
  AND2_X1 U10272 ( .A1(n10321), .A2(n10397), .ZN(n10395) );
  OR2_X1 U10273 ( .A1(n10323), .A2(n10324), .ZN(n10397) );
  OR2_X1 U10274 ( .A1(n8762), .A2(n8838), .ZN(n10324) );
  OR2_X1 U10275 ( .A1(n10398), .A2(n10399), .ZN(n10323) );
  AND2_X1 U10276 ( .A1(n10320), .A2(n10319), .ZN(n10399) );
  AND2_X1 U10277 ( .A1(n10317), .A2(n10400), .ZN(n10398) );
  OR2_X1 U10278 ( .A1(n10319), .A2(n10320), .ZN(n10400) );
  OR2_X1 U10279 ( .A1(n8766), .A2(n8838), .ZN(n10320) );
  OR2_X1 U10280 ( .A1(n10401), .A2(n10402), .ZN(n10319) );
  AND2_X1 U10281 ( .A1(n10316), .A2(n10315), .ZN(n10402) );
  AND2_X1 U10282 ( .A1(n10313), .A2(n10403), .ZN(n10401) );
  OR2_X1 U10283 ( .A1(n10315), .A2(n10316), .ZN(n10403) );
  OR2_X1 U10284 ( .A1(n8770), .A2(n8838), .ZN(n10316) );
  OR2_X1 U10285 ( .A1(n10404), .A2(n10405), .ZN(n10315) );
  AND2_X1 U10286 ( .A1(n10312), .A2(n10311), .ZN(n10405) );
  AND2_X1 U10287 ( .A1(n10309), .A2(n10406), .ZN(n10404) );
  OR2_X1 U10288 ( .A1(n10311), .A2(n10312), .ZN(n10406) );
  OR2_X1 U10289 ( .A1(n8774), .A2(n8838), .ZN(n10312) );
  OR2_X1 U10290 ( .A1(n10407), .A2(n10408), .ZN(n10311) );
  AND2_X1 U10291 ( .A1(n10308), .A2(n10307), .ZN(n10408) );
  AND2_X1 U10292 ( .A1(n10305), .A2(n10409), .ZN(n10407) );
  OR2_X1 U10293 ( .A1(n10307), .A2(n10308), .ZN(n10409) );
  OR2_X1 U10294 ( .A1(n8778), .A2(n8838), .ZN(n10308) );
  OR2_X1 U10295 ( .A1(n10410), .A2(n10411), .ZN(n10307) );
  AND2_X1 U10296 ( .A1(n10304), .A2(n10303), .ZN(n10411) );
  AND2_X1 U10297 ( .A1(n10301), .A2(n10412), .ZN(n10410) );
  OR2_X1 U10298 ( .A1(n10303), .A2(n10304), .ZN(n10412) );
  OR2_X1 U10299 ( .A1(n8782), .A2(n8838), .ZN(n10304) );
  OR2_X1 U10300 ( .A1(n10413), .A2(n10414), .ZN(n10303) );
  AND2_X1 U10301 ( .A1(n10300), .A2(n10299), .ZN(n10414) );
  AND2_X1 U10302 ( .A1(n10297), .A2(n10415), .ZN(n10413) );
  OR2_X1 U10303 ( .A1(n10299), .A2(n10300), .ZN(n10415) );
  OR2_X1 U10304 ( .A1(n8786), .A2(n8838), .ZN(n10300) );
  OR2_X1 U10305 ( .A1(n10416), .A2(n10417), .ZN(n10299) );
  AND2_X1 U10306 ( .A1(n10296), .A2(n10295), .ZN(n10417) );
  AND2_X1 U10307 ( .A1(n10293), .A2(n10418), .ZN(n10416) );
  OR2_X1 U10308 ( .A1(n10295), .A2(n10296), .ZN(n10418) );
  OR2_X1 U10309 ( .A1(n8790), .A2(n8838), .ZN(n10296) );
  OR2_X1 U10310 ( .A1(n10419), .A2(n10420), .ZN(n10295) );
  AND2_X1 U10311 ( .A1(n10292), .A2(n10291), .ZN(n10420) );
  AND2_X1 U10312 ( .A1(n10289), .A2(n10421), .ZN(n10419) );
  OR2_X1 U10313 ( .A1(n10291), .A2(n10292), .ZN(n10421) );
  OR2_X1 U10314 ( .A1(n8794), .A2(n8838), .ZN(n10292) );
  OR2_X1 U10315 ( .A1(n10422), .A2(n10423), .ZN(n10291) );
  AND2_X1 U10316 ( .A1(n10288), .A2(n10287), .ZN(n10423) );
  AND2_X1 U10317 ( .A1(n10285), .A2(n10424), .ZN(n10422) );
  OR2_X1 U10318 ( .A1(n10287), .A2(n10288), .ZN(n10424) );
  OR2_X1 U10319 ( .A1(n8798), .A2(n8838), .ZN(n10288) );
  OR2_X1 U10320 ( .A1(n10425), .A2(n10426), .ZN(n10287) );
  AND2_X1 U10321 ( .A1(n10284), .A2(n10283), .ZN(n10426) );
  AND2_X1 U10322 ( .A1(n10281), .A2(n10427), .ZN(n10425) );
  OR2_X1 U10323 ( .A1(n10283), .A2(n10284), .ZN(n10427) );
  OR2_X1 U10324 ( .A1(n8802), .A2(n8838), .ZN(n10284) );
  OR2_X1 U10325 ( .A1(n10428), .A2(n10429), .ZN(n10283) );
  AND2_X1 U10326 ( .A1(n10280), .A2(n10279), .ZN(n10429) );
  AND2_X1 U10327 ( .A1(n10277), .A2(n10430), .ZN(n10428) );
  OR2_X1 U10328 ( .A1(n10279), .A2(n10280), .ZN(n10430) );
  OR2_X1 U10329 ( .A1(n8806), .A2(n8838), .ZN(n10280) );
  OR2_X1 U10330 ( .A1(n10431), .A2(n10432), .ZN(n10279) );
  AND2_X1 U10331 ( .A1(n10276), .A2(n10275), .ZN(n10432) );
  AND2_X1 U10332 ( .A1(n10273), .A2(n10433), .ZN(n10431) );
  OR2_X1 U10333 ( .A1(n10275), .A2(n10276), .ZN(n10433) );
  OR2_X1 U10334 ( .A1(n8810), .A2(n8838), .ZN(n10276) );
  OR2_X1 U10335 ( .A1(n10434), .A2(n10435), .ZN(n10275) );
  AND2_X1 U10336 ( .A1(n10272), .A2(n10271), .ZN(n10435) );
  AND2_X1 U10337 ( .A1(n10269), .A2(n10436), .ZN(n10434) );
  OR2_X1 U10338 ( .A1(n10271), .A2(n10272), .ZN(n10436) );
  OR2_X1 U10339 ( .A1(n8140), .A2(n8838), .ZN(n10272) );
  OR2_X1 U10340 ( .A1(n10437), .A2(n10438), .ZN(n10271) );
  AND2_X1 U10341 ( .A1(n10268), .A2(n10267), .ZN(n10438) );
  AND2_X1 U10342 ( .A1(n10265), .A2(n10439), .ZN(n10437) );
  OR2_X1 U10343 ( .A1(n10267), .A2(n10268), .ZN(n10439) );
  OR2_X1 U10344 ( .A1(n8115), .A2(n8838), .ZN(n10268) );
  OR2_X1 U10345 ( .A1(n10440), .A2(n10441), .ZN(n10267) );
  AND2_X1 U10346 ( .A1(n10264), .A2(n10263), .ZN(n10441) );
  AND2_X1 U10347 ( .A1(n10261), .A2(n10442), .ZN(n10440) );
  OR2_X1 U10348 ( .A1(n10263), .A2(n10264), .ZN(n10442) );
  OR2_X1 U10349 ( .A1(n8090), .A2(n8838), .ZN(n10264) );
  OR2_X1 U10350 ( .A1(n10443), .A2(n10444), .ZN(n10263) );
  AND2_X1 U10351 ( .A1(n10260), .A2(n10259), .ZN(n10444) );
  AND2_X1 U10352 ( .A1(n10257), .A2(n10445), .ZN(n10443) );
  OR2_X1 U10353 ( .A1(n10259), .A2(n10260), .ZN(n10445) );
  OR2_X1 U10354 ( .A1(n8065), .A2(n8838), .ZN(n10260) );
  OR2_X1 U10355 ( .A1(n10446), .A2(n10447), .ZN(n10259) );
  AND2_X1 U10356 ( .A1(n10256), .A2(n10255), .ZN(n10447) );
  AND2_X1 U10357 ( .A1(n10253), .A2(n10448), .ZN(n10446) );
  OR2_X1 U10358 ( .A1(n10255), .A2(n10256), .ZN(n10448) );
  OR2_X1 U10359 ( .A1(n8040), .A2(n8838), .ZN(n10256) );
  OR2_X1 U10360 ( .A1(n10449), .A2(n10450), .ZN(n10255) );
  AND2_X1 U10361 ( .A1(n10252), .A2(n10251), .ZN(n10450) );
  AND2_X1 U10362 ( .A1(n10249), .A2(n10451), .ZN(n10449) );
  OR2_X1 U10363 ( .A1(n10251), .A2(n10252), .ZN(n10451) );
  OR2_X1 U10364 ( .A1(n8015), .A2(n8838), .ZN(n10252) );
  OR2_X1 U10365 ( .A1(n10452), .A2(n10453), .ZN(n10251) );
  AND2_X1 U10366 ( .A1(n8839), .A2(n10248), .ZN(n10453) );
  AND2_X1 U10367 ( .A1(n10246), .A2(n10454), .ZN(n10452) );
  OR2_X1 U10368 ( .A1(n10248), .A2(n8839), .ZN(n10454) );
  OR2_X1 U10369 ( .A1(n7979), .A2(n8838), .ZN(n8839) );
  OR2_X1 U10370 ( .A1(n10455), .A2(n10456), .ZN(n10248) );
  AND2_X1 U10371 ( .A1(n10242), .A2(n10245), .ZN(n10456) );
  AND2_X1 U10372 ( .A1(n10457), .A2(n10458), .ZN(n10455) );
  OR2_X1 U10373 ( .A1(n10245), .A2(n10242), .ZN(n10458) );
  OR2_X1 U10374 ( .A1(n7954), .A2(n8838), .ZN(n10242) );
  OR3_X1 U10375 ( .A1(n8838), .A2(n8834), .A3(n9796), .ZN(n10245) );
  INV_X1 U10376 ( .A(n10244), .ZN(n10457) );
  OR2_X1 U10377 ( .A1(n10459), .A2(n10460), .ZN(n10244) );
  AND2_X1 U10378 ( .A1(b_27_), .A2(n10461), .ZN(n10460) );
  OR2_X1 U10379 ( .A1(n10462), .A2(n9801), .ZN(n10461) );
  AND2_X1 U10380 ( .A1(a_30_), .A2(n8830), .ZN(n10462) );
  AND2_X1 U10381 ( .A1(b_26_), .A2(n10463), .ZN(n10459) );
  OR2_X1 U10382 ( .A1(n10464), .A2(n7920), .ZN(n10463) );
  AND2_X1 U10383 ( .A1(a_31_), .A2(n8834), .ZN(n10464) );
  XNOR2_X1 U10384 ( .A(n10465), .B(n10466), .ZN(n10246) );
  XOR2_X1 U10385 ( .A(n10467), .B(n10468), .Z(n10466) );
  XOR2_X1 U10386 ( .A(n10469), .B(n10470), .Z(n10249) );
  XOR2_X1 U10387 ( .A(n10471), .B(n10472), .Z(n10470) );
  XOR2_X1 U10388 ( .A(n10473), .B(n10474), .Z(n10253) );
  XOR2_X1 U10389 ( .A(n10475), .B(n8835), .Z(n10474) );
  XOR2_X1 U10390 ( .A(n10476), .B(n10477), .Z(n10257) );
  XOR2_X1 U10391 ( .A(n10478), .B(n10479), .Z(n10477) );
  XOR2_X1 U10392 ( .A(n10480), .B(n10481), .Z(n10261) );
  XOR2_X1 U10393 ( .A(n10482), .B(n10483), .Z(n10481) );
  XOR2_X1 U10394 ( .A(n10484), .B(n10485), .Z(n10265) );
  XOR2_X1 U10395 ( .A(n10486), .B(n10487), .Z(n10485) );
  XOR2_X1 U10396 ( .A(n10488), .B(n10489), .Z(n10269) );
  XOR2_X1 U10397 ( .A(n10490), .B(n10491), .Z(n10489) );
  XOR2_X1 U10398 ( .A(n10492), .B(n10493), .Z(n10273) );
  XOR2_X1 U10399 ( .A(n10494), .B(n10495), .Z(n10493) );
  XOR2_X1 U10400 ( .A(n10496), .B(n10497), .Z(n10277) );
  XOR2_X1 U10401 ( .A(n10498), .B(n10499), .Z(n10497) );
  XOR2_X1 U10402 ( .A(n10500), .B(n10501), .Z(n10281) );
  XOR2_X1 U10403 ( .A(n10502), .B(n10503), .Z(n10501) );
  XOR2_X1 U10404 ( .A(n10504), .B(n10505), .Z(n10285) );
  XOR2_X1 U10405 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR2_X1 U10406 ( .A(n10508), .B(n10509), .Z(n10289) );
  XOR2_X1 U10407 ( .A(n10510), .B(n10511), .Z(n10509) );
  XOR2_X1 U10408 ( .A(n10512), .B(n10513), .Z(n10293) );
  XOR2_X1 U10409 ( .A(n10514), .B(n10515), .Z(n10513) );
  XOR2_X1 U10410 ( .A(n10516), .B(n10517), .Z(n10297) );
  XOR2_X1 U10411 ( .A(n10518), .B(n10519), .Z(n10517) );
  XOR2_X1 U10412 ( .A(n10520), .B(n10521), .Z(n10301) );
  XOR2_X1 U10413 ( .A(n10522), .B(n10523), .Z(n10521) );
  XOR2_X1 U10414 ( .A(n10524), .B(n10525), .Z(n10305) );
  XOR2_X1 U10415 ( .A(n10526), .B(n10527), .Z(n10525) );
  XOR2_X1 U10416 ( .A(n10528), .B(n10529), .Z(n10309) );
  XOR2_X1 U10417 ( .A(n10530), .B(n10531), .Z(n10529) );
  XOR2_X1 U10418 ( .A(n10532), .B(n10533), .Z(n10313) );
  XOR2_X1 U10419 ( .A(n10534), .B(n10535), .Z(n10533) );
  XOR2_X1 U10420 ( .A(n10536), .B(n10537), .Z(n10317) );
  XOR2_X1 U10421 ( .A(n10538), .B(n10539), .Z(n10537) );
  XOR2_X1 U10422 ( .A(n10540), .B(n10541), .Z(n10321) );
  XOR2_X1 U10423 ( .A(n10542), .B(n10543), .Z(n10541) );
  XOR2_X1 U10424 ( .A(n10544), .B(n10545), .Z(n10325) );
  XOR2_X1 U10425 ( .A(n10546), .B(n10547), .Z(n10545) );
  XOR2_X1 U10426 ( .A(n10548), .B(n10549), .Z(n10329) );
  XOR2_X1 U10427 ( .A(n10550), .B(n10551), .Z(n10549) );
  XOR2_X1 U10428 ( .A(n10552), .B(n10553), .Z(n10333) );
  XOR2_X1 U10429 ( .A(n10554), .B(n10555), .Z(n10553) );
  XNOR2_X1 U10430 ( .A(n10556), .B(n10557), .ZN(n10337) );
  XNOR2_X1 U10431 ( .A(n10558), .B(n10559), .ZN(n10556) );
  XOR2_X1 U10432 ( .A(n10560), .B(n10561), .Z(n10341) );
  XOR2_X1 U10433 ( .A(n10562), .B(n10563), .Z(n10561) );
  XOR2_X1 U10434 ( .A(n10564), .B(n10565), .Z(n10345) );
  XOR2_X1 U10435 ( .A(n10566), .B(n10567), .Z(n10565) );
  OR2_X1 U10436 ( .A1(n8734), .A2(n8838), .ZN(n10351) );
  XOR2_X1 U10437 ( .A(n10568), .B(n10569), .Z(n10350) );
  XOR2_X1 U10438 ( .A(n10570), .B(n10571), .Z(n10569) );
  XNOR2_X1 U10439 ( .A(n10572), .B(n10573), .ZN(n10353) );
  XNOR2_X1 U10440 ( .A(n10574), .B(n10575), .ZN(n10572) );
  XOR2_X1 U10441 ( .A(n10576), .B(n10577), .Z(n10141) );
  XOR2_X1 U10442 ( .A(n10578), .B(n10579), .Z(n10577) );
  OR2_X1 U10443 ( .A1(n9688), .A2(n9687), .ZN(n8892) );
  XOR2_X1 U10444 ( .A(n9683), .B(n9685), .Z(n9687) );
  INV_X1 U10445 ( .A(n10359), .ZN(n9688) );
  OR2_X1 U10446 ( .A1(n10361), .A2(n10362), .ZN(n10359) );
  OR2_X1 U10447 ( .A1(n10580), .A2(n10581), .ZN(n10362) );
  AND2_X1 U10448 ( .A1(n10363), .A2(n10366), .ZN(n10581) );
  AND2_X1 U10449 ( .A1(n10582), .A2(n10365), .ZN(n10580) );
  OR2_X1 U10450 ( .A1(n10583), .A2(n10584), .ZN(n10365) );
  AND2_X1 U10451 ( .A1(n10576), .A2(n10579), .ZN(n10584) );
  AND2_X1 U10452 ( .A1(n10585), .A2(n10578), .ZN(n10583) );
  OR2_X1 U10453 ( .A1(n10586), .A2(n10587), .ZN(n10578) );
  AND2_X1 U10454 ( .A1(n10575), .A2(n10574), .ZN(n10587) );
  AND2_X1 U10455 ( .A1(n10573), .A2(n10588), .ZN(n10586) );
  OR2_X1 U10456 ( .A1(n10574), .A2(n10575), .ZN(n10588) );
  OR2_X1 U10457 ( .A1(n10589), .A2(n10590), .ZN(n10575) );
  AND2_X1 U10458 ( .A1(n10571), .A2(n10570), .ZN(n10590) );
  AND2_X1 U10459 ( .A1(n10568), .A2(n10591), .ZN(n10589) );
  OR2_X1 U10460 ( .A1(n10570), .A2(n10571), .ZN(n10591) );
  OR2_X1 U10461 ( .A1(n8738), .A2(n8834), .ZN(n10571) );
  OR2_X1 U10462 ( .A1(n10592), .A2(n10593), .ZN(n10570) );
  AND2_X1 U10463 ( .A1(n10567), .A2(n10566), .ZN(n10593) );
  AND2_X1 U10464 ( .A1(n10564), .A2(n10594), .ZN(n10592) );
  OR2_X1 U10465 ( .A1(n10566), .A2(n10567), .ZN(n10594) );
  OR2_X1 U10466 ( .A1(n8742), .A2(n8834), .ZN(n10567) );
  OR2_X1 U10467 ( .A1(n10595), .A2(n10596), .ZN(n10566) );
  AND2_X1 U10468 ( .A1(n10563), .A2(n10562), .ZN(n10596) );
  AND2_X1 U10469 ( .A1(n10560), .A2(n10597), .ZN(n10595) );
  OR2_X1 U10470 ( .A1(n10562), .A2(n10563), .ZN(n10597) );
  OR2_X1 U10471 ( .A1(n8746), .A2(n8834), .ZN(n10563) );
  OR2_X1 U10472 ( .A1(n10598), .A2(n10599), .ZN(n10562) );
  AND2_X1 U10473 ( .A1(n10559), .A2(n10558), .ZN(n10599) );
  AND2_X1 U10474 ( .A1(n10557), .A2(n10600), .ZN(n10598) );
  OR2_X1 U10475 ( .A1(n10558), .A2(n10559), .ZN(n10600) );
  OR2_X1 U10476 ( .A1(n10601), .A2(n10602), .ZN(n10559) );
  AND2_X1 U10477 ( .A1(n10555), .A2(n10554), .ZN(n10602) );
  AND2_X1 U10478 ( .A1(n10552), .A2(n10603), .ZN(n10601) );
  OR2_X1 U10479 ( .A1(n10554), .A2(n10555), .ZN(n10603) );
  OR2_X1 U10480 ( .A1(n8754), .A2(n8834), .ZN(n10555) );
  OR2_X1 U10481 ( .A1(n10604), .A2(n10605), .ZN(n10554) );
  AND2_X1 U10482 ( .A1(n10551), .A2(n10550), .ZN(n10605) );
  AND2_X1 U10483 ( .A1(n10548), .A2(n10606), .ZN(n10604) );
  OR2_X1 U10484 ( .A1(n10550), .A2(n10551), .ZN(n10606) );
  OR2_X1 U10485 ( .A1(n8758), .A2(n8834), .ZN(n10551) );
  OR2_X1 U10486 ( .A1(n10607), .A2(n10608), .ZN(n10550) );
  AND2_X1 U10487 ( .A1(n10547), .A2(n10546), .ZN(n10608) );
  AND2_X1 U10488 ( .A1(n10544), .A2(n10609), .ZN(n10607) );
  OR2_X1 U10489 ( .A1(n10546), .A2(n10547), .ZN(n10609) );
  OR2_X1 U10490 ( .A1(n8762), .A2(n8834), .ZN(n10547) );
  OR2_X1 U10491 ( .A1(n10610), .A2(n10611), .ZN(n10546) );
  AND2_X1 U10492 ( .A1(n10543), .A2(n10542), .ZN(n10611) );
  AND2_X1 U10493 ( .A1(n10540), .A2(n10612), .ZN(n10610) );
  OR2_X1 U10494 ( .A1(n10542), .A2(n10543), .ZN(n10612) );
  OR2_X1 U10495 ( .A1(n8766), .A2(n8834), .ZN(n10543) );
  OR2_X1 U10496 ( .A1(n10613), .A2(n10614), .ZN(n10542) );
  AND2_X1 U10497 ( .A1(n10539), .A2(n10538), .ZN(n10614) );
  AND2_X1 U10498 ( .A1(n10536), .A2(n10615), .ZN(n10613) );
  OR2_X1 U10499 ( .A1(n10538), .A2(n10539), .ZN(n10615) );
  OR2_X1 U10500 ( .A1(n8770), .A2(n8834), .ZN(n10539) );
  OR2_X1 U10501 ( .A1(n10616), .A2(n10617), .ZN(n10538) );
  AND2_X1 U10502 ( .A1(n10535), .A2(n10534), .ZN(n10617) );
  AND2_X1 U10503 ( .A1(n10532), .A2(n10618), .ZN(n10616) );
  OR2_X1 U10504 ( .A1(n10534), .A2(n10535), .ZN(n10618) );
  OR2_X1 U10505 ( .A1(n8774), .A2(n8834), .ZN(n10535) );
  OR2_X1 U10506 ( .A1(n10619), .A2(n10620), .ZN(n10534) );
  AND2_X1 U10507 ( .A1(n10531), .A2(n10530), .ZN(n10620) );
  AND2_X1 U10508 ( .A1(n10528), .A2(n10621), .ZN(n10619) );
  OR2_X1 U10509 ( .A1(n10530), .A2(n10531), .ZN(n10621) );
  OR2_X1 U10510 ( .A1(n8778), .A2(n8834), .ZN(n10531) );
  OR2_X1 U10511 ( .A1(n10622), .A2(n10623), .ZN(n10530) );
  AND2_X1 U10512 ( .A1(n10527), .A2(n10526), .ZN(n10623) );
  AND2_X1 U10513 ( .A1(n10524), .A2(n10624), .ZN(n10622) );
  OR2_X1 U10514 ( .A1(n10526), .A2(n10527), .ZN(n10624) );
  OR2_X1 U10515 ( .A1(n8782), .A2(n8834), .ZN(n10527) );
  OR2_X1 U10516 ( .A1(n10625), .A2(n10626), .ZN(n10526) );
  AND2_X1 U10517 ( .A1(n10523), .A2(n10522), .ZN(n10626) );
  AND2_X1 U10518 ( .A1(n10520), .A2(n10627), .ZN(n10625) );
  OR2_X1 U10519 ( .A1(n10522), .A2(n10523), .ZN(n10627) );
  OR2_X1 U10520 ( .A1(n8786), .A2(n8834), .ZN(n10523) );
  OR2_X1 U10521 ( .A1(n10628), .A2(n10629), .ZN(n10522) );
  AND2_X1 U10522 ( .A1(n10519), .A2(n10518), .ZN(n10629) );
  AND2_X1 U10523 ( .A1(n10516), .A2(n10630), .ZN(n10628) );
  OR2_X1 U10524 ( .A1(n10518), .A2(n10519), .ZN(n10630) );
  OR2_X1 U10525 ( .A1(n8790), .A2(n8834), .ZN(n10519) );
  OR2_X1 U10526 ( .A1(n10631), .A2(n10632), .ZN(n10518) );
  AND2_X1 U10527 ( .A1(n10515), .A2(n10514), .ZN(n10632) );
  AND2_X1 U10528 ( .A1(n10512), .A2(n10633), .ZN(n10631) );
  OR2_X1 U10529 ( .A1(n10514), .A2(n10515), .ZN(n10633) );
  OR2_X1 U10530 ( .A1(n8794), .A2(n8834), .ZN(n10515) );
  OR2_X1 U10531 ( .A1(n10634), .A2(n10635), .ZN(n10514) );
  AND2_X1 U10532 ( .A1(n10511), .A2(n10510), .ZN(n10635) );
  AND2_X1 U10533 ( .A1(n10508), .A2(n10636), .ZN(n10634) );
  OR2_X1 U10534 ( .A1(n10510), .A2(n10511), .ZN(n10636) );
  OR2_X1 U10535 ( .A1(n8798), .A2(n8834), .ZN(n10511) );
  OR2_X1 U10536 ( .A1(n10637), .A2(n10638), .ZN(n10510) );
  AND2_X1 U10537 ( .A1(n10507), .A2(n10506), .ZN(n10638) );
  AND2_X1 U10538 ( .A1(n10504), .A2(n10639), .ZN(n10637) );
  OR2_X1 U10539 ( .A1(n10506), .A2(n10507), .ZN(n10639) );
  OR2_X1 U10540 ( .A1(n8802), .A2(n8834), .ZN(n10507) );
  OR2_X1 U10541 ( .A1(n10640), .A2(n10641), .ZN(n10506) );
  AND2_X1 U10542 ( .A1(n10503), .A2(n10502), .ZN(n10641) );
  AND2_X1 U10543 ( .A1(n10500), .A2(n10642), .ZN(n10640) );
  OR2_X1 U10544 ( .A1(n10502), .A2(n10503), .ZN(n10642) );
  OR2_X1 U10545 ( .A1(n8806), .A2(n8834), .ZN(n10503) );
  OR2_X1 U10546 ( .A1(n10643), .A2(n10644), .ZN(n10502) );
  AND2_X1 U10547 ( .A1(n10499), .A2(n10498), .ZN(n10644) );
  AND2_X1 U10548 ( .A1(n10496), .A2(n10645), .ZN(n10643) );
  OR2_X1 U10549 ( .A1(n10498), .A2(n10499), .ZN(n10645) );
  OR2_X1 U10550 ( .A1(n8810), .A2(n8834), .ZN(n10499) );
  OR2_X1 U10551 ( .A1(n10646), .A2(n10647), .ZN(n10498) );
  AND2_X1 U10552 ( .A1(n10495), .A2(n10494), .ZN(n10647) );
  AND2_X1 U10553 ( .A1(n10492), .A2(n10648), .ZN(n10646) );
  OR2_X1 U10554 ( .A1(n10494), .A2(n10495), .ZN(n10648) );
  OR2_X1 U10555 ( .A1(n8140), .A2(n8834), .ZN(n10495) );
  OR2_X1 U10556 ( .A1(n10649), .A2(n10650), .ZN(n10494) );
  AND2_X1 U10557 ( .A1(n10491), .A2(n10490), .ZN(n10650) );
  AND2_X1 U10558 ( .A1(n10488), .A2(n10651), .ZN(n10649) );
  OR2_X1 U10559 ( .A1(n10490), .A2(n10491), .ZN(n10651) );
  OR2_X1 U10560 ( .A1(n8115), .A2(n8834), .ZN(n10491) );
  OR2_X1 U10561 ( .A1(n10652), .A2(n10653), .ZN(n10490) );
  AND2_X1 U10562 ( .A1(n10487), .A2(n10486), .ZN(n10653) );
  AND2_X1 U10563 ( .A1(n10484), .A2(n10654), .ZN(n10652) );
  OR2_X1 U10564 ( .A1(n10486), .A2(n10487), .ZN(n10654) );
  OR2_X1 U10565 ( .A1(n8090), .A2(n8834), .ZN(n10487) );
  OR2_X1 U10566 ( .A1(n10655), .A2(n10656), .ZN(n10486) );
  AND2_X1 U10567 ( .A1(n10483), .A2(n10482), .ZN(n10656) );
  AND2_X1 U10568 ( .A1(n10480), .A2(n10657), .ZN(n10655) );
  OR2_X1 U10569 ( .A1(n10482), .A2(n10483), .ZN(n10657) );
  OR2_X1 U10570 ( .A1(n8065), .A2(n8834), .ZN(n10483) );
  OR2_X1 U10571 ( .A1(n10658), .A2(n10659), .ZN(n10482) );
  AND2_X1 U10572 ( .A1(n10479), .A2(n10478), .ZN(n10659) );
  AND2_X1 U10573 ( .A1(n10476), .A2(n10660), .ZN(n10658) );
  OR2_X1 U10574 ( .A1(n10478), .A2(n10479), .ZN(n10660) );
  OR2_X1 U10575 ( .A1(n8040), .A2(n8834), .ZN(n10479) );
  OR2_X1 U10576 ( .A1(n10661), .A2(n10662), .ZN(n10478) );
  AND2_X1 U10577 ( .A1(n8835), .A2(n10475), .ZN(n10662) );
  AND2_X1 U10578 ( .A1(n10473), .A2(n10663), .ZN(n10661) );
  OR2_X1 U10579 ( .A1(n10475), .A2(n8835), .ZN(n10663) );
  OR2_X1 U10580 ( .A1(n8015), .A2(n8834), .ZN(n8835) );
  OR2_X1 U10581 ( .A1(n10664), .A2(n10665), .ZN(n10475) );
  AND2_X1 U10582 ( .A1(n10472), .A2(n10471), .ZN(n10665) );
  AND2_X1 U10583 ( .A1(n10469), .A2(n10666), .ZN(n10664) );
  OR2_X1 U10584 ( .A1(n10471), .A2(n10472), .ZN(n10666) );
  OR2_X1 U10585 ( .A1(n7979), .A2(n8834), .ZN(n10472) );
  OR2_X1 U10586 ( .A1(n10667), .A2(n10668), .ZN(n10471) );
  AND2_X1 U10587 ( .A1(n10465), .A2(n10468), .ZN(n10668) );
  AND2_X1 U10588 ( .A1(n10669), .A2(n10670), .ZN(n10667) );
  OR2_X1 U10589 ( .A1(n10468), .A2(n10465), .ZN(n10670) );
  OR2_X1 U10590 ( .A1(n7954), .A2(n8834), .ZN(n10465) );
  OR3_X1 U10591 ( .A1(n8834), .A2(n8830), .A3(n9796), .ZN(n10468) );
  INV_X1 U10592 ( .A(n10467), .ZN(n10669) );
  OR2_X1 U10593 ( .A1(n10671), .A2(n10672), .ZN(n10467) );
  AND2_X1 U10594 ( .A1(b_26_), .A2(n10673), .ZN(n10672) );
  OR2_X1 U10595 ( .A1(n10674), .A2(n9801), .ZN(n10673) );
  AND2_X1 U10596 ( .A1(a_30_), .A2(n8826), .ZN(n10674) );
  AND2_X1 U10597 ( .A1(b_25_), .A2(n10675), .ZN(n10671) );
  OR2_X1 U10598 ( .A1(n10676), .A2(n7920), .ZN(n10675) );
  AND2_X1 U10599 ( .A1(a_31_), .A2(n8830), .ZN(n10676) );
  XNOR2_X1 U10600 ( .A(n10677), .B(n10678), .ZN(n10469) );
  XOR2_X1 U10601 ( .A(n10679), .B(n10680), .Z(n10678) );
  XOR2_X1 U10602 ( .A(n10681), .B(n10682), .Z(n10473) );
  XOR2_X1 U10603 ( .A(n10683), .B(n10684), .Z(n10682) );
  XOR2_X1 U10604 ( .A(n10685), .B(n10686), .Z(n10476) );
  XOR2_X1 U10605 ( .A(n10687), .B(n10688), .Z(n10686) );
  XOR2_X1 U10606 ( .A(n10689), .B(n10690), .Z(n10480) );
  XOR2_X1 U10607 ( .A(n10691), .B(n8831), .Z(n10690) );
  XOR2_X1 U10608 ( .A(n10692), .B(n10693), .Z(n10484) );
  XOR2_X1 U10609 ( .A(n10694), .B(n10695), .Z(n10693) );
  XOR2_X1 U10610 ( .A(n10696), .B(n10697), .Z(n10488) );
  XOR2_X1 U10611 ( .A(n10698), .B(n10699), .Z(n10697) );
  XOR2_X1 U10612 ( .A(n10700), .B(n10701), .Z(n10492) );
  XOR2_X1 U10613 ( .A(n10702), .B(n10703), .Z(n10701) );
  XOR2_X1 U10614 ( .A(n10704), .B(n10705), .Z(n10496) );
  XOR2_X1 U10615 ( .A(n10706), .B(n10707), .Z(n10705) );
  XOR2_X1 U10616 ( .A(n10708), .B(n10709), .Z(n10500) );
  XOR2_X1 U10617 ( .A(n10710), .B(n10711), .Z(n10709) );
  XOR2_X1 U10618 ( .A(n10712), .B(n10713), .Z(n10504) );
  XOR2_X1 U10619 ( .A(n10714), .B(n10715), .Z(n10713) );
  XOR2_X1 U10620 ( .A(n10716), .B(n10717), .Z(n10508) );
  XOR2_X1 U10621 ( .A(n10718), .B(n10719), .Z(n10717) );
  XOR2_X1 U10622 ( .A(n10720), .B(n10721), .Z(n10512) );
  XOR2_X1 U10623 ( .A(n10722), .B(n10723), .Z(n10721) );
  XOR2_X1 U10624 ( .A(n10724), .B(n10725), .Z(n10516) );
  XOR2_X1 U10625 ( .A(n10726), .B(n10727), .Z(n10725) );
  XOR2_X1 U10626 ( .A(n10728), .B(n10729), .Z(n10520) );
  XOR2_X1 U10627 ( .A(n10730), .B(n10731), .Z(n10729) );
  XOR2_X1 U10628 ( .A(n10732), .B(n10733), .Z(n10524) );
  XOR2_X1 U10629 ( .A(n10734), .B(n10735), .Z(n10733) );
  XOR2_X1 U10630 ( .A(n10736), .B(n10737), .Z(n10528) );
  XOR2_X1 U10631 ( .A(n10738), .B(n10739), .Z(n10737) );
  XOR2_X1 U10632 ( .A(n10740), .B(n10741), .Z(n10532) );
  XOR2_X1 U10633 ( .A(n10742), .B(n10743), .Z(n10741) );
  XOR2_X1 U10634 ( .A(n10744), .B(n10745), .Z(n10536) );
  XOR2_X1 U10635 ( .A(n10746), .B(n10747), .Z(n10745) );
  XOR2_X1 U10636 ( .A(n10748), .B(n10749), .Z(n10540) );
  XOR2_X1 U10637 ( .A(n10750), .B(n10751), .Z(n10749) );
  XOR2_X1 U10638 ( .A(n10752), .B(n10753), .Z(n10544) );
  XOR2_X1 U10639 ( .A(n10754), .B(n10755), .Z(n10753) );
  XOR2_X1 U10640 ( .A(n10756), .B(n10757), .Z(n10548) );
  XOR2_X1 U10641 ( .A(n10758), .B(n10759), .Z(n10757) );
  XOR2_X1 U10642 ( .A(n10760), .B(n10761), .Z(n10552) );
  XOR2_X1 U10643 ( .A(n10762), .B(n10763), .Z(n10761) );
  OR2_X1 U10644 ( .A1(n8750), .A2(n8834), .ZN(n10558) );
  XOR2_X1 U10645 ( .A(n10764), .B(n10765), .Z(n10557) );
  XOR2_X1 U10646 ( .A(n10766), .B(n10767), .Z(n10765) );
  XNOR2_X1 U10647 ( .A(n10768), .B(n10769), .ZN(n10560) );
  XNOR2_X1 U10648 ( .A(n10770), .B(n10771), .ZN(n10768) );
  XOR2_X1 U10649 ( .A(n10772), .B(n10773), .Z(n10564) );
  XOR2_X1 U10650 ( .A(n10774), .B(n10775), .Z(n10773) );
  XOR2_X1 U10651 ( .A(n10776), .B(n10777), .Z(n10568) );
  XOR2_X1 U10652 ( .A(n10778), .B(n10779), .Z(n10777) );
  OR2_X1 U10653 ( .A1(n8734), .A2(n8834), .ZN(n10574) );
  XOR2_X1 U10654 ( .A(n10780), .B(n10781), .Z(n10573) );
  XOR2_X1 U10655 ( .A(n10782), .B(n10783), .Z(n10781) );
  OR2_X1 U10656 ( .A1(n10576), .A2(n10579), .ZN(n10585) );
  OR2_X1 U10657 ( .A1(n8730), .A2(n8834), .ZN(n10579) );
  XOR2_X1 U10658 ( .A(n10784), .B(n10785), .Z(n10576) );
  XOR2_X1 U10659 ( .A(n10786), .B(n10787), .Z(n10785) );
  OR2_X1 U10660 ( .A1(n10363), .A2(n10366), .ZN(n10582) );
  OR2_X1 U10661 ( .A1(n9248), .A2(n8834), .ZN(n10366) );
  XOR2_X1 U10662 ( .A(n10788), .B(n10789), .Z(n10363) );
  XOR2_X1 U10663 ( .A(n10790), .B(n10791), .Z(n10789) );
  XOR2_X1 U10664 ( .A(n10792), .B(n10793), .Z(n10361) );
  XOR2_X1 U10665 ( .A(n10794), .B(n10795), .Z(n10793) );
  OR2_X1 U10666 ( .A1(n10796), .A2(n9684), .ZN(n8900) );
  XOR2_X1 U10667 ( .A(n9660), .B(n9662), .Z(n9684) );
  OR2_X1 U10668 ( .A1(n10797), .A2(n10798), .ZN(n9662) );
  AND2_X1 U10669 ( .A1(n10799), .A2(n10800), .ZN(n10798) );
  AND2_X1 U10670 ( .A1(n10801), .A2(n10802), .ZN(n10797) );
  OR2_X1 U10671 ( .A1(n10799), .A2(n10800), .ZN(n10802) );
  XOR2_X1 U10672 ( .A(n9669), .B(n10803), .Z(n9660) );
  XOR2_X1 U10673 ( .A(n9668), .B(n9667), .Z(n10803) );
  OR2_X1 U10674 ( .A1(n9248), .A2(n8822), .ZN(n9667) );
  OR2_X1 U10675 ( .A1(n10804), .A2(n10805), .ZN(n9668) );
  AND2_X1 U10676 ( .A1(n10806), .A2(n10807), .ZN(n10805) );
  AND2_X1 U10677 ( .A1(n10808), .A2(n10809), .ZN(n10804) );
  OR2_X1 U10678 ( .A1(n10806), .A2(n10807), .ZN(n10809) );
  XOR2_X1 U10679 ( .A(n9676), .B(n10810), .Z(n9669) );
  XOR2_X1 U10680 ( .A(n9675), .B(n9674), .Z(n10810) );
  OR2_X1 U10681 ( .A1(n8730), .A2(n8818), .ZN(n9674) );
  OR2_X1 U10682 ( .A1(n10811), .A2(n10812), .ZN(n9675) );
  AND2_X1 U10683 ( .A1(n10813), .A2(n10814), .ZN(n10812) );
  AND2_X1 U10684 ( .A1(n10815), .A2(n10816), .ZN(n10811) );
  OR2_X1 U10685 ( .A1(n10813), .A2(n10814), .ZN(n10816) );
  XOR2_X1 U10686 ( .A(n10817), .B(n10818), .Z(n9676) );
  XOR2_X1 U10687 ( .A(n10819), .B(n10820), .Z(n10818) );
  AND2_X1 U10688 ( .A1(n9685), .A2(n9683), .ZN(n10796) );
  XNOR2_X1 U10689 ( .A(n10801), .B(n10821), .ZN(n9683) );
  XOR2_X1 U10690 ( .A(n10800), .B(n10799), .Z(n10821) );
  OR2_X1 U10691 ( .A1(n9248), .A2(n8826), .ZN(n10799) );
  OR2_X1 U10692 ( .A1(n10822), .A2(n10823), .ZN(n10800) );
  AND2_X1 U10693 ( .A1(n10824), .A2(n10825), .ZN(n10823) );
  AND2_X1 U10694 ( .A1(n10826), .A2(n10827), .ZN(n10822) );
  OR2_X1 U10695 ( .A1(n10824), .A2(n10825), .ZN(n10827) );
  XNOR2_X1 U10696 ( .A(n10828), .B(n10808), .ZN(n10801) );
  XOR2_X1 U10697 ( .A(n10815), .B(n10829), .Z(n10808) );
  XOR2_X1 U10698 ( .A(n10814), .B(n10813), .Z(n10829) );
  OR2_X1 U10699 ( .A1(n8734), .A2(n8818), .ZN(n10813) );
  OR2_X1 U10700 ( .A1(n10830), .A2(n10831), .ZN(n10814) );
  AND2_X1 U10701 ( .A1(n10832), .A2(n10833), .ZN(n10831) );
  AND2_X1 U10702 ( .A1(n10834), .A2(n10835), .ZN(n10830) );
  OR2_X1 U10703 ( .A1(n10832), .A2(n10833), .ZN(n10835) );
  XOR2_X1 U10704 ( .A(n10836), .B(n10837), .Z(n10815) );
  XOR2_X1 U10705 ( .A(n10838), .B(n10839), .Z(n10837) );
  XNOR2_X1 U10706 ( .A(n10807), .B(n10806), .ZN(n10828) );
  OR2_X1 U10707 ( .A1(n10840), .A2(n10841), .ZN(n10806) );
  AND2_X1 U10708 ( .A1(n10842), .A2(n10843), .ZN(n10841) );
  AND2_X1 U10709 ( .A1(n10844), .A2(n10845), .ZN(n10840) );
  OR2_X1 U10710 ( .A1(n10842), .A2(n10843), .ZN(n10845) );
  OR2_X1 U10711 ( .A1(n8730), .A2(n8822), .ZN(n10807) );
  INV_X1 U10712 ( .A(n10846), .ZN(n9685) );
  OR2_X1 U10713 ( .A1(n10847), .A2(n10848), .ZN(n10846) );
  AND2_X1 U10714 ( .A1(n10795), .A2(n10794), .ZN(n10848) );
  AND2_X1 U10715 ( .A1(n10792), .A2(n10849), .ZN(n10847) );
  OR2_X1 U10716 ( .A1(n10794), .A2(n10795), .ZN(n10849) );
  OR2_X1 U10717 ( .A1(n9248), .A2(n8830), .ZN(n10795) );
  OR2_X1 U10718 ( .A1(n10850), .A2(n10851), .ZN(n10794) );
  AND2_X1 U10719 ( .A1(n10791), .A2(n10790), .ZN(n10851) );
  AND2_X1 U10720 ( .A1(n10788), .A2(n10852), .ZN(n10850) );
  OR2_X1 U10721 ( .A1(n10790), .A2(n10791), .ZN(n10852) );
  OR2_X1 U10722 ( .A1(n8730), .A2(n8830), .ZN(n10791) );
  OR2_X1 U10723 ( .A1(n10853), .A2(n10854), .ZN(n10790) );
  AND2_X1 U10724 ( .A1(n10787), .A2(n10786), .ZN(n10854) );
  AND2_X1 U10725 ( .A1(n10784), .A2(n10855), .ZN(n10853) );
  OR2_X1 U10726 ( .A1(n10786), .A2(n10787), .ZN(n10855) );
  OR2_X1 U10727 ( .A1(n8734), .A2(n8830), .ZN(n10787) );
  OR2_X1 U10728 ( .A1(n10856), .A2(n10857), .ZN(n10786) );
  AND2_X1 U10729 ( .A1(n10783), .A2(n10782), .ZN(n10857) );
  AND2_X1 U10730 ( .A1(n10780), .A2(n10858), .ZN(n10856) );
  OR2_X1 U10731 ( .A1(n10782), .A2(n10783), .ZN(n10858) );
  OR2_X1 U10732 ( .A1(n8738), .A2(n8830), .ZN(n10783) );
  OR2_X1 U10733 ( .A1(n10859), .A2(n10860), .ZN(n10782) );
  AND2_X1 U10734 ( .A1(n10779), .A2(n10778), .ZN(n10860) );
  AND2_X1 U10735 ( .A1(n10776), .A2(n10861), .ZN(n10859) );
  OR2_X1 U10736 ( .A1(n10778), .A2(n10779), .ZN(n10861) );
  OR2_X1 U10737 ( .A1(n8742), .A2(n8830), .ZN(n10779) );
  OR2_X1 U10738 ( .A1(n10862), .A2(n10863), .ZN(n10778) );
  AND2_X1 U10739 ( .A1(n10775), .A2(n10774), .ZN(n10863) );
  AND2_X1 U10740 ( .A1(n10772), .A2(n10864), .ZN(n10862) );
  OR2_X1 U10741 ( .A1(n10774), .A2(n10775), .ZN(n10864) );
  OR2_X1 U10742 ( .A1(n8746), .A2(n8830), .ZN(n10775) );
  OR2_X1 U10743 ( .A1(n10865), .A2(n10866), .ZN(n10774) );
  AND2_X1 U10744 ( .A1(n10771), .A2(n10770), .ZN(n10866) );
  AND2_X1 U10745 ( .A1(n10769), .A2(n10867), .ZN(n10865) );
  OR2_X1 U10746 ( .A1(n10770), .A2(n10771), .ZN(n10867) );
  OR2_X1 U10747 ( .A1(n10868), .A2(n10869), .ZN(n10771) );
  AND2_X1 U10748 ( .A1(n10767), .A2(n10766), .ZN(n10869) );
  AND2_X1 U10749 ( .A1(n10764), .A2(n10870), .ZN(n10868) );
  OR2_X1 U10750 ( .A1(n10766), .A2(n10767), .ZN(n10870) );
  OR2_X1 U10751 ( .A1(n8754), .A2(n8830), .ZN(n10767) );
  OR2_X1 U10752 ( .A1(n10871), .A2(n10872), .ZN(n10766) );
  AND2_X1 U10753 ( .A1(n10763), .A2(n10762), .ZN(n10872) );
  AND2_X1 U10754 ( .A1(n10760), .A2(n10873), .ZN(n10871) );
  OR2_X1 U10755 ( .A1(n10762), .A2(n10763), .ZN(n10873) );
  OR2_X1 U10756 ( .A1(n8758), .A2(n8830), .ZN(n10763) );
  OR2_X1 U10757 ( .A1(n10874), .A2(n10875), .ZN(n10762) );
  AND2_X1 U10758 ( .A1(n10759), .A2(n10758), .ZN(n10875) );
  AND2_X1 U10759 ( .A1(n10756), .A2(n10876), .ZN(n10874) );
  OR2_X1 U10760 ( .A1(n10758), .A2(n10759), .ZN(n10876) );
  OR2_X1 U10761 ( .A1(n8762), .A2(n8830), .ZN(n10759) );
  OR2_X1 U10762 ( .A1(n10877), .A2(n10878), .ZN(n10758) );
  AND2_X1 U10763 ( .A1(n10755), .A2(n10754), .ZN(n10878) );
  AND2_X1 U10764 ( .A1(n10752), .A2(n10879), .ZN(n10877) );
  OR2_X1 U10765 ( .A1(n10754), .A2(n10755), .ZN(n10879) );
  OR2_X1 U10766 ( .A1(n8766), .A2(n8830), .ZN(n10755) );
  OR2_X1 U10767 ( .A1(n10880), .A2(n10881), .ZN(n10754) );
  AND2_X1 U10768 ( .A1(n10751), .A2(n10750), .ZN(n10881) );
  AND2_X1 U10769 ( .A1(n10748), .A2(n10882), .ZN(n10880) );
  OR2_X1 U10770 ( .A1(n10750), .A2(n10751), .ZN(n10882) );
  OR2_X1 U10771 ( .A1(n8770), .A2(n8830), .ZN(n10751) );
  OR2_X1 U10772 ( .A1(n10883), .A2(n10884), .ZN(n10750) );
  AND2_X1 U10773 ( .A1(n10747), .A2(n10746), .ZN(n10884) );
  AND2_X1 U10774 ( .A1(n10744), .A2(n10885), .ZN(n10883) );
  OR2_X1 U10775 ( .A1(n10746), .A2(n10747), .ZN(n10885) );
  OR2_X1 U10776 ( .A1(n8774), .A2(n8830), .ZN(n10747) );
  OR2_X1 U10777 ( .A1(n10886), .A2(n10887), .ZN(n10746) );
  AND2_X1 U10778 ( .A1(n10743), .A2(n10742), .ZN(n10887) );
  AND2_X1 U10779 ( .A1(n10740), .A2(n10888), .ZN(n10886) );
  OR2_X1 U10780 ( .A1(n10742), .A2(n10743), .ZN(n10888) );
  OR2_X1 U10781 ( .A1(n8778), .A2(n8830), .ZN(n10743) );
  OR2_X1 U10782 ( .A1(n10889), .A2(n10890), .ZN(n10742) );
  AND2_X1 U10783 ( .A1(n10739), .A2(n10738), .ZN(n10890) );
  AND2_X1 U10784 ( .A1(n10736), .A2(n10891), .ZN(n10889) );
  OR2_X1 U10785 ( .A1(n10738), .A2(n10739), .ZN(n10891) );
  OR2_X1 U10786 ( .A1(n8782), .A2(n8830), .ZN(n10739) );
  OR2_X1 U10787 ( .A1(n10892), .A2(n10893), .ZN(n10738) );
  AND2_X1 U10788 ( .A1(n10735), .A2(n10734), .ZN(n10893) );
  AND2_X1 U10789 ( .A1(n10732), .A2(n10894), .ZN(n10892) );
  OR2_X1 U10790 ( .A1(n10734), .A2(n10735), .ZN(n10894) );
  OR2_X1 U10791 ( .A1(n8786), .A2(n8830), .ZN(n10735) );
  OR2_X1 U10792 ( .A1(n10895), .A2(n10896), .ZN(n10734) );
  AND2_X1 U10793 ( .A1(n10731), .A2(n10730), .ZN(n10896) );
  AND2_X1 U10794 ( .A1(n10728), .A2(n10897), .ZN(n10895) );
  OR2_X1 U10795 ( .A1(n10730), .A2(n10731), .ZN(n10897) );
  OR2_X1 U10796 ( .A1(n8790), .A2(n8830), .ZN(n10731) );
  OR2_X1 U10797 ( .A1(n10898), .A2(n10899), .ZN(n10730) );
  AND2_X1 U10798 ( .A1(n10727), .A2(n10726), .ZN(n10899) );
  AND2_X1 U10799 ( .A1(n10724), .A2(n10900), .ZN(n10898) );
  OR2_X1 U10800 ( .A1(n10726), .A2(n10727), .ZN(n10900) );
  OR2_X1 U10801 ( .A1(n8794), .A2(n8830), .ZN(n10727) );
  OR2_X1 U10802 ( .A1(n10901), .A2(n10902), .ZN(n10726) );
  AND2_X1 U10803 ( .A1(n10723), .A2(n10722), .ZN(n10902) );
  AND2_X1 U10804 ( .A1(n10720), .A2(n10903), .ZN(n10901) );
  OR2_X1 U10805 ( .A1(n10722), .A2(n10723), .ZN(n10903) );
  OR2_X1 U10806 ( .A1(n8798), .A2(n8830), .ZN(n10723) );
  OR2_X1 U10807 ( .A1(n10904), .A2(n10905), .ZN(n10722) );
  AND2_X1 U10808 ( .A1(n10719), .A2(n10718), .ZN(n10905) );
  AND2_X1 U10809 ( .A1(n10716), .A2(n10906), .ZN(n10904) );
  OR2_X1 U10810 ( .A1(n10718), .A2(n10719), .ZN(n10906) );
  OR2_X1 U10811 ( .A1(n8802), .A2(n8830), .ZN(n10719) );
  OR2_X1 U10812 ( .A1(n10907), .A2(n10908), .ZN(n10718) );
  AND2_X1 U10813 ( .A1(n10715), .A2(n10714), .ZN(n10908) );
  AND2_X1 U10814 ( .A1(n10712), .A2(n10909), .ZN(n10907) );
  OR2_X1 U10815 ( .A1(n10714), .A2(n10715), .ZN(n10909) );
  OR2_X1 U10816 ( .A1(n8806), .A2(n8830), .ZN(n10715) );
  OR2_X1 U10817 ( .A1(n10910), .A2(n10911), .ZN(n10714) );
  AND2_X1 U10818 ( .A1(n10711), .A2(n10710), .ZN(n10911) );
  AND2_X1 U10819 ( .A1(n10708), .A2(n10912), .ZN(n10910) );
  OR2_X1 U10820 ( .A1(n10710), .A2(n10711), .ZN(n10912) );
  OR2_X1 U10821 ( .A1(n8810), .A2(n8830), .ZN(n10711) );
  OR2_X1 U10822 ( .A1(n10913), .A2(n10914), .ZN(n10710) );
  AND2_X1 U10823 ( .A1(n10707), .A2(n10706), .ZN(n10914) );
  AND2_X1 U10824 ( .A1(n10704), .A2(n10915), .ZN(n10913) );
  OR2_X1 U10825 ( .A1(n10706), .A2(n10707), .ZN(n10915) );
  OR2_X1 U10826 ( .A1(n8140), .A2(n8830), .ZN(n10707) );
  OR2_X1 U10827 ( .A1(n10916), .A2(n10917), .ZN(n10706) );
  AND2_X1 U10828 ( .A1(n10703), .A2(n10702), .ZN(n10917) );
  AND2_X1 U10829 ( .A1(n10700), .A2(n10918), .ZN(n10916) );
  OR2_X1 U10830 ( .A1(n10702), .A2(n10703), .ZN(n10918) );
  OR2_X1 U10831 ( .A1(n8115), .A2(n8830), .ZN(n10703) );
  OR2_X1 U10832 ( .A1(n10919), .A2(n10920), .ZN(n10702) );
  AND2_X1 U10833 ( .A1(n10699), .A2(n10698), .ZN(n10920) );
  AND2_X1 U10834 ( .A1(n10696), .A2(n10921), .ZN(n10919) );
  OR2_X1 U10835 ( .A1(n10698), .A2(n10699), .ZN(n10921) );
  OR2_X1 U10836 ( .A1(n8090), .A2(n8830), .ZN(n10699) );
  OR2_X1 U10837 ( .A1(n10922), .A2(n10923), .ZN(n10698) );
  AND2_X1 U10838 ( .A1(n10695), .A2(n10694), .ZN(n10923) );
  AND2_X1 U10839 ( .A1(n10692), .A2(n10924), .ZN(n10922) );
  OR2_X1 U10840 ( .A1(n10694), .A2(n10695), .ZN(n10924) );
  OR2_X1 U10841 ( .A1(n8065), .A2(n8830), .ZN(n10695) );
  OR2_X1 U10842 ( .A1(n10925), .A2(n10926), .ZN(n10694) );
  AND2_X1 U10843 ( .A1(n8831), .A2(n10691), .ZN(n10926) );
  AND2_X1 U10844 ( .A1(n10689), .A2(n10927), .ZN(n10925) );
  OR2_X1 U10845 ( .A1(n10691), .A2(n8831), .ZN(n10927) );
  OR2_X1 U10846 ( .A1(n8040), .A2(n8830), .ZN(n8831) );
  OR2_X1 U10847 ( .A1(n10928), .A2(n10929), .ZN(n10691) );
  AND2_X1 U10848 ( .A1(n10688), .A2(n10687), .ZN(n10929) );
  AND2_X1 U10849 ( .A1(n10685), .A2(n10930), .ZN(n10928) );
  OR2_X1 U10850 ( .A1(n10687), .A2(n10688), .ZN(n10930) );
  OR2_X1 U10851 ( .A1(n8015), .A2(n8830), .ZN(n10688) );
  OR2_X1 U10852 ( .A1(n10931), .A2(n10932), .ZN(n10687) );
  AND2_X1 U10853 ( .A1(n10684), .A2(n10683), .ZN(n10932) );
  AND2_X1 U10854 ( .A1(n10681), .A2(n10933), .ZN(n10931) );
  OR2_X1 U10855 ( .A1(n10683), .A2(n10684), .ZN(n10933) );
  OR2_X1 U10856 ( .A1(n7979), .A2(n8830), .ZN(n10684) );
  OR2_X1 U10857 ( .A1(n10934), .A2(n10935), .ZN(n10683) );
  AND2_X1 U10858 ( .A1(n10677), .A2(n10680), .ZN(n10935) );
  AND2_X1 U10859 ( .A1(n10936), .A2(n10937), .ZN(n10934) );
  OR2_X1 U10860 ( .A1(n10680), .A2(n10677), .ZN(n10937) );
  OR2_X1 U10861 ( .A1(n7954), .A2(n8830), .ZN(n10677) );
  OR3_X1 U10862 ( .A1(n8830), .A2(n8826), .A3(n9796), .ZN(n10680) );
  INV_X1 U10863 ( .A(n10679), .ZN(n10936) );
  OR2_X1 U10864 ( .A1(n10938), .A2(n10939), .ZN(n10679) );
  AND2_X1 U10865 ( .A1(b_25_), .A2(n10940), .ZN(n10939) );
  OR2_X1 U10866 ( .A1(n10941), .A2(n9801), .ZN(n10940) );
  AND2_X1 U10867 ( .A1(a_30_), .A2(n8822), .ZN(n10941) );
  AND2_X1 U10868 ( .A1(b_24_), .A2(n10942), .ZN(n10938) );
  OR2_X1 U10869 ( .A1(n10943), .A2(n7920), .ZN(n10942) );
  AND2_X1 U10870 ( .A1(a_31_), .A2(n8826), .ZN(n10943) );
  XNOR2_X1 U10871 ( .A(n10944), .B(n10945), .ZN(n10681) );
  XOR2_X1 U10872 ( .A(n10946), .B(n10947), .Z(n10945) );
  XOR2_X1 U10873 ( .A(n10948), .B(n10949), .Z(n10685) );
  XOR2_X1 U10874 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR2_X1 U10875 ( .A(n10952), .B(n10953), .Z(n10689) );
  XOR2_X1 U10876 ( .A(n10954), .B(n10955), .Z(n10953) );
  XOR2_X1 U10877 ( .A(n10956), .B(n10957), .Z(n10692) );
  XOR2_X1 U10878 ( .A(n10958), .B(n10959), .Z(n10957) );
  XOR2_X1 U10879 ( .A(n10960), .B(n10961), .Z(n10696) );
  XOR2_X1 U10880 ( .A(n10962), .B(n8827), .Z(n10961) );
  XOR2_X1 U10881 ( .A(n10963), .B(n10964), .Z(n10700) );
  XOR2_X1 U10882 ( .A(n10965), .B(n10966), .Z(n10964) );
  XOR2_X1 U10883 ( .A(n10967), .B(n10968), .Z(n10704) );
  XOR2_X1 U10884 ( .A(n10969), .B(n10970), .Z(n10968) );
  XOR2_X1 U10885 ( .A(n10971), .B(n10972), .Z(n10708) );
  XOR2_X1 U10886 ( .A(n10973), .B(n10974), .Z(n10972) );
  XOR2_X1 U10887 ( .A(n10975), .B(n10976), .Z(n10712) );
  XOR2_X1 U10888 ( .A(n10977), .B(n10978), .Z(n10976) );
  XOR2_X1 U10889 ( .A(n10979), .B(n10980), .Z(n10716) );
  XOR2_X1 U10890 ( .A(n10981), .B(n10982), .Z(n10980) );
  XOR2_X1 U10891 ( .A(n10983), .B(n10984), .Z(n10720) );
  XOR2_X1 U10892 ( .A(n10985), .B(n10986), .Z(n10984) );
  XOR2_X1 U10893 ( .A(n10987), .B(n10988), .Z(n10724) );
  XOR2_X1 U10894 ( .A(n10989), .B(n10990), .Z(n10988) );
  XOR2_X1 U10895 ( .A(n10991), .B(n10992), .Z(n10728) );
  XOR2_X1 U10896 ( .A(n10993), .B(n10994), .Z(n10992) );
  XOR2_X1 U10897 ( .A(n10995), .B(n10996), .Z(n10732) );
  XOR2_X1 U10898 ( .A(n10997), .B(n10998), .Z(n10996) );
  XOR2_X1 U10899 ( .A(n10999), .B(n11000), .Z(n10736) );
  XOR2_X1 U10900 ( .A(n11001), .B(n11002), .Z(n11000) );
  XOR2_X1 U10901 ( .A(n11003), .B(n11004), .Z(n10740) );
  XOR2_X1 U10902 ( .A(n11005), .B(n11006), .Z(n11004) );
  XOR2_X1 U10903 ( .A(n11007), .B(n11008), .Z(n10744) );
  XOR2_X1 U10904 ( .A(n11009), .B(n11010), .Z(n11008) );
  XOR2_X1 U10905 ( .A(n11011), .B(n11012), .Z(n10748) );
  XOR2_X1 U10906 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR2_X1 U10907 ( .A(n11015), .B(n11016), .Z(n10752) );
  XOR2_X1 U10908 ( .A(n11017), .B(n11018), .Z(n11016) );
  XNOR2_X1 U10909 ( .A(n11019), .B(n11020), .ZN(n10756) );
  XNOR2_X1 U10910 ( .A(n11021), .B(n11022), .ZN(n11019) );
  XOR2_X1 U10911 ( .A(n11023), .B(n11024), .Z(n10760) );
  XOR2_X1 U10912 ( .A(n11025), .B(n11026), .Z(n11024) );
  XOR2_X1 U10913 ( .A(n11027), .B(n11028), .Z(n10764) );
  XOR2_X1 U10914 ( .A(n11029), .B(n11030), .Z(n11028) );
  OR2_X1 U10915 ( .A1(n8750), .A2(n8830), .ZN(n10770) );
  XOR2_X1 U10916 ( .A(n11031), .B(n11032), .Z(n10769) );
  XOR2_X1 U10917 ( .A(n11033), .B(n11034), .Z(n11032) );
  XNOR2_X1 U10918 ( .A(n11035), .B(n11036), .ZN(n10772) );
  XNOR2_X1 U10919 ( .A(n11037), .B(n11038), .ZN(n11035) );
  XOR2_X1 U10920 ( .A(n11039), .B(n11040), .Z(n10776) );
  XOR2_X1 U10921 ( .A(n11041), .B(n11042), .Z(n11040) );
  XOR2_X1 U10922 ( .A(n11043), .B(n11044), .Z(n10780) );
  XOR2_X1 U10923 ( .A(n11045), .B(n11046), .Z(n11044) );
  XOR2_X1 U10924 ( .A(n11047), .B(n11048), .Z(n10784) );
  XOR2_X1 U10925 ( .A(n11049), .B(n11050), .Z(n11048) );
  XOR2_X1 U10926 ( .A(n11051), .B(n11052), .Z(n10788) );
  XOR2_X1 U10927 ( .A(n11053), .B(n11054), .Z(n11052) );
  XOR2_X1 U10928 ( .A(n10826), .B(n11055), .Z(n10792) );
  XOR2_X1 U10929 ( .A(n10825), .B(n10824), .Z(n11055) );
  OR2_X1 U10930 ( .A1(n8730), .A2(n8826), .ZN(n10824) );
  OR2_X1 U10931 ( .A1(n11056), .A2(n11057), .ZN(n10825) );
  AND2_X1 U10932 ( .A1(n11054), .A2(n11053), .ZN(n11057) );
  AND2_X1 U10933 ( .A1(n11051), .A2(n11058), .ZN(n11056) );
  OR2_X1 U10934 ( .A1(n11054), .A2(n11053), .ZN(n11058) );
  OR2_X1 U10935 ( .A1(n11059), .A2(n11060), .ZN(n11053) );
  AND2_X1 U10936 ( .A1(n11050), .A2(n11049), .ZN(n11060) );
  AND2_X1 U10937 ( .A1(n11047), .A2(n11061), .ZN(n11059) );
  OR2_X1 U10938 ( .A1(n11050), .A2(n11049), .ZN(n11061) );
  OR2_X1 U10939 ( .A1(n11062), .A2(n11063), .ZN(n11049) );
  AND2_X1 U10940 ( .A1(n11046), .A2(n11045), .ZN(n11063) );
  AND2_X1 U10941 ( .A1(n11043), .A2(n11064), .ZN(n11062) );
  OR2_X1 U10942 ( .A1(n11046), .A2(n11045), .ZN(n11064) );
  OR2_X1 U10943 ( .A1(n11065), .A2(n11066), .ZN(n11045) );
  AND2_X1 U10944 ( .A1(n11042), .A2(n11041), .ZN(n11066) );
  AND2_X1 U10945 ( .A1(n11039), .A2(n11067), .ZN(n11065) );
  OR2_X1 U10946 ( .A1(n11042), .A2(n11041), .ZN(n11067) );
  OR2_X1 U10947 ( .A1(n11068), .A2(n11069), .ZN(n11041) );
  AND2_X1 U10948 ( .A1(n11038), .A2(n11037), .ZN(n11069) );
  AND2_X1 U10949 ( .A1(n11036), .A2(n11070), .ZN(n11068) );
  OR2_X1 U10950 ( .A1(n11038), .A2(n11037), .ZN(n11070) );
  OR2_X1 U10951 ( .A1(n8750), .A2(n8826), .ZN(n11037) );
  OR2_X1 U10952 ( .A1(n11071), .A2(n11072), .ZN(n11038) );
  AND2_X1 U10953 ( .A1(n11034), .A2(n11033), .ZN(n11072) );
  AND2_X1 U10954 ( .A1(n11031), .A2(n11073), .ZN(n11071) );
  OR2_X1 U10955 ( .A1(n11034), .A2(n11033), .ZN(n11073) );
  OR2_X1 U10956 ( .A1(n11074), .A2(n11075), .ZN(n11033) );
  AND2_X1 U10957 ( .A1(n11030), .A2(n11029), .ZN(n11075) );
  AND2_X1 U10958 ( .A1(n11027), .A2(n11076), .ZN(n11074) );
  OR2_X1 U10959 ( .A1(n11030), .A2(n11029), .ZN(n11076) );
  OR2_X1 U10960 ( .A1(n11077), .A2(n11078), .ZN(n11029) );
  AND2_X1 U10961 ( .A1(n11026), .A2(n11025), .ZN(n11078) );
  AND2_X1 U10962 ( .A1(n11023), .A2(n11079), .ZN(n11077) );
  OR2_X1 U10963 ( .A1(n11026), .A2(n11025), .ZN(n11079) );
  OR2_X1 U10964 ( .A1(n11080), .A2(n11081), .ZN(n11025) );
  AND2_X1 U10965 ( .A1(n11022), .A2(n11021), .ZN(n11081) );
  AND2_X1 U10966 ( .A1(n11020), .A2(n11082), .ZN(n11080) );
  OR2_X1 U10967 ( .A1(n11022), .A2(n11021), .ZN(n11082) );
  OR2_X1 U10968 ( .A1(n8766), .A2(n8826), .ZN(n11021) );
  OR2_X1 U10969 ( .A1(n11083), .A2(n11084), .ZN(n11022) );
  AND2_X1 U10970 ( .A1(n11018), .A2(n11017), .ZN(n11084) );
  AND2_X1 U10971 ( .A1(n11015), .A2(n11085), .ZN(n11083) );
  OR2_X1 U10972 ( .A1(n11018), .A2(n11017), .ZN(n11085) );
  OR2_X1 U10973 ( .A1(n11086), .A2(n11087), .ZN(n11017) );
  AND2_X1 U10974 ( .A1(n11014), .A2(n11013), .ZN(n11087) );
  AND2_X1 U10975 ( .A1(n11011), .A2(n11088), .ZN(n11086) );
  OR2_X1 U10976 ( .A1(n11014), .A2(n11013), .ZN(n11088) );
  OR2_X1 U10977 ( .A1(n11089), .A2(n11090), .ZN(n11013) );
  AND2_X1 U10978 ( .A1(n11010), .A2(n11009), .ZN(n11090) );
  AND2_X1 U10979 ( .A1(n11007), .A2(n11091), .ZN(n11089) );
  OR2_X1 U10980 ( .A1(n11010), .A2(n11009), .ZN(n11091) );
  OR2_X1 U10981 ( .A1(n11092), .A2(n11093), .ZN(n11009) );
  AND2_X1 U10982 ( .A1(n11006), .A2(n11005), .ZN(n11093) );
  AND2_X1 U10983 ( .A1(n11003), .A2(n11094), .ZN(n11092) );
  OR2_X1 U10984 ( .A1(n11006), .A2(n11005), .ZN(n11094) );
  OR2_X1 U10985 ( .A1(n11095), .A2(n11096), .ZN(n11005) );
  AND2_X1 U10986 ( .A1(n11002), .A2(n11001), .ZN(n11096) );
  AND2_X1 U10987 ( .A1(n10999), .A2(n11097), .ZN(n11095) );
  OR2_X1 U10988 ( .A1(n11002), .A2(n11001), .ZN(n11097) );
  OR2_X1 U10989 ( .A1(n11098), .A2(n11099), .ZN(n11001) );
  AND2_X1 U10990 ( .A1(n10998), .A2(n10997), .ZN(n11099) );
  AND2_X1 U10991 ( .A1(n10995), .A2(n11100), .ZN(n11098) );
  OR2_X1 U10992 ( .A1(n10998), .A2(n10997), .ZN(n11100) );
  OR2_X1 U10993 ( .A1(n11101), .A2(n11102), .ZN(n10997) );
  AND2_X1 U10994 ( .A1(n10994), .A2(n10993), .ZN(n11102) );
  AND2_X1 U10995 ( .A1(n10991), .A2(n11103), .ZN(n11101) );
  OR2_X1 U10996 ( .A1(n10994), .A2(n10993), .ZN(n11103) );
  OR2_X1 U10997 ( .A1(n11104), .A2(n11105), .ZN(n10993) );
  AND2_X1 U10998 ( .A1(n10990), .A2(n10989), .ZN(n11105) );
  AND2_X1 U10999 ( .A1(n10987), .A2(n11106), .ZN(n11104) );
  OR2_X1 U11000 ( .A1(n10990), .A2(n10989), .ZN(n11106) );
  OR2_X1 U11001 ( .A1(n11107), .A2(n11108), .ZN(n10989) );
  AND2_X1 U11002 ( .A1(n10986), .A2(n10985), .ZN(n11108) );
  AND2_X1 U11003 ( .A1(n10983), .A2(n11109), .ZN(n11107) );
  OR2_X1 U11004 ( .A1(n10986), .A2(n10985), .ZN(n11109) );
  OR2_X1 U11005 ( .A1(n11110), .A2(n11111), .ZN(n10985) );
  AND2_X1 U11006 ( .A1(n10982), .A2(n10981), .ZN(n11111) );
  AND2_X1 U11007 ( .A1(n10979), .A2(n11112), .ZN(n11110) );
  OR2_X1 U11008 ( .A1(n10982), .A2(n10981), .ZN(n11112) );
  OR2_X1 U11009 ( .A1(n11113), .A2(n11114), .ZN(n10981) );
  AND2_X1 U11010 ( .A1(n10978), .A2(n10977), .ZN(n11114) );
  AND2_X1 U11011 ( .A1(n10975), .A2(n11115), .ZN(n11113) );
  OR2_X1 U11012 ( .A1(n10978), .A2(n10977), .ZN(n11115) );
  OR2_X1 U11013 ( .A1(n11116), .A2(n11117), .ZN(n10977) );
  AND2_X1 U11014 ( .A1(n10974), .A2(n10973), .ZN(n11117) );
  AND2_X1 U11015 ( .A1(n10971), .A2(n11118), .ZN(n11116) );
  OR2_X1 U11016 ( .A1(n10974), .A2(n10973), .ZN(n11118) );
  OR2_X1 U11017 ( .A1(n11119), .A2(n11120), .ZN(n10973) );
  AND2_X1 U11018 ( .A1(n10970), .A2(n10969), .ZN(n11120) );
  AND2_X1 U11019 ( .A1(n10967), .A2(n11121), .ZN(n11119) );
  OR2_X1 U11020 ( .A1(n10970), .A2(n10969), .ZN(n11121) );
  OR2_X1 U11021 ( .A1(n11122), .A2(n11123), .ZN(n10969) );
  AND2_X1 U11022 ( .A1(n10966), .A2(n10965), .ZN(n11123) );
  AND2_X1 U11023 ( .A1(n10963), .A2(n11124), .ZN(n11122) );
  OR2_X1 U11024 ( .A1(n10966), .A2(n10965), .ZN(n11124) );
  OR2_X1 U11025 ( .A1(n11125), .A2(n11126), .ZN(n10965) );
  AND2_X1 U11026 ( .A1(n8827), .A2(n10962), .ZN(n11126) );
  AND2_X1 U11027 ( .A1(n10960), .A2(n11127), .ZN(n11125) );
  OR2_X1 U11028 ( .A1(n8827), .A2(n10962), .ZN(n11127) );
  OR2_X1 U11029 ( .A1(n11128), .A2(n11129), .ZN(n10962) );
  AND2_X1 U11030 ( .A1(n10959), .A2(n10958), .ZN(n11129) );
  AND2_X1 U11031 ( .A1(n10956), .A2(n11130), .ZN(n11128) );
  OR2_X1 U11032 ( .A1(n10959), .A2(n10958), .ZN(n11130) );
  OR2_X1 U11033 ( .A1(n11131), .A2(n11132), .ZN(n10958) );
  AND2_X1 U11034 ( .A1(n10955), .A2(n10954), .ZN(n11132) );
  AND2_X1 U11035 ( .A1(n10952), .A2(n11133), .ZN(n11131) );
  OR2_X1 U11036 ( .A1(n10955), .A2(n10954), .ZN(n11133) );
  OR2_X1 U11037 ( .A1(n11134), .A2(n11135), .ZN(n10954) );
  AND2_X1 U11038 ( .A1(n10951), .A2(n10950), .ZN(n11135) );
  AND2_X1 U11039 ( .A1(n10948), .A2(n11136), .ZN(n11134) );
  OR2_X1 U11040 ( .A1(n10951), .A2(n10950), .ZN(n11136) );
  OR2_X1 U11041 ( .A1(n11137), .A2(n11138), .ZN(n10950) );
  AND2_X1 U11042 ( .A1(n10944), .A2(n10947), .ZN(n11138) );
  AND2_X1 U11043 ( .A1(n11139), .A2(n11140), .ZN(n11137) );
  OR2_X1 U11044 ( .A1(n10944), .A2(n10947), .ZN(n11140) );
  OR3_X1 U11045 ( .A1(n8826), .A2(n8822), .A3(n9796), .ZN(n10947) );
  OR2_X1 U11046 ( .A1(n7954), .A2(n8826), .ZN(n10944) );
  INV_X1 U11047 ( .A(n10946), .ZN(n11139) );
  OR2_X1 U11048 ( .A1(n11141), .A2(n11142), .ZN(n10946) );
  AND2_X1 U11049 ( .A1(b_24_), .A2(n11143), .ZN(n11142) );
  OR2_X1 U11050 ( .A1(n11144), .A2(n9801), .ZN(n11143) );
  AND2_X1 U11051 ( .A1(a_30_), .A2(n8818), .ZN(n11144) );
  AND2_X1 U11052 ( .A1(b_23_), .A2(n11145), .ZN(n11141) );
  OR2_X1 U11053 ( .A1(n11146), .A2(n7920), .ZN(n11145) );
  AND2_X1 U11054 ( .A1(a_31_), .A2(n8822), .ZN(n11146) );
  OR2_X1 U11055 ( .A1(n7979), .A2(n8826), .ZN(n10951) );
  XNOR2_X1 U11056 ( .A(n11147), .B(n11148), .ZN(n10948) );
  XOR2_X1 U11057 ( .A(n11149), .B(n11150), .Z(n11148) );
  OR2_X1 U11058 ( .A1(n8015), .A2(n8826), .ZN(n10955) );
  XOR2_X1 U11059 ( .A(n11151), .B(n11152), .Z(n10952) );
  XOR2_X1 U11060 ( .A(n11153), .B(n11154), .Z(n11152) );
  OR2_X1 U11061 ( .A1(n8040), .A2(n8826), .ZN(n10959) );
  XOR2_X1 U11062 ( .A(n11155), .B(n11156), .Z(n10956) );
  XOR2_X1 U11063 ( .A(n11157), .B(n11158), .Z(n11156) );
  OR2_X1 U11064 ( .A1(n8065), .A2(n8826), .ZN(n8827) );
  XOR2_X1 U11065 ( .A(n11159), .B(n11160), .Z(n10960) );
  XOR2_X1 U11066 ( .A(n11161), .B(n11162), .Z(n11160) );
  OR2_X1 U11067 ( .A1(n8090), .A2(n8826), .ZN(n10966) );
  XOR2_X1 U11068 ( .A(n11163), .B(n11164), .Z(n10963) );
  XOR2_X1 U11069 ( .A(n11165), .B(n11166), .Z(n11164) );
  OR2_X1 U11070 ( .A1(n8115), .A2(n8826), .ZN(n10970) );
  XOR2_X1 U11071 ( .A(n11167), .B(n11168), .Z(n10967) );
  XOR2_X1 U11072 ( .A(n11169), .B(n8823), .Z(n11168) );
  OR2_X1 U11073 ( .A1(n8140), .A2(n8826), .ZN(n10974) );
  XOR2_X1 U11074 ( .A(n11170), .B(n11171), .Z(n10971) );
  XOR2_X1 U11075 ( .A(n11172), .B(n11173), .Z(n11171) );
  OR2_X1 U11076 ( .A1(n8810), .A2(n8826), .ZN(n10978) );
  XOR2_X1 U11077 ( .A(n11174), .B(n11175), .Z(n10975) );
  XOR2_X1 U11078 ( .A(n11176), .B(n11177), .Z(n11175) );
  OR2_X1 U11079 ( .A1(n8806), .A2(n8826), .ZN(n10982) );
  XOR2_X1 U11080 ( .A(n11178), .B(n11179), .Z(n10979) );
  XOR2_X1 U11081 ( .A(n11180), .B(n11181), .Z(n11179) );
  OR2_X1 U11082 ( .A1(n8802), .A2(n8826), .ZN(n10986) );
  XOR2_X1 U11083 ( .A(n11182), .B(n11183), .Z(n10983) );
  XOR2_X1 U11084 ( .A(n11184), .B(n11185), .Z(n11183) );
  OR2_X1 U11085 ( .A1(n8798), .A2(n8826), .ZN(n10990) );
  XOR2_X1 U11086 ( .A(n11186), .B(n11187), .Z(n10987) );
  XOR2_X1 U11087 ( .A(n11188), .B(n11189), .Z(n11187) );
  OR2_X1 U11088 ( .A1(n8794), .A2(n8826), .ZN(n10994) );
  XOR2_X1 U11089 ( .A(n11190), .B(n11191), .Z(n10991) );
  XOR2_X1 U11090 ( .A(n11192), .B(n11193), .Z(n11191) );
  OR2_X1 U11091 ( .A1(n8790), .A2(n8826), .ZN(n10998) );
  XOR2_X1 U11092 ( .A(n11194), .B(n11195), .Z(n10995) );
  XOR2_X1 U11093 ( .A(n11196), .B(n11197), .Z(n11195) );
  OR2_X1 U11094 ( .A1(n8786), .A2(n8826), .ZN(n11002) );
  XOR2_X1 U11095 ( .A(n11198), .B(n11199), .Z(n10999) );
  XOR2_X1 U11096 ( .A(n11200), .B(n11201), .Z(n11199) );
  OR2_X1 U11097 ( .A1(n8782), .A2(n8826), .ZN(n11006) );
  XOR2_X1 U11098 ( .A(n11202), .B(n11203), .Z(n11003) );
  XOR2_X1 U11099 ( .A(n11204), .B(n11205), .Z(n11203) );
  OR2_X1 U11100 ( .A1(n8778), .A2(n8826), .ZN(n11010) );
  XOR2_X1 U11101 ( .A(n11206), .B(n11207), .Z(n11007) );
  XOR2_X1 U11102 ( .A(n11208), .B(n11209), .Z(n11207) );
  OR2_X1 U11103 ( .A1(n8774), .A2(n8826), .ZN(n11014) );
  XOR2_X1 U11104 ( .A(n11210), .B(n11211), .Z(n11011) );
  XOR2_X1 U11105 ( .A(n11212), .B(n11213), .Z(n11211) );
  OR2_X1 U11106 ( .A1(n8770), .A2(n8826), .ZN(n11018) );
  XOR2_X1 U11107 ( .A(n11214), .B(n11215), .Z(n11015) );
  XOR2_X1 U11108 ( .A(n11216), .B(n11217), .Z(n11215) );
  XOR2_X1 U11109 ( .A(n11218), .B(n11219), .Z(n11020) );
  XOR2_X1 U11110 ( .A(n11220), .B(n11221), .Z(n11219) );
  OR2_X1 U11111 ( .A1(n8762), .A2(n8826), .ZN(n11026) );
  XNOR2_X1 U11112 ( .A(n11222), .B(n11223), .ZN(n11023) );
  XNOR2_X1 U11113 ( .A(n11224), .B(n11225), .ZN(n11222) );
  OR2_X1 U11114 ( .A1(n8758), .A2(n8826), .ZN(n11030) );
  XOR2_X1 U11115 ( .A(n11226), .B(n11227), .Z(n11027) );
  XOR2_X1 U11116 ( .A(n11228), .B(n11229), .Z(n11227) );
  OR2_X1 U11117 ( .A1(n8754), .A2(n8826), .ZN(n11034) );
  XOR2_X1 U11118 ( .A(n11230), .B(n11231), .Z(n11031) );
  XOR2_X1 U11119 ( .A(n11232), .B(n11233), .Z(n11231) );
  XOR2_X1 U11120 ( .A(n11234), .B(n11235), .Z(n11036) );
  XOR2_X1 U11121 ( .A(n11236), .B(n11237), .Z(n11235) );
  OR2_X1 U11122 ( .A1(n8746), .A2(n8826), .ZN(n11042) );
  XNOR2_X1 U11123 ( .A(n11238), .B(n11239), .ZN(n11039) );
  XNOR2_X1 U11124 ( .A(n11240), .B(n11241), .ZN(n11238) );
  OR2_X1 U11125 ( .A1(n8742), .A2(n8826), .ZN(n11046) );
  XOR2_X1 U11126 ( .A(n11242), .B(n11243), .Z(n11043) );
  XOR2_X1 U11127 ( .A(n11244), .B(n11245), .Z(n11243) );
  OR2_X1 U11128 ( .A1(n8738), .A2(n8826), .ZN(n11050) );
  XOR2_X1 U11129 ( .A(n11246), .B(n11247), .Z(n11047) );
  XOR2_X1 U11130 ( .A(n11248), .B(n11249), .Z(n11247) );
  OR2_X1 U11131 ( .A1(n8734), .A2(n8826), .ZN(n11054) );
  XNOR2_X1 U11132 ( .A(n11250), .B(n11251), .ZN(n11051) );
  XNOR2_X1 U11133 ( .A(n11252), .B(n11253), .ZN(n11250) );
  XOR2_X1 U11134 ( .A(n10844), .B(n11254), .Z(n10826) );
  XOR2_X1 U11135 ( .A(n10843), .B(n10842), .Z(n11254) );
  OR2_X1 U11136 ( .A1(n8734), .A2(n8822), .ZN(n10842) );
  OR2_X1 U11137 ( .A1(n11255), .A2(n11256), .ZN(n10843) );
  AND2_X1 U11138 ( .A1(n11253), .A2(n11252), .ZN(n11256) );
  AND2_X1 U11139 ( .A1(n11251), .A2(n11257), .ZN(n11255) );
  OR2_X1 U11140 ( .A1(n11253), .A2(n11252), .ZN(n11257) );
  OR2_X1 U11141 ( .A1(n8738), .A2(n8822), .ZN(n11252) );
  OR2_X1 U11142 ( .A1(n11258), .A2(n11259), .ZN(n11253) );
  AND2_X1 U11143 ( .A1(n11249), .A2(n11248), .ZN(n11259) );
  AND2_X1 U11144 ( .A1(n11246), .A2(n11260), .ZN(n11258) );
  OR2_X1 U11145 ( .A1(n11249), .A2(n11248), .ZN(n11260) );
  OR2_X1 U11146 ( .A1(n11261), .A2(n11262), .ZN(n11248) );
  AND2_X1 U11147 ( .A1(n11245), .A2(n11244), .ZN(n11262) );
  AND2_X1 U11148 ( .A1(n11242), .A2(n11263), .ZN(n11261) );
  OR2_X1 U11149 ( .A1(n11245), .A2(n11244), .ZN(n11263) );
  OR2_X1 U11150 ( .A1(n11264), .A2(n11265), .ZN(n11244) );
  AND2_X1 U11151 ( .A1(n11241), .A2(n11240), .ZN(n11265) );
  AND2_X1 U11152 ( .A1(n11239), .A2(n11266), .ZN(n11264) );
  OR2_X1 U11153 ( .A1(n11241), .A2(n11240), .ZN(n11266) );
  OR2_X1 U11154 ( .A1(n8750), .A2(n8822), .ZN(n11240) );
  OR2_X1 U11155 ( .A1(n11267), .A2(n11268), .ZN(n11241) );
  AND2_X1 U11156 ( .A1(n11237), .A2(n11236), .ZN(n11268) );
  AND2_X1 U11157 ( .A1(n11234), .A2(n11269), .ZN(n11267) );
  OR2_X1 U11158 ( .A1(n11237), .A2(n11236), .ZN(n11269) );
  OR2_X1 U11159 ( .A1(n11270), .A2(n11271), .ZN(n11236) );
  AND2_X1 U11160 ( .A1(n11233), .A2(n11232), .ZN(n11271) );
  AND2_X1 U11161 ( .A1(n11230), .A2(n11272), .ZN(n11270) );
  OR2_X1 U11162 ( .A1(n11233), .A2(n11232), .ZN(n11272) );
  OR2_X1 U11163 ( .A1(n11273), .A2(n11274), .ZN(n11232) );
  AND2_X1 U11164 ( .A1(n11229), .A2(n11228), .ZN(n11274) );
  AND2_X1 U11165 ( .A1(n11226), .A2(n11275), .ZN(n11273) );
  OR2_X1 U11166 ( .A1(n11229), .A2(n11228), .ZN(n11275) );
  OR2_X1 U11167 ( .A1(n11276), .A2(n11277), .ZN(n11228) );
  AND2_X1 U11168 ( .A1(n11225), .A2(n11224), .ZN(n11277) );
  AND2_X1 U11169 ( .A1(n11223), .A2(n11278), .ZN(n11276) );
  OR2_X1 U11170 ( .A1(n11225), .A2(n11224), .ZN(n11278) );
  OR2_X1 U11171 ( .A1(n8766), .A2(n8822), .ZN(n11224) );
  OR2_X1 U11172 ( .A1(n11279), .A2(n11280), .ZN(n11225) );
  AND2_X1 U11173 ( .A1(n11221), .A2(n11220), .ZN(n11280) );
  AND2_X1 U11174 ( .A1(n11218), .A2(n11281), .ZN(n11279) );
  OR2_X1 U11175 ( .A1(n11221), .A2(n11220), .ZN(n11281) );
  OR2_X1 U11176 ( .A1(n11282), .A2(n11283), .ZN(n11220) );
  AND2_X1 U11177 ( .A1(n11217), .A2(n11216), .ZN(n11283) );
  AND2_X1 U11178 ( .A1(n11214), .A2(n11284), .ZN(n11282) );
  OR2_X1 U11179 ( .A1(n11217), .A2(n11216), .ZN(n11284) );
  OR2_X1 U11180 ( .A1(n11285), .A2(n11286), .ZN(n11216) );
  AND2_X1 U11181 ( .A1(n11213), .A2(n11212), .ZN(n11286) );
  AND2_X1 U11182 ( .A1(n11210), .A2(n11287), .ZN(n11285) );
  OR2_X1 U11183 ( .A1(n11213), .A2(n11212), .ZN(n11287) );
  OR2_X1 U11184 ( .A1(n11288), .A2(n11289), .ZN(n11212) );
  AND2_X1 U11185 ( .A1(n11209), .A2(n11208), .ZN(n11289) );
  AND2_X1 U11186 ( .A1(n11206), .A2(n11290), .ZN(n11288) );
  OR2_X1 U11187 ( .A1(n11209), .A2(n11208), .ZN(n11290) );
  OR2_X1 U11188 ( .A1(n11291), .A2(n11292), .ZN(n11208) );
  AND2_X1 U11189 ( .A1(n11205), .A2(n11204), .ZN(n11292) );
  AND2_X1 U11190 ( .A1(n11202), .A2(n11293), .ZN(n11291) );
  OR2_X1 U11191 ( .A1(n11205), .A2(n11204), .ZN(n11293) );
  OR2_X1 U11192 ( .A1(n11294), .A2(n11295), .ZN(n11204) );
  AND2_X1 U11193 ( .A1(n11201), .A2(n11200), .ZN(n11295) );
  AND2_X1 U11194 ( .A1(n11198), .A2(n11296), .ZN(n11294) );
  OR2_X1 U11195 ( .A1(n11201), .A2(n11200), .ZN(n11296) );
  OR2_X1 U11196 ( .A1(n11297), .A2(n11298), .ZN(n11200) );
  AND2_X1 U11197 ( .A1(n11197), .A2(n11196), .ZN(n11298) );
  AND2_X1 U11198 ( .A1(n11194), .A2(n11299), .ZN(n11297) );
  OR2_X1 U11199 ( .A1(n11197), .A2(n11196), .ZN(n11299) );
  OR2_X1 U11200 ( .A1(n11300), .A2(n11301), .ZN(n11196) );
  AND2_X1 U11201 ( .A1(n11193), .A2(n11192), .ZN(n11301) );
  AND2_X1 U11202 ( .A1(n11190), .A2(n11302), .ZN(n11300) );
  OR2_X1 U11203 ( .A1(n11193), .A2(n11192), .ZN(n11302) );
  OR2_X1 U11204 ( .A1(n11303), .A2(n11304), .ZN(n11192) );
  AND2_X1 U11205 ( .A1(n11189), .A2(n11188), .ZN(n11304) );
  AND2_X1 U11206 ( .A1(n11186), .A2(n11305), .ZN(n11303) );
  OR2_X1 U11207 ( .A1(n11189), .A2(n11188), .ZN(n11305) );
  OR2_X1 U11208 ( .A1(n11306), .A2(n11307), .ZN(n11188) );
  AND2_X1 U11209 ( .A1(n11185), .A2(n11184), .ZN(n11307) );
  AND2_X1 U11210 ( .A1(n11182), .A2(n11308), .ZN(n11306) );
  OR2_X1 U11211 ( .A1(n11185), .A2(n11184), .ZN(n11308) );
  OR2_X1 U11212 ( .A1(n11309), .A2(n11310), .ZN(n11184) );
  AND2_X1 U11213 ( .A1(n11181), .A2(n11180), .ZN(n11310) );
  AND2_X1 U11214 ( .A1(n11178), .A2(n11311), .ZN(n11309) );
  OR2_X1 U11215 ( .A1(n11181), .A2(n11180), .ZN(n11311) );
  OR2_X1 U11216 ( .A1(n11312), .A2(n11313), .ZN(n11180) );
  AND2_X1 U11217 ( .A1(n11177), .A2(n11176), .ZN(n11313) );
  AND2_X1 U11218 ( .A1(n11174), .A2(n11314), .ZN(n11312) );
  OR2_X1 U11219 ( .A1(n11177), .A2(n11176), .ZN(n11314) );
  OR2_X1 U11220 ( .A1(n11315), .A2(n11316), .ZN(n11176) );
  AND2_X1 U11221 ( .A1(n11173), .A2(n11172), .ZN(n11316) );
  AND2_X1 U11222 ( .A1(n11170), .A2(n11317), .ZN(n11315) );
  OR2_X1 U11223 ( .A1(n11173), .A2(n11172), .ZN(n11317) );
  OR2_X1 U11224 ( .A1(n11318), .A2(n11319), .ZN(n11172) );
  AND2_X1 U11225 ( .A1(n8823), .A2(n11169), .ZN(n11319) );
  AND2_X1 U11226 ( .A1(n11167), .A2(n11320), .ZN(n11318) );
  OR2_X1 U11227 ( .A1(n8823), .A2(n11169), .ZN(n11320) );
  OR2_X1 U11228 ( .A1(n11321), .A2(n11322), .ZN(n11169) );
  AND2_X1 U11229 ( .A1(n11166), .A2(n11165), .ZN(n11322) );
  AND2_X1 U11230 ( .A1(n11163), .A2(n11323), .ZN(n11321) );
  OR2_X1 U11231 ( .A1(n11166), .A2(n11165), .ZN(n11323) );
  OR2_X1 U11232 ( .A1(n11324), .A2(n11325), .ZN(n11165) );
  AND2_X1 U11233 ( .A1(n11162), .A2(n11161), .ZN(n11325) );
  AND2_X1 U11234 ( .A1(n11159), .A2(n11326), .ZN(n11324) );
  OR2_X1 U11235 ( .A1(n11162), .A2(n11161), .ZN(n11326) );
  OR2_X1 U11236 ( .A1(n11327), .A2(n11328), .ZN(n11161) );
  AND2_X1 U11237 ( .A1(n11158), .A2(n11157), .ZN(n11328) );
  AND2_X1 U11238 ( .A1(n11155), .A2(n11329), .ZN(n11327) );
  OR2_X1 U11239 ( .A1(n11158), .A2(n11157), .ZN(n11329) );
  OR2_X1 U11240 ( .A1(n11330), .A2(n11331), .ZN(n11157) );
  AND2_X1 U11241 ( .A1(n11154), .A2(n11153), .ZN(n11331) );
  AND2_X1 U11242 ( .A1(n11151), .A2(n11332), .ZN(n11330) );
  OR2_X1 U11243 ( .A1(n11154), .A2(n11153), .ZN(n11332) );
  OR2_X1 U11244 ( .A1(n11333), .A2(n11334), .ZN(n11153) );
  AND2_X1 U11245 ( .A1(n11147), .A2(n11150), .ZN(n11334) );
  AND2_X1 U11246 ( .A1(n11335), .A2(n11336), .ZN(n11333) );
  OR2_X1 U11247 ( .A1(n11147), .A2(n11150), .ZN(n11336) );
  OR3_X1 U11248 ( .A1(n8822), .A2(n8818), .A3(n9796), .ZN(n11150) );
  OR2_X1 U11249 ( .A1(n7954), .A2(n8822), .ZN(n11147) );
  INV_X1 U11250 ( .A(n11149), .ZN(n11335) );
  OR2_X1 U11251 ( .A1(n11337), .A2(n11338), .ZN(n11149) );
  AND2_X1 U11252 ( .A1(b_23_), .A2(n11339), .ZN(n11338) );
  OR2_X1 U11253 ( .A1(n11340), .A2(n9801), .ZN(n11339) );
  AND2_X1 U11254 ( .A1(a_30_), .A2(n8814), .ZN(n11340) );
  AND2_X1 U11255 ( .A1(b_22_), .A2(n11341), .ZN(n11337) );
  OR2_X1 U11256 ( .A1(n11342), .A2(n7920), .ZN(n11341) );
  AND2_X1 U11257 ( .A1(a_31_), .A2(n8818), .ZN(n11342) );
  OR2_X1 U11258 ( .A1(n7979), .A2(n8822), .ZN(n11154) );
  XNOR2_X1 U11259 ( .A(n11343), .B(n11344), .ZN(n11151) );
  XOR2_X1 U11260 ( .A(n11345), .B(n11346), .Z(n11344) );
  OR2_X1 U11261 ( .A1(n8015), .A2(n8822), .ZN(n11158) );
  XOR2_X1 U11262 ( .A(n11347), .B(n11348), .Z(n11155) );
  XOR2_X1 U11263 ( .A(n11349), .B(n11350), .Z(n11348) );
  OR2_X1 U11264 ( .A1(n8040), .A2(n8822), .ZN(n11162) );
  XOR2_X1 U11265 ( .A(n11351), .B(n11352), .Z(n11159) );
  XOR2_X1 U11266 ( .A(n11353), .B(n11354), .Z(n11352) );
  OR2_X1 U11267 ( .A1(n8065), .A2(n8822), .ZN(n11166) );
  XOR2_X1 U11268 ( .A(n11355), .B(n11356), .Z(n11163) );
  XOR2_X1 U11269 ( .A(n11357), .B(n11358), .Z(n11356) );
  OR2_X1 U11270 ( .A1(n8090), .A2(n8822), .ZN(n8823) );
  XOR2_X1 U11271 ( .A(n11359), .B(n11360), .Z(n11167) );
  XOR2_X1 U11272 ( .A(n11361), .B(n11362), .Z(n11360) );
  OR2_X1 U11273 ( .A1(n8115), .A2(n8822), .ZN(n11173) );
  XOR2_X1 U11274 ( .A(n11363), .B(n11364), .Z(n11170) );
  XOR2_X1 U11275 ( .A(n11365), .B(n11366), .Z(n11364) );
  OR2_X1 U11276 ( .A1(n8140), .A2(n8822), .ZN(n11177) );
  XOR2_X1 U11277 ( .A(n11367), .B(n11368), .Z(n11174) );
  XOR2_X1 U11278 ( .A(n11369), .B(n8819), .Z(n11368) );
  OR2_X1 U11279 ( .A1(n8810), .A2(n8822), .ZN(n11181) );
  XOR2_X1 U11280 ( .A(n11370), .B(n11371), .Z(n11178) );
  XOR2_X1 U11281 ( .A(n11372), .B(n11373), .Z(n11371) );
  OR2_X1 U11282 ( .A1(n8806), .A2(n8822), .ZN(n11185) );
  XOR2_X1 U11283 ( .A(n11374), .B(n11375), .Z(n11182) );
  XOR2_X1 U11284 ( .A(n11376), .B(n11377), .Z(n11375) );
  OR2_X1 U11285 ( .A1(n8802), .A2(n8822), .ZN(n11189) );
  XOR2_X1 U11286 ( .A(n11378), .B(n11379), .Z(n11186) );
  XOR2_X1 U11287 ( .A(n11380), .B(n11381), .Z(n11379) );
  OR2_X1 U11288 ( .A1(n8798), .A2(n8822), .ZN(n11193) );
  XOR2_X1 U11289 ( .A(n11382), .B(n11383), .Z(n11190) );
  XOR2_X1 U11290 ( .A(n11384), .B(n11385), .Z(n11383) );
  OR2_X1 U11291 ( .A1(n8794), .A2(n8822), .ZN(n11197) );
  XOR2_X1 U11292 ( .A(n11386), .B(n11387), .Z(n11194) );
  XOR2_X1 U11293 ( .A(n11388), .B(n11389), .Z(n11387) );
  OR2_X1 U11294 ( .A1(n8790), .A2(n8822), .ZN(n11201) );
  XOR2_X1 U11295 ( .A(n11390), .B(n11391), .Z(n11198) );
  XOR2_X1 U11296 ( .A(n11392), .B(n11393), .Z(n11391) );
  OR2_X1 U11297 ( .A1(n8786), .A2(n8822), .ZN(n11205) );
  XOR2_X1 U11298 ( .A(n11394), .B(n11395), .Z(n11202) );
  XOR2_X1 U11299 ( .A(n11396), .B(n11397), .Z(n11395) );
  OR2_X1 U11300 ( .A1(n8782), .A2(n8822), .ZN(n11209) );
  XOR2_X1 U11301 ( .A(n11398), .B(n11399), .Z(n11206) );
  XOR2_X1 U11302 ( .A(n11400), .B(n11401), .Z(n11399) );
  OR2_X1 U11303 ( .A1(n8778), .A2(n8822), .ZN(n11213) );
  XNOR2_X1 U11304 ( .A(n11402), .B(n11403), .ZN(n11210) );
  XNOR2_X1 U11305 ( .A(n11404), .B(n11405), .ZN(n11402) );
  OR2_X1 U11306 ( .A1(n8774), .A2(n8822), .ZN(n11217) );
  XOR2_X1 U11307 ( .A(n11406), .B(n11407), .Z(n11214) );
  XOR2_X1 U11308 ( .A(n11408), .B(n11409), .Z(n11407) );
  OR2_X1 U11309 ( .A1(n8770), .A2(n8822), .ZN(n11221) );
  XOR2_X1 U11310 ( .A(n11410), .B(n11411), .Z(n11218) );
  XOR2_X1 U11311 ( .A(n11412), .B(n11413), .Z(n11411) );
  XOR2_X1 U11312 ( .A(n11414), .B(n11415), .Z(n11223) );
  XOR2_X1 U11313 ( .A(n11416), .B(n11417), .Z(n11415) );
  OR2_X1 U11314 ( .A1(n8762), .A2(n8822), .ZN(n11229) );
  XNOR2_X1 U11315 ( .A(n11418), .B(n11419), .ZN(n11226) );
  XNOR2_X1 U11316 ( .A(n11420), .B(n11421), .ZN(n11418) );
  OR2_X1 U11317 ( .A1(n8758), .A2(n8822), .ZN(n11233) );
  XOR2_X1 U11318 ( .A(n11422), .B(n11423), .Z(n11230) );
  XOR2_X1 U11319 ( .A(n11424), .B(n11425), .Z(n11423) );
  OR2_X1 U11320 ( .A1(n8754), .A2(n8822), .ZN(n11237) );
  XOR2_X1 U11321 ( .A(n11426), .B(n11427), .Z(n11234) );
  XOR2_X1 U11322 ( .A(n11428), .B(n11429), .Z(n11427) );
  XOR2_X1 U11323 ( .A(n11430), .B(n11431), .Z(n11239) );
  XOR2_X1 U11324 ( .A(n11432), .B(n11433), .Z(n11431) );
  OR2_X1 U11325 ( .A1(n8746), .A2(n8822), .ZN(n11245) );
  XNOR2_X1 U11326 ( .A(n11434), .B(n11435), .ZN(n11242) );
  XNOR2_X1 U11327 ( .A(n11436), .B(n11437), .ZN(n11434) );
  OR2_X1 U11328 ( .A1(n8742), .A2(n8822), .ZN(n11249) );
  XOR2_X1 U11329 ( .A(n11438), .B(n11439), .Z(n11246) );
  XOR2_X1 U11330 ( .A(n11440), .B(n11441), .Z(n11439) );
  XOR2_X1 U11331 ( .A(n11442), .B(n11443), .Z(n11251) );
  XOR2_X1 U11332 ( .A(n11444), .B(n11445), .Z(n11443) );
  XOR2_X1 U11333 ( .A(n10834), .B(n11446), .Z(n10844) );
  XOR2_X1 U11334 ( .A(n10833), .B(n10832), .Z(n11446) );
  OR2_X1 U11335 ( .A1(n8738), .A2(n8818), .ZN(n10832) );
  OR2_X1 U11336 ( .A1(n11447), .A2(n11448), .ZN(n10833) );
  AND2_X1 U11337 ( .A1(n11445), .A2(n11444), .ZN(n11448) );
  AND2_X1 U11338 ( .A1(n11442), .A2(n11449), .ZN(n11447) );
  OR2_X1 U11339 ( .A1(n11445), .A2(n11444), .ZN(n11449) );
  OR2_X1 U11340 ( .A1(n11450), .A2(n11451), .ZN(n11444) );
  AND2_X1 U11341 ( .A1(n11441), .A2(n11440), .ZN(n11451) );
  AND2_X1 U11342 ( .A1(n11438), .A2(n11452), .ZN(n11450) );
  OR2_X1 U11343 ( .A1(n11441), .A2(n11440), .ZN(n11452) );
  OR2_X1 U11344 ( .A1(n11453), .A2(n11454), .ZN(n11440) );
  AND2_X1 U11345 ( .A1(n11437), .A2(n11436), .ZN(n11454) );
  AND2_X1 U11346 ( .A1(n11435), .A2(n11455), .ZN(n11453) );
  OR2_X1 U11347 ( .A1(n11437), .A2(n11436), .ZN(n11455) );
  OR2_X1 U11348 ( .A1(n8750), .A2(n8818), .ZN(n11436) );
  OR2_X1 U11349 ( .A1(n11456), .A2(n11457), .ZN(n11437) );
  AND2_X1 U11350 ( .A1(n11433), .A2(n11432), .ZN(n11457) );
  AND2_X1 U11351 ( .A1(n11430), .A2(n11458), .ZN(n11456) );
  OR2_X1 U11352 ( .A1(n11433), .A2(n11432), .ZN(n11458) );
  OR2_X1 U11353 ( .A1(n11459), .A2(n11460), .ZN(n11432) );
  AND2_X1 U11354 ( .A1(n11429), .A2(n11428), .ZN(n11460) );
  AND2_X1 U11355 ( .A1(n11426), .A2(n11461), .ZN(n11459) );
  OR2_X1 U11356 ( .A1(n11429), .A2(n11428), .ZN(n11461) );
  OR2_X1 U11357 ( .A1(n11462), .A2(n11463), .ZN(n11428) );
  AND2_X1 U11358 ( .A1(n11425), .A2(n11424), .ZN(n11463) );
  AND2_X1 U11359 ( .A1(n11422), .A2(n11464), .ZN(n11462) );
  OR2_X1 U11360 ( .A1(n11425), .A2(n11424), .ZN(n11464) );
  OR2_X1 U11361 ( .A1(n11465), .A2(n11466), .ZN(n11424) );
  AND2_X1 U11362 ( .A1(n11421), .A2(n11420), .ZN(n11466) );
  AND2_X1 U11363 ( .A1(n11419), .A2(n11467), .ZN(n11465) );
  OR2_X1 U11364 ( .A1(n11421), .A2(n11420), .ZN(n11467) );
  OR2_X1 U11365 ( .A1(n8766), .A2(n8818), .ZN(n11420) );
  OR2_X1 U11366 ( .A1(n11468), .A2(n11469), .ZN(n11421) );
  AND2_X1 U11367 ( .A1(n11417), .A2(n11416), .ZN(n11469) );
  AND2_X1 U11368 ( .A1(n11414), .A2(n11470), .ZN(n11468) );
  OR2_X1 U11369 ( .A1(n11417), .A2(n11416), .ZN(n11470) );
  OR2_X1 U11370 ( .A1(n11471), .A2(n11472), .ZN(n11416) );
  AND2_X1 U11371 ( .A1(n11413), .A2(n11412), .ZN(n11472) );
  AND2_X1 U11372 ( .A1(n11410), .A2(n11473), .ZN(n11471) );
  OR2_X1 U11373 ( .A1(n11413), .A2(n11412), .ZN(n11473) );
  OR2_X1 U11374 ( .A1(n11474), .A2(n11475), .ZN(n11412) );
  AND2_X1 U11375 ( .A1(n11409), .A2(n11408), .ZN(n11475) );
  AND2_X1 U11376 ( .A1(n11406), .A2(n11476), .ZN(n11474) );
  OR2_X1 U11377 ( .A1(n11409), .A2(n11408), .ZN(n11476) );
  OR2_X1 U11378 ( .A1(n11477), .A2(n11478), .ZN(n11408) );
  AND2_X1 U11379 ( .A1(n11405), .A2(n11404), .ZN(n11478) );
  AND2_X1 U11380 ( .A1(n11403), .A2(n11479), .ZN(n11477) );
  OR2_X1 U11381 ( .A1(n11405), .A2(n11404), .ZN(n11479) );
  OR2_X1 U11382 ( .A1(n8782), .A2(n8818), .ZN(n11404) );
  OR2_X1 U11383 ( .A1(n11480), .A2(n11481), .ZN(n11405) );
  AND2_X1 U11384 ( .A1(n11401), .A2(n11400), .ZN(n11481) );
  AND2_X1 U11385 ( .A1(n11398), .A2(n11482), .ZN(n11480) );
  OR2_X1 U11386 ( .A1(n11401), .A2(n11400), .ZN(n11482) );
  OR2_X1 U11387 ( .A1(n11483), .A2(n11484), .ZN(n11400) );
  AND2_X1 U11388 ( .A1(n11397), .A2(n11396), .ZN(n11484) );
  AND2_X1 U11389 ( .A1(n11394), .A2(n11485), .ZN(n11483) );
  OR2_X1 U11390 ( .A1(n11397), .A2(n11396), .ZN(n11485) );
  OR2_X1 U11391 ( .A1(n11486), .A2(n11487), .ZN(n11396) );
  AND2_X1 U11392 ( .A1(n11393), .A2(n11392), .ZN(n11487) );
  AND2_X1 U11393 ( .A1(n11390), .A2(n11488), .ZN(n11486) );
  OR2_X1 U11394 ( .A1(n11393), .A2(n11392), .ZN(n11488) );
  OR2_X1 U11395 ( .A1(n11489), .A2(n11490), .ZN(n11392) );
  AND2_X1 U11396 ( .A1(n11389), .A2(n11388), .ZN(n11490) );
  AND2_X1 U11397 ( .A1(n11386), .A2(n11491), .ZN(n11489) );
  OR2_X1 U11398 ( .A1(n11389), .A2(n11388), .ZN(n11491) );
  OR2_X1 U11399 ( .A1(n11492), .A2(n11493), .ZN(n11388) );
  AND2_X1 U11400 ( .A1(n11385), .A2(n11384), .ZN(n11493) );
  AND2_X1 U11401 ( .A1(n11382), .A2(n11494), .ZN(n11492) );
  OR2_X1 U11402 ( .A1(n11385), .A2(n11384), .ZN(n11494) );
  OR2_X1 U11403 ( .A1(n11495), .A2(n11496), .ZN(n11384) );
  AND2_X1 U11404 ( .A1(n11381), .A2(n11380), .ZN(n11496) );
  AND2_X1 U11405 ( .A1(n11378), .A2(n11497), .ZN(n11495) );
  OR2_X1 U11406 ( .A1(n11381), .A2(n11380), .ZN(n11497) );
  OR2_X1 U11407 ( .A1(n11498), .A2(n11499), .ZN(n11380) );
  AND2_X1 U11408 ( .A1(n11377), .A2(n11376), .ZN(n11499) );
  AND2_X1 U11409 ( .A1(n11374), .A2(n11500), .ZN(n11498) );
  OR2_X1 U11410 ( .A1(n11377), .A2(n11376), .ZN(n11500) );
  OR2_X1 U11411 ( .A1(n11501), .A2(n11502), .ZN(n11376) );
  AND2_X1 U11412 ( .A1(n11373), .A2(n11372), .ZN(n11502) );
  AND2_X1 U11413 ( .A1(n11370), .A2(n11503), .ZN(n11501) );
  OR2_X1 U11414 ( .A1(n11373), .A2(n11372), .ZN(n11503) );
  OR2_X1 U11415 ( .A1(n11504), .A2(n11505), .ZN(n11372) );
  AND2_X1 U11416 ( .A1(n8819), .A2(n11369), .ZN(n11505) );
  AND2_X1 U11417 ( .A1(n11367), .A2(n11506), .ZN(n11504) );
  OR2_X1 U11418 ( .A1(n8819), .A2(n11369), .ZN(n11506) );
  OR2_X1 U11419 ( .A1(n11507), .A2(n11508), .ZN(n11369) );
  AND2_X1 U11420 ( .A1(n11366), .A2(n11365), .ZN(n11508) );
  AND2_X1 U11421 ( .A1(n11363), .A2(n11509), .ZN(n11507) );
  OR2_X1 U11422 ( .A1(n11366), .A2(n11365), .ZN(n11509) );
  OR2_X1 U11423 ( .A1(n11510), .A2(n11511), .ZN(n11365) );
  AND2_X1 U11424 ( .A1(n11362), .A2(n11361), .ZN(n11511) );
  AND2_X1 U11425 ( .A1(n11359), .A2(n11512), .ZN(n11510) );
  OR2_X1 U11426 ( .A1(n11362), .A2(n11361), .ZN(n11512) );
  OR2_X1 U11427 ( .A1(n11513), .A2(n11514), .ZN(n11361) );
  AND2_X1 U11428 ( .A1(n11358), .A2(n11357), .ZN(n11514) );
  AND2_X1 U11429 ( .A1(n11355), .A2(n11515), .ZN(n11513) );
  OR2_X1 U11430 ( .A1(n11358), .A2(n11357), .ZN(n11515) );
  OR2_X1 U11431 ( .A1(n11516), .A2(n11517), .ZN(n11357) );
  AND2_X1 U11432 ( .A1(n11354), .A2(n11353), .ZN(n11517) );
  AND2_X1 U11433 ( .A1(n11351), .A2(n11518), .ZN(n11516) );
  OR2_X1 U11434 ( .A1(n11354), .A2(n11353), .ZN(n11518) );
  OR2_X1 U11435 ( .A1(n11519), .A2(n11520), .ZN(n11353) );
  AND2_X1 U11436 ( .A1(n11350), .A2(n11349), .ZN(n11520) );
  AND2_X1 U11437 ( .A1(n11347), .A2(n11521), .ZN(n11519) );
  OR2_X1 U11438 ( .A1(n11350), .A2(n11349), .ZN(n11521) );
  OR2_X1 U11439 ( .A1(n11522), .A2(n11523), .ZN(n11349) );
  AND2_X1 U11440 ( .A1(n11343), .A2(n11346), .ZN(n11523) );
  AND2_X1 U11441 ( .A1(n11524), .A2(n11525), .ZN(n11522) );
  OR2_X1 U11442 ( .A1(n11343), .A2(n11346), .ZN(n11525) );
  OR3_X1 U11443 ( .A1(n8818), .A2(n8814), .A3(n9796), .ZN(n11346) );
  OR2_X1 U11444 ( .A1(n7954), .A2(n8818), .ZN(n11343) );
  INV_X1 U11445 ( .A(n11345), .ZN(n11524) );
  OR2_X1 U11446 ( .A1(n11526), .A2(n11527), .ZN(n11345) );
  AND2_X1 U11447 ( .A1(b_22_), .A2(n11528), .ZN(n11527) );
  OR2_X1 U11448 ( .A1(n11529), .A2(n9801), .ZN(n11528) );
  AND2_X1 U11449 ( .A1(a_30_), .A2(n8811), .ZN(n11529) );
  AND2_X1 U11450 ( .A1(b_21_), .A2(n11530), .ZN(n11526) );
  OR2_X1 U11451 ( .A1(n11531), .A2(n7920), .ZN(n11530) );
  AND2_X1 U11452 ( .A1(a_31_), .A2(n8814), .ZN(n11531) );
  OR2_X1 U11453 ( .A1(n7979), .A2(n8818), .ZN(n11350) );
  XNOR2_X1 U11454 ( .A(n11532), .B(n11533), .ZN(n11347) );
  XOR2_X1 U11455 ( .A(n11534), .B(n11535), .Z(n11533) );
  OR2_X1 U11456 ( .A1(n8015), .A2(n8818), .ZN(n11354) );
  XOR2_X1 U11457 ( .A(n11536), .B(n11537), .Z(n11351) );
  XOR2_X1 U11458 ( .A(n11538), .B(n11539), .Z(n11537) );
  OR2_X1 U11459 ( .A1(n8040), .A2(n8818), .ZN(n11358) );
  XOR2_X1 U11460 ( .A(n11540), .B(n11541), .Z(n11355) );
  XOR2_X1 U11461 ( .A(n11542), .B(n11543), .Z(n11541) );
  OR2_X1 U11462 ( .A1(n8065), .A2(n8818), .ZN(n11362) );
  XOR2_X1 U11463 ( .A(n11544), .B(n11545), .Z(n11359) );
  XOR2_X1 U11464 ( .A(n11546), .B(n11547), .Z(n11545) );
  OR2_X1 U11465 ( .A1(n8090), .A2(n8818), .ZN(n11366) );
  XOR2_X1 U11466 ( .A(n11548), .B(n11549), .Z(n11363) );
  XOR2_X1 U11467 ( .A(n11550), .B(n11551), .Z(n11549) );
  OR2_X1 U11468 ( .A1(n8115), .A2(n8818), .ZN(n8819) );
  XOR2_X1 U11469 ( .A(n11552), .B(n11553), .Z(n11367) );
  XOR2_X1 U11470 ( .A(n11554), .B(n11555), .Z(n11553) );
  OR2_X1 U11471 ( .A1(n8140), .A2(n8818), .ZN(n11373) );
  XOR2_X1 U11472 ( .A(n11556), .B(n11557), .Z(n11370) );
  XOR2_X1 U11473 ( .A(n11558), .B(n11559), .Z(n11557) );
  OR2_X1 U11474 ( .A1(n8810), .A2(n8818), .ZN(n11377) );
  XOR2_X1 U11475 ( .A(n11560), .B(n11561), .Z(n11374) );
  XOR2_X1 U11476 ( .A(n11562), .B(n8815), .Z(n11561) );
  OR2_X1 U11477 ( .A1(n8806), .A2(n8818), .ZN(n11381) );
  XOR2_X1 U11478 ( .A(n11563), .B(n11564), .Z(n11378) );
  XOR2_X1 U11479 ( .A(n11565), .B(n11566), .Z(n11564) );
  OR2_X1 U11480 ( .A1(n8802), .A2(n8818), .ZN(n11385) );
  XOR2_X1 U11481 ( .A(n11567), .B(n11568), .Z(n11382) );
  XOR2_X1 U11482 ( .A(n11569), .B(n11570), .Z(n11568) );
  OR2_X1 U11483 ( .A1(n8798), .A2(n8818), .ZN(n11389) );
  XOR2_X1 U11484 ( .A(n11571), .B(n11572), .Z(n11386) );
  XOR2_X1 U11485 ( .A(n11573), .B(n11574), .Z(n11572) );
  OR2_X1 U11486 ( .A1(n8794), .A2(n8818), .ZN(n11393) );
  XOR2_X1 U11487 ( .A(n11575), .B(n11576), .Z(n11390) );
  XOR2_X1 U11488 ( .A(n11577), .B(n11578), .Z(n11576) );
  OR2_X1 U11489 ( .A1(n8790), .A2(n8818), .ZN(n11397) );
  XOR2_X1 U11490 ( .A(n11579), .B(n11580), .Z(n11394) );
  XOR2_X1 U11491 ( .A(n11581), .B(n11582), .Z(n11580) );
  OR2_X1 U11492 ( .A1(n8786), .A2(n8818), .ZN(n11401) );
  XOR2_X1 U11493 ( .A(n11583), .B(n11584), .Z(n11398) );
  XOR2_X1 U11494 ( .A(n11585), .B(n11586), .Z(n11584) );
  XOR2_X1 U11495 ( .A(n11587), .B(n11588), .Z(n11403) );
  XOR2_X1 U11496 ( .A(n11589), .B(n11590), .Z(n11588) );
  OR2_X1 U11497 ( .A1(n8778), .A2(n8818), .ZN(n11409) );
  XOR2_X1 U11498 ( .A(n11591), .B(n11592), .Z(n11406) );
  XOR2_X1 U11499 ( .A(n11593), .B(n11594), .Z(n11592) );
  OR2_X1 U11500 ( .A1(n8774), .A2(n8818), .ZN(n11413) );
  XOR2_X1 U11501 ( .A(n11595), .B(n11596), .Z(n11410) );
  XOR2_X1 U11502 ( .A(n11597), .B(n11598), .Z(n11596) );
  OR2_X1 U11503 ( .A1(n8770), .A2(n8818), .ZN(n11417) );
  XOR2_X1 U11504 ( .A(n11599), .B(n11600), .Z(n11414) );
  XOR2_X1 U11505 ( .A(n11601), .B(n11602), .Z(n11600) );
  XOR2_X1 U11506 ( .A(n11603), .B(n11604), .Z(n11419) );
  XOR2_X1 U11507 ( .A(n11605), .B(n11606), .Z(n11604) );
  OR2_X1 U11508 ( .A1(n8762), .A2(n8818), .ZN(n11425) );
  XOR2_X1 U11509 ( .A(n11607), .B(n11608), .Z(n11422) );
  XOR2_X1 U11510 ( .A(n11609), .B(n11610), .Z(n11608) );
  OR2_X1 U11511 ( .A1(n8758), .A2(n8818), .ZN(n11429) );
  XOR2_X1 U11512 ( .A(n11611), .B(n11612), .Z(n11426) );
  XOR2_X1 U11513 ( .A(n11613), .B(n11614), .Z(n11612) );
  OR2_X1 U11514 ( .A1(n8754), .A2(n8818), .ZN(n11433) );
  XOR2_X1 U11515 ( .A(n11615), .B(n11616), .Z(n11430) );
  XOR2_X1 U11516 ( .A(n11617), .B(n11618), .Z(n11616) );
  XOR2_X1 U11517 ( .A(n11619), .B(n11620), .Z(n11435) );
  XOR2_X1 U11518 ( .A(n11621), .B(n11622), .Z(n11620) );
  OR2_X1 U11519 ( .A1(n8746), .A2(n8818), .ZN(n11441) );
  XOR2_X1 U11520 ( .A(n11623), .B(n11624), .Z(n11438) );
  XOR2_X1 U11521 ( .A(n11625), .B(n11626), .Z(n11624) );
  OR2_X1 U11522 ( .A1(n8742), .A2(n8818), .ZN(n11445) );
  XOR2_X1 U11523 ( .A(n11627), .B(n11628), .Z(n11442) );
  XOR2_X1 U11524 ( .A(n11629), .B(n11630), .Z(n11628) );
  XOR2_X1 U11525 ( .A(n11631), .B(n11632), .Z(n10834) );
  XOR2_X1 U11526 ( .A(n11633), .B(n11634), .Z(n11632) );
  OR2_X1 U11527 ( .A1(n11635), .A2(n9631), .ZN(n8925) );
  XOR2_X1 U11528 ( .A(n9579), .B(n9581), .Z(n9631) );
  OR2_X1 U11529 ( .A1(n11636), .A2(n11637), .ZN(n9581) );
  AND2_X1 U11530 ( .A1(n11638), .A2(n11639), .ZN(n11637) );
  AND2_X1 U11531 ( .A1(n11640), .A2(n11641), .ZN(n11636) );
  OR2_X1 U11532 ( .A1(n11638), .A2(n11639), .ZN(n11641) );
  XOR2_X1 U11533 ( .A(n9588), .B(n11642), .Z(n9579) );
  XOR2_X1 U11534 ( .A(n9587), .B(n9586), .Z(n11642) );
  OR2_X1 U11535 ( .A1(n9248), .A2(n8807), .ZN(n9586) );
  OR2_X1 U11536 ( .A1(n11643), .A2(n11644), .ZN(n9587) );
  AND2_X1 U11537 ( .A1(n11645), .A2(n11646), .ZN(n11644) );
  AND2_X1 U11538 ( .A1(n11647), .A2(n11648), .ZN(n11643) );
  OR2_X1 U11539 ( .A1(n11645), .A2(n11646), .ZN(n11648) );
  XOR2_X1 U11540 ( .A(n9595), .B(n11649), .Z(n9588) );
  XOR2_X1 U11541 ( .A(n9594), .B(n9593), .Z(n11649) );
  OR2_X1 U11542 ( .A1(n8730), .A2(n8803), .ZN(n9593) );
  OR2_X1 U11543 ( .A1(n11650), .A2(n11651), .ZN(n9594) );
  AND2_X1 U11544 ( .A1(n11652), .A2(n11653), .ZN(n11651) );
  AND2_X1 U11545 ( .A1(n11654), .A2(n11655), .ZN(n11650) );
  OR2_X1 U11546 ( .A1(n11652), .A2(n11653), .ZN(n11655) );
  XOR2_X1 U11547 ( .A(n9602), .B(n11656), .Z(n9595) );
  XOR2_X1 U11548 ( .A(n9601), .B(n9600), .Z(n11656) );
  OR2_X1 U11549 ( .A1(n8734), .A2(n8799), .ZN(n9600) );
  OR2_X1 U11550 ( .A1(n11657), .A2(n11658), .ZN(n9601) );
  AND2_X1 U11551 ( .A1(n11659), .A2(n11660), .ZN(n11658) );
  AND2_X1 U11552 ( .A1(n11661), .A2(n11662), .ZN(n11657) );
  OR2_X1 U11553 ( .A1(n11659), .A2(n11660), .ZN(n11662) );
  XOR2_X1 U11554 ( .A(n9609), .B(n11663), .Z(n9602) );
  XOR2_X1 U11555 ( .A(n9608), .B(n9607), .Z(n11663) );
  OR2_X1 U11556 ( .A1(n8738), .A2(n8795), .ZN(n9607) );
  OR2_X1 U11557 ( .A1(n11664), .A2(n11665), .ZN(n9608) );
  AND2_X1 U11558 ( .A1(n11666), .A2(n11667), .ZN(n11665) );
  AND2_X1 U11559 ( .A1(n11668), .A2(n11669), .ZN(n11664) );
  OR2_X1 U11560 ( .A1(n11666), .A2(n11667), .ZN(n11669) );
  XOR2_X1 U11561 ( .A(n9616), .B(n11670), .Z(n9609) );
  XOR2_X1 U11562 ( .A(n9615), .B(n9614), .Z(n11670) );
  OR2_X1 U11563 ( .A1(n8742), .A2(n8791), .ZN(n9614) );
  OR2_X1 U11564 ( .A1(n11671), .A2(n11672), .ZN(n9615) );
  AND2_X1 U11565 ( .A1(n11673), .A2(n11674), .ZN(n11672) );
  AND2_X1 U11566 ( .A1(n11675), .A2(n11676), .ZN(n11671) );
  OR2_X1 U11567 ( .A1(n11673), .A2(n11674), .ZN(n11676) );
  XOR2_X1 U11568 ( .A(n9623), .B(n11677), .Z(n9616) );
  XOR2_X1 U11569 ( .A(n9622), .B(n9621), .Z(n11677) );
  OR2_X1 U11570 ( .A1(n8746), .A2(n8787), .ZN(n9621) );
  OR2_X1 U11571 ( .A1(n11678), .A2(n11679), .ZN(n9622) );
  AND2_X1 U11572 ( .A1(n11680), .A2(n11681), .ZN(n11679) );
  AND2_X1 U11573 ( .A1(n11682), .A2(n11683), .ZN(n11678) );
  OR2_X1 U11574 ( .A1(n11681), .A2(n11680), .ZN(n11683) );
  XOR2_X1 U11575 ( .A(n11684), .B(n11685), .Z(n9623) );
  XOR2_X1 U11576 ( .A(n11686), .B(n11687), .Z(n11685) );
  AND2_X1 U11577 ( .A1(n9632), .A2(n9630), .ZN(n11635) );
  XNOR2_X1 U11578 ( .A(n11640), .B(n11688), .ZN(n9630) );
  XOR2_X1 U11579 ( .A(n11639), .B(n11638), .Z(n11688) );
  OR2_X1 U11580 ( .A1(n9248), .A2(n8811), .ZN(n11638) );
  OR2_X1 U11581 ( .A1(n11689), .A2(n11690), .ZN(n11639) );
  AND2_X1 U11582 ( .A1(n11691), .A2(n11692), .ZN(n11690) );
  AND2_X1 U11583 ( .A1(n11693), .A2(n11694), .ZN(n11689) );
  OR2_X1 U11584 ( .A1(n11691), .A2(n11692), .ZN(n11694) );
  XOR2_X1 U11585 ( .A(n11647), .B(n11695), .Z(n11640) );
  XOR2_X1 U11586 ( .A(n11646), .B(n11645), .Z(n11695) );
  OR2_X1 U11587 ( .A1(n8730), .A2(n8807), .ZN(n11645) );
  OR2_X1 U11588 ( .A1(n11696), .A2(n11697), .ZN(n11646) );
  AND2_X1 U11589 ( .A1(n11698), .A2(n11699), .ZN(n11697) );
  AND2_X1 U11590 ( .A1(n11700), .A2(n11701), .ZN(n11696) );
  OR2_X1 U11591 ( .A1(n11698), .A2(n11699), .ZN(n11701) );
  XOR2_X1 U11592 ( .A(n11654), .B(n11702), .Z(n11647) );
  XOR2_X1 U11593 ( .A(n11653), .B(n11652), .Z(n11702) );
  OR2_X1 U11594 ( .A1(n8734), .A2(n8803), .ZN(n11652) );
  OR2_X1 U11595 ( .A1(n11703), .A2(n11704), .ZN(n11653) );
  AND2_X1 U11596 ( .A1(n11705), .A2(n11706), .ZN(n11704) );
  AND2_X1 U11597 ( .A1(n11707), .A2(n11708), .ZN(n11703) );
  OR2_X1 U11598 ( .A1(n11705), .A2(n11706), .ZN(n11708) );
  XOR2_X1 U11599 ( .A(n11661), .B(n11709), .Z(n11654) );
  XOR2_X1 U11600 ( .A(n11660), .B(n11659), .Z(n11709) );
  OR2_X1 U11601 ( .A1(n8738), .A2(n8799), .ZN(n11659) );
  OR2_X1 U11602 ( .A1(n11710), .A2(n11711), .ZN(n11660) );
  AND2_X1 U11603 ( .A1(n11712), .A2(n11713), .ZN(n11711) );
  AND2_X1 U11604 ( .A1(n11714), .A2(n11715), .ZN(n11710) );
  OR2_X1 U11605 ( .A1(n11712), .A2(n11713), .ZN(n11715) );
  XOR2_X1 U11606 ( .A(n11668), .B(n11716), .Z(n11661) );
  XOR2_X1 U11607 ( .A(n11667), .B(n11666), .Z(n11716) );
  OR2_X1 U11608 ( .A1(n8742), .A2(n8795), .ZN(n11666) );
  OR2_X1 U11609 ( .A1(n11717), .A2(n11718), .ZN(n11667) );
  AND2_X1 U11610 ( .A1(n11719), .A2(n11720), .ZN(n11718) );
  AND2_X1 U11611 ( .A1(n11721), .A2(n11722), .ZN(n11717) );
  OR2_X1 U11612 ( .A1(n11719), .A2(n11720), .ZN(n11722) );
  XOR2_X1 U11613 ( .A(n11675), .B(n11723), .Z(n11668) );
  XOR2_X1 U11614 ( .A(n11674), .B(n11673), .Z(n11723) );
  OR2_X1 U11615 ( .A1(n8746), .A2(n8791), .ZN(n11673) );
  OR2_X1 U11616 ( .A1(n11724), .A2(n11725), .ZN(n11674) );
  AND2_X1 U11617 ( .A1(n11726), .A2(n11727), .ZN(n11725) );
  AND2_X1 U11618 ( .A1(n11728), .A2(n11729), .ZN(n11724) );
  OR2_X1 U11619 ( .A1(n11726), .A2(n11727), .ZN(n11729) );
  XOR2_X1 U11620 ( .A(n11682), .B(n11730), .Z(n11675) );
  XOR2_X1 U11621 ( .A(n11681), .B(n11680), .Z(n11730) );
  OR2_X1 U11622 ( .A1(n8750), .A2(n8787), .ZN(n11680) );
  OR2_X1 U11623 ( .A1(n11731), .A2(n11732), .ZN(n11681) );
  AND2_X1 U11624 ( .A1(n11733), .A2(n11734), .ZN(n11732) );
  AND2_X1 U11625 ( .A1(n11735), .A2(n11736), .ZN(n11731) );
  OR2_X1 U11626 ( .A1(n11734), .A2(n11733), .ZN(n11736) );
  XOR2_X1 U11627 ( .A(n11737), .B(n11738), .Z(n11682) );
  XOR2_X1 U11628 ( .A(n11739), .B(n11740), .Z(n11738) );
  INV_X1 U11629 ( .A(n9640), .ZN(n9632) );
  OR2_X1 U11630 ( .A1(n11741), .A2(n11742), .ZN(n9640) );
  AND2_X1 U11631 ( .A1(n9657), .A2(n9656), .ZN(n11742) );
  AND2_X1 U11632 ( .A1(n9654), .A2(n11743), .ZN(n11741) );
  OR2_X1 U11633 ( .A1(n9656), .A2(n9657), .ZN(n11743) );
  OR2_X1 U11634 ( .A1(n9248), .A2(n8814), .ZN(n9657) );
  OR2_X1 U11635 ( .A1(n11744), .A2(n11745), .ZN(n9656) );
  AND2_X1 U11636 ( .A1(n9681), .A2(n9680), .ZN(n11745) );
  AND2_X1 U11637 ( .A1(n9678), .A2(n11746), .ZN(n11744) );
  OR2_X1 U11638 ( .A1(n9680), .A2(n9681), .ZN(n11746) );
  OR2_X1 U11639 ( .A1(n8730), .A2(n8814), .ZN(n9681) );
  OR2_X1 U11640 ( .A1(n11747), .A2(n11748), .ZN(n9680) );
  AND2_X1 U11641 ( .A1(n10820), .A2(n10819), .ZN(n11748) );
  AND2_X1 U11642 ( .A1(n10817), .A2(n11749), .ZN(n11747) );
  OR2_X1 U11643 ( .A1(n10819), .A2(n10820), .ZN(n11749) );
  OR2_X1 U11644 ( .A1(n8734), .A2(n8814), .ZN(n10820) );
  OR2_X1 U11645 ( .A1(n11750), .A2(n11751), .ZN(n10819) );
  AND2_X1 U11646 ( .A1(n10839), .A2(n10838), .ZN(n11751) );
  AND2_X1 U11647 ( .A1(n10836), .A2(n11752), .ZN(n11750) );
  OR2_X1 U11648 ( .A1(n10838), .A2(n10839), .ZN(n11752) );
  OR2_X1 U11649 ( .A1(n8738), .A2(n8814), .ZN(n10839) );
  OR2_X1 U11650 ( .A1(n11753), .A2(n11754), .ZN(n10838) );
  AND2_X1 U11651 ( .A1(n11634), .A2(n11633), .ZN(n11754) );
  AND2_X1 U11652 ( .A1(n11631), .A2(n11755), .ZN(n11753) );
  OR2_X1 U11653 ( .A1(n11633), .A2(n11634), .ZN(n11755) );
  OR2_X1 U11654 ( .A1(n8742), .A2(n8814), .ZN(n11634) );
  OR2_X1 U11655 ( .A1(n11756), .A2(n11757), .ZN(n11633) );
  AND2_X1 U11656 ( .A1(n11630), .A2(n11629), .ZN(n11757) );
  AND2_X1 U11657 ( .A1(n11627), .A2(n11758), .ZN(n11756) );
  OR2_X1 U11658 ( .A1(n11629), .A2(n11630), .ZN(n11758) );
  OR2_X1 U11659 ( .A1(n8746), .A2(n8814), .ZN(n11630) );
  OR2_X1 U11660 ( .A1(n11759), .A2(n11760), .ZN(n11629) );
  AND2_X1 U11661 ( .A1(n11626), .A2(n11625), .ZN(n11760) );
  AND2_X1 U11662 ( .A1(n11623), .A2(n11761), .ZN(n11759) );
  OR2_X1 U11663 ( .A1(n11625), .A2(n11626), .ZN(n11761) );
  OR2_X1 U11664 ( .A1(n8750), .A2(n8814), .ZN(n11626) );
  OR2_X1 U11665 ( .A1(n11762), .A2(n11763), .ZN(n11625) );
  AND2_X1 U11666 ( .A1(n11622), .A2(n11621), .ZN(n11763) );
  AND2_X1 U11667 ( .A1(n11619), .A2(n11764), .ZN(n11762) );
  OR2_X1 U11668 ( .A1(n11621), .A2(n11622), .ZN(n11764) );
  OR2_X1 U11669 ( .A1(n8754), .A2(n8814), .ZN(n11622) );
  OR2_X1 U11670 ( .A1(n11765), .A2(n11766), .ZN(n11621) );
  AND2_X1 U11671 ( .A1(n11618), .A2(n11617), .ZN(n11766) );
  AND2_X1 U11672 ( .A1(n11615), .A2(n11767), .ZN(n11765) );
  OR2_X1 U11673 ( .A1(n11617), .A2(n11618), .ZN(n11767) );
  OR2_X1 U11674 ( .A1(n8758), .A2(n8814), .ZN(n11618) );
  OR2_X1 U11675 ( .A1(n11768), .A2(n11769), .ZN(n11617) );
  AND2_X1 U11676 ( .A1(n11614), .A2(n11613), .ZN(n11769) );
  AND2_X1 U11677 ( .A1(n11611), .A2(n11770), .ZN(n11768) );
  OR2_X1 U11678 ( .A1(n11613), .A2(n11614), .ZN(n11770) );
  OR2_X1 U11679 ( .A1(n8762), .A2(n8814), .ZN(n11614) );
  OR2_X1 U11680 ( .A1(n11771), .A2(n11772), .ZN(n11613) );
  AND2_X1 U11681 ( .A1(n11610), .A2(n11609), .ZN(n11772) );
  AND2_X1 U11682 ( .A1(n11607), .A2(n11773), .ZN(n11771) );
  OR2_X1 U11683 ( .A1(n11609), .A2(n11610), .ZN(n11773) );
  OR2_X1 U11684 ( .A1(n8766), .A2(n8814), .ZN(n11610) );
  OR2_X1 U11685 ( .A1(n11774), .A2(n11775), .ZN(n11609) );
  AND2_X1 U11686 ( .A1(n11606), .A2(n11605), .ZN(n11775) );
  AND2_X1 U11687 ( .A1(n11603), .A2(n11776), .ZN(n11774) );
  OR2_X1 U11688 ( .A1(n11605), .A2(n11606), .ZN(n11776) );
  OR2_X1 U11689 ( .A1(n8770), .A2(n8814), .ZN(n11606) );
  OR2_X1 U11690 ( .A1(n11777), .A2(n11778), .ZN(n11605) );
  AND2_X1 U11691 ( .A1(n11602), .A2(n11601), .ZN(n11778) );
  AND2_X1 U11692 ( .A1(n11599), .A2(n11779), .ZN(n11777) );
  OR2_X1 U11693 ( .A1(n11601), .A2(n11602), .ZN(n11779) );
  OR2_X1 U11694 ( .A1(n8774), .A2(n8814), .ZN(n11602) );
  OR2_X1 U11695 ( .A1(n11780), .A2(n11781), .ZN(n11601) );
  AND2_X1 U11696 ( .A1(n11598), .A2(n11597), .ZN(n11781) );
  AND2_X1 U11697 ( .A1(n11595), .A2(n11782), .ZN(n11780) );
  OR2_X1 U11698 ( .A1(n11597), .A2(n11598), .ZN(n11782) );
  OR2_X1 U11699 ( .A1(n8778), .A2(n8814), .ZN(n11598) );
  OR2_X1 U11700 ( .A1(n11783), .A2(n11784), .ZN(n11597) );
  AND2_X1 U11701 ( .A1(n11594), .A2(n11593), .ZN(n11784) );
  AND2_X1 U11702 ( .A1(n11591), .A2(n11785), .ZN(n11783) );
  OR2_X1 U11703 ( .A1(n11593), .A2(n11594), .ZN(n11785) );
  OR2_X1 U11704 ( .A1(n8782), .A2(n8814), .ZN(n11594) );
  OR2_X1 U11705 ( .A1(n11786), .A2(n11787), .ZN(n11593) );
  AND2_X1 U11706 ( .A1(n11590), .A2(n11589), .ZN(n11787) );
  AND2_X1 U11707 ( .A1(n11587), .A2(n11788), .ZN(n11786) );
  OR2_X1 U11708 ( .A1(n11589), .A2(n11590), .ZN(n11788) );
  OR2_X1 U11709 ( .A1(n8786), .A2(n8814), .ZN(n11590) );
  OR2_X1 U11710 ( .A1(n11789), .A2(n11790), .ZN(n11589) );
  AND2_X1 U11711 ( .A1(n11586), .A2(n11585), .ZN(n11790) );
  AND2_X1 U11712 ( .A1(n11583), .A2(n11791), .ZN(n11789) );
  OR2_X1 U11713 ( .A1(n11585), .A2(n11586), .ZN(n11791) );
  OR2_X1 U11714 ( .A1(n8790), .A2(n8814), .ZN(n11586) );
  OR2_X1 U11715 ( .A1(n11792), .A2(n11793), .ZN(n11585) );
  AND2_X1 U11716 ( .A1(n11582), .A2(n11581), .ZN(n11793) );
  AND2_X1 U11717 ( .A1(n11579), .A2(n11794), .ZN(n11792) );
  OR2_X1 U11718 ( .A1(n11581), .A2(n11582), .ZN(n11794) );
  OR2_X1 U11719 ( .A1(n8794), .A2(n8814), .ZN(n11582) );
  OR2_X1 U11720 ( .A1(n11795), .A2(n11796), .ZN(n11581) );
  AND2_X1 U11721 ( .A1(n11578), .A2(n11577), .ZN(n11796) );
  AND2_X1 U11722 ( .A1(n11575), .A2(n11797), .ZN(n11795) );
  OR2_X1 U11723 ( .A1(n11577), .A2(n11578), .ZN(n11797) );
  OR2_X1 U11724 ( .A1(n8798), .A2(n8814), .ZN(n11578) );
  OR2_X1 U11725 ( .A1(n11798), .A2(n11799), .ZN(n11577) );
  AND2_X1 U11726 ( .A1(n11574), .A2(n11573), .ZN(n11799) );
  AND2_X1 U11727 ( .A1(n11571), .A2(n11800), .ZN(n11798) );
  OR2_X1 U11728 ( .A1(n11573), .A2(n11574), .ZN(n11800) );
  OR2_X1 U11729 ( .A1(n8802), .A2(n8814), .ZN(n11574) );
  OR2_X1 U11730 ( .A1(n11801), .A2(n11802), .ZN(n11573) );
  AND2_X1 U11731 ( .A1(n11570), .A2(n11569), .ZN(n11802) );
  AND2_X1 U11732 ( .A1(n11567), .A2(n11803), .ZN(n11801) );
  OR2_X1 U11733 ( .A1(n11569), .A2(n11570), .ZN(n11803) );
  OR2_X1 U11734 ( .A1(n8806), .A2(n8814), .ZN(n11570) );
  OR2_X1 U11735 ( .A1(n11804), .A2(n11805), .ZN(n11569) );
  AND2_X1 U11736 ( .A1(n11566), .A2(n11565), .ZN(n11805) );
  AND2_X1 U11737 ( .A1(n11563), .A2(n11806), .ZN(n11804) );
  OR2_X1 U11738 ( .A1(n11565), .A2(n11566), .ZN(n11806) );
  OR2_X1 U11739 ( .A1(n8810), .A2(n8814), .ZN(n11566) );
  OR2_X1 U11740 ( .A1(n11807), .A2(n11808), .ZN(n11565) );
  AND2_X1 U11741 ( .A1(n8815), .A2(n11562), .ZN(n11808) );
  AND2_X1 U11742 ( .A1(n11560), .A2(n11809), .ZN(n11807) );
  OR2_X1 U11743 ( .A1(n11562), .A2(n8815), .ZN(n11809) );
  OR2_X1 U11744 ( .A1(n8140), .A2(n8814), .ZN(n8815) );
  OR2_X1 U11745 ( .A1(n11810), .A2(n11811), .ZN(n11562) );
  AND2_X1 U11746 ( .A1(n11559), .A2(n11558), .ZN(n11811) );
  AND2_X1 U11747 ( .A1(n11556), .A2(n11812), .ZN(n11810) );
  OR2_X1 U11748 ( .A1(n11558), .A2(n11559), .ZN(n11812) );
  OR2_X1 U11749 ( .A1(n8115), .A2(n8814), .ZN(n11559) );
  OR2_X1 U11750 ( .A1(n11813), .A2(n11814), .ZN(n11558) );
  AND2_X1 U11751 ( .A1(n11555), .A2(n11554), .ZN(n11814) );
  AND2_X1 U11752 ( .A1(n11552), .A2(n11815), .ZN(n11813) );
  OR2_X1 U11753 ( .A1(n11554), .A2(n11555), .ZN(n11815) );
  OR2_X1 U11754 ( .A1(n8090), .A2(n8814), .ZN(n11555) );
  OR2_X1 U11755 ( .A1(n11816), .A2(n11817), .ZN(n11554) );
  AND2_X1 U11756 ( .A1(n11551), .A2(n11550), .ZN(n11817) );
  AND2_X1 U11757 ( .A1(n11548), .A2(n11818), .ZN(n11816) );
  OR2_X1 U11758 ( .A1(n11550), .A2(n11551), .ZN(n11818) );
  OR2_X1 U11759 ( .A1(n8065), .A2(n8814), .ZN(n11551) );
  OR2_X1 U11760 ( .A1(n11819), .A2(n11820), .ZN(n11550) );
  AND2_X1 U11761 ( .A1(n11547), .A2(n11546), .ZN(n11820) );
  AND2_X1 U11762 ( .A1(n11544), .A2(n11821), .ZN(n11819) );
  OR2_X1 U11763 ( .A1(n11546), .A2(n11547), .ZN(n11821) );
  OR2_X1 U11764 ( .A1(n8040), .A2(n8814), .ZN(n11547) );
  OR2_X1 U11765 ( .A1(n11822), .A2(n11823), .ZN(n11546) );
  AND2_X1 U11766 ( .A1(n11543), .A2(n11542), .ZN(n11823) );
  AND2_X1 U11767 ( .A1(n11540), .A2(n11824), .ZN(n11822) );
  OR2_X1 U11768 ( .A1(n11542), .A2(n11543), .ZN(n11824) );
  OR2_X1 U11769 ( .A1(n8015), .A2(n8814), .ZN(n11543) );
  OR2_X1 U11770 ( .A1(n11825), .A2(n11826), .ZN(n11542) );
  AND2_X1 U11771 ( .A1(n11539), .A2(n11538), .ZN(n11826) );
  AND2_X1 U11772 ( .A1(n11536), .A2(n11827), .ZN(n11825) );
  OR2_X1 U11773 ( .A1(n11538), .A2(n11539), .ZN(n11827) );
  OR2_X1 U11774 ( .A1(n7979), .A2(n8814), .ZN(n11539) );
  OR2_X1 U11775 ( .A1(n11828), .A2(n11829), .ZN(n11538) );
  AND2_X1 U11776 ( .A1(n11532), .A2(n11535), .ZN(n11829) );
  AND2_X1 U11777 ( .A1(n11830), .A2(n11831), .ZN(n11828) );
  OR2_X1 U11778 ( .A1(n11535), .A2(n11532), .ZN(n11831) );
  OR2_X1 U11779 ( .A1(n7954), .A2(n8814), .ZN(n11532) );
  OR3_X1 U11780 ( .A1(n8814), .A2(n8811), .A3(n9796), .ZN(n11535) );
  INV_X1 U11781 ( .A(n11534), .ZN(n11830) );
  OR2_X1 U11782 ( .A1(n11832), .A2(n11833), .ZN(n11534) );
  AND2_X1 U11783 ( .A1(b_21_), .A2(n11834), .ZN(n11833) );
  OR2_X1 U11784 ( .A1(n11835), .A2(n9801), .ZN(n11834) );
  AND2_X1 U11785 ( .A1(a_30_), .A2(n8807), .ZN(n11835) );
  AND2_X1 U11786 ( .A1(b_20_), .A2(n11836), .ZN(n11832) );
  OR2_X1 U11787 ( .A1(n11837), .A2(n7920), .ZN(n11836) );
  AND2_X1 U11788 ( .A1(a_31_), .A2(n8811), .ZN(n11837) );
  XNOR2_X1 U11789 ( .A(n11838), .B(n11839), .ZN(n11536) );
  XOR2_X1 U11790 ( .A(n11840), .B(n11841), .Z(n11839) );
  XOR2_X1 U11791 ( .A(n11842), .B(n11843), .Z(n11540) );
  XOR2_X1 U11792 ( .A(n11844), .B(n11845), .Z(n11843) );
  XOR2_X1 U11793 ( .A(n11846), .B(n11847), .Z(n11544) );
  XOR2_X1 U11794 ( .A(n11848), .B(n11849), .Z(n11847) );
  XOR2_X1 U11795 ( .A(n11850), .B(n11851), .Z(n11548) );
  XOR2_X1 U11796 ( .A(n11852), .B(n11853), .Z(n11851) );
  XOR2_X1 U11797 ( .A(n11854), .B(n11855), .Z(n11552) );
  XOR2_X1 U11798 ( .A(n11856), .B(n11857), .Z(n11855) );
  XOR2_X1 U11799 ( .A(n11858), .B(n11859), .Z(n11556) );
  XOR2_X1 U11800 ( .A(n11860), .B(n11861), .Z(n11859) );
  XOR2_X1 U11801 ( .A(n11862), .B(n11863), .Z(n11560) );
  XOR2_X1 U11802 ( .A(n11864), .B(n11865), .Z(n11863) );
  XOR2_X1 U11803 ( .A(n11866), .B(n11867), .Z(n11563) );
  XOR2_X1 U11804 ( .A(n11868), .B(n11869), .Z(n11867) );
  XOR2_X1 U11805 ( .A(n11870), .B(n11871), .Z(n11567) );
  XOR2_X1 U11806 ( .A(n11872), .B(n8162), .Z(n11871) );
  XOR2_X1 U11807 ( .A(n11873), .B(n11874), .Z(n11571) );
  XOR2_X1 U11808 ( .A(n11875), .B(n11876), .Z(n11874) );
  XOR2_X1 U11809 ( .A(n11877), .B(n11878), .Z(n11575) );
  XOR2_X1 U11810 ( .A(n11879), .B(n11880), .Z(n11878) );
  XOR2_X1 U11811 ( .A(n11881), .B(n11882), .Z(n11579) );
  XOR2_X1 U11812 ( .A(n11883), .B(n11884), .Z(n11882) );
  XOR2_X1 U11813 ( .A(n11885), .B(n11886), .Z(n11583) );
  XOR2_X1 U11814 ( .A(n11887), .B(n11888), .Z(n11886) );
  XOR2_X1 U11815 ( .A(n11889), .B(n11890), .Z(n11587) );
  XOR2_X1 U11816 ( .A(n11891), .B(n11892), .Z(n11890) );
  XOR2_X1 U11817 ( .A(n11893), .B(n11894), .Z(n11591) );
  XOR2_X1 U11818 ( .A(n11895), .B(n11896), .Z(n11894) );
  XOR2_X1 U11819 ( .A(n11897), .B(n11898), .Z(n11595) );
  XOR2_X1 U11820 ( .A(n11899), .B(n11900), .Z(n11898) );
  XOR2_X1 U11821 ( .A(n11901), .B(n11902), .Z(n11599) );
  XOR2_X1 U11822 ( .A(n11903), .B(n11904), .Z(n11902) );
  XOR2_X1 U11823 ( .A(n11905), .B(n11906), .Z(n11603) );
  XOR2_X1 U11824 ( .A(n11907), .B(n11908), .Z(n11906) );
  XOR2_X1 U11825 ( .A(n11909), .B(n11910), .Z(n11607) );
  XOR2_X1 U11826 ( .A(n11911), .B(n11912), .Z(n11910) );
  XOR2_X1 U11827 ( .A(n11913), .B(n11914), .Z(n11611) );
  XOR2_X1 U11828 ( .A(n11915), .B(n11916), .Z(n11914) );
  XOR2_X1 U11829 ( .A(n11917), .B(n11918), .Z(n11615) );
  XOR2_X1 U11830 ( .A(n11919), .B(n11920), .Z(n11918) );
  XOR2_X1 U11831 ( .A(n11921), .B(n11922), .Z(n11619) );
  XOR2_X1 U11832 ( .A(n11923), .B(n11924), .Z(n11922) );
  XOR2_X1 U11833 ( .A(n11925), .B(n11926), .Z(n11623) );
  XOR2_X1 U11834 ( .A(n11927), .B(n11928), .Z(n11926) );
  XOR2_X1 U11835 ( .A(n11929), .B(n11930), .Z(n11627) );
  XOR2_X1 U11836 ( .A(n11931), .B(n11932), .Z(n11930) );
  XOR2_X1 U11837 ( .A(n11933), .B(n11934), .Z(n11631) );
  XOR2_X1 U11838 ( .A(n11935), .B(n11936), .Z(n11934) );
  XOR2_X1 U11839 ( .A(n11937), .B(n11938), .Z(n10836) );
  XOR2_X1 U11840 ( .A(n11939), .B(n11940), .Z(n11938) );
  XOR2_X1 U11841 ( .A(n11941), .B(n11942), .Z(n10817) );
  XOR2_X1 U11842 ( .A(n11943), .B(n11944), .Z(n11942) );
  XOR2_X1 U11843 ( .A(n11945), .B(n11946), .Z(n9678) );
  XOR2_X1 U11844 ( .A(n11947), .B(n11948), .Z(n11946) );
  XOR2_X1 U11845 ( .A(n11693), .B(n11949), .Z(n9654) );
  XOR2_X1 U11846 ( .A(n11692), .B(n11691), .Z(n11949) );
  OR2_X1 U11847 ( .A1(n8730), .A2(n8811), .ZN(n11691) );
  OR2_X1 U11848 ( .A1(n11950), .A2(n11951), .ZN(n11692) );
  AND2_X1 U11849 ( .A1(n11948), .A2(n11947), .ZN(n11951) );
  AND2_X1 U11850 ( .A1(n11945), .A2(n11952), .ZN(n11950) );
  OR2_X1 U11851 ( .A1(n11948), .A2(n11947), .ZN(n11952) );
  OR2_X1 U11852 ( .A1(n11953), .A2(n11954), .ZN(n11947) );
  AND2_X1 U11853 ( .A1(n11944), .A2(n11943), .ZN(n11954) );
  AND2_X1 U11854 ( .A1(n11941), .A2(n11955), .ZN(n11953) );
  OR2_X1 U11855 ( .A1(n11944), .A2(n11943), .ZN(n11955) );
  OR2_X1 U11856 ( .A1(n11956), .A2(n11957), .ZN(n11943) );
  AND2_X1 U11857 ( .A1(n11940), .A2(n11939), .ZN(n11957) );
  AND2_X1 U11858 ( .A1(n11937), .A2(n11958), .ZN(n11956) );
  OR2_X1 U11859 ( .A1(n11940), .A2(n11939), .ZN(n11958) );
  OR2_X1 U11860 ( .A1(n11959), .A2(n11960), .ZN(n11939) );
  AND2_X1 U11861 ( .A1(n11936), .A2(n11935), .ZN(n11960) );
  AND2_X1 U11862 ( .A1(n11933), .A2(n11961), .ZN(n11959) );
  OR2_X1 U11863 ( .A1(n11936), .A2(n11935), .ZN(n11961) );
  OR2_X1 U11864 ( .A1(n11962), .A2(n11963), .ZN(n11935) );
  AND2_X1 U11865 ( .A1(n11932), .A2(n11931), .ZN(n11963) );
  AND2_X1 U11866 ( .A1(n11929), .A2(n11964), .ZN(n11962) );
  OR2_X1 U11867 ( .A1(n11932), .A2(n11931), .ZN(n11964) );
  OR2_X1 U11868 ( .A1(n11965), .A2(n11966), .ZN(n11931) );
  AND2_X1 U11869 ( .A1(n11928), .A2(n11927), .ZN(n11966) );
  AND2_X1 U11870 ( .A1(n11925), .A2(n11967), .ZN(n11965) );
  OR2_X1 U11871 ( .A1(n11928), .A2(n11927), .ZN(n11967) );
  OR2_X1 U11872 ( .A1(n11968), .A2(n11969), .ZN(n11927) );
  AND2_X1 U11873 ( .A1(n11924), .A2(n11923), .ZN(n11969) );
  AND2_X1 U11874 ( .A1(n11921), .A2(n11970), .ZN(n11968) );
  OR2_X1 U11875 ( .A1(n11924), .A2(n11923), .ZN(n11970) );
  OR2_X1 U11876 ( .A1(n11971), .A2(n11972), .ZN(n11923) );
  AND2_X1 U11877 ( .A1(n11920), .A2(n11919), .ZN(n11972) );
  AND2_X1 U11878 ( .A1(n11917), .A2(n11973), .ZN(n11971) );
  OR2_X1 U11879 ( .A1(n11920), .A2(n11919), .ZN(n11973) );
  OR2_X1 U11880 ( .A1(n11974), .A2(n11975), .ZN(n11919) );
  AND2_X1 U11881 ( .A1(n11916), .A2(n11915), .ZN(n11975) );
  AND2_X1 U11882 ( .A1(n11913), .A2(n11976), .ZN(n11974) );
  OR2_X1 U11883 ( .A1(n11916), .A2(n11915), .ZN(n11976) );
  OR2_X1 U11884 ( .A1(n11977), .A2(n11978), .ZN(n11915) );
  AND2_X1 U11885 ( .A1(n11912), .A2(n11911), .ZN(n11978) );
  AND2_X1 U11886 ( .A1(n11909), .A2(n11979), .ZN(n11977) );
  OR2_X1 U11887 ( .A1(n11912), .A2(n11911), .ZN(n11979) );
  OR2_X1 U11888 ( .A1(n11980), .A2(n11981), .ZN(n11911) );
  AND2_X1 U11889 ( .A1(n11908), .A2(n11907), .ZN(n11981) );
  AND2_X1 U11890 ( .A1(n11905), .A2(n11982), .ZN(n11980) );
  OR2_X1 U11891 ( .A1(n11908), .A2(n11907), .ZN(n11982) );
  OR2_X1 U11892 ( .A1(n11983), .A2(n11984), .ZN(n11907) );
  AND2_X1 U11893 ( .A1(n11904), .A2(n11903), .ZN(n11984) );
  AND2_X1 U11894 ( .A1(n11901), .A2(n11985), .ZN(n11983) );
  OR2_X1 U11895 ( .A1(n11904), .A2(n11903), .ZN(n11985) );
  OR2_X1 U11896 ( .A1(n11986), .A2(n11987), .ZN(n11903) );
  AND2_X1 U11897 ( .A1(n11900), .A2(n11899), .ZN(n11987) );
  AND2_X1 U11898 ( .A1(n11897), .A2(n11988), .ZN(n11986) );
  OR2_X1 U11899 ( .A1(n11900), .A2(n11899), .ZN(n11988) );
  OR2_X1 U11900 ( .A1(n11989), .A2(n11990), .ZN(n11899) );
  AND2_X1 U11901 ( .A1(n11896), .A2(n11895), .ZN(n11990) );
  AND2_X1 U11902 ( .A1(n11893), .A2(n11991), .ZN(n11989) );
  OR2_X1 U11903 ( .A1(n11896), .A2(n11895), .ZN(n11991) );
  OR2_X1 U11904 ( .A1(n11992), .A2(n11993), .ZN(n11895) );
  AND2_X1 U11905 ( .A1(n11892), .A2(n11891), .ZN(n11993) );
  AND2_X1 U11906 ( .A1(n11889), .A2(n11994), .ZN(n11992) );
  OR2_X1 U11907 ( .A1(n11892), .A2(n11891), .ZN(n11994) );
  OR2_X1 U11908 ( .A1(n11995), .A2(n11996), .ZN(n11891) );
  AND2_X1 U11909 ( .A1(n11888), .A2(n11887), .ZN(n11996) );
  AND2_X1 U11910 ( .A1(n11885), .A2(n11997), .ZN(n11995) );
  OR2_X1 U11911 ( .A1(n11888), .A2(n11887), .ZN(n11997) );
  OR2_X1 U11912 ( .A1(n11998), .A2(n11999), .ZN(n11887) );
  AND2_X1 U11913 ( .A1(n11884), .A2(n11883), .ZN(n11999) );
  AND2_X1 U11914 ( .A1(n11881), .A2(n12000), .ZN(n11998) );
  OR2_X1 U11915 ( .A1(n11884), .A2(n11883), .ZN(n12000) );
  OR2_X1 U11916 ( .A1(n12001), .A2(n12002), .ZN(n11883) );
  AND2_X1 U11917 ( .A1(n11880), .A2(n11879), .ZN(n12002) );
  AND2_X1 U11918 ( .A1(n11877), .A2(n12003), .ZN(n12001) );
  OR2_X1 U11919 ( .A1(n11880), .A2(n11879), .ZN(n12003) );
  OR2_X1 U11920 ( .A1(n12004), .A2(n12005), .ZN(n11879) );
  AND2_X1 U11921 ( .A1(n11876), .A2(n11875), .ZN(n12005) );
  AND2_X1 U11922 ( .A1(n11873), .A2(n12006), .ZN(n12004) );
  OR2_X1 U11923 ( .A1(n11876), .A2(n11875), .ZN(n12006) );
  OR2_X1 U11924 ( .A1(n12007), .A2(n12008), .ZN(n11875) );
  AND2_X1 U11925 ( .A1(n8162), .A2(n11872), .ZN(n12008) );
  AND2_X1 U11926 ( .A1(n11870), .A2(n12009), .ZN(n12007) );
  OR2_X1 U11927 ( .A1(n8162), .A2(n11872), .ZN(n12009) );
  OR2_X1 U11928 ( .A1(n12010), .A2(n12011), .ZN(n11872) );
  AND2_X1 U11929 ( .A1(n11869), .A2(n11868), .ZN(n12011) );
  AND2_X1 U11930 ( .A1(n11866), .A2(n12012), .ZN(n12010) );
  OR2_X1 U11931 ( .A1(n11869), .A2(n11868), .ZN(n12012) );
  OR2_X1 U11932 ( .A1(n12013), .A2(n12014), .ZN(n11868) );
  AND2_X1 U11933 ( .A1(n11865), .A2(n11864), .ZN(n12014) );
  AND2_X1 U11934 ( .A1(n11862), .A2(n12015), .ZN(n12013) );
  OR2_X1 U11935 ( .A1(n11865), .A2(n11864), .ZN(n12015) );
  OR2_X1 U11936 ( .A1(n12016), .A2(n12017), .ZN(n11864) );
  AND2_X1 U11937 ( .A1(n11861), .A2(n11860), .ZN(n12017) );
  AND2_X1 U11938 ( .A1(n11858), .A2(n12018), .ZN(n12016) );
  OR2_X1 U11939 ( .A1(n11861), .A2(n11860), .ZN(n12018) );
  OR2_X1 U11940 ( .A1(n12019), .A2(n12020), .ZN(n11860) );
  AND2_X1 U11941 ( .A1(n11857), .A2(n11856), .ZN(n12020) );
  AND2_X1 U11942 ( .A1(n11854), .A2(n12021), .ZN(n12019) );
  OR2_X1 U11943 ( .A1(n11857), .A2(n11856), .ZN(n12021) );
  OR2_X1 U11944 ( .A1(n12022), .A2(n12023), .ZN(n11856) );
  AND2_X1 U11945 ( .A1(n11853), .A2(n11852), .ZN(n12023) );
  AND2_X1 U11946 ( .A1(n11850), .A2(n12024), .ZN(n12022) );
  OR2_X1 U11947 ( .A1(n11853), .A2(n11852), .ZN(n12024) );
  OR2_X1 U11948 ( .A1(n12025), .A2(n12026), .ZN(n11852) );
  AND2_X1 U11949 ( .A1(n11849), .A2(n11848), .ZN(n12026) );
  AND2_X1 U11950 ( .A1(n11846), .A2(n12027), .ZN(n12025) );
  OR2_X1 U11951 ( .A1(n11849), .A2(n11848), .ZN(n12027) );
  OR2_X1 U11952 ( .A1(n12028), .A2(n12029), .ZN(n11848) );
  AND2_X1 U11953 ( .A1(n11845), .A2(n11844), .ZN(n12029) );
  AND2_X1 U11954 ( .A1(n11842), .A2(n12030), .ZN(n12028) );
  OR2_X1 U11955 ( .A1(n11845), .A2(n11844), .ZN(n12030) );
  OR2_X1 U11956 ( .A1(n12031), .A2(n12032), .ZN(n11844) );
  AND2_X1 U11957 ( .A1(n11838), .A2(n11841), .ZN(n12032) );
  AND2_X1 U11958 ( .A1(n12033), .A2(n12034), .ZN(n12031) );
  OR2_X1 U11959 ( .A1(n11838), .A2(n11841), .ZN(n12034) );
  OR3_X1 U11960 ( .A1(n8811), .A2(n8807), .A3(n9796), .ZN(n11841) );
  OR2_X1 U11961 ( .A1(n7954), .A2(n8811), .ZN(n11838) );
  INV_X1 U11962 ( .A(n11840), .ZN(n12033) );
  OR2_X1 U11963 ( .A1(n12035), .A2(n12036), .ZN(n11840) );
  AND2_X1 U11964 ( .A1(b_20_), .A2(n12037), .ZN(n12036) );
  OR2_X1 U11965 ( .A1(n12038), .A2(n9801), .ZN(n12037) );
  AND2_X1 U11966 ( .A1(a_30_), .A2(n8803), .ZN(n12038) );
  AND2_X1 U11967 ( .A1(b_19_), .A2(n12039), .ZN(n12035) );
  OR2_X1 U11968 ( .A1(n12040), .A2(n7920), .ZN(n12039) );
  AND2_X1 U11969 ( .A1(a_31_), .A2(n8807), .ZN(n12040) );
  OR2_X1 U11970 ( .A1(n7979), .A2(n8811), .ZN(n11845) );
  XNOR2_X1 U11971 ( .A(n12041), .B(n12042), .ZN(n11842) );
  XOR2_X1 U11972 ( .A(n12043), .B(n12044), .Z(n12042) );
  OR2_X1 U11973 ( .A1(n8015), .A2(n8811), .ZN(n11849) );
  XOR2_X1 U11974 ( .A(n12045), .B(n12046), .Z(n11846) );
  XOR2_X1 U11975 ( .A(n12047), .B(n12048), .Z(n12046) );
  OR2_X1 U11976 ( .A1(n8040), .A2(n8811), .ZN(n11853) );
  XOR2_X1 U11977 ( .A(n12049), .B(n12050), .Z(n11850) );
  XOR2_X1 U11978 ( .A(n12051), .B(n12052), .Z(n12050) );
  OR2_X1 U11979 ( .A1(n8065), .A2(n8811), .ZN(n11857) );
  XOR2_X1 U11980 ( .A(n12053), .B(n12054), .Z(n11854) );
  XOR2_X1 U11981 ( .A(n12055), .B(n12056), .Z(n12054) );
  OR2_X1 U11982 ( .A1(n8090), .A2(n8811), .ZN(n11861) );
  XOR2_X1 U11983 ( .A(n12057), .B(n12058), .Z(n11858) );
  XOR2_X1 U11984 ( .A(n12059), .B(n12060), .Z(n12058) );
  OR2_X1 U11985 ( .A1(n8115), .A2(n8811), .ZN(n11865) );
  XOR2_X1 U11986 ( .A(n12061), .B(n12062), .Z(n11862) );
  XOR2_X1 U11987 ( .A(n12063), .B(n12064), .Z(n12062) );
  OR2_X1 U11988 ( .A1(n8140), .A2(n8811), .ZN(n11869) );
  XOR2_X1 U11989 ( .A(n12065), .B(n12066), .Z(n11866) );
  XOR2_X1 U11990 ( .A(n12067), .B(n12068), .Z(n12066) );
  OR2_X1 U11991 ( .A1(n8810), .A2(n8811), .ZN(n8162) );
  XOR2_X1 U11992 ( .A(n12069), .B(n12070), .Z(n11870) );
  XOR2_X1 U11993 ( .A(n12071), .B(n12072), .Z(n12070) );
  OR2_X1 U11994 ( .A1(n8806), .A2(n8811), .ZN(n11876) );
  XOR2_X1 U11995 ( .A(n12073), .B(n12074), .Z(n11873) );
  XOR2_X1 U11996 ( .A(n12075), .B(n12076), .Z(n12074) );
  OR2_X1 U11997 ( .A1(n8802), .A2(n8811), .ZN(n11880) );
  XOR2_X1 U11998 ( .A(n12077), .B(n12078), .Z(n11877) );
  XOR2_X1 U11999 ( .A(n12079), .B(n8188), .Z(n12078) );
  OR2_X1 U12000 ( .A1(n8798), .A2(n8811), .ZN(n11884) );
  XOR2_X1 U12001 ( .A(n12080), .B(n12081), .Z(n11881) );
  XOR2_X1 U12002 ( .A(n12082), .B(n12083), .Z(n12081) );
  OR2_X1 U12003 ( .A1(n8794), .A2(n8811), .ZN(n11888) );
  XOR2_X1 U12004 ( .A(n12084), .B(n12085), .Z(n11885) );
  XOR2_X1 U12005 ( .A(n12086), .B(n12087), .Z(n12085) );
  OR2_X1 U12006 ( .A1(n8790), .A2(n8811), .ZN(n11892) );
  XOR2_X1 U12007 ( .A(n12088), .B(n12089), .Z(n11889) );
  XOR2_X1 U12008 ( .A(n12090), .B(n12091), .Z(n12089) );
  OR2_X1 U12009 ( .A1(n8786), .A2(n8811), .ZN(n11896) );
  XOR2_X1 U12010 ( .A(n12092), .B(n12093), .Z(n11893) );
  XOR2_X1 U12011 ( .A(n12094), .B(n12095), .Z(n12093) );
  OR2_X1 U12012 ( .A1(n8782), .A2(n8811), .ZN(n11900) );
  XOR2_X1 U12013 ( .A(n12096), .B(n12097), .Z(n11897) );
  XOR2_X1 U12014 ( .A(n12098), .B(n12099), .Z(n12097) );
  OR2_X1 U12015 ( .A1(n8778), .A2(n8811), .ZN(n11904) );
  XOR2_X1 U12016 ( .A(n12100), .B(n12101), .Z(n11901) );
  XOR2_X1 U12017 ( .A(n12102), .B(n12103), .Z(n12101) );
  OR2_X1 U12018 ( .A1(n8774), .A2(n8811), .ZN(n11908) );
  XOR2_X1 U12019 ( .A(n12104), .B(n12105), .Z(n11905) );
  XOR2_X1 U12020 ( .A(n12106), .B(n12107), .Z(n12105) );
  OR2_X1 U12021 ( .A1(n8770), .A2(n8811), .ZN(n11912) );
  XOR2_X1 U12022 ( .A(n12108), .B(n12109), .Z(n11909) );
  XOR2_X1 U12023 ( .A(n12110), .B(n12111), .Z(n12109) );
  OR2_X1 U12024 ( .A1(n8766), .A2(n8811), .ZN(n11916) );
  XOR2_X1 U12025 ( .A(n12112), .B(n12113), .Z(n11913) );
  XOR2_X1 U12026 ( .A(n12114), .B(n12115), .Z(n12113) );
  OR2_X1 U12027 ( .A1(n8762), .A2(n8811), .ZN(n11920) );
  XOR2_X1 U12028 ( .A(n12116), .B(n12117), .Z(n11917) );
  XOR2_X1 U12029 ( .A(n12118), .B(n12119), .Z(n12117) );
  OR2_X1 U12030 ( .A1(n8758), .A2(n8811), .ZN(n11924) );
  XOR2_X1 U12031 ( .A(n12120), .B(n12121), .Z(n11921) );
  XOR2_X1 U12032 ( .A(n12122), .B(n12123), .Z(n12121) );
  OR2_X1 U12033 ( .A1(n8754), .A2(n8811), .ZN(n11928) );
  XOR2_X1 U12034 ( .A(n12124), .B(n12125), .Z(n11925) );
  XOR2_X1 U12035 ( .A(n12126), .B(n12127), .Z(n12125) );
  OR2_X1 U12036 ( .A1(n8750), .A2(n8811), .ZN(n11932) );
  XOR2_X1 U12037 ( .A(n12128), .B(n12129), .Z(n11929) );
  XOR2_X1 U12038 ( .A(n12130), .B(n12131), .Z(n12129) );
  OR2_X1 U12039 ( .A1(n8746), .A2(n8811), .ZN(n11936) );
  XOR2_X1 U12040 ( .A(n12132), .B(n12133), .Z(n11933) );
  XOR2_X1 U12041 ( .A(n12134), .B(n12135), .Z(n12133) );
  OR2_X1 U12042 ( .A1(n8742), .A2(n8811), .ZN(n11940) );
  XOR2_X1 U12043 ( .A(n12136), .B(n12137), .Z(n11937) );
  XOR2_X1 U12044 ( .A(n12138), .B(n12139), .Z(n12137) );
  OR2_X1 U12045 ( .A1(n8738), .A2(n8811), .ZN(n11944) );
  XOR2_X1 U12046 ( .A(n12140), .B(n12141), .Z(n11941) );
  XOR2_X1 U12047 ( .A(n12142), .B(n12143), .Z(n12141) );
  OR2_X1 U12048 ( .A1(n8734), .A2(n8811), .ZN(n11948) );
  XOR2_X1 U12049 ( .A(n12144), .B(n12145), .Z(n11945) );
  XOR2_X1 U12050 ( .A(n12146), .B(n12147), .Z(n12145) );
  XOR2_X1 U12051 ( .A(n11700), .B(n12148), .Z(n11693) );
  XOR2_X1 U12052 ( .A(n11699), .B(n11698), .Z(n12148) );
  OR2_X1 U12053 ( .A1(n8734), .A2(n8807), .ZN(n11698) );
  OR2_X1 U12054 ( .A1(n12149), .A2(n12150), .ZN(n11699) );
  AND2_X1 U12055 ( .A1(n12147), .A2(n12146), .ZN(n12150) );
  AND2_X1 U12056 ( .A1(n12144), .A2(n12151), .ZN(n12149) );
  OR2_X1 U12057 ( .A1(n12147), .A2(n12146), .ZN(n12151) );
  OR2_X1 U12058 ( .A1(n12152), .A2(n12153), .ZN(n12146) );
  AND2_X1 U12059 ( .A1(n12143), .A2(n12142), .ZN(n12153) );
  AND2_X1 U12060 ( .A1(n12140), .A2(n12154), .ZN(n12152) );
  OR2_X1 U12061 ( .A1(n12143), .A2(n12142), .ZN(n12154) );
  OR2_X1 U12062 ( .A1(n12155), .A2(n12156), .ZN(n12142) );
  AND2_X1 U12063 ( .A1(n12139), .A2(n12138), .ZN(n12156) );
  AND2_X1 U12064 ( .A1(n12136), .A2(n12157), .ZN(n12155) );
  OR2_X1 U12065 ( .A1(n12139), .A2(n12138), .ZN(n12157) );
  OR2_X1 U12066 ( .A1(n12158), .A2(n12159), .ZN(n12138) );
  AND2_X1 U12067 ( .A1(n12135), .A2(n12134), .ZN(n12159) );
  AND2_X1 U12068 ( .A1(n12132), .A2(n12160), .ZN(n12158) );
  OR2_X1 U12069 ( .A1(n12135), .A2(n12134), .ZN(n12160) );
  OR2_X1 U12070 ( .A1(n12161), .A2(n12162), .ZN(n12134) );
  AND2_X1 U12071 ( .A1(n12131), .A2(n12130), .ZN(n12162) );
  AND2_X1 U12072 ( .A1(n12128), .A2(n12163), .ZN(n12161) );
  OR2_X1 U12073 ( .A1(n12131), .A2(n12130), .ZN(n12163) );
  OR2_X1 U12074 ( .A1(n12164), .A2(n12165), .ZN(n12130) );
  AND2_X1 U12075 ( .A1(n12127), .A2(n12126), .ZN(n12165) );
  AND2_X1 U12076 ( .A1(n12124), .A2(n12166), .ZN(n12164) );
  OR2_X1 U12077 ( .A1(n12127), .A2(n12126), .ZN(n12166) );
  OR2_X1 U12078 ( .A1(n12167), .A2(n12168), .ZN(n12126) );
  AND2_X1 U12079 ( .A1(n12123), .A2(n12122), .ZN(n12168) );
  AND2_X1 U12080 ( .A1(n12120), .A2(n12169), .ZN(n12167) );
  OR2_X1 U12081 ( .A1(n12123), .A2(n12122), .ZN(n12169) );
  OR2_X1 U12082 ( .A1(n12170), .A2(n12171), .ZN(n12122) );
  AND2_X1 U12083 ( .A1(n12119), .A2(n12118), .ZN(n12171) );
  AND2_X1 U12084 ( .A1(n12116), .A2(n12172), .ZN(n12170) );
  OR2_X1 U12085 ( .A1(n12119), .A2(n12118), .ZN(n12172) );
  OR2_X1 U12086 ( .A1(n12173), .A2(n12174), .ZN(n12118) );
  AND2_X1 U12087 ( .A1(n12115), .A2(n12114), .ZN(n12174) );
  AND2_X1 U12088 ( .A1(n12112), .A2(n12175), .ZN(n12173) );
  OR2_X1 U12089 ( .A1(n12115), .A2(n12114), .ZN(n12175) );
  OR2_X1 U12090 ( .A1(n12176), .A2(n12177), .ZN(n12114) );
  AND2_X1 U12091 ( .A1(n12111), .A2(n12110), .ZN(n12177) );
  AND2_X1 U12092 ( .A1(n12108), .A2(n12178), .ZN(n12176) );
  OR2_X1 U12093 ( .A1(n12111), .A2(n12110), .ZN(n12178) );
  OR2_X1 U12094 ( .A1(n12179), .A2(n12180), .ZN(n12110) );
  AND2_X1 U12095 ( .A1(n12107), .A2(n12106), .ZN(n12180) );
  AND2_X1 U12096 ( .A1(n12104), .A2(n12181), .ZN(n12179) );
  OR2_X1 U12097 ( .A1(n12107), .A2(n12106), .ZN(n12181) );
  OR2_X1 U12098 ( .A1(n12182), .A2(n12183), .ZN(n12106) );
  AND2_X1 U12099 ( .A1(n12103), .A2(n12102), .ZN(n12183) );
  AND2_X1 U12100 ( .A1(n12100), .A2(n12184), .ZN(n12182) );
  OR2_X1 U12101 ( .A1(n12103), .A2(n12102), .ZN(n12184) );
  OR2_X1 U12102 ( .A1(n12185), .A2(n12186), .ZN(n12102) );
  AND2_X1 U12103 ( .A1(n12099), .A2(n12098), .ZN(n12186) );
  AND2_X1 U12104 ( .A1(n12096), .A2(n12187), .ZN(n12185) );
  OR2_X1 U12105 ( .A1(n12099), .A2(n12098), .ZN(n12187) );
  OR2_X1 U12106 ( .A1(n12188), .A2(n12189), .ZN(n12098) );
  AND2_X1 U12107 ( .A1(n12095), .A2(n12094), .ZN(n12189) );
  AND2_X1 U12108 ( .A1(n12092), .A2(n12190), .ZN(n12188) );
  OR2_X1 U12109 ( .A1(n12095), .A2(n12094), .ZN(n12190) );
  OR2_X1 U12110 ( .A1(n12191), .A2(n12192), .ZN(n12094) );
  AND2_X1 U12111 ( .A1(n12091), .A2(n12090), .ZN(n12192) );
  AND2_X1 U12112 ( .A1(n12088), .A2(n12193), .ZN(n12191) );
  OR2_X1 U12113 ( .A1(n12091), .A2(n12090), .ZN(n12193) );
  OR2_X1 U12114 ( .A1(n12194), .A2(n12195), .ZN(n12090) );
  AND2_X1 U12115 ( .A1(n12087), .A2(n12086), .ZN(n12195) );
  AND2_X1 U12116 ( .A1(n12084), .A2(n12196), .ZN(n12194) );
  OR2_X1 U12117 ( .A1(n12087), .A2(n12086), .ZN(n12196) );
  OR2_X1 U12118 ( .A1(n12197), .A2(n12198), .ZN(n12086) );
  AND2_X1 U12119 ( .A1(n12083), .A2(n12082), .ZN(n12198) );
  AND2_X1 U12120 ( .A1(n12080), .A2(n12199), .ZN(n12197) );
  OR2_X1 U12121 ( .A1(n12083), .A2(n12082), .ZN(n12199) );
  OR2_X1 U12122 ( .A1(n12200), .A2(n12201), .ZN(n12082) );
  AND2_X1 U12123 ( .A1(n8188), .A2(n12079), .ZN(n12201) );
  AND2_X1 U12124 ( .A1(n12077), .A2(n12202), .ZN(n12200) );
  OR2_X1 U12125 ( .A1(n8188), .A2(n12079), .ZN(n12202) );
  OR2_X1 U12126 ( .A1(n12203), .A2(n12204), .ZN(n12079) );
  AND2_X1 U12127 ( .A1(n12076), .A2(n12075), .ZN(n12204) );
  AND2_X1 U12128 ( .A1(n12073), .A2(n12205), .ZN(n12203) );
  OR2_X1 U12129 ( .A1(n12076), .A2(n12075), .ZN(n12205) );
  OR2_X1 U12130 ( .A1(n12206), .A2(n12207), .ZN(n12075) );
  AND2_X1 U12131 ( .A1(n12072), .A2(n12071), .ZN(n12207) );
  AND2_X1 U12132 ( .A1(n12069), .A2(n12208), .ZN(n12206) );
  OR2_X1 U12133 ( .A1(n12072), .A2(n12071), .ZN(n12208) );
  OR2_X1 U12134 ( .A1(n12209), .A2(n12210), .ZN(n12071) );
  AND2_X1 U12135 ( .A1(n12068), .A2(n12067), .ZN(n12210) );
  AND2_X1 U12136 ( .A1(n12065), .A2(n12211), .ZN(n12209) );
  OR2_X1 U12137 ( .A1(n12068), .A2(n12067), .ZN(n12211) );
  OR2_X1 U12138 ( .A1(n12212), .A2(n12213), .ZN(n12067) );
  AND2_X1 U12139 ( .A1(n12064), .A2(n12063), .ZN(n12213) );
  AND2_X1 U12140 ( .A1(n12061), .A2(n12214), .ZN(n12212) );
  OR2_X1 U12141 ( .A1(n12064), .A2(n12063), .ZN(n12214) );
  OR2_X1 U12142 ( .A1(n12215), .A2(n12216), .ZN(n12063) );
  AND2_X1 U12143 ( .A1(n12060), .A2(n12059), .ZN(n12216) );
  AND2_X1 U12144 ( .A1(n12057), .A2(n12217), .ZN(n12215) );
  OR2_X1 U12145 ( .A1(n12060), .A2(n12059), .ZN(n12217) );
  OR2_X1 U12146 ( .A1(n12218), .A2(n12219), .ZN(n12059) );
  AND2_X1 U12147 ( .A1(n12056), .A2(n12055), .ZN(n12219) );
  AND2_X1 U12148 ( .A1(n12053), .A2(n12220), .ZN(n12218) );
  OR2_X1 U12149 ( .A1(n12056), .A2(n12055), .ZN(n12220) );
  OR2_X1 U12150 ( .A1(n12221), .A2(n12222), .ZN(n12055) );
  AND2_X1 U12151 ( .A1(n12052), .A2(n12051), .ZN(n12222) );
  AND2_X1 U12152 ( .A1(n12049), .A2(n12223), .ZN(n12221) );
  OR2_X1 U12153 ( .A1(n12052), .A2(n12051), .ZN(n12223) );
  OR2_X1 U12154 ( .A1(n12224), .A2(n12225), .ZN(n12051) );
  AND2_X1 U12155 ( .A1(n12048), .A2(n12047), .ZN(n12225) );
  AND2_X1 U12156 ( .A1(n12045), .A2(n12226), .ZN(n12224) );
  OR2_X1 U12157 ( .A1(n12048), .A2(n12047), .ZN(n12226) );
  OR2_X1 U12158 ( .A1(n12227), .A2(n12228), .ZN(n12047) );
  AND2_X1 U12159 ( .A1(n12041), .A2(n12044), .ZN(n12228) );
  AND2_X1 U12160 ( .A1(n12229), .A2(n12230), .ZN(n12227) );
  OR2_X1 U12161 ( .A1(n12041), .A2(n12044), .ZN(n12230) );
  OR3_X1 U12162 ( .A1(n8807), .A2(n8803), .A3(n9796), .ZN(n12044) );
  OR2_X1 U12163 ( .A1(n7954), .A2(n8807), .ZN(n12041) );
  INV_X1 U12164 ( .A(n12043), .ZN(n12229) );
  OR2_X1 U12165 ( .A1(n12231), .A2(n12232), .ZN(n12043) );
  AND2_X1 U12166 ( .A1(b_19_), .A2(n12233), .ZN(n12232) );
  OR2_X1 U12167 ( .A1(n12234), .A2(n9801), .ZN(n12233) );
  AND2_X1 U12168 ( .A1(a_30_), .A2(n8799), .ZN(n12234) );
  AND2_X1 U12169 ( .A1(b_18_), .A2(n12235), .ZN(n12231) );
  OR2_X1 U12170 ( .A1(n12236), .A2(n7920), .ZN(n12235) );
  AND2_X1 U12171 ( .A1(a_31_), .A2(n8803), .ZN(n12236) );
  OR2_X1 U12172 ( .A1(n7979), .A2(n8807), .ZN(n12048) );
  XNOR2_X1 U12173 ( .A(n12237), .B(n12238), .ZN(n12045) );
  XOR2_X1 U12174 ( .A(n12239), .B(n12240), .Z(n12238) );
  OR2_X1 U12175 ( .A1(n8015), .A2(n8807), .ZN(n12052) );
  XOR2_X1 U12176 ( .A(n12241), .B(n12242), .Z(n12049) );
  XOR2_X1 U12177 ( .A(n12243), .B(n12244), .Z(n12242) );
  OR2_X1 U12178 ( .A1(n8040), .A2(n8807), .ZN(n12056) );
  XOR2_X1 U12179 ( .A(n12245), .B(n12246), .Z(n12053) );
  XOR2_X1 U12180 ( .A(n12247), .B(n12248), .Z(n12246) );
  OR2_X1 U12181 ( .A1(n8065), .A2(n8807), .ZN(n12060) );
  XOR2_X1 U12182 ( .A(n12249), .B(n12250), .Z(n12057) );
  XOR2_X1 U12183 ( .A(n12251), .B(n12252), .Z(n12250) );
  OR2_X1 U12184 ( .A1(n8090), .A2(n8807), .ZN(n12064) );
  XOR2_X1 U12185 ( .A(n12253), .B(n12254), .Z(n12061) );
  XOR2_X1 U12186 ( .A(n12255), .B(n12256), .Z(n12254) );
  OR2_X1 U12187 ( .A1(n8115), .A2(n8807), .ZN(n12068) );
  XOR2_X1 U12188 ( .A(n12257), .B(n12258), .Z(n12065) );
  XOR2_X1 U12189 ( .A(n12259), .B(n12260), .Z(n12258) );
  OR2_X1 U12190 ( .A1(n8140), .A2(n8807), .ZN(n12072) );
  XOR2_X1 U12191 ( .A(n12261), .B(n12262), .Z(n12069) );
  XOR2_X1 U12192 ( .A(n12263), .B(n12264), .Z(n12262) );
  OR2_X1 U12193 ( .A1(n8810), .A2(n8807), .ZN(n12076) );
  XOR2_X1 U12194 ( .A(n12265), .B(n12266), .Z(n12073) );
  XOR2_X1 U12195 ( .A(n12267), .B(n12268), .Z(n12266) );
  OR2_X1 U12196 ( .A1(n8806), .A2(n8807), .ZN(n8188) );
  XOR2_X1 U12197 ( .A(n12269), .B(n12270), .Z(n12077) );
  XOR2_X1 U12198 ( .A(n12271), .B(n12272), .Z(n12270) );
  OR2_X1 U12199 ( .A1(n8802), .A2(n8807), .ZN(n12083) );
  XOR2_X1 U12200 ( .A(n12273), .B(n12274), .Z(n12080) );
  XOR2_X1 U12201 ( .A(n12275), .B(n12276), .Z(n12274) );
  OR2_X1 U12202 ( .A1(n8798), .A2(n8807), .ZN(n12087) );
  XOR2_X1 U12203 ( .A(n12277), .B(n12278), .Z(n12084) );
  XOR2_X1 U12204 ( .A(n12279), .B(n8214), .Z(n12278) );
  OR2_X1 U12205 ( .A1(n8794), .A2(n8807), .ZN(n12091) );
  XOR2_X1 U12206 ( .A(n12280), .B(n12281), .Z(n12088) );
  XOR2_X1 U12207 ( .A(n12282), .B(n12283), .Z(n12281) );
  OR2_X1 U12208 ( .A1(n8790), .A2(n8807), .ZN(n12095) );
  XOR2_X1 U12209 ( .A(n12284), .B(n12285), .Z(n12092) );
  XOR2_X1 U12210 ( .A(n12286), .B(n12287), .Z(n12285) );
  OR2_X1 U12211 ( .A1(n8786), .A2(n8807), .ZN(n12099) );
  XOR2_X1 U12212 ( .A(n12288), .B(n12289), .Z(n12096) );
  XOR2_X1 U12213 ( .A(n12290), .B(n12291), .Z(n12289) );
  OR2_X1 U12214 ( .A1(n8782), .A2(n8807), .ZN(n12103) );
  XOR2_X1 U12215 ( .A(n12292), .B(n12293), .Z(n12100) );
  XOR2_X1 U12216 ( .A(n12294), .B(n12295), .Z(n12293) );
  OR2_X1 U12217 ( .A1(n8778), .A2(n8807), .ZN(n12107) );
  XOR2_X1 U12218 ( .A(n12296), .B(n12297), .Z(n12104) );
  XOR2_X1 U12219 ( .A(n12298), .B(n12299), .Z(n12297) );
  OR2_X1 U12220 ( .A1(n8774), .A2(n8807), .ZN(n12111) );
  XOR2_X1 U12221 ( .A(n12300), .B(n12301), .Z(n12108) );
  XOR2_X1 U12222 ( .A(n12302), .B(n12303), .Z(n12301) );
  OR2_X1 U12223 ( .A1(n8770), .A2(n8807), .ZN(n12115) );
  XOR2_X1 U12224 ( .A(n12304), .B(n12305), .Z(n12112) );
  XOR2_X1 U12225 ( .A(n12306), .B(n12307), .Z(n12305) );
  OR2_X1 U12226 ( .A1(n8766), .A2(n8807), .ZN(n12119) );
  XOR2_X1 U12227 ( .A(n12308), .B(n12309), .Z(n12116) );
  XOR2_X1 U12228 ( .A(n12310), .B(n12311), .Z(n12309) );
  OR2_X1 U12229 ( .A1(n8762), .A2(n8807), .ZN(n12123) );
  XOR2_X1 U12230 ( .A(n12312), .B(n12313), .Z(n12120) );
  XOR2_X1 U12231 ( .A(n12314), .B(n12315), .Z(n12313) );
  OR2_X1 U12232 ( .A1(n8758), .A2(n8807), .ZN(n12127) );
  XOR2_X1 U12233 ( .A(n12316), .B(n12317), .Z(n12124) );
  XOR2_X1 U12234 ( .A(n12318), .B(n12319), .Z(n12317) );
  OR2_X1 U12235 ( .A1(n8754), .A2(n8807), .ZN(n12131) );
  XOR2_X1 U12236 ( .A(n12320), .B(n12321), .Z(n12128) );
  XOR2_X1 U12237 ( .A(n12322), .B(n12323), .Z(n12321) );
  OR2_X1 U12238 ( .A1(n8750), .A2(n8807), .ZN(n12135) );
  XOR2_X1 U12239 ( .A(n12324), .B(n12325), .Z(n12132) );
  XOR2_X1 U12240 ( .A(n12326), .B(n12327), .Z(n12325) );
  OR2_X1 U12241 ( .A1(n8746), .A2(n8807), .ZN(n12139) );
  XOR2_X1 U12242 ( .A(n12328), .B(n12329), .Z(n12136) );
  XOR2_X1 U12243 ( .A(n12330), .B(n12331), .Z(n12329) );
  OR2_X1 U12244 ( .A1(n8742), .A2(n8807), .ZN(n12143) );
  XOR2_X1 U12245 ( .A(n12332), .B(n12333), .Z(n12140) );
  XOR2_X1 U12246 ( .A(n12334), .B(n12335), .Z(n12333) );
  OR2_X1 U12247 ( .A1(n8738), .A2(n8807), .ZN(n12147) );
  XOR2_X1 U12248 ( .A(n12336), .B(n12337), .Z(n12144) );
  XOR2_X1 U12249 ( .A(n12338), .B(n12339), .Z(n12337) );
  XOR2_X1 U12250 ( .A(n11707), .B(n12340), .Z(n11700) );
  XOR2_X1 U12251 ( .A(n11706), .B(n11705), .Z(n12340) );
  OR2_X1 U12252 ( .A1(n8738), .A2(n8803), .ZN(n11705) );
  OR2_X1 U12253 ( .A1(n12341), .A2(n12342), .ZN(n11706) );
  AND2_X1 U12254 ( .A1(n12339), .A2(n12338), .ZN(n12342) );
  AND2_X1 U12255 ( .A1(n12336), .A2(n12343), .ZN(n12341) );
  OR2_X1 U12256 ( .A1(n12339), .A2(n12338), .ZN(n12343) );
  OR2_X1 U12257 ( .A1(n12344), .A2(n12345), .ZN(n12338) );
  AND2_X1 U12258 ( .A1(n12335), .A2(n12334), .ZN(n12345) );
  AND2_X1 U12259 ( .A1(n12332), .A2(n12346), .ZN(n12344) );
  OR2_X1 U12260 ( .A1(n12335), .A2(n12334), .ZN(n12346) );
  OR2_X1 U12261 ( .A1(n12347), .A2(n12348), .ZN(n12334) );
  AND2_X1 U12262 ( .A1(n12331), .A2(n12330), .ZN(n12348) );
  AND2_X1 U12263 ( .A1(n12328), .A2(n12349), .ZN(n12347) );
  OR2_X1 U12264 ( .A1(n12331), .A2(n12330), .ZN(n12349) );
  OR2_X1 U12265 ( .A1(n12350), .A2(n12351), .ZN(n12330) );
  AND2_X1 U12266 ( .A1(n12327), .A2(n12326), .ZN(n12351) );
  AND2_X1 U12267 ( .A1(n12324), .A2(n12352), .ZN(n12350) );
  OR2_X1 U12268 ( .A1(n12327), .A2(n12326), .ZN(n12352) );
  OR2_X1 U12269 ( .A1(n12353), .A2(n12354), .ZN(n12326) );
  AND2_X1 U12270 ( .A1(n12323), .A2(n12322), .ZN(n12354) );
  AND2_X1 U12271 ( .A1(n12320), .A2(n12355), .ZN(n12353) );
  OR2_X1 U12272 ( .A1(n12323), .A2(n12322), .ZN(n12355) );
  OR2_X1 U12273 ( .A1(n12356), .A2(n12357), .ZN(n12322) );
  AND2_X1 U12274 ( .A1(n12319), .A2(n12318), .ZN(n12357) );
  AND2_X1 U12275 ( .A1(n12316), .A2(n12358), .ZN(n12356) );
  OR2_X1 U12276 ( .A1(n12319), .A2(n12318), .ZN(n12358) );
  OR2_X1 U12277 ( .A1(n12359), .A2(n12360), .ZN(n12318) );
  AND2_X1 U12278 ( .A1(n12315), .A2(n12314), .ZN(n12360) );
  AND2_X1 U12279 ( .A1(n12312), .A2(n12361), .ZN(n12359) );
  OR2_X1 U12280 ( .A1(n12315), .A2(n12314), .ZN(n12361) );
  OR2_X1 U12281 ( .A1(n12362), .A2(n12363), .ZN(n12314) );
  AND2_X1 U12282 ( .A1(n12311), .A2(n12310), .ZN(n12363) );
  AND2_X1 U12283 ( .A1(n12308), .A2(n12364), .ZN(n12362) );
  OR2_X1 U12284 ( .A1(n12311), .A2(n12310), .ZN(n12364) );
  OR2_X1 U12285 ( .A1(n12365), .A2(n12366), .ZN(n12310) );
  AND2_X1 U12286 ( .A1(n12307), .A2(n12306), .ZN(n12366) );
  AND2_X1 U12287 ( .A1(n12304), .A2(n12367), .ZN(n12365) );
  OR2_X1 U12288 ( .A1(n12307), .A2(n12306), .ZN(n12367) );
  OR2_X1 U12289 ( .A1(n12368), .A2(n12369), .ZN(n12306) );
  AND2_X1 U12290 ( .A1(n12303), .A2(n12302), .ZN(n12369) );
  AND2_X1 U12291 ( .A1(n12300), .A2(n12370), .ZN(n12368) );
  OR2_X1 U12292 ( .A1(n12303), .A2(n12302), .ZN(n12370) );
  OR2_X1 U12293 ( .A1(n12371), .A2(n12372), .ZN(n12302) );
  AND2_X1 U12294 ( .A1(n12299), .A2(n12298), .ZN(n12372) );
  AND2_X1 U12295 ( .A1(n12296), .A2(n12373), .ZN(n12371) );
  OR2_X1 U12296 ( .A1(n12299), .A2(n12298), .ZN(n12373) );
  OR2_X1 U12297 ( .A1(n12374), .A2(n12375), .ZN(n12298) );
  AND2_X1 U12298 ( .A1(n12295), .A2(n12294), .ZN(n12375) );
  AND2_X1 U12299 ( .A1(n12292), .A2(n12376), .ZN(n12374) );
  OR2_X1 U12300 ( .A1(n12295), .A2(n12294), .ZN(n12376) );
  OR2_X1 U12301 ( .A1(n12377), .A2(n12378), .ZN(n12294) );
  AND2_X1 U12302 ( .A1(n12291), .A2(n12290), .ZN(n12378) );
  AND2_X1 U12303 ( .A1(n12288), .A2(n12379), .ZN(n12377) );
  OR2_X1 U12304 ( .A1(n12291), .A2(n12290), .ZN(n12379) );
  OR2_X1 U12305 ( .A1(n12380), .A2(n12381), .ZN(n12290) );
  AND2_X1 U12306 ( .A1(n12287), .A2(n12286), .ZN(n12381) );
  AND2_X1 U12307 ( .A1(n12284), .A2(n12382), .ZN(n12380) );
  OR2_X1 U12308 ( .A1(n12287), .A2(n12286), .ZN(n12382) );
  OR2_X1 U12309 ( .A1(n12383), .A2(n12384), .ZN(n12286) );
  AND2_X1 U12310 ( .A1(n12283), .A2(n12282), .ZN(n12384) );
  AND2_X1 U12311 ( .A1(n12280), .A2(n12385), .ZN(n12383) );
  OR2_X1 U12312 ( .A1(n12283), .A2(n12282), .ZN(n12385) );
  OR2_X1 U12313 ( .A1(n12386), .A2(n12387), .ZN(n12282) );
  AND2_X1 U12314 ( .A1(n8214), .A2(n12279), .ZN(n12387) );
  AND2_X1 U12315 ( .A1(n12277), .A2(n12388), .ZN(n12386) );
  OR2_X1 U12316 ( .A1(n8214), .A2(n12279), .ZN(n12388) );
  OR2_X1 U12317 ( .A1(n12389), .A2(n12390), .ZN(n12279) );
  AND2_X1 U12318 ( .A1(n12276), .A2(n12275), .ZN(n12390) );
  AND2_X1 U12319 ( .A1(n12273), .A2(n12391), .ZN(n12389) );
  OR2_X1 U12320 ( .A1(n12276), .A2(n12275), .ZN(n12391) );
  OR2_X1 U12321 ( .A1(n12392), .A2(n12393), .ZN(n12275) );
  AND2_X1 U12322 ( .A1(n12272), .A2(n12271), .ZN(n12393) );
  AND2_X1 U12323 ( .A1(n12269), .A2(n12394), .ZN(n12392) );
  OR2_X1 U12324 ( .A1(n12272), .A2(n12271), .ZN(n12394) );
  OR2_X1 U12325 ( .A1(n12395), .A2(n12396), .ZN(n12271) );
  AND2_X1 U12326 ( .A1(n12268), .A2(n12267), .ZN(n12396) );
  AND2_X1 U12327 ( .A1(n12265), .A2(n12397), .ZN(n12395) );
  OR2_X1 U12328 ( .A1(n12268), .A2(n12267), .ZN(n12397) );
  OR2_X1 U12329 ( .A1(n12398), .A2(n12399), .ZN(n12267) );
  AND2_X1 U12330 ( .A1(n12264), .A2(n12263), .ZN(n12399) );
  AND2_X1 U12331 ( .A1(n12261), .A2(n12400), .ZN(n12398) );
  OR2_X1 U12332 ( .A1(n12264), .A2(n12263), .ZN(n12400) );
  OR2_X1 U12333 ( .A1(n12401), .A2(n12402), .ZN(n12263) );
  AND2_X1 U12334 ( .A1(n12260), .A2(n12259), .ZN(n12402) );
  AND2_X1 U12335 ( .A1(n12257), .A2(n12403), .ZN(n12401) );
  OR2_X1 U12336 ( .A1(n12260), .A2(n12259), .ZN(n12403) );
  OR2_X1 U12337 ( .A1(n12404), .A2(n12405), .ZN(n12259) );
  AND2_X1 U12338 ( .A1(n12256), .A2(n12255), .ZN(n12405) );
  AND2_X1 U12339 ( .A1(n12253), .A2(n12406), .ZN(n12404) );
  OR2_X1 U12340 ( .A1(n12256), .A2(n12255), .ZN(n12406) );
  OR2_X1 U12341 ( .A1(n12407), .A2(n12408), .ZN(n12255) );
  AND2_X1 U12342 ( .A1(n12252), .A2(n12251), .ZN(n12408) );
  AND2_X1 U12343 ( .A1(n12249), .A2(n12409), .ZN(n12407) );
  OR2_X1 U12344 ( .A1(n12252), .A2(n12251), .ZN(n12409) );
  OR2_X1 U12345 ( .A1(n12410), .A2(n12411), .ZN(n12251) );
  AND2_X1 U12346 ( .A1(n12248), .A2(n12247), .ZN(n12411) );
  AND2_X1 U12347 ( .A1(n12245), .A2(n12412), .ZN(n12410) );
  OR2_X1 U12348 ( .A1(n12248), .A2(n12247), .ZN(n12412) );
  OR2_X1 U12349 ( .A1(n12413), .A2(n12414), .ZN(n12247) );
  AND2_X1 U12350 ( .A1(n12244), .A2(n12243), .ZN(n12414) );
  AND2_X1 U12351 ( .A1(n12241), .A2(n12415), .ZN(n12413) );
  OR2_X1 U12352 ( .A1(n12244), .A2(n12243), .ZN(n12415) );
  OR2_X1 U12353 ( .A1(n12416), .A2(n12417), .ZN(n12243) );
  AND2_X1 U12354 ( .A1(n12237), .A2(n12240), .ZN(n12417) );
  AND2_X1 U12355 ( .A1(n12418), .A2(n12419), .ZN(n12416) );
  OR2_X1 U12356 ( .A1(n12237), .A2(n12240), .ZN(n12419) );
  OR3_X1 U12357 ( .A1(n8803), .A2(n8799), .A3(n9796), .ZN(n12240) );
  OR2_X1 U12358 ( .A1(n7954), .A2(n8803), .ZN(n12237) );
  INV_X1 U12359 ( .A(n12239), .ZN(n12418) );
  OR2_X1 U12360 ( .A1(n12420), .A2(n12421), .ZN(n12239) );
  AND2_X1 U12361 ( .A1(b_18_), .A2(n12422), .ZN(n12421) );
  OR2_X1 U12362 ( .A1(n12423), .A2(n9801), .ZN(n12422) );
  AND2_X1 U12363 ( .A1(a_30_), .A2(n8795), .ZN(n12423) );
  AND2_X1 U12364 ( .A1(b_17_), .A2(n12424), .ZN(n12420) );
  OR2_X1 U12365 ( .A1(n12425), .A2(n7920), .ZN(n12424) );
  AND2_X1 U12366 ( .A1(a_31_), .A2(n8799), .ZN(n12425) );
  OR2_X1 U12367 ( .A1(n7979), .A2(n8803), .ZN(n12244) );
  XNOR2_X1 U12368 ( .A(n12426), .B(n12427), .ZN(n12241) );
  XOR2_X1 U12369 ( .A(n12428), .B(n12429), .Z(n12427) );
  OR2_X1 U12370 ( .A1(n8015), .A2(n8803), .ZN(n12248) );
  XOR2_X1 U12371 ( .A(n12430), .B(n12431), .Z(n12245) );
  XOR2_X1 U12372 ( .A(n12432), .B(n12433), .Z(n12431) );
  OR2_X1 U12373 ( .A1(n8040), .A2(n8803), .ZN(n12252) );
  XOR2_X1 U12374 ( .A(n12434), .B(n12435), .Z(n12249) );
  XOR2_X1 U12375 ( .A(n12436), .B(n12437), .Z(n12435) );
  OR2_X1 U12376 ( .A1(n8065), .A2(n8803), .ZN(n12256) );
  XOR2_X1 U12377 ( .A(n12438), .B(n12439), .Z(n12253) );
  XOR2_X1 U12378 ( .A(n12440), .B(n12441), .Z(n12439) );
  OR2_X1 U12379 ( .A1(n8090), .A2(n8803), .ZN(n12260) );
  XOR2_X1 U12380 ( .A(n12442), .B(n12443), .Z(n12257) );
  XOR2_X1 U12381 ( .A(n12444), .B(n12445), .Z(n12443) );
  OR2_X1 U12382 ( .A1(n8115), .A2(n8803), .ZN(n12264) );
  XOR2_X1 U12383 ( .A(n12446), .B(n12447), .Z(n12261) );
  XOR2_X1 U12384 ( .A(n12448), .B(n12449), .Z(n12447) );
  OR2_X1 U12385 ( .A1(n8140), .A2(n8803), .ZN(n12268) );
  XOR2_X1 U12386 ( .A(n12450), .B(n12451), .Z(n12265) );
  XOR2_X1 U12387 ( .A(n12452), .B(n12453), .Z(n12451) );
  OR2_X1 U12388 ( .A1(n8810), .A2(n8803), .ZN(n12272) );
  XOR2_X1 U12389 ( .A(n12454), .B(n12455), .Z(n12269) );
  XOR2_X1 U12390 ( .A(n12456), .B(n12457), .Z(n12455) );
  OR2_X1 U12391 ( .A1(n8806), .A2(n8803), .ZN(n12276) );
  XOR2_X1 U12392 ( .A(n12458), .B(n12459), .Z(n12273) );
  XOR2_X1 U12393 ( .A(n12460), .B(n12461), .Z(n12459) );
  OR2_X1 U12394 ( .A1(n8802), .A2(n8803), .ZN(n8214) );
  XOR2_X1 U12395 ( .A(n12462), .B(n12463), .Z(n12277) );
  XOR2_X1 U12396 ( .A(n12464), .B(n12465), .Z(n12463) );
  OR2_X1 U12397 ( .A1(n8798), .A2(n8803), .ZN(n12283) );
  XOR2_X1 U12398 ( .A(n12466), .B(n12467), .Z(n12280) );
  XOR2_X1 U12399 ( .A(n12468), .B(n12469), .Z(n12467) );
  OR2_X1 U12400 ( .A1(n8794), .A2(n8803), .ZN(n12287) );
  XOR2_X1 U12401 ( .A(n12470), .B(n12471), .Z(n12284) );
  XOR2_X1 U12402 ( .A(n12472), .B(n8240), .Z(n12471) );
  OR2_X1 U12403 ( .A1(n8790), .A2(n8803), .ZN(n12291) );
  XOR2_X1 U12404 ( .A(n12473), .B(n12474), .Z(n12288) );
  XOR2_X1 U12405 ( .A(n12475), .B(n12476), .Z(n12474) );
  OR2_X1 U12406 ( .A1(n8786), .A2(n8803), .ZN(n12295) );
  XOR2_X1 U12407 ( .A(n12477), .B(n12478), .Z(n12292) );
  XOR2_X1 U12408 ( .A(n12479), .B(n12480), .Z(n12478) );
  OR2_X1 U12409 ( .A1(n8782), .A2(n8803), .ZN(n12299) );
  XOR2_X1 U12410 ( .A(n12481), .B(n12482), .Z(n12296) );
  XOR2_X1 U12411 ( .A(n12483), .B(n12484), .Z(n12482) );
  OR2_X1 U12412 ( .A1(n8778), .A2(n8803), .ZN(n12303) );
  XOR2_X1 U12413 ( .A(n12485), .B(n12486), .Z(n12300) );
  XOR2_X1 U12414 ( .A(n12487), .B(n12488), .Z(n12486) );
  OR2_X1 U12415 ( .A1(n8774), .A2(n8803), .ZN(n12307) );
  XOR2_X1 U12416 ( .A(n12489), .B(n12490), .Z(n12304) );
  XOR2_X1 U12417 ( .A(n12491), .B(n12492), .Z(n12490) );
  OR2_X1 U12418 ( .A1(n8770), .A2(n8803), .ZN(n12311) );
  XOR2_X1 U12419 ( .A(n12493), .B(n12494), .Z(n12308) );
  XOR2_X1 U12420 ( .A(n12495), .B(n12496), .Z(n12494) );
  OR2_X1 U12421 ( .A1(n8766), .A2(n8803), .ZN(n12315) );
  XOR2_X1 U12422 ( .A(n12497), .B(n12498), .Z(n12312) );
  XOR2_X1 U12423 ( .A(n12499), .B(n12500), .Z(n12498) );
  OR2_X1 U12424 ( .A1(n8762), .A2(n8803), .ZN(n12319) );
  XOR2_X1 U12425 ( .A(n12501), .B(n12502), .Z(n12316) );
  XOR2_X1 U12426 ( .A(n12503), .B(n12504), .Z(n12502) );
  OR2_X1 U12427 ( .A1(n8758), .A2(n8803), .ZN(n12323) );
  XOR2_X1 U12428 ( .A(n12505), .B(n12506), .Z(n12320) );
  XOR2_X1 U12429 ( .A(n12507), .B(n12508), .Z(n12506) );
  OR2_X1 U12430 ( .A1(n8754), .A2(n8803), .ZN(n12327) );
  XOR2_X1 U12431 ( .A(n12509), .B(n12510), .Z(n12324) );
  XOR2_X1 U12432 ( .A(n12511), .B(n12512), .Z(n12510) );
  OR2_X1 U12433 ( .A1(n8750), .A2(n8803), .ZN(n12331) );
  XOR2_X1 U12434 ( .A(n12513), .B(n12514), .Z(n12328) );
  XOR2_X1 U12435 ( .A(n12515), .B(n12516), .Z(n12514) );
  OR2_X1 U12436 ( .A1(n8746), .A2(n8803), .ZN(n12335) );
  XOR2_X1 U12437 ( .A(n12517), .B(n12518), .Z(n12332) );
  XOR2_X1 U12438 ( .A(n12519), .B(n12520), .Z(n12518) );
  OR2_X1 U12439 ( .A1(n8742), .A2(n8803), .ZN(n12339) );
  XOR2_X1 U12440 ( .A(n12521), .B(n12522), .Z(n12336) );
  XOR2_X1 U12441 ( .A(n12523), .B(n12524), .Z(n12522) );
  XOR2_X1 U12442 ( .A(n11714), .B(n12525), .Z(n11707) );
  XOR2_X1 U12443 ( .A(n11713), .B(n11712), .Z(n12525) );
  OR2_X1 U12444 ( .A1(n8742), .A2(n8799), .ZN(n11712) );
  OR2_X1 U12445 ( .A1(n12526), .A2(n12527), .ZN(n11713) );
  AND2_X1 U12446 ( .A1(n12524), .A2(n12523), .ZN(n12527) );
  AND2_X1 U12447 ( .A1(n12521), .A2(n12528), .ZN(n12526) );
  OR2_X1 U12448 ( .A1(n12524), .A2(n12523), .ZN(n12528) );
  OR2_X1 U12449 ( .A1(n12529), .A2(n12530), .ZN(n12523) );
  AND2_X1 U12450 ( .A1(n12520), .A2(n12519), .ZN(n12530) );
  AND2_X1 U12451 ( .A1(n12517), .A2(n12531), .ZN(n12529) );
  OR2_X1 U12452 ( .A1(n12520), .A2(n12519), .ZN(n12531) );
  OR2_X1 U12453 ( .A1(n12532), .A2(n12533), .ZN(n12519) );
  AND2_X1 U12454 ( .A1(n12516), .A2(n12515), .ZN(n12533) );
  AND2_X1 U12455 ( .A1(n12513), .A2(n12534), .ZN(n12532) );
  OR2_X1 U12456 ( .A1(n12516), .A2(n12515), .ZN(n12534) );
  OR2_X1 U12457 ( .A1(n12535), .A2(n12536), .ZN(n12515) );
  AND2_X1 U12458 ( .A1(n12512), .A2(n12511), .ZN(n12536) );
  AND2_X1 U12459 ( .A1(n12509), .A2(n12537), .ZN(n12535) );
  OR2_X1 U12460 ( .A1(n12512), .A2(n12511), .ZN(n12537) );
  OR2_X1 U12461 ( .A1(n12538), .A2(n12539), .ZN(n12511) );
  AND2_X1 U12462 ( .A1(n12508), .A2(n12507), .ZN(n12539) );
  AND2_X1 U12463 ( .A1(n12505), .A2(n12540), .ZN(n12538) );
  OR2_X1 U12464 ( .A1(n12508), .A2(n12507), .ZN(n12540) );
  OR2_X1 U12465 ( .A1(n12541), .A2(n12542), .ZN(n12507) );
  AND2_X1 U12466 ( .A1(n12504), .A2(n12503), .ZN(n12542) );
  AND2_X1 U12467 ( .A1(n12501), .A2(n12543), .ZN(n12541) );
  OR2_X1 U12468 ( .A1(n12504), .A2(n12503), .ZN(n12543) );
  OR2_X1 U12469 ( .A1(n12544), .A2(n12545), .ZN(n12503) );
  AND2_X1 U12470 ( .A1(n12500), .A2(n12499), .ZN(n12545) );
  AND2_X1 U12471 ( .A1(n12497), .A2(n12546), .ZN(n12544) );
  OR2_X1 U12472 ( .A1(n12500), .A2(n12499), .ZN(n12546) );
  OR2_X1 U12473 ( .A1(n12547), .A2(n12548), .ZN(n12499) );
  AND2_X1 U12474 ( .A1(n12496), .A2(n12495), .ZN(n12548) );
  AND2_X1 U12475 ( .A1(n12493), .A2(n12549), .ZN(n12547) );
  OR2_X1 U12476 ( .A1(n12496), .A2(n12495), .ZN(n12549) );
  OR2_X1 U12477 ( .A1(n12550), .A2(n12551), .ZN(n12495) );
  AND2_X1 U12478 ( .A1(n12492), .A2(n12491), .ZN(n12551) );
  AND2_X1 U12479 ( .A1(n12489), .A2(n12552), .ZN(n12550) );
  OR2_X1 U12480 ( .A1(n12492), .A2(n12491), .ZN(n12552) );
  OR2_X1 U12481 ( .A1(n12553), .A2(n12554), .ZN(n12491) );
  AND2_X1 U12482 ( .A1(n12488), .A2(n12487), .ZN(n12554) );
  AND2_X1 U12483 ( .A1(n12485), .A2(n12555), .ZN(n12553) );
  OR2_X1 U12484 ( .A1(n12488), .A2(n12487), .ZN(n12555) );
  OR2_X1 U12485 ( .A1(n12556), .A2(n12557), .ZN(n12487) );
  AND2_X1 U12486 ( .A1(n12484), .A2(n12483), .ZN(n12557) );
  AND2_X1 U12487 ( .A1(n12481), .A2(n12558), .ZN(n12556) );
  OR2_X1 U12488 ( .A1(n12484), .A2(n12483), .ZN(n12558) );
  OR2_X1 U12489 ( .A1(n12559), .A2(n12560), .ZN(n12483) );
  AND2_X1 U12490 ( .A1(n12480), .A2(n12479), .ZN(n12560) );
  AND2_X1 U12491 ( .A1(n12477), .A2(n12561), .ZN(n12559) );
  OR2_X1 U12492 ( .A1(n12480), .A2(n12479), .ZN(n12561) );
  OR2_X1 U12493 ( .A1(n12562), .A2(n12563), .ZN(n12479) );
  AND2_X1 U12494 ( .A1(n12476), .A2(n12475), .ZN(n12563) );
  AND2_X1 U12495 ( .A1(n12473), .A2(n12564), .ZN(n12562) );
  OR2_X1 U12496 ( .A1(n12476), .A2(n12475), .ZN(n12564) );
  OR2_X1 U12497 ( .A1(n12565), .A2(n12566), .ZN(n12475) );
  AND2_X1 U12498 ( .A1(n8240), .A2(n12472), .ZN(n12566) );
  AND2_X1 U12499 ( .A1(n12470), .A2(n12567), .ZN(n12565) );
  OR2_X1 U12500 ( .A1(n8240), .A2(n12472), .ZN(n12567) );
  OR2_X1 U12501 ( .A1(n12568), .A2(n12569), .ZN(n12472) );
  AND2_X1 U12502 ( .A1(n12469), .A2(n12468), .ZN(n12569) );
  AND2_X1 U12503 ( .A1(n12466), .A2(n12570), .ZN(n12568) );
  OR2_X1 U12504 ( .A1(n12469), .A2(n12468), .ZN(n12570) );
  OR2_X1 U12505 ( .A1(n12571), .A2(n12572), .ZN(n12468) );
  AND2_X1 U12506 ( .A1(n12465), .A2(n12464), .ZN(n12572) );
  AND2_X1 U12507 ( .A1(n12462), .A2(n12573), .ZN(n12571) );
  OR2_X1 U12508 ( .A1(n12465), .A2(n12464), .ZN(n12573) );
  OR2_X1 U12509 ( .A1(n12574), .A2(n12575), .ZN(n12464) );
  AND2_X1 U12510 ( .A1(n12461), .A2(n12460), .ZN(n12575) );
  AND2_X1 U12511 ( .A1(n12458), .A2(n12576), .ZN(n12574) );
  OR2_X1 U12512 ( .A1(n12461), .A2(n12460), .ZN(n12576) );
  OR2_X1 U12513 ( .A1(n12577), .A2(n12578), .ZN(n12460) );
  AND2_X1 U12514 ( .A1(n12457), .A2(n12456), .ZN(n12578) );
  AND2_X1 U12515 ( .A1(n12454), .A2(n12579), .ZN(n12577) );
  OR2_X1 U12516 ( .A1(n12457), .A2(n12456), .ZN(n12579) );
  OR2_X1 U12517 ( .A1(n12580), .A2(n12581), .ZN(n12456) );
  AND2_X1 U12518 ( .A1(n12453), .A2(n12452), .ZN(n12581) );
  AND2_X1 U12519 ( .A1(n12450), .A2(n12582), .ZN(n12580) );
  OR2_X1 U12520 ( .A1(n12453), .A2(n12452), .ZN(n12582) );
  OR2_X1 U12521 ( .A1(n12583), .A2(n12584), .ZN(n12452) );
  AND2_X1 U12522 ( .A1(n12449), .A2(n12448), .ZN(n12584) );
  AND2_X1 U12523 ( .A1(n12446), .A2(n12585), .ZN(n12583) );
  OR2_X1 U12524 ( .A1(n12449), .A2(n12448), .ZN(n12585) );
  OR2_X1 U12525 ( .A1(n12586), .A2(n12587), .ZN(n12448) );
  AND2_X1 U12526 ( .A1(n12445), .A2(n12444), .ZN(n12587) );
  AND2_X1 U12527 ( .A1(n12442), .A2(n12588), .ZN(n12586) );
  OR2_X1 U12528 ( .A1(n12445), .A2(n12444), .ZN(n12588) );
  OR2_X1 U12529 ( .A1(n12589), .A2(n12590), .ZN(n12444) );
  AND2_X1 U12530 ( .A1(n12441), .A2(n12440), .ZN(n12590) );
  AND2_X1 U12531 ( .A1(n12438), .A2(n12591), .ZN(n12589) );
  OR2_X1 U12532 ( .A1(n12441), .A2(n12440), .ZN(n12591) );
  OR2_X1 U12533 ( .A1(n12592), .A2(n12593), .ZN(n12440) );
  AND2_X1 U12534 ( .A1(n12437), .A2(n12436), .ZN(n12593) );
  AND2_X1 U12535 ( .A1(n12434), .A2(n12594), .ZN(n12592) );
  OR2_X1 U12536 ( .A1(n12437), .A2(n12436), .ZN(n12594) );
  OR2_X1 U12537 ( .A1(n12595), .A2(n12596), .ZN(n12436) );
  AND2_X1 U12538 ( .A1(n12433), .A2(n12432), .ZN(n12596) );
  AND2_X1 U12539 ( .A1(n12430), .A2(n12597), .ZN(n12595) );
  OR2_X1 U12540 ( .A1(n12433), .A2(n12432), .ZN(n12597) );
  OR2_X1 U12541 ( .A1(n12598), .A2(n12599), .ZN(n12432) );
  AND2_X1 U12542 ( .A1(n12426), .A2(n12429), .ZN(n12599) );
  AND2_X1 U12543 ( .A1(n12600), .A2(n12601), .ZN(n12598) );
  OR2_X1 U12544 ( .A1(n12426), .A2(n12429), .ZN(n12601) );
  OR3_X1 U12545 ( .A1(n8799), .A2(n8795), .A3(n9796), .ZN(n12429) );
  OR2_X1 U12546 ( .A1(n7954), .A2(n8799), .ZN(n12426) );
  INV_X1 U12547 ( .A(n12428), .ZN(n12600) );
  OR2_X1 U12548 ( .A1(n12602), .A2(n12603), .ZN(n12428) );
  AND2_X1 U12549 ( .A1(b_17_), .A2(n12604), .ZN(n12603) );
  OR2_X1 U12550 ( .A1(n12605), .A2(n9801), .ZN(n12604) );
  AND2_X1 U12551 ( .A1(a_30_), .A2(n8791), .ZN(n12605) );
  AND2_X1 U12552 ( .A1(b_16_), .A2(n12606), .ZN(n12602) );
  OR2_X1 U12553 ( .A1(n12607), .A2(n7920), .ZN(n12606) );
  AND2_X1 U12554 ( .A1(a_31_), .A2(n8795), .ZN(n12607) );
  OR2_X1 U12555 ( .A1(n7979), .A2(n8799), .ZN(n12433) );
  XNOR2_X1 U12556 ( .A(n12608), .B(n12609), .ZN(n12430) );
  XOR2_X1 U12557 ( .A(n12610), .B(n12611), .Z(n12609) );
  OR2_X1 U12558 ( .A1(n8015), .A2(n8799), .ZN(n12437) );
  XOR2_X1 U12559 ( .A(n12612), .B(n12613), .Z(n12434) );
  XOR2_X1 U12560 ( .A(n12614), .B(n12615), .Z(n12613) );
  OR2_X1 U12561 ( .A1(n8040), .A2(n8799), .ZN(n12441) );
  XOR2_X1 U12562 ( .A(n12616), .B(n12617), .Z(n12438) );
  XOR2_X1 U12563 ( .A(n12618), .B(n12619), .Z(n12617) );
  OR2_X1 U12564 ( .A1(n8065), .A2(n8799), .ZN(n12445) );
  XOR2_X1 U12565 ( .A(n12620), .B(n12621), .Z(n12442) );
  XOR2_X1 U12566 ( .A(n12622), .B(n12623), .Z(n12621) );
  OR2_X1 U12567 ( .A1(n8090), .A2(n8799), .ZN(n12449) );
  XOR2_X1 U12568 ( .A(n12624), .B(n12625), .Z(n12446) );
  XOR2_X1 U12569 ( .A(n12626), .B(n12627), .Z(n12625) );
  OR2_X1 U12570 ( .A1(n8115), .A2(n8799), .ZN(n12453) );
  XOR2_X1 U12571 ( .A(n12628), .B(n12629), .Z(n12450) );
  XOR2_X1 U12572 ( .A(n12630), .B(n12631), .Z(n12629) );
  OR2_X1 U12573 ( .A1(n8140), .A2(n8799), .ZN(n12457) );
  XOR2_X1 U12574 ( .A(n12632), .B(n12633), .Z(n12454) );
  XOR2_X1 U12575 ( .A(n12634), .B(n12635), .Z(n12633) );
  OR2_X1 U12576 ( .A1(n8810), .A2(n8799), .ZN(n12461) );
  XOR2_X1 U12577 ( .A(n12636), .B(n12637), .Z(n12458) );
  XOR2_X1 U12578 ( .A(n12638), .B(n12639), .Z(n12637) );
  OR2_X1 U12579 ( .A1(n8806), .A2(n8799), .ZN(n12465) );
  XOR2_X1 U12580 ( .A(n12640), .B(n12641), .Z(n12462) );
  XOR2_X1 U12581 ( .A(n12642), .B(n12643), .Z(n12641) );
  OR2_X1 U12582 ( .A1(n8802), .A2(n8799), .ZN(n12469) );
  XOR2_X1 U12583 ( .A(n12644), .B(n12645), .Z(n12466) );
  XOR2_X1 U12584 ( .A(n12646), .B(n12647), .Z(n12645) );
  OR2_X1 U12585 ( .A1(n8798), .A2(n8799), .ZN(n8240) );
  XOR2_X1 U12586 ( .A(n12648), .B(n12649), .Z(n12470) );
  XOR2_X1 U12587 ( .A(n12650), .B(n12651), .Z(n12649) );
  OR2_X1 U12588 ( .A1(n8794), .A2(n8799), .ZN(n12476) );
  XOR2_X1 U12589 ( .A(n12652), .B(n12653), .Z(n12473) );
  XOR2_X1 U12590 ( .A(n12654), .B(n12655), .Z(n12653) );
  OR2_X1 U12591 ( .A1(n8790), .A2(n8799), .ZN(n12480) );
  XOR2_X1 U12592 ( .A(n12656), .B(n12657), .Z(n12477) );
  XOR2_X1 U12593 ( .A(n12658), .B(n8270), .Z(n12657) );
  OR2_X1 U12594 ( .A1(n8786), .A2(n8799), .ZN(n12484) );
  XOR2_X1 U12595 ( .A(n12659), .B(n12660), .Z(n12481) );
  XOR2_X1 U12596 ( .A(n12661), .B(n12662), .Z(n12660) );
  OR2_X1 U12597 ( .A1(n8782), .A2(n8799), .ZN(n12488) );
  XOR2_X1 U12598 ( .A(n12663), .B(n12664), .Z(n12485) );
  XOR2_X1 U12599 ( .A(n12665), .B(n12666), .Z(n12664) );
  OR2_X1 U12600 ( .A1(n8778), .A2(n8799), .ZN(n12492) );
  XOR2_X1 U12601 ( .A(n12667), .B(n12668), .Z(n12489) );
  XOR2_X1 U12602 ( .A(n12669), .B(n12670), .Z(n12668) );
  OR2_X1 U12603 ( .A1(n8774), .A2(n8799), .ZN(n12496) );
  XOR2_X1 U12604 ( .A(n12671), .B(n12672), .Z(n12493) );
  XOR2_X1 U12605 ( .A(n12673), .B(n12674), .Z(n12672) );
  OR2_X1 U12606 ( .A1(n8770), .A2(n8799), .ZN(n12500) );
  XOR2_X1 U12607 ( .A(n12675), .B(n12676), .Z(n12497) );
  XOR2_X1 U12608 ( .A(n12677), .B(n12678), .Z(n12676) );
  OR2_X1 U12609 ( .A1(n8766), .A2(n8799), .ZN(n12504) );
  XOR2_X1 U12610 ( .A(n12679), .B(n12680), .Z(n12501) );
  XOR2_X1 U12611 ( .A(n12681), .B(n12682), .Z(n12680) );
  OR2_X1 U12612 ( .A1(n8762), .A2(n8799), .ZN(n12508) );
  XOR2_X1 U12613 ( .A(n12683), .B(n12684), .Z(n12505) );
  XOR2_X1 U12614 ( .A(n12685), .B(n12686), .Z(n12684) );
  OR2_X1 U12615 ( .A1(n8758), .A2(n8799), .ZN(n12512) );
  XOR2_X1 U12616 ( .A(n12687), .B(n12688), .Z(n12509) );
  XOR2_X1 U12617 ( .A(n12689), .B(n12690), .Z(n12688) );
  OR2_X1 U12618 ( .A1(n8754), .A2(n8799), .ZN(n12516) );
  XOR2_X1 U12619 ( .A(n12691), .B(n12692), .Z(n12513) );
  XOR2_X1 U12620 ( .A(n12693), .B(n12694), .Z(n12692) );
  OR2_X1 U12621 ( .A1(n8750), .A2(n8799), .ZN(n12520) );
  XOR2_X1 U12622 ( .A(n12695), .B(n12696), .Z(n12517) );
  XOR2_X1 U12623 ( .A(n12697), .B(n12698), .Z(n12696) );
  OR2_X1 U12624 ( .A1(n8746), .A2(n8799), .ZN(n12524) );
  XOR2_X1 U12625 ( .A(n12699), .B(n12700), .Z(n12521) );
  XOR2_X1 U12626 ( .A(n12701), .B(n12702), .Z(n12700) );
  XOR2_X1 U12627 ( .A(n11721), .B(n12703), .Z(n11714) );
  XOR2_X1 U12628 ( .A(n11720), .B(n11719), .Z(n12703) );
  OR2_X1 U12629 ( .A1(n8746), .A2(n8795), .ZN(n11719) );
  OR2_X1 U12630 ( .A1(n12704), .A2(n12705), .ZN(n11720) );
  AND2_X1 U12631 ( .A1(n12702), .A2(n12701), .ZN(n12705) );
  AND2_X1 U12632 ( .A1(n12699), .A2(n12706), .ZN(n12704) );
  OR2_X1 U12633 ( .A1(n12702), .A2(n12701), .ZN(n12706) );
  OR2_X1 U12634 ( .A1(n12707), .A2(n12708), .ZN(n12701) );
  AND2_X1 U12635 ( .A1(n12698), .A2(n12697), .ZN(n12708) );
  AND2_X1 U12636 ( .A1(n12695), .A2(n12709), .ZN(n12707) );
  OR2_X1 U12637 ( .A1(n12698), .A2(n12697), .ZN(n12709) );
  OR2_X1 U12638 ( .A1(n12710), .A2(n12711), .ZN(n12697) );
  AND2_X1 U12639 ( .A1(n12694), .A2(n12693), .ZN(n12711) );
  AND2_X1 U12640 ( .A1(n12691), .A2(n12712), .ZN(n12710) );
  OR2_X1 U12641 ( .A1(n12694), .A2(n12693), .ZN(n12712) );
  OR2_X1 U12642 ( .A1(n12713), .A2(n12714), .ZN(n12693) );
  AND2_X1 U12643 ( .A1(n12690), .A2(n12689), .ZN(n12714) );
  AND2_X1 U12644 ( .A1(n12687), .A2(n12715), .ZN(n12713) );
  OR2_X1 U12645 ( .A1(n12690), .A2(n12689), .ZN(n12715) );
  OR2_X1 U12646 ( .A1(n12716), .A2(n12717), .ZN(n12689) );
  AND2_X1 U12647 ( .A1(n12686), .A2(n12685), .ZN(n12717) );
  AND2_X1 U12648 ( .A1(n12683), .A2(n12718), .ZN(n12716) );
  OR2_X1 U12649 ( .A1(n12686), .A2(n12685), .ZN(n12718) );
  OR2_X1 U12650 ( .A1(n12719), .A2(n12720), .ZN(n12685) );
  AND2_X1 U12651 ( .A1(n12682), .A2(n12681), .ZN(n12720) );
  AND2_X1 U12652 ( .A1(n12679), .A2(n12721), .ZN(n12719) );
  OR2_X1 U12653 ( .A1(n12682), .A2(n12681), .ZN(n12721) );
  OR2_X1 U12654 ( .A1(n12722), .A2(n12723), .ZN(n12681) );
  AND2_X1 U12655 ( .A1(n12678), .A2(n12677), .ZN(n12723) );
  AND2_X1 U12656 ( .A1(n12675), .A2(n12724), .ZN(n12722) );
  OR2_X1 U12657 ( .A1(n12678), .A2(n12677), .ZN(n12724) );
  OR2_X1 U12658 ( .A1(n12725), .A2(n12726), .ZN(n12677) );
  AND2_X1 U12659 ( .A1(n12674), .A2(n12673), .ZN(n12726) );
  AND2_X1 U12660 ( .A1(n12671), .A2(n12727), .ZN(n12725) );
  OR2_X1 U12661 ( .A1(n12674), .A2(n12673), .ZN(n12727) );
  OR2_X1 U12662 ( .A1(n12728), .A2(n12729), .ZN(n12673) );
  AND2_X1 U12663 ( .A1(n12670), .A2(n12669), .ZN(n12729) );
  AND2_X1 U12664 ( .A1(n12667), .A2(n12730), .ZN(n12728) );
  OR2_X1 U12665 ( .A1(n12670), .A2(n12669), .ZN(n12730) );
  OR2_X1 U12666 ( .A1(n12731), .A2(n12732), .ZN(n12669) );
  AND2_X1 U12667 ( .A1(n12666), .A2(n12665), .ZN(n12732) );
  AND2_X1 U12668 ( .A1(n12663), .A2(n12733), .ZN(n12731) );
  OR2_X1 U12669 ( .A1(n12666), .A2(n12665), .ZN(n12733) );
  OR2_X1 U12670 ( .A1(n12734), .A2(n12735), .ZN(n12665) );
  AND2_X1 U12671 ( .A1(n12662), .A2(n12661), .ZN(n12735) );
  AND2_X1 U12672 ( .A1(n12659), .A2(n12736), .ZN(n12734) );
  OR2_X1 U12673 ( .A1(n12662), .A2(n12661), .ZN(n12736) );
  OR2_X1 U12674 ( .A1(n12737), .A2(n12738), .ZN(n12661) );
  AND2_X1 U12675 ( .A1(n8270), .A2(n12658), .ZN(n12738) );
  AND2_X1 U12676 ( .A1(n12656), .A2(n12739), .ZN(n12737) );
  OR2_X1 U12677 ( .A1(n8270), .A2(n12658), .ZN(n12739) );
  OR2_X1 U12678 ( .A1(n12740), .A2(n12741), .ZN(n12658) );
  AND2_X1 U12679 ( .A1(n12655), .A2(n12654), .ZN(n12741) );
  AND2_X1 U12680 ( .A1(n12652), .A2(n12742), .ZN(n12740) );
  OR2_X1 U12681 ( .A1(n12655), .A2(n12654), .ZN(n12742) );
  OR2_X1 U12682 ( .A1(n12743), .A2(n12744), .ZN(n12654) );
  AND2_X1 U12683 ( .A1(n12651), .A2(n12650), .ZN(n12744) );
  AND2_X1 U12684 ( .A1(n12648), .A2(n12745), .ZN(n12743) );
  OR2_X1 U12685 ( .A1(n12651), .A2(n12650), .ZN(n12745) );
  OR2_X1 U12686 ( .A1(n12746), .A2(n12747), .ZN(n12650) );
  AND2_X1 U12687 ( .A1(n12647), .A2(n12646), .ZN(n12747) );
  AND2_X1 U12688 ( .A1(n12644), .A2(n12748), .ZN(n12746) );
  OR2_X1 U12689 ( .A1(n12647), .A2(n12646), .ZN(n12748) );
  OR2_X1 U12690 ( .A1(n12749), .A2(n12750), .ZN(n12646) );
  AND2_X1 U12691 ( .A1(n12643), .A2(n12642), .ZN(n12750) );
  AND2_X1 U12692 ( .A1(n12640), .A2(n12751), .ZN(n12749) );
  OR2_X1 U12693 ( .A1(n12643), .A2(n12642), .ZN(n12751) );
  OR2_X1 U12694 ( .A1(n12752), .A2(n12753), .ZN(n12642) );
  AND2_X1 U12695 ( .A1(n12639), .A2(n12638), .ZN(n12753) );
  AND2_X1 U12696 ( .A1(n12636), .A2(n12754), .ZN(n12752) );
  OR2_X1 U12697 ( .A1(n12639), .A2(n12638), .ZN(n12754) );
  OR2_X1 U12698 ( .A1(n12755), .A2(n12756), .ZN(n12638) );
  AND2_X1 U12699 ( .A1(n12635), .A2(n12634), .ZN(n12756) );
  AND2_X1 U12700 ( .A1(n12632), .A2(n12757), .ZN(n12755) );
  OR2_X1 U12701 ( .A1(n12635), .A2(n12634), .ZN(n12757) );
  OR2_X1 U12702 ( .A1(n12758), .A2(n12759), .ZN(n12634) );
  AND2_X1 U12703 ( .A1(n12631), .A2(n12630), .ZN(n12759) );
  AND2_X1 U12704 ( .A1(n12628), .A2(n12760), .ZN(n12758) );
  OR2_X1 U12705 ( .A1(n12631), .A2(n12630), .ZN(n12760) );
  OR2_X1 U12706 ( .A1(n12761), .A2(n12762), .ZN(n12630) );
  AND2_X1 U12707 ( .A1(n12627), .A2(n12626), .ZN(n12762) );
  AND2_X1 U12708 ( .A1(n12624), .A2(n12763), .ZN(n12761) );
  OR2_X1 U12709 ( .A1(n12627), .A2(n12626), .ZN(n12763) );
  OR2_X1 U12710 ( .A1(n12764), .A2(n12765), .ZN(n12626) );
  AND2_X1 U12711 ( .A1(n12623), .A2(n12622), .ZN(n12765) );
  AND2_X1 U12712 ( .A1(n12620), .A2(n12766), .ZN(n12764) );
  OR2_X1 U12713 ( .A1(n12623), .A2(n12622), .ZN(n12766) );
  OR2_X1 U12714 ( .A1(n12767), .A2(n12768), .ZN(n12622) );
  AND2_X1 U12715 ( .A1(n12619), .A2(n12618), .ZN(n12768) );
  AND2_X1 U12716 ( .A1(n12616), .A2(n12769), .ZN(n12767) );
  OR2_X1 U12717 ( .A1(n12619), .A2(n12618), .ZN(n12769) );
  OR2_X1 U12718 ( .A1(n12770), .A2(n12771), .ZN(n12618) );
  AND2_X1 U12719 ( .A1(n12615), .A2(n12614), .ZN(n12771) );
  AND2_X1 U12720 ( .A1(n12612), .A2(n12772), .ZN(n12770) );
  OR2_X1 U12721 ( .A1(n12615), .A2(n12614), .ZN(n12772) );
  OR2_X1 U12722 ( .A1(n12773), .A2(n12774), .ZN(n12614) );
  AND2_X1 U12723 ( .A1(n12608), .A2(n12611), .ZN(n12774) );
  AND2_X1 U12724 ( .A1(n12775), .A2(n12776), .ZN(n12773) );
  OR2_X1 U12725 ( .A1(n12608), .A2(n12611), .ZN(n12776) );
  OR3_X1 U12726 ( .A1(n8795), .A2(n8791), .A3(n9796), .ZN(n12611) );
  OR2_X1 U12727 ( .A1(n7954), .A2(n8795), .ZN(n12608) );
  INV_X1 U12728 ( .A(n12610), .ZN(n12775) );
  OR2_X1 U12729 ( .A1(n12777), .A2(n12778), .ZN(n12610) );
  AND2_X1 U12730 ( .A1(b_16_), .A2(n12779), .ZN(n12778) );
  OR2_X1 U12731 ( .A1(n12780), .A2(n9801), .ZN(n12779) );
  AND2_X1 U12732 ( .A1(a_30_), .A2(n8787), .ZN(n12780) );
  AND2_X1 U12733 ( .A1(b_15_), .A2(n12781), .ZN(n12777) );
  OR2_X1 U12734 ( .A1(n12782), .A2(n7920), .ZN(n12781) );
  AND2_X1 U12735 ( .A1(a_31_), .A2(n8791), .ZN(n12782) );
  OR2_X1 U12736 ( .A1(n7979), .A2(n8795), .ZN(n12615) );
  XNOR2_X1 U12737 ( .A(n12783), .B(n12784), .ZN(n12612) );
  XOR2_X1 U12738 ( .A(n12785), .B(n12786), .Z(n12784) );
  OR2_X1 U12739 ( .A1(n8015), .A2(n8795), .ZN(n12619) );
  XOR2_X1 U12740 ( .A(n12787), .B(n12788), .Z(n12616) );
  XOR2_X1 U12741 ( .A(n12789), .B(n12790), .Z(n12788) );
  OR2_X1 U12742 ( .A1(n8040), .A2(n8795), .ZN(n12623) );
  XOR2_X1 U12743 ( .A(n12791), .B(n12792), .Z(n12620) );
  XOR2_X1 U12744 ( .A(n12793), .B(n12794), .Z(n12792) );
  OR2_X1 U12745 ( .A1(n8065), .A2(n8795), .ZN(n12627) );
  XOR2_X1 U12746 ( .A(n12795), .B(n12796), .Z(n12624) );
  XOR2_X1 U12747 ( .A(n12797), .B(n12798), .Z(n12796) );
  OR2_X1 U12748 ( .A1(n8090), .A2(n8795), .ZN(n12631) );
  XOR2_X1 U12749 ( .A(n12799), .B(n12800), .Z(n12628) );
  XOR2_X1 U12750 ( .A(n12801), .B(n12802), .Z(n12800) );
  OR2_X1 U12751 ( .A1(n8115), .A2(n8795), .ZN(n12635) );
  XOR2_X1 U12752 ( .A(n12803), .B(n12804), .Z(n12632) );
  XOR2_X1 U12753 ( .A(n12805), .B(n12806), .Z(n12804) );
  OR2_X1 U12754 ( .A1(n8140), .A2(n8795), .ZN(n12639) );
  XOR2_X1 U12755 ( .A(n12807), .B(n12808), .Z(n12636) );
  XOR2_X1 U12756 ( .A(n12809), .B(n12810), .Z(n12808) );
  OR2_X1 U12757 ( .A1(n8810), .A2(n8795), .ZN(n12643) );
  XOR2_X1 U12758 ( .A(n12811), .B(n12812), .Z(n12640) );
  XOR2_X1 U12759 ( .A(n12813), .B(n12814), .Z(n12812) );
  OR2_X1 U12760 ( .A1(n8806), .A2(n8795), .ZN(n12647) );
  XOR2_X1 U12761 ( .A(n12815), .B(n12816), .Z(n12644) );
  XOR2_X1 U12762 ( .A(n12817), .B(n12818), .Z(n12816) );
  OR2_X1 U12763 ( .A1(n8802), .A2(n8795), .ZN(n12651) );
  XOR2_X1 U12764 ( .A(n12819), .B(n12820), .Z(n12648) );
  XOR2_X1 U12765 ( .A(n12821), .B(n12822), .Z(n12820) );
  OR2_X1 U12766 ( .A1(n8798), .A2(n8795), .ZN(n12655) );
  XOR2_X1 U12767 ( .A(n12823), .B(n12824), .Z(n12652) );
  XOR2_X1 U12768 ( .A(n12825), .B(n12826), .Z(n12824) );
  OR2_X1 U12769 ( .A1(n8794), .A2(n8795), .ZN(n8270) );
  XOR2_X1 U12770 ( .A(n12827), .B(n12828), .Z(n12656) );
  XOR2_X1 U12771 ( .A(n12829), .B(n12830), .Z(n12828) );
  OR2_X1 U12772 ( .A1(n8790), .A2(n8795), .ZN(n12662) );
  XOR2_X1 U12773 ( .A(n12831), .B(n12832), .Z(n12659) );
  XOR2_X1 U12774 ( .A(n12833), .B(n12834), .Z(n12832) );
  OR2_X1 U12775 ( .A1(n8786), .A2(n8795), .ZN(n12666) );
  XOR2_X1 U12776 ( .A(n12835), .B(n12836), .Z(n12663) );
  XOR2_X1 U12777 ( .A(n12837), .B(n8296), .Z(n12836) );
  OR2_X1 U12778 ( .A1(n8782), .A2(n8795), .ZN(n12670) );
  XOR2_X1 U12779 ( .A(n12838), .B(n12839), .Z(n12667) );
  XOR2_X1 U12780 ( .A(n12840), .B(n12841), .Z(n12839) );
  OR2_X1 U12781 ( .A1(n8778), .A2(n8795), .ZN(n12674) );
  XOR2_X1 U12782 ( .A(n12842), .B(n12843), .Z(n12671) );
  XOR2_X1 U12783 ( .A(n12844), .B(n12845), .Z(n12843) );
  OR2_X1 U12784 ( .A1(n8774), .A2(n8795), .ZN(n12678) );
  XOR2_X1 U12785 ( .A(n12846), .B(n12847), .Z(n12675) );
  XOR2_X1 U12786 ( .A(n12848), .B(n12849), .Z(n12847) );
  OR2_X1 U12787 ( .A1(n8770), .A2(n8795), .ZN(n12682) );
  XOR2_X1 U12788 ( .A(n12850), .B(n12851), .Z(n12679) );
  XOR2_X1 U12789 ( .A(n12852), .B(n12853), .Z(n12851) );
  OR2_X1 U12790 ( .A1(n8766), .A2(n8795), .ZN(n12686) );
  XOR2_X1 U12791 ( .A(n12854), .B(n12855), .Z(n12683) );
  XOR2_X1 U12792 ( .A(n12856), .B(n12857), .Z(n12855) );
  OR2_X1 U12793 ( .A1(n8762), .A2(n8795), .ZN(n12690) );
  XOR2_X1 U12794 ( .A(n12858), .B(n12859), .Z(n12687) );
  XOR2_X1 U12795 ( .A(n12860), .B(n12861), .Z(n12859) );
  OR2_X1 U12796 ( .A1(n8758), .A2(n8795), .ZN(n12694) );
  XOR2_X1 U12797 ( .A(n12862), .B(n12863), .Z(n12691) );
  XOR2_X1 U12798 ( .A(n12864), .B(n12865), .Z(n12863) );
  OR2_X1 U12799 ( .A1(n8754), .A2(n8795), .ZN(n12698) );
  XOR2_X1 U12800 ( .A(n12866), .B(n12867), .Z(n12695) );
  XOR2_X1 U12801 ( .A(n12868), .B(n12869), .Z(n12867) );
  OR2_X1 U12802 ( .A1(n8750), .A2(n8795), .ZN(n12702) );
  XOR2_X1 U12803 ( .A(n12870), .B(n12871), .Z(n12699) );
  XOR2_X1 U12804 ( .A(n12872), .B(n12873), .Z(n12871) );
  XOR2_X1 U12805 ( .A(n11728), .B(n12874), .Z(n11721) );
  XOR2_X1 U12806 ( .A(n11727), .B(n11726), .Z(n12874) );
  OR2_X1 U12807 ( .A1(n8750), .A2(n8791), .ZN(n11726) );
  OR2_X1 U12808 ( .A1(n12875), .A2(n12876), .ZN(n11727) );
  AND2_X1 U12809 ( .A1(n12873), .A2(n12872), .ZN(n12876) );
  AND2_X1 U12810 ( .A1(n12870), .A2(n12877), .ZN(n12875) );
  OR2_X1 U12811 ( .A1(n12873), .A2(n12872), .ZN(n12877) );
  OR2_X1 U12812 ( .A1(n12878), .A2(n12879), .ZN(n12872) );
  AND2_X1 U12813 ( .A1(n12869), .A2(n12868), .ZN(n12879) );
  AND2_X1 U12814 ( .A1(n12866), .A2(n12880), .ZN(n12878) );
  OR2_X1 U12815 ( .A1(n12869), .A2(n12868), .ZN(n12880) );
  OR2_X1 U12816 ( .A1(n12881), .A2(n12882), .ZN(n12868) );
  AND2_X1 U12817 ( .A1(n12865), .A2(n12864), .ZN(n12882) );
  AND2_X1 U12818 ( .A1(n12862), .A2(n12883), .ZN(n12881) );
  OR2_X1 U12819 ( .A1(n12865), .A2(n12864), .ZN(n12883) );
  OR2_X1 U12820 ( .A1(n12884), .A2(n12885), .ZN(n12864) );
  AND2_X1 U12821 ( .A1(n12861), .A2(n12860), .ZN(n12885) );
  AND2_X1 U12822 ( .A1(n12858), .A2(n12886), .ZN(n12884) );
  OR2_X1 U12823 ( .A1(n12861), .A2(n12860), .ZN(n12886) );
  OR2_X1 U12824 ( .A1(n12887), .A2(n12888), .ZN(n12860) );
  AND2_X1 U12825 ( .A1(n12857), .A2(n12856), .ZN(n12888) );
  AND2_X1 U12826 ( .A1(n12854), .A2(n12889), .ZN(n12887) );
  OR2_X1 U12827 ( .A1(n12857), .A2(n12856), .ZN(n12889) );
  OR2_X1 U12828 ( .A1(n12890), .A2(n12891), .ZN(n12856) );
  AND2_X1 U12829 ( .A1(n12853), .A2(n12852), .ZN(n12891) );
  AND2_X1 U12830 ( .A1(n12850), .A2(n12892), .ZN(n12890) );
  OR2_X1 U12831 ( .A1(n12853), .A2(n12852), .ZN(n12892) );
  OR2_X1 U12832 ( .A1(n12893), .A2(n12894), .ZN(n12852) );
  AND2_X1 U12833 ( .A1(n12846), .A2(n12849), .ZN(n12894) );
  AND2_X1 U12834 ( .A1(n12895), .A2(n12848), .ZN(n12893) );
  OR2_X1 U12835 ( .A1(n12896), .A2(n12897), .ZN(n12848) );
  AND2_X1 U12836 ( .A1(n12845), .A2(n12844), .ZN(n12897) );
  AND2_X1 U12837 ( .A1(n12842), .A2(n12898), .ZN(n12896) );
  OR2_X1 U12838 ( .A1(n12845), .A2(n12844), .ZN(n12898) );
  OR2_X1 U12839 ( .A1(n12899), .A2(n12900), .ZN(n12844) );
  AND2_X1 U12840 ( .A1(n12838), .A2(n12841), .ZN(n12900) );
  AND2_X1 U12841 ( .A1(n12901), .A2(n12840), .ZN(n12899) );
  OR2_X1 U12842 ( .A1(n12902), .A2(n12903), .ZN(n12840) );
  AND2_X1 U12843 ( .A1(n12835), .A2(n8296), .ZN(n12903) );
  AND2_X1 U12844 ( .A1(n12904), .A2(n12837), .ZN(n12902) );
  OR2_X1 U12845 ( .A1(n12905), .A2(n12906), .ZN(n12837) );
  AND2_X1 U12846 ( .A1(n12831), .A2(n12834), .ZN(n12906) );
  AND2_X1 U12847 ( .A1(n12907), .A2(n12833), .ZN(n12905) );
  OR2_X1 U12848 ( .A1(n12908), .A2(n12909), .ZN(n12833) );
  AND2_X1 U12849 ( .A1(n12827), .A2(n12830), .ZN(n12909) );
  AND2_X1 U12850 ( .A1(n12910), .A2(n12829), .ZN(n12908) );
  OR2_X1 U12851 ( .A1(n12911), .A2(n12912), .ZN(n12829) );
  AND2_X1 U12852 ( .A1(n12823), .A2(n12826), .ZN(n12912) );
  AND2_X1 U12853 ( .A1(n12913), .A2(n12825), .ZN(n12911) );
  OR2_X1 U12854 ( .A1(n12914), .A2(n12915), .ZN(n12825) );
  AND2_X1 U12855 ( .A1(n12819), .A2(n12822), .ZN(n12915) );
  AND2_X1 U12856 ( .A1(n12916), .A2(n12821), .ZN(n12914) );
  OR2_X1 U12857 ( .A1(n12917), .A2(n12918), .ZN(n12821) );
  AND2_X1 U12858 ( .A1(n12815), .A2(n12818), .ZN(n12918) );
  AND2_X1 U12859 ( .A1(n12919), .A2(n12817), .ZN(n12917) );
  OR2_X1 U12860 ( .A1(n12920), .A2(n12921), .ZN(n12817) );
  AND2_X1 U12861 ( .A1(n12811), .A2(n12814), .ZN(n12921) );
  AND2_X1 U12862 ( .A1(n12922), .A2(n12813), .ZN(n12920) );
  OR2_X1 U12863 ( .A1(n12923), .A2(n12924), .ZN(n12813) );
  AND2_X1 U12864 ( .A1(n12807), .A2(n12810), .ZN(n12924) );
  AND2_X1 U12865 ( .A1(n12925), .A2(n12809), .ZN(n12923) );
  OR2_X1 U12866 ( .A1(n12926), .A2(n12927), .ZN(n12809) );
  AND2_X1 U12867 ( .A1(n12803), .A2(n12806), .ZN(n12927) );
  AND2_X1 U12868 ( .A1(n12928), .A2(n12805), .ZN(n12926) );
  OR2_X1 U12869 ( .A1(n12929), .A2(n12930), .ZN(n12805) );
  AND2_X1 U12870 ( .A1(n12799), .A2(n12802), .ZN(n12930) );
  AND2_X1 U12871 ( .A1(n12931), .A2(n12801), .ZN(n12929) );
  OR2_X1 U12872 ( .A1(n12932), .A2(n12933), .ZN(n12801) );
  AND2_X1 U12873 ( .A1(n12795), .A2(n12798), .ZN(n12933) );
  AND2_X1 U12874 ( .A1(n12934), .A2(n12797), .ZN(n12932) );
  OR2_X1 U12875 ( .A1(n12935), .A2(n12936), .ZN(n12797) );
  AND2_X1 U12876 ( .A1(n12791), .A2(n12794), .ZN(n12936) );
  AND2_X1 U12877 ( .A1(n12937), .A2(n12793), .ZN(n12935) );
  OR2_X1 U12878 ( .A1(n12938), .A2(n12939), .ZN(n12793) );
  AND2_X1 U12879 ( .A1(n12787), .A2(n12790), .ZN(n12939) );
  AND2_X1 U12880 ( .A1(n12940), .A2(n12789), .ZN(n12938) );
  OR2_X1 U12881 ( .A1(n12941), .A2(n12942), .ZN(n12789) );
  AND2_X1 U12882 ( .A1(n12783), .A2(n12786), .ZN(n12942) );
  AND2_X1 U12883 ( .A1(n12943), .A2(n12944), .ZN(n12941) );
  OR2_X1 U12884 ( .A1(n12783), .A2(n12786), .ZN(n12944) );
  OR3_X1 U12885 ( .A1(n8791), .A2(n8787), .A3(n9796), .ZN(n12786) );
  OR2_X1 U12886 ( .A1(n7954), .A2(n8791), .ZN(n12783) );
  INV_X1 U12887 ( .A(n12785), .ZN(n12943) );
  OR2_X1 U12888 ( .A1(n12945), .A2(n12946), .ZN(n12785) );
  AND2_X1 U12889 ( .A1(b_15_), .A2(n12947), .ZN(n12946) );
  OR2_X1 U12890 ( .A1(n12948), .A2(n9801), .ZN(n12947) );
  AND2_X1 U12891 ( .A1(a_30_), .A2(n8783), .ZN(n12948) );
  AND2_X1 U12892 ( .A1(b_14_), .A2(n12949), .ZN(n12945) );
  OR2_X1 U12893 ( .A1(n12950), .A2(n7920), .ZN(n12949) );
  AND2_X1 U12894 ( .A1(a_31_), .A2(n8787), .ZN(n12950) );
  OR2_X1 U12895 ( .A1(n12787), .A2(n12790), .ZN(n12940) );
  OR2_X1 U12896 ( .A1(n7979), .A2(n8791), .ZN(n12790) );
  XNOR2_X1 U12897 ( .A(n12951), .B(n12952), .ZN(n12787) );
  XOR2_X1 U12898 ( .A(n12953), .B(n12954), .Z(n12952) );
  OR2_X1 U12899 ( .A1(n12791), .A2(n12794), .ZN(n12937) );
  OR2_X1 U12900 ( .A1(n8015), .A2(n8791), .ZN(n12794) );
  XOR2_X1 U12901 ( .A(n12955), .B(n12956), .Z(n12791) );
  XOR2_X1 U12902 ( .A(n12957), .B(n12958), .Z(n12956) );
  OR2_X1 U12903 ( .A1(n12795), .A2(n12798), .ZN(n12934) );
  OR2_X1 U12904 ( .A1(n8040), .A2(n8791), .ZN(n12798) );
  XOR2_X1 U12905 ( .A(n12959), .B(n12960), .Z(n12795) );
  XOR2_X1 U12906 ( .A(n12961), .B(n12962), .Z(n12960) );
  OR2_X1 U12907 ( .A1(n12799), .A2(n12802), .ZN(n12931) );
  OR2_X1 U12908 ( .A1(n8065), .A2(n8791), .ZN(n12802) );
  XOR2_X1 U12909 ( .A(n12963), .B(n12964), .Z(n12799) );
  XOR2_X1 U12910 ( .A(n12965), .B(n12966), .Z(n12964) );
  OR2_X1 U12911 ( .A1(n12803), .A2(n12806), .ZN(n12928) );
  OR2_X1 U12912 ( .A1(n8090), .A2(n8791), .ZN(n12806) );
  XOR2_X1 U12913 ( .A(n12967), .B(n12968), .Z(n12803) );
  XOR2_X1 U12914 ( .A(n12969), .B(n12970), .Z(n12968) );
  OR2_X1 U12915 ( .A1(n12807), .A2(n12810), .ZN(n12925) );
  OR2_X1 U12916 ( .A1(n8115), .A2(n8791), .ZN(n12810) );
  XOR2_X1 U12917 ( .A(n12971), .B(n12972), .Z(n12807) );
  XOR2_X1 U12918 ( .A(n12973), .B(n12974), .Z(n12972) );
  OR2_X1 U12919 ( .A1(n12811), .A2(n12814), .ZN(n12922) );
  OR2_X1 U12920 ( .A1(n8140), .A2(n8791), .ZN(n12814) );
  XOR2_X1 U12921 ( .A(n12975), .B(n12976), .Z(n12811) );
  XOR2_X1 U12922 ( .A(n12977), .B(n12978), .Z(n12976) );
  OR2_X1 U12923 ( .A1(n12815), .A2(n12818), .ZN(n12919) );
  OR2_X1 U12924 ( .A1(n8810), .A2(n8791), .ZN(n12818) );
  XOR2_X1 U12925 ( .A(n12979), .B(n12980), .Z(n12815) );
  XOR2_X1 U12926 ( .A(n12981), .B(n12982), .Z(n12980) );
  OR2_X1 U12927 ( .A1(n12819), .A2(n12822), .ZN(n12916) );
  OR2_X1 U12928 ( .A1(n8806), .A2(n8791), .ZN(n12822) );
  XOR2_X1 U12929 ( .A(n12983), .B(n12984), .Z(n12819) );
  XOR2_X1 U12930 ( .A(n12985), .B(n12986), .Z(n12984) );
  OR2_X1 U12931 ( .A1(n12823), .A2(n12826), .ZN(n12913) );
  OR2_X1 U12932 ( .A1(n8802), .A2(n8791), .ZN(n12826) );
  XOR2_X1 U12933 ( .A(n12987), .B(n12988), .Z(n12823) );
  XOR2_X1 U12934 ( .A(n12989), .B(n12990), .Z(n12988) );
  OR2_X1 U12935 ( .A1(n12827), .A2(n12830), .ZN(n12910) );
  OR2_X1 U12936 ( .A1(n8798), .A2(n8791), .ZN(n12830) );
  XOR2_X1 U12937 ( .A(n12991), .B(n12992), .Z(n12827) );
  XOR2_X1 U12938 ( .A(n12993), .B(n12994), .Z(n12992) );
  OR2_X1 U12939 ( .A1(n12831), .A2(n12834), .ZN(n12907) );
  OR2_X1 U12940 ( .A1(n8794), .A2(n8791), .ZN(n12834) );
  XOR2_X1 U12941 ( .A(n12995), .B(n12996), .Z(n12831) );
  XOR2_X1 U12942 ( .A(n12997), .B(n12998), .Z(n12996) );
  OR2_X1 U12943 ( .A1(n12835), .A2(n8296), .ZN(n12904) );
  OR2_X1 U12944 ( .A1(n8790), .A2(n8791), .ZN(n8296) );
  XOR2_X1 U12945 ( .A(n12999), .B(n13000), .Z(n12835) );
  XOR2_X1 U12946 ( .A(n13001), .B(n13002), .Z(n13000) );
  OR2_X1 U12947 ( .A1(n12838), .A2(n12841), .ZN(n12901) );
  OR2_X1 U12948 ( .A1(n8786), .A2(n8791), .ZN(n12841) );
  XOR2_X1 U12949 ( .A(n13003), .B(n13004), .Z(n12838) );
  XOR2_X1 U12950 ( .A(n13005), .B(n13006), .Z(n13004) );
  OR2_X1 U12951 ( .A1(n8782), .A2(n8791), .ZN(n12845) );
  XOR2_X1 U12952 ( .A(n13007), .B(n13008), .Z(n12842) );
  XOR2_X1 U12953 ( .A(n13009), .B(n8322), .Z(n13008) );
  OR2_X1 U12954 ( .A1(n12846), .A2(n12849), .ZN(n12895) );
  OR2_X1 U12955 ( .A1(n8778), .A2(n8791), .ZN(n12849) );
  XOR2_X1 U12956 ( .A(n13010), .B(n13011), .Z(n12846) );
  XOR2_X1 U12957 ( .A(n13012), .B(n13013), .Z(n13011) );
  OR2_X1 U12958 ( .A1(n8774), .A2(n8791), .ZN(n12853) );
  XOR2_X1 U12959 ( .A(n13014), .B(n13015), .Z(n12850) );
  XOR2_X1 U12960 ( .A(n13016), .B(n13017), .Z(n13015) );
  OR2_X1 U12961 ( .A1(n8770), .A2(n8791), .ZN(n12857) );
  XOR2_X1 U12962 ( .A(n13018), .B(n13019), .Z(n12854) );
  XOR2_X1 U12963 ( .A(n13020), .B(n13021), .Z(n13019) );
  OR2_X1 U12964 ( .A1(n8766), .A2(n8791), .ZN(n12861) );
  XOR2_X1 U12965 ( .A(n13022), .B(n13023), .Z(n12858) );
  XOR2_X1 U12966 ( .A(n13024), .B(n13025), .Z(n13023) );
  OR2_X1 U12967 ( .A1(n8762), .A2(n8791), .ZN(n12865) );
  XOR2_X1 U12968 ( .A(n13026), .B(n13027), .Z(n12862) );
  XOR2_X1 U12969 ( .A(n13028), .B(n13029), .Z(n13027) );
  OR2_X1 U12970 ( .A1(n8758), .A2(n8791), .ZN(n12869) );
  XOR2_X1 U12971 ( .A(n13030), .B(n13031), .Z(n12866) );
  XOR2_X1 U12972 ( .A(n13032), .B(n13033), .Z(n13031) );
  OR2_X1 U12973 ( .A1(n8754), .A2(n8791), .ZN(n12873) );
  XOR2_X1 U12974 ( .A(n13034), .B(n13035), .Z(n12870) );
  XOR2_X1 U12975 ( .A(n13036), .B(n13037), .Z(n13035) );
  XOR2_X1 U12976 ( .A(n11735), .B(n13038), .Z(n11728) );
  XOR2_X1 U12977 ( .A(n11734), .B(n11733), .Z(n13038) );
  OR2_X1 U12978 ( .A1(n8754), .A2(n8787), .ZN(n11733) );
  OR2_X1 U12979 ( .A1(n13039), .A2(n13040), .ZN(n11734) );
  AND2_X1 U12980 ( .A1(n13037), .A2(n13036), .ZN(n13040) );
  AND2_X1 U12981 ( .A1(n13034), .A2(n13041), .ZN(n13039) );
  OR2_X1 U12982 ( .A1(n13036), .A2(n13037), .ZN(n13041) );
  OR2_X1 U12983 ( .A1(n8758), .A2(n8787), .ZN(n13037) );
  OR2_X1 U12984 ( .A1(n13042), .A2(n13043), .ZN(n13036) );
  AND2_X1 U12985 ( .A1(n13033), .A2(n13032), .ZN(n13043) );
  AND2_X1 U12986 ( .A1(n13030), .A2(n13044), .ZN(n13042) );
  OR2_X1 U12987 ( .A1(n13032), .A2(n13033), .ZN(n13044) );
  OR2_X1 U12988 ( .A1(n8762), .A2(n8787), .ZN(n13033) );
  OR2_X1 U12989 ( .A1(n13045), .A2(n13046), .ZN(n13032) );
  AND2_X1 U12990 ( .A1(n13029), .A2(n13028), .ZN(n13046) );
  AND2_X1 U12991 ( .A1(n13026), .A2(n13047), .ZN(n13045) );
  OR2_X1 U12992 ( .A1(n13028), .A2(n13029), .ZN(n13047) );
  OR2_X1 U12993 ( .A1(n8766), .A2(n8787), .ZN(n13029) );
  OR2_X1 U12994 ( .A1(n13048), .A2(n13049), .ZN(n13028) );
  AND2_X1 U12995 ( .A1(n13025), .A2(n13024), .ZN(n13049) );
  AND2_X1 U12996 ( .A1(n13022), .A2(n13050), .ZN(n13048) );
  OR2_X1 U12997 ( .A1(n13024), .A2(n13025), .ZN(n13050) );
  OR2_X1 U12998 ( .A1(n8770), .A2(n8787), .ZN(n13025) );
  OR2_X1 U12999 ( .A1(n13051), .A2(n13052), .ZN(n13024) );
  AND2_X1 U13000 ( .A1(n13021), .A2(n13020), .ZN(n13052) );
  AND2_X1 U13001 ( .A1(n13018), .A2(n13053), .ZN(n13051) );
  OR2_X1 U13002 ( .A1(n13020), .A2(n13021), .ZN(n13053) );
  OR2_X1 U13003 ( .A1(n8774), .A2(n8787), .ZN(n13021) );
  OR2_X1 U13004 ( .A1(n13054), .A2(n13055), .ZN(n13020) );
  AND2_X1 U13005 ( .A1(n13017), .A2(n13016), .ZN(n13055) );
  AND2_X1 U13006 ( .A1(n13014), .A2(n13056), .ZN(n13054) );
  OR2_X1 U13007 ( .A1(n13016), .A2(n13017), .ZN(n13056) );
  OR2_X1 U13008 ( .A1(n8778), .A2(n8787), .ZN(n13017) );
  OR2_X1 U13009 ( .A1(n13057), .A2(n13058), .ZN(n13016) );
  AND2_X1 U13010 ( .A1(n13013), .A2(n13012), .ZN(n13058) );
  AND2_X1 U13011 ( .A1(n13010), .A2(n13059), .ZN(n13057) );
  OR2_X1 U13012 ( .A1(n13012), .A2(n13013), .ZN(n13059) );
  OR2_X1 U13013 ( .A1(n8782), .A2(n8787), .ZN(n13013) );
  OR2_X1 U13014 ( .A1(n13060), .A2(n13061), .ZN(n13012) );
  AND2_X1 U13015 ( .A1(n8322), .A2(n13009), .ZN(n13061) );
  AND2_X1 U13016 ( .A1(n13007), .A2(n13062), .ZN(n13060) );
  OR2_X1 U13017 ( .A1(n13009), .A2(n8322), .ZN(n13062) );
  OR2_X1 U13018 ( .A1(n8786), .A2(n8787), .ZN(n8322) );
  OR2_X1 U13019 ( .A1(n13063), .A2(n13064), .ZN(n13009) );
  AND2_X1 U13020 ( .A1(n13006), .A2(n13005), .ZN(n13064) );
  AND2_X1 U13021 ( .A1(n13003), .A2(n13065), .ZN(n13063) );
  OR2_X1 U13022 ( .A1(n13005), .A2(n13006), .ZN(n13065) );
  OR2_X1 U13023 ( .A1(n8790), .A2(n8787), .ZN(n13006) );
  OR2_X1 U13024 ( .A1(n13066), .A2(n13067), .ZN(n13005) );
  AND2_X1 U13025 ( .A1(n13002), .A2(n13001), .ZN(n13067) );
  AND2_X1 U13026 ( .A1(n12999), .A2(n13068), .ZN(n13066) );
  OR2_X1 U13027 ( .A1(n13001), .A2(n13002), .ZN(n13068) );
  OR2_X1 U13028 ( .A1(n8794), .A2(n8787), .ZN(n13002) );
  OR2_X1 U13029 ( .A1(n13069), .A2(n13070), .ZN(n13001) );
  AND2_X1 U13030 ( .A1(n12998), .A2(n12997), .ZN(n13070) );
  AND2_X1 U13031 ( .A1(n12995), .A2(n13071), .ZN(n13069) );
  OR2_X1 U13032 ( .A1(n12997), .A2(n12998), .ZN(n13071) );
  OR2_X1 U13033 ( .A1(n8798), .A2(n8787), .ZN(n12998) );
  OR2_X1 U13034 ( .A1(n13072), .A2(n13073), .ZN(n12997) );
  AND2_X1 U13035 ( .A1(n12994), .A2(n12993), .ZN(n13073) );
  AND2_X1 U13036 ( .A1(n12991), .A2(n13074), .ZN(n13072) );
  OR2_X1 U13037 ( .A1(n12993), .A2(n12994), .ZN(n13074) );
  OR2_X1 U13038 ( .A1(n8802), .A2(n8787), .ZN(n12994) );
  OR2_X1 U13039 ( .A1(n13075), .A2(n13076), .ZN(n12993) );
  AND2_X1 U13040 ( .A1(n12990), .A2(n12989), .ZN(n13076) );
  AND2_X1 U13041 ( .A1(n12987), .A2(n13077), .ZN(n13075) );
  OR2_X1 U13042 ( .A1(n12989), .A2(n12990), .ZN(n13077) );
  OR2_X1 U13043 ( .A1(n8806), .A2(n8787), .ZN(n12990) );
  OR2_X1 U13044 ( .A1(n13078), .A2(n13079), .ZN(n12989) );
  AND2_X1 U13045 ( .A1(n12986), .A2(n12985), .ZN(n13079) );
  AND2_X1 U13046 ( .A1(n12983), .A2(n13080), .ZN(n13078) );
  OR2_X1 U13047 ( .A1(n12985), .A2(n12986), .ZN(n13080) );
  OR2_X1 U13048 ( .A1(n8810), .A2(n8787), .ZN(n12986) );
  OR2_X1 U13049 ( .A1(n13081), .A2(n13082), .ZN(n12985) );
  AND2_X1 U13050 ( .A1(n12982), .A2(n12981), .ZN(n13082) );
  AND2_X1 U13051 ( .A1(n12979), .A2(n13083), .ZN(n13081) );
  OR2_X1 U13052 ( .A1(n12981), .A2(n12982), .ZN(n13083) );
  OR2_X1 U13053 ( .A1(n8140), .A2(n8787), .ZN(n12982) );
  OR2_X1 U13054 ( .A1(n13084), .A2(n13085), .ZN(n12981) );
  AND2_X1 U13055 ( .A1(n12978), .A2(n12977), .ZN(n13085) );
  AND2_X1 U13056 ( .A1(n12975), .A2(n13086), .ZN(n13084) );
  OR2_X1 U13057 ( .A1(n12977), .A2(n12978), .ZN(n13086) );
  OR2_X1 U13058 ( .A1(n8115), .A2(n8787), .ZN(n12978) );
  OR2_X1 U13059 ( .A1(n13087), .A2(n13088), .ZN(n12977) );
  AND2_X1 U13060 ( .A1(n12974), .A2(n12973), .ZN(n13088) );
  AND2_X1 U13061 ( .A1(n12971), .A2(n13089), .ZN(n13087) );
  OR2_X1 U13062 ( .A1(n12973), .A2(n12974), .ZN(n13089) );
  OR2_X1 U13063 ( .A1(n8090), .A2(n8787), .ZN(n12974) );
  OR2_X1 U13064 ( .A1(n13090), .A2(n13091), .ZN(n12973) );
  AND2_X1 U13065 ( .A1(n12970), .A2(n12969), .ZN(n13091) );
  AND2_X1 U13066 ( .A1(n12967), .A2(n13092), .ZN(n13090) );
  OR2_X1 U13067 ( .A1(n12969), .A2(n12970), .ZN(n13092) );
  OR2_X1 U13068 ( .A1(n8065), .A2(n8787), .ZN(n12970) );
  OR2_X1 U13069 ( .A1(n13093), .A2(n13094), .ZN(n12969) );
  AND2_X1 U13070 ( .A1(n12966), .A2(n12965), .ZN(n13094) );
  AND2_X1 U13071 ( .A1(n12963), .A2(n13095), .ZN(n13093) );
  OR2_X1 U13072 ( .A1(n12965), .A2(n12966), .ZN(n13095) );
  OR2_X1 U13073 ( .A1(n8040), .A2(n8787), .ZN(n12966) );
  OR2_X1 U13074 ( .A1(n13096), .A2(n13097), .ZN(n12965) );
  AND2_X1 U13075 ( .A1(n12962), .A2(n12961), .ZN(n13097) );
  AND2_X1 U13076 ( .A1(n12959), .A2(n13098), .ZN(n13096) );
  OR2_X1 U13077 ( .A1(n12961), .A2(n12962), .ZN(n13098) );
  OR2_X1 U13078 ( .A1(n8015), .A2(n8787), .ZN(n12962) );
  OR2_X1 U13079 ( .A1(n13099), .A2(n13100), .ZN(n12961) );
  AND2_X1 U13080 ( .A1(n12958), .A2(n12957), .ZN(n13100) );
  AND2_X1 U13081 ( .A1(n12955), .A2(n13101), .ZN(n13099) );
  OR2_X1 U13082 ( .A1(n12957), .A2(n12958), .ZN(n13101) );
  OR2_X1 U13083 ( .A1(n7979), .A2(n8787), .ZN(n12958) );
  OR2_X1 U13084 ( .A1(n13102), .A2(n13103), .ZN(n12957) );
  AND2_X1 U13085 ( .A1(n12951), .A2(n12954), .ZN(n13103) );
  AND2_X1 U13086 ( .A1(n13104), .A2(n13105), .ZN(n13102) );
  OR2_X1 U13087 ( .A1(n12954), .A2(n12951), .ZN(n13105) );
  OR2_X1 U13088 ( .A1(n7954), .A2(n8787), .ZN(n12951) );
  OR3_X1 U13089 ( .A1(n8787), .A2(n8783), .A3(n9796), .ZN(n12954) );
  INV_X1 U13090 ( .A(n12953), .ZN(n13104) );
  OR2_X1 U13091 ( .A1(n13106), .A2(n13107), .ZN(n12953) );
  AND2_X1 U13092 ( .A1(b_14_), .A2(n13108), .ZN(n13107) );
  OR2_X1 U13093 ( .A1(n13109), .A2(n9801), .ZN(n13108) );
  AND2_X1 U13094 ( .A1(a_30_), .A2(n8779), .ZN(n13109) );
  AND2_X1 U13095 ( .A1(b_13_), .A2(n13110), .ZN(n13106) );
  OR2_X1 U13096 ( .A1(n13111), .A2(n7920), .ZN(n13110) );
  AND2_X1 U13097 ( .A1(a_31_), .A2(n8783), .ZN(n13111) );
  XNOR2_X1 U13098 ( .A(n13112), .B(n13113), .ZN(n12955) );
  XOR2_X1 U13099 ( .A(n13114), .B(n13115), .Z(n13113) );
  XOR2_X1 U13100 ( .A(n13116), .B(n13117), .Z(n12959) );
  XOR2_X1 U13101 ( .A(n13118), .B(n13119), .Z(n13117) );
  XOR2_X1 U13102 ( .A(n13120), .B(n13121), .Z(n12963) );
  XOR2_X1 U13103 ( .A(n13122), .B(n13123), .Z(n13121) );
  XOR2_X1 U13104 ( .A(n13124), .B(n13125), .Z(n12967) );
  XOR2_X1 U13105 ( .A(n13126), .B(n13127), .Z(n13125) );
  XOR2_X1 U13106 ( .A(n13128), .B(n13129), .Z(n12971) );
  XOR2_X1 U13107 ( .A(n13130), .B(n13131), .Z(n13129) );
  XOR2_X1 U13108 ( .A(n13132), .B(n13133), .Z(n12975) );
  XOR2_X1 U13109 ( .A(n13134), .B(n13135), .Z(n13133) );
  XOR2_X1 U13110 ( .A(n13136), .B(n13137), .Z(n12979) );
  XOR2_X1 U13111 ( .A(n13138), .B(n13139), .Z(n13137) );
  XOR2_X1 U13112 ( .A(n13140), .B(n13141), .Z(n12983) );
  XOR2_X1 U13113 ( .A(n13142), .B(n13143), .Z(n13141) );
  XOR2_X1 U13114 ( .A(n13144), .B(n13145), .Z(n12987) );
  XOR2_X1 U13115 ( .A(n13146), .B(n13147), .Z(n13145) );
  XOR2_X1 U13116 ( .A(n13148), .B(n13149), .Z(n12991) );
  XOR2_X1 U13117 ( .A(n13150), .B(n13151), .Z(n13149) );
  XOR2_X1 U13118 ( .A(n13152), .B(n13153), .Z(n12995) );
  XOR2_X1 U13119 ( .A(n13154), .B(n13155), .Z(n13153) );
  XOR2_X1 U13120 ( .A(n13156), .B(n13157), .Z(n12999) );
  XOR2_X1 U13121 ( .A(n13158), .B(n13159), .Z(n13157) );
  XOR2_X1 U13122 ( .A(n13160), .B(n13161), .Z(n13003) );
  XOR2_X1 U13123 ( .A(n13162), .B(n13163), .Z(n13161) );
  XOR2_X1 U13124 ( .A(n13164), .B(n13165), .Z(n13007) );
  XOR2_X1 U13125 ( .A(n13166), .B(n13167), .Z(n13165) );
  XOR2_X1 U13126 ( .A(n13168), .B(n13169), .Z(n13010) );
  XOR2_X1 U13127 ( .A(n13170), .B(n13171), .Z(n13169) );
  XOR2_X1 U13128 ( .A(n13172), .B(n13173), .Z(n13014) );
  XOR2_X1 U13129 ( .A(n13174), .B(n8348), .Z(n13173) );
  XOR2_X1 U13130 ( .A(n13175), .B(n13176), .Z(n13018) );
  XOR2_X1 U13131 ( .A(n13177), .B(n13178), .Z(n13176) );
  XOR2_X1 U13132 ( .A(n13179), .B(n13180), .Z(n13022) );
  XOR2_X1 U13133 ( .A(n13181), .B(n13182), .Z(n13180) );
  XOR2_X1 U13134 ( .A(n13183), .B(n13184), .Z(n13026) );
  XOR2_X1 U13135 ( .A(n13185), .B(n13186), .Z(n13184) );
  XOR2_X1 U13136 ( .A(n13187), .B(n13188), .Z(n13030) );
  XOR2_X1 U13137 ( .A(n13189), .B(n13190), .Z(n13188) );
  XOR2_X1 U13138 ( .A(n13191), .B(n13192), .Z(n13034) );
  XOR2_X1 U13139 ( .A(n13193), .B(n13194), .Z(n13192) );
  XOR2_X1 U13140 ( .A(n13195), .B(n13196), .Z(n11735) );
  XOR2_X1 U13141 ( .A(n13197), .B(n13198), .Z(n13196) );
  XOR2_X1 U13142 ( .A(n8995), .B(n8994), .Z(n8982) );
  INV_X1 U13143 ( .A(n13199), .ZN(n8994) );
  OR2_X1 U13144 ( .A1(n13200), .A2(n13201), .ZN(n13199) );
  AND2_X1 U13145 ( .A1(n9438), .A2(n9437), .ZN(n13201) );
  AND2_X1 U13146 ( .A1(n9435), .A2(n13202), .ZN(n13200) );
  OR2_X1 U13147 ( .A1(n9437), .A2(n9438), .ZN(n13202) );
  OR2_X1 U13148 ( .A1(n9248), .A2(n8783), .ZN(n9438) );
  OR2_X1 U13149 ( .A1(n13203), .A2(n13204), .ZN(n9437) );
  AND2_X1 U13150 ( .A1(n9462), .A2(n9461), .ZN(n13204) );
  AND2_X1 U13151 ( .A1(n9459), .A2(n13205), .ZN(n13203) );
  OR2_X1 U13152 ( .A1(n9461), .A2(n9462), .ZN(n13205) );
  OR2_X1 U13153 ( .A1(n8730), .A2(n8783), .ZN(n9462) );
  OR2_X1 U13154 ( .A1(n13206), .A2(n13207), .ZN(n9461) );
  AND2_X1 U13155 ( .A1(n9493), .A2(n9492), .ZN(n13207) );
  AND2_X1 U13156 ( .A1(n9490), .A2(n13208), .ZN(n13206) );
  OR2_X1 U13157 ( .A1(n9492), .A2(n9493), .ZN(n13208) );
  OR2_X1 U13158 ( .A1(n8734), .A2(n8783), .ZN(n9493) );
  OR2_X1 U13159 ( .A1(n13209), .A2(n13210), .ZN(n9492) );
  AND2_X1 U13160 ( .A1(n9531), .A2(n9530), .ZN(n13210) );
  AND2_X1 U13161 ( .A1(n9528), .A2(n13211), .ZN(n13209) );
  OR2_X1 U13162 ( .A1(n9530), .A2(n9531), .ZN(n13211) );
  OR2_X1 U13163 ( .A1(n8738), .A2(n8783), .ZN(n9531) );
  OR2_X1 U13164 ( .A1(n13212), .A2(n13213), .ZN(n9530) );
  AND2_X1 U13165 ( .A1(n9576), .A2(n9575), .ZN(n13213) );
  AND2_X1 U13166 ( .A1(n9573), .A2(n13214), .ZN(n13212) );
  OR2_X1 U13167 ( .A1(n9575), .A2(n9576), .ZN(n13214) );
  OR2_X1 U13168 ( .A1(n8742), .A2(n8783), .ZN(n9576) );
  OR2_X1 U13169 ( .A1(n13215), .A2(n13216), .ZN(n9575) );
  AND2_X1 U13170 ( .A1(n9628), .A2(n9627), .ZN(n13216) );
  AND2_X1 U13171 ( .A1(n9625), .A2(n13217), .ZN(n13215) );
  OR2_X1 U13172 ( .A1(n9627), .A2(n9628), .ZN(n13217) );
  OR2_X1 U13173 ( .A1(n8746), .A2(n8783), .ZN(n9628) );
  OR2_X1 U13174 ( .A1(n13218), .A2(n13219), .ZN(n9627) );
  AND2_X1 U13175 ( .A1(n11687), .A2(n11686), .ZN(n13219) );
  AND2_X1 U13176 ( .A1(n11684), .A2(n13220), .ZN(n13218) );
  OR2_X1 U13177 ( .A1(n11686), .A2(n11687), .ZN(n13220) );
  OR2_X1 U13178 ( .A1(n8750), .A2(n8783), .ZN(n11687) );
  OR2_X1 U13179 ( .A1(n13221), .A2(n13222), .ZN(n11686) );
  AND2_X1 U13180 ( .A1(n11740), .A2(n11739), .ZN(n13222) );
  AND2_X1 U13181 ( .A1(n11737), .A2(n13223), .ZN(n13221) );
  OR2_X1 U13182 ( .A1(n11739), .A2(n11740), .ZN(n13223) );
  OR2_X1 U13183 ( .A1(n8754), .A2(n8783), .ZN(n11740) );
  OR2_X1 U13184 ( .A1(n13224), .A2(n13225), .ZN(n11739) );
  AND2_X1 U13185 ( .A1(n13198), .A2(n13197), .ZN(n13225) );
  AND2_X1 U13186 ( .A1(n13195), .A2(n13226), .ZN(n13224) );
  OR2_X1 U13187 ( .A1(n13197), .A2(n13198), .ZN(n13226) );
  OR2_X1 U13188 ( .A1(n8758), .A2(n8783), .ZN(n13198) );
  OR2_X1 U13189 ( .A1(n13227), .A2(n13228), .ZN(n13197) );
  AND2_X1 U13190 ( .A1(n13194), .A2(n13193), .ZN(n13228) );
  AND2_X1 U13191 ( .A1(n13191), .A2(n13229), .ZN(n13227) );
  OR2_X1 U13192 ( .A1(n13193), .A2(n13194), .ZN(n13229) );
  OR2_X1 U13193 ( .A1(n8762), .A2(n8783), .ZN(n13194) );
  OR2_X1 U13194 ( .A1(n13230), .A2(n13231), .ZN(n13193) );
  AND2_X1 U13195 ( .A1(n13190), .A2(n13189), .ZN(n13231) );
  AND2_X1 U13196 ( .A1(n13187), .A2(n13232), .ZN(n13230) );
  OR2_X1 U13197 ( .A1(n13189), .A2(n13190), .ZN(n13232) );
  OR2_X1 U13198 ( .A1(n8766), .A2(n8783), .ZN(n13190) );
  OR2_X1 U13199 ( .A1(n13233), .A2(n13234), .ZN(n13189) );
  AND2_X1 U13200 ( .A1(n13186), .A2(n13185), .ZN(n13234) );
  AND2_X1 U13201 ( .A1(n13183), .A2(n13235), .ZN(n13233) );
  OR2_X1 U13202 ( .A1(n13185), .A2(n13186), .ZN(n13235) );
  OR2_X1 U13203 ( .A1(n8770), .A2(n8783), .ZN(n13186) );
  OR2_X1 U13204 ( .A1(n13236), .A2(n13237), .ZN(n13185) );
  AND2_X1 U13205 ( .A1(n13182), .A2(n13181), .ZN(n13237) );
  AND2_X1 U13206 ( .A1(n13179), .A2(n13238), .ZN(n13236) );
  OR2_X1 U13207 ( .A1(n13181), .A2(n13182), .ZN(n13238) );
  OR2_X1 U13208 ( .A1(n8774), .A2(n8783), .ZN(n13182) );
  OR2_X1 U13209 ( .A1(n13239), .A2(n13240), .ZN(n13181) );
  AND2_X1 U13210 ( .A1(n13178), .A2(n13177), .ZN(n13240) );
  AND2_X1 U13211 ( .A1(n13175), .A2(n13241), .ZN(n13239) );
  OR2_X1 U13212 ( .A1(n13177), .A2(n13178), .ZN(n13241) );
  OR2_X1 U13213 ( .A1(n8778), .A2(n8783), .ZN(n13178) );
  OR2_X1 U13214 ( .A1(n13242), .A2(n13243), .ZN(n13177) );
  AND2_X1 U13215 ( .A1(n8348), .A2(n13174), .ZN(n13243) );
  AND2_X1 U13216 ( .A1(n13172), .A2(n13244), .ZN(n13242) );
  OR2_X1 U13217 ( .A1(n13174), .A2(n8348), .ZN(n13244) );
  OR2_X1 U13218 ( .A1(n8782), .A2(n8783), .ZN(n8348) );
  OR2_X1 U13219 ( .A1(n13245), .A2(n13246), .ZN(n13174) );
  AND2_X1 U13220 ( .A1(n13171), .A2(n13170), .ZN(n13246) );
  AND2_X1 U13221 ( .A1(n13168), .A2(n13247), .ZN(n13245) );
  OR2_X1 U13222 ( .A1(n13170), .A2(n13171), .ZN(n13247) );
  OR2_X1 U13223 ( .A1(n8786), .A2(n8783), .ZN(n13171) );
  OR2_X1 U13224 ( .A1(n13248), .A2(n13249), .ZN(n13170) );
  AND2_X1 U13225 ( .A1(n13167), .A2(n13166), .ZN(n13249) );
  AND2_X1 U13226 ( .A1(n13164), .A2(n13250), .ZN(n13248) );
  OR2_X1 U13227 ( .A1(n13166), .A2(n13167), .ZN(n13250) );
  OR2_X1 U13228 ( .A1(n8790), .A2(n8783), .ZN(n13167) );
  OR2_X1 U13229 ( .A1(n13251), .A2(n13252), .ZN(n13166) );
  AND2_X1 U13230 ( .A1(n13163), .A2(n13162), .ZN(n13252) );
  AND2_X1 U13231 ( .A1(n13160), .A2(n13253), .ZN(n13251) );
  OR2_X1 U13232 ( .A1(n13162), .A2(n13163), .ZN(n13253) );
  OR2_X1 U13233 ( .A1(n8794), .A2(n8783), .ZN(n13163) );
  OR2_X1 U13234 ( .A1(n13254), .A2(n13255), .ZN(n13162) );
  AND2_X1 U13235 ( .A1(n13159), .A2(n13158), .ZN(n13255) );
  AND2_X1 U13236 ( .A1(n13156), .A2(n13256), .ZN(n13254) );
  OR2_X1 U13237 ( .A1(n13158), .A2(n13159), .ZN(n13256) );
  OR2_X1 U13238 ( .A1(n8798), .A2(n8783), .ZN(n13159) );
  OR2_X1 U13239 ( .A1(n13257), .A2(n13258), .ZN(n13158) );
  AND2_X1 U13240 ( .A1(n13155), .A2(n13154), .ZN(n13258) );
  AND2_X1 U13241 ( .A1(n13152), .A2(n13259), .ZN(n13257) );
  OR2_X1 U13242 ( .A1(n13154), .A2(n13155), .ZN(n13259) );
  OR2_X1 U13243 ( .A1(n8802), .A2(n8783), .ZN(n13155) );
  OR2_X1 U13244 ( .A1(n13260), .A2(n13261), .ZN(n13154) );
  AND2_X1 U13245 ( .A1(n13151), .A2(n13150), .ZN(n13261) );
  AND2_X1 U13246 ( .A1(n13148), .A2(n13262), .ZN(n13260) );
  OR2_X1 U13247 ( .A1(n13150), .A2(n13151), .ZN(n13262) );
  OR2_X1 U13248 ( .A1(n8806), .A2(n8783), .ZN(n13151) );
  OR2_X1 U13249 ( .A1(n13263), .A2(n13264), .ZN(n13150) );
  AND2_X1 U13250 ( .A1(n13147), .A2(n13146), .ZN(n13264) );
  AND2_X1 U13251 ( .A1(n13144), .A2(n13265), .ZN(n13263) );
  OR2_X1 U13252 ( .A1(n13146), .A2(n13147), .ZN(n13265) );
  OR2_X1 U13253 ( .A1(n8810), .A2(n8783), .ZN(n13147) );
  OR2_X1 U13254 ( .A1(n13266), .A2(n13267), .ZN(n13146) );
  AND2_X1 U13255 ( .A1(n13143), .A2(n13142), .ZN(n13267) );
  AND2_X1 U13256 ( .A1(n13140), .A2(n13268), .ZN(n13266) );
  OR2_X1 U13257 ( .A1(n13142), .A2(n13143), .ZN(n13268) );
  OR2_X1 U13258 ( .A1(n8140), .A2(n8783), .ZN(n13143) );
  OR2_X1 U13259 ( .A1(n13269), .A2(n13270), .ZN(n13142) );
  AND2_X1 U13260 ( .A1(n13139), .A2(n13138), .ZN(n13270) );
  AND2_X1 U13261 ( .A1(n13136), .A2(n13271), .ZN(n13269) );
  OR2_X1 U13262 ( .A1(n13138), .A2(n13139), .ZN(n13271) );
  OR2_X1 U13263 ( .A1(n8115), .A2(n8783), .ZN(n13139) );
  OR2_X1 U13264 ( .A1(n13272), .A2(n13273), .ZN(n13138) );
  AND2_X1 U13265 ( .A1(n13135), .A2(n13134), .ZN(n13273) );
  AND2_X1 U13266 ( .A1(n13132), .A2(n13274), .ZN(n13272) );
  OR2_X1 U13267 ( .A1(n13134), .A2(n13135), .ZN(n13274) );
  OR2_X1 U13268 ( .A1(n8090), .A2(n8783), .ZN(n13135) );
  OR2_X1 U13269 ( .A1(n13275), .A2(n13276), .ZN(n13134) );
  AND2_X1 U13270 ( .A1(n13131), .A2(n13130), .ZN(n13276) );
  AND2_X1 U13271 ( .A1(n13128), .A2(n13277), .ZN(n13275) );
  OR2_X1 U13272 ( .A1(n13130), .A2(n13131), .ZN(n13277) );
  OR2_X1 U13273 ( .A1(n8065), .A2(n8783), .ZN(n13131) );
  OR2_X1 U13274 ( .A1(n13278), .A2(n13279), .ZN(n13130) );
  AND2_X1 U13275 ( .A1(n13127), .A2(n13126), .ZN(n13279) );
  AND2_X1 U13276 ( .A1(n13124), .A2(n13280), .ZN(n13278) );
  OR2_X1 U13277 ( .A1(n13126), .A2(n13127), .ZN(n13280) );
  OR2_X1 U13278 ( .A1(n8040), .A2(n8783), .ZN(n13127) );
  OR2_X1 U13279 ( .A1(n13281), .A2(n13282), .ZN(n13126) );
  AND2_X1 U13280 ( .A1(n13123), .A2(n13122), .ZN(n13282) );
  AND2_X1 U13281 ( .A1(n13120), .A2(n13283), .ZN(n13281) );
  OR2_X1 U13282 ( .A1(n13122), .A2(n13123), .ZN(n13283) );
  OR2_X1 U13283 ( .A1(n8015), .A2(n8783), .ZN(n13123) );
  OR2_X1 U13284 ( .A1(n13284), .A2(n13285), .ZN(n13122) );
  AND2_X1 U13285 ( .A1(n13119), .A2(n13118), .ZN(n13285) );
  AND2_X1 U13286 ( .A1(n13116), .A2(n13286), .ZN(n13284) );
  OR2_X1 U13287 ( .A1(n13118), .A2(n13119), .ZN(n13286) );
  OR2_X1 U13288 ( .A1(n7979), .A2(n8783), .ZN(n13119) );
  OR2_X1 U13289 ( .A1(n13287), .A2(n13288), .ZN(n13118) );
  AND2_X1 U13290 ( .A1(n13112), .A2(n13115), .ZN(n13288) );
  AND2_X1 U13291 ( .A1(n13289), .A2(n13290), .ZN(n13287) );
  OR2_X1 U13292 ( .A1(n13115), .A2(n13112), .ZN(n13290) );
  OR2_X1 U13293 ( .A1(n7954), .A2(n8783), .ZN(n13112) );
  OR3_X1 U13294 ( .A1(n8783), .A2(n8779), .A3(n9796), .ZN(n13115) );
  INV_X1 U13295 ( .A(n13114), .ZN(n13289) );
  OR2_X1 U13296 ( .A1(n13291), .A2(n13292), .ZN(n13114) );
  AND2_X1 U13297 ( .A1(b_13_), .A2(n13293), .ZN(n13292) );
  OR2_X1 U13298 ( .A1(n13294), .A2(n9801), .ZN(n13293) );
  AND2_X1 U13299 ( .A1(a_30_), .A2(n8775), .ZN(n13294) );
  AND2_X1 U13300 ( .A1(b_12_), .A2(n13295), .ZN(n13291) );
  OR2_X1 U13301 ( .A1(n13296), .A2(n7920), .ZN(n13295) );
  AND2_X1 U13302 ( .A1(a_31_), .A2(n8779), .ZN(n13296) );
  XNOR2_X1 U13303 ( .A(n13297), .B(n13298), .ZN(n13116) );
  XOR2_X1 U13304 ( .A(n13299), .B(n13300), .Z(n13298) );
  XOR2_X1 U13305 ( .A(n13301), .B(n13302), .Z(n13120) );
  XOR2_X1 U13306 ( .A(n13303), .B(n13304), .Z(n13302) );
  XOR2_X1 U13307 ( .A(n13305), .B(n13306), .Z(n13124) );
  XOR2_X1 U13308 ( .A(n13307), .B(n13308), .Z(n13306) );
  XOR2_X1 U13309 ( .A(n13309), .B(n13310), .Z(n13128) );
  XOR2_X1 U13310 ( .A(n13311), .B(n13312), .Z(n13310) );
  XOR2_X1 U13311 ( .A(n13313), .B(n13314), .Z(n13132) );
  XOR2_X1 U13312 ( .A(n13315), .B(n13316), .Z(n13314) );
  XOR2_X1 U13313 ( .A(n13317), .B(n13318), .Z(n13136) );
  XOR2_X1 U13314 ( .A(n13319), .B(n13320), .Z(n13318) );
  XOR2_X1 U13315 ( .A(n13321), .B(n13322), .Z(n13140) );
  XOR2_X1 U13316 ( .A(n13323), .B(n13324), .Z(n13322) );
  XOR2_X1 U13317 ( .A(n13325), .B(n13326), .Z(n13144) );
  XOR2_X1 U13318 ( .A(n13327), .B(n13328), .Z(n13326) );
  XOR2_X1 U13319 ( .A(n13329), .B(n13330), .Z(n13148) );
  XOR2_X1 U13320 ( .A(n13331), .B(n13332), .Z(n13330) );
  XOR2_X1 U13321 ( .A(n13333), .B(n13334), .Z(n13152) );
  XOR2_X1 U13322 ( .A(n13335), .B(n13336), .Z(n13334) );
  XOR2_X1 U13323 ( .A(n13337), .B(n13338), .Z(n13156) );
  XOR2_X1 U13324 ( .A(n13339), .B(n13340), .Z(n13338) );
  XOR2_X1 U13325 ( .A(n13341), .B(n13342), .Z(n13160) );
  XOR2_X1 U13326 ( .A(n13343), .B(n13344), .Z(n13342) );
  XOR2_X1 U13327 ( .A(n13345), .B(n13346), .Z(n13164) );
  XOR2_X1 U13328 ( .A(n13347), .B(n13348), .Z(n13346) );
  XOR2_X1 U13329 ( .A(n13349), .B(n13350), .Z(n13168) );
  XOR2_X1 U13330 ( .A(n13351), .B(n13352), .Z(n13350) );
  XOR2_X1 U13331 ( .A(n13353), .B(n13354), .Z(n13172) );
  XOR2_X1 U13332 ( .A(n13355), .B(n13356), .Z(n13354) );
  XOR2_X1 U13333 ( .A(n13357), .B(n13358), .Z(n13175) );
  XOR2_X1 U13334 ( .A(n13359), .B(n13360), .Z(n13358) );
  XOR2_X1 U13335 ( .A(n13361), .B(n13362), .Z(n13179) );
  XOR2_X1 U13336 ( .A(n13363), .B(n8374), .Z(n13362) );
  XOR2_X1 U13337 ( .A(n13364), .B(n13365), .Z(n13183) );
  XOR2_X1 U13338 ( .A(n13366), .B(n13367), .Z(n13365) );
  XOR2_X1 U13339 ( .A(n13368), .B(n13369), .Z(n13187) );
  XOR2_X1 U13340 ( .A(n13370), .B(n13371), .Z(n13369) );
  XOR2_X1 U13341 ( .A(n13372), .B(n13373), .Z(n13191) );
  XOR2_X1 U13342 ( .A(n13374), .B(n13375), .Z(n13373) );
  XOR2_X1 U13343 ( .A(n13376), .B(n13377), .Z(n13195) );
  XOR2_X1 U13344 ( .A(n13378), .B(n13379), .Z(n13377) );
  XOR2_X1 U13345 ( .A(n13380), .B(n13381), .Z(n11737) );
  XOR2_X1 U13346 ( .A(n13382), .B(n13383), .Z(n13381) );
  XOR2_X1 U13347 ( .A(n13384), .B(n13385), .Z(n11684) );
  XOR2_X1 U13348 ( .A(n13386), .B(n13387), .Z(n13385) );
  XOR2_X1 U13349 ( .A(n13388), .B(n13389), .Z(n9625) );
  XOR2_X1 U13350 ( .A(n13390), .B(n13391), .Z(n13389) );
  XOR2_X1 U13351 ( .A(n13392), .B(n13393), .Z(n9573) );
  XOR2_X1 U13352 ( .A(n13394), .B(n13395), .Z(n13393) );
  XOR2_X1 U13353 ( .A(n13396), .B(n13397), .Z(n9528) );
  XOR2_X1 U13354 ( .A(n13398), .B(n13399), .Z(n13397) );
  XOR2_X1 U13355 ( .A(n13400), .B(n13401), .Z(n9490) );
  XOR2_X1 U13356 ( .A(n13402), .B(n13403), .Z(n13401) );
  XOR2_X1 U13357 ( .A(n13404), .B(n13405), .Z(n9459) );
  XOR2_X1 U13358 ( .A(n13406), .B(n13407), .Z(n13405) );
  XOR2_X1 U13359 ( .A(n13408), .B(n13409), .Z(n9435) );
  XOR2_X1 U13360 ( .A(n13410), .B(n13411), .Z(n13409) );
  XNOR2_X1 U13361 ( .A(n13412), .B(n13413), .ZN(n8995) );
  XOR2_X1 U13362 ( .A(n13414), .B(n13415), .Z(n13413) );
  XOR2_X1 U13363 ( .A(n9006), .B(n9005), .Z(n8993) );
  INV_X1 U13364 ( .A(n13416), .ZN(n9005) );
  OR2_X1 U13365 ( .A1(n13417), .A2(n13418), .ZN(n13416) );
  AND2_X1 U13366 ( .A1(n13415), .A2(n13414), .ZN(n13418) );
  AND2_X1 U13367 ( .A1(n13412), .A2(n13419), .ZN(n13417) );
  OR2_X1 U13368 ( .A1(n13414), .A2(n13415), .ZN(n13419) );
  OR2_X1 U13369 ( .A1(n9248), .A2(n8779), .ZN(n13415) );
  OR2_X1 U13370 ( .A1(n13420), .A2(n13421), .ZN(n13414) );
  AND2_X1 U13371 ( .A1(n13411), .A2(n13410), .ZN(n13421) );
  AND2_X1 U13372 ( .A1(n13408), .A2(n13422), .ZN(n13420) );
  OR2_X1 U13373 ( .A1(n13410), .A2(n13411), .ZN(n13422) );
  OR2_X1 U13374 ( .A1(n8730), .A2(n8779), .ZN(n13411) );
  OR2_X1 U13375 ( .A1(n13423), .A2(n13424), .ZN(n13410) );
  AND2_X1 U13376 ( .A1(n13407), .A2(n13406), .ZN(n13424) );
  AND2_X1 U13377 ( .A1(n13404), .A2(n13425), .ZN(n13423) );
  OR2_X1 U13378 ( .A1(n13406), .A2(n13407), .ZN(n13425) );
  OR2_X1 U13379 ( .A1(n8734), .A2(n8779), .ZN(n13407) );
  OR2_X1 U13380 ( .A1(n13426), .A2(n13427), .ZN(n13406) );
  AND2_X1 U13381 ( .A1(n13403), .A2(n13402), .ZN(n13427) );
  AND2_X1 U13382 ( .A1(n13400), .A2(n13428), .ZN(n13426) );
  OR2_X1 U13383 ( .A1(n13402), .A2(n13403), .ZN(n13428) );
  OR2_X1 U13384 ( .A1(n8738), .A2(n8779), .ZN(n13403) );
  OR2_X1 U13385 ( .A1(n13429), .A2(n13430), .ZN(n13402) );
  AND2_X1 U13386 ( .A1(n13399), .A2(n13398), .ZN(n13430) );
  AND2_X1 U13387 ( .A1(n13396), .A2(n13431), .ZN(n13429) );
  OR2_X1 U13388 ( .A1(n13398), .A2(n13399), .ZN(n13431) );
  OR2_X1 U13389 ( .A1(n8742), .A2(n8779), .ZN(n13399) );
  OR2_X1 U13390 ( .A1(n13432), .A2(n13433), .ZN(n13398) );
  AND2_X1 U13391 ( .A1(n13395), .A2(n13394), .ZN(n13433) );
  AND2_X1 U13392 ( .A1(n13392), .A2(n13434), .ZN(n13432) );
  OR2_X1 U13393 ( .A1(n13394), .A2(n13395), .ZN(n13434) );
  OR2_X1 U13394 ( .A1(n8746), .A2(n8779), .ZN(n13395) );
  OR2_X1 U13395 ( .A1(n13435), .A2(n13436), .ZN(n13394) );
  AND2_X1 U13396 ( .A1(n13391), .A2(n13390), .ZN(n13436) );
  AND2_X1 U13397 ( .A1(n13388), .A2(n13437), .ZN(n13435) );
  OR2_X1 U13398 ( .A1(n13390), .A2(n13391), .ZN(n13437) );
  OR2_X1 U13399 ( .A1(n8750), .A2(n8779), .ZN(n13391) );
  OR2_X1 U13400 ( .A1(n13438), .A2(n13439), .ZN(n13390) );
  AND2_X1 U13401 ( .A1(n13387), .A2(n13386), .ZN(n13439) );
  AND2_X1 U13402 ( .A1(n13384), .A2(n13440), .ZN(n13438) );
  OR2_X1 U13403 ( .A1(n13386), .A2(n13387), .ZN(n13440) );
  OR2_X1 U13404 ( .A1(n8754), .A2(n8779), .ZN(n13387) );
  OR2_X1 U13405 ( .A1(n13441), .A2(n13442), .ZN(n13386) );
  AND2_X1 U13406 ( .A1(n13383), .A2(n13382), .ZN(n13442) );
  AND2_X1 U13407 ( .A1(n13380), .A2(n13443), .ZN(n13441) );
  OR2_X1 U13408 ( .A1(n13382), .A2(n13383), .ZN(n13443) );
  OR2_X1 U13409 ( .A1(n8758), .A2(n8779), .ZN(n13383) );
  OR2_X1 U13410 ( .A1(n13444), .A2(n13445), .ZN(n13382) );
  AND2_X1 U13411 ( .A1(n13379), .A2(n13378), .ZN(n13445) );
  AND2_X1 U13412 ( .A1(n13376), .A2(n13446), .ZN(n13444) );
  OR2_X1 U13413 ( .A1(n13378), .A2(n13379), .ZN(n13446) );
  OR2_X1 U13414 ( .A1(n8762), .A2(n8779), .ZN(n13379) );
  OR2_X1 U13415 ( .A1(n13447), .A2(n13448), .ZN(n13378) );
  AND2_X1 U13416 ( .A1(n13375), .A2(n13374), .ZN(n13448) );
  AND2_X1 U13417 ( .A1(n13372), .A2(n13449), .ZN(n13447) );
  OR2_X1 U13418 ( .A1(n13374), .A2(n13375), .ZN(n13449) );
  OR2_X1 U13419 ( .A1(n8766), .A2(n8779), .ZN(n13375) );
  OR2_X1 U13420 ( .A1(n13450), .A2(n13451), .ZN(n13374) );
  AND2_X1 U13421 ( .A1(n13371), .A2(n13370), .ZN(n13451) );
  AND2_X1 U13422 ( .A1(n13368), .A2(n13452), .ZN(n13450) );
  OR2_X1 U13423 ( .A1(n13370), .A2(n13371), .ZN(n13452) );
  OR2_X1 U13424 ( .A1(n8770), .A2(n8779), .ZN(n13371) );
  OR2_X1 U13425 ( .A1(n13453), .A2(n13454), .ZN(n13370) );
  AND2_X1 U13426 ( .A1(n13367), .A2(n13366), .ZN(n13454) );
  AND2_X1 U13427 ( .A1(n13364), .A2(n13455), .ZN(n13453) );
  OR2_X1 U13428 ( .A1(n13366), .A2(n13367), .ZN(n13455) );
  OR2_X1 U13429 ( .A1(n8774), .A2(n8779), .ZN(n13367) );
  OR2_X1 U13430 ( .A1(n13456), .A2(n13457), .ZN(n13366) );
  AND2_X1 U13431 ( .A1(n8374), .A2(n13363), .ZN(n13457) );
  AND2_X1 U13432 ( .A1(n13361), .A2(n13458), .ZN(n13456) );
  OR2_X1 U13433 ( .A1(n13363), .A2(n8374), .ZN(n13458) );
  OR2_X1 U13434 ( .A1(n8778), .A2(n8779), .ZN(n8374) );
  OR2_X1 U13435 ( .A1(n13459), .A2(n13460), .ZN(n13363) );
  AND2_X1 U13436 ( .A1(n13360), .A2(n13359), .ZN(n13460) );
  AND2_X1 U13437 ( .A1(n13357), .A2(n13461), .ZN(n13459) );
  OR2_X1 U13438 ( .A1(n13359), .A2(n13360), .ZN(n13461) );
  OR2_X1 U13439 ( .A1(n8782), .A2(n8779), .ZN(n13360) );
  OR2_X1 U13440 ( .A1(n13462), .A2(n13463), .ZN(n13359) );
  AND2_X1 U13441 ( .A1(n13356), .A2(n13355), .ZN(n13463) );
  AND2_X1 U13442 ( .A1(n13353), .A2(n13464), .ZN(n13462) );
  OR2_X1 U13443 ( .A1(n13355), .A2(n13356), .ZN(n13464) );
  OR2_X1 U13444 ( .A1(n8786), .A2(n8779), .ZN(n13356) );
  OR2_X1 U13445 ( .A1(n13465), .A2(n13466), .ZN(n13355) );
  AND2_X1 U13446 ( .A1(n13352), .A2(n13351), .ZN(n13466) );
  AND2_X1 U13447 ( .A1(n13349), .A2(n13467), .ZN(n13465) );
  OR2_X1 U13448 ( .A1(n13351), .A2(n13352), .ZN(n13467) );
  OR2_X1 U13449 ( .A1(n8790), .A2(n8779), .ZN(n13352) );
  OR2_X1 U13450 ( .A1(n13468), .A2(n13469), .ZN(n13351) );
  AND2_X1 U13451 ( .A1(n13348), .A2(n13347), .ZN(n13469) );
  AND2_X1 U13452 ( .A1(n13345), .A2(n13470), .ZN(n13468) );
  OR2_X1 U13453 ( .A1(n13347), .A2(n13348), .ZN(n13470) );
  OR2_X1 U13454 ( .A1(n8794), .A2(n8779), .ZN(n13348) );
  OR2_X1 U13455 ( .A1(n13471), .A2(n13472), .ZN(n13347) );
  AND2_X1 U13456 ( .A1(n13344), .A2(n13343), .ZN(n13472) );
  AND2_X1 U13457 ( .A1(n13341), .A2(n13473), .ZN(n13471) );
  OR2_X1 U13458 ( .A1(n13343), .A2(n13344), .ZN(n13473) );
  OR2_X1 U13459 ( .A1(n8798), .A2(n8779), .ZN(n13344) );
  OR2_X1 U13460 ( .A1(n13474), .A2(n13475), .ZN(n13343) );
  AND2_X1 U13461 ( .A1(n13340), .A2(n13339), .ZN(n13475) );
  AND2_X1 U13462 ( .A1(n13337), .A2(n13476), .ZN(n13474) );
  OR2_X1 U13463 ( .A1(n13339), .A2(n13340), .ZN(n13476) );
  OR2_X1 U13464 ( .A1(n8802), .A2(n8779), .ZN(n13340) );
  OR2_X1 U13465 ( .A1(n13477), .A2(n13478), .ZN(n13339) );
  AND2_X1 U13466 ( .A1(n13336), .A2(n13335), .ZN(n13478) );
  AND2_X1 U13467 ( .A1(n13333), .A2(n13479), .ZN(n13477) );
  OR2_X1 U13468 ( .A1(n13335), .A2(n13336), .ZN(n13479) );
  OR2_X1 U13469 ( .A1(n8806), .A2(n8779), .ZN(n13336) );
  OR2_X1 U13470 ( .A1(n13480), .A2(n13481), .ZN(n13335) );
  AND2_X1 U13471 ( .A1(n13332), .A2(n13331), .ZN(n13481) );
  AND2_X1 U13472 ( .A1(n13329), .A2(n13482), .ZN(n13480) );
  OR2_X1 U13473 ( .A1(n13331), .A2(n13332), .ZN(n13482) );
  OR2_X1 U13474 ( .A1(n8810), .A2(n8779), .ZN(n13332) );
  OR2_X1 U13475 ( .A1(n13483), .A2(n13484), .ZN(n13331) );
  AND2_X1 U13476 ( .A1(n13328), .A2(n13327), .ZN(n13484) );
  AND2_X1 U13477 ( .A1(n13325), .A2(n13485), .ZN(n13483) );
  OR2_X1 U13478 ( .A1(n13327), .A2(n13328), .ZN(n13485) );
  OR2_X1 U13479 ( .A1(n8140), .A2(n8779), .ZN(n13328) );
  OR2_X1 U13480 ( .A1(n13486), .A2(n13487), .ZN(n13327) );
  AND2_X1 U13481 ( .A1(n13324), .A2(n13323), .ZN(n13487) );
  AND2_X1 U13482 ( .A1(n13321), .A2(n13488), .ZN(n13486) );
  OR2_X1 U13483 ( .A1(n13323), .A2(n13324), .ZN(n13488) );
  OR2_X1 U13484 ( .A1(n8115), .A2(n8779), .ZN(n13324) );
  OR2_X1 U13485 ( .A1(n13489), .A2(n13490), .ZN(n13323) );
  AND2_X1 U13486 ( .A1(n13320), .A2(n13319), .ZN(n13490) );
  AND2_X1 U13487 ( .A1(n13317), .A2(n13491), .ZN(n13489) );
  OR2_X1 U13488 ( .A1(n13319), .A2(n13320), .ZN(n13491) );
  OR2_X1 U13489 ( .A1(n8090), .A2(n8779), .ZN(n13320) );
  OR2_X1 U13490 ( .A1(n13492), .A2(n13493), .ZN(n13319) );
  AND2_X1 U13491 ( .A1(n13316), .A2(n13315), .ZN(n13493) );
  AND2_X1 U13492 ( .A1(n13313), .A2(n13494), .ZN(n13492) );
  OR2_X1 U13493 ( .A1(n13315), .A2(n13316), .ZN(n13494) );
  OR2_X1 U13494 ( .A1(n8065), .A2(n8779), .ZN(n13316) );
  OR2_X1 U13495 ( .A1(n13495), .A2(n13496), .ZN(n13315) );
  AND2_X1 U13496 ( .A1(n13312), .A2(n13311), .ZN(n13496) );
  AND2_X1 U13497 ( .A1(n13309), .A2(n13497), .ZN(n13495) );
  OR2_X1 U13498 ( .A1(n13311), .A2(n13312), .ZN(n13497) );
  OR2_X1 U13499 ( .A1(n8040), .A2(n8779), .ZN(n13312) );
  OR2_X1 U13500 ( .A1(n13498), .A2(n13499), .ZN(n13311) );
  AND2_X1 U13501 ( .A1(n13308), .A2(n13307), .ZN(n13499) );
  AND2_X1 U13502 ( .A1(n13305), .A2(n13500), .ZN(n13498) );
  OR2_X1 U13503 ( .A1(n13307), .A2(n13308), .ZN(n13500) );
  OR2_X1 U13504 ( .A1(n8015), .A2(n8779), .ZN(n13308) );
  OR2_X1 U13505 ( .A1(n13501), .A2(n13502), .ZN(n13307) );
  AND2_X1 U13506 ( .A1(n13304), .A2(n13303), .ZN(n13502) );
  AND2_X1 U13507 ( .A1(n13301), .A2(n13503), .ZN(n13501) );
  OR2_X1 U13508 ( .A1(n13303), .A2(n13304), .ZN(n13503) );
  OR2_X1 U13509 ( .A1(n7979), .A2(n8779), .ZN(n13304) );
  OR2_X1 U13510 ( .A1(n13504), .A2(n13505), .ZN(n13303) );
  AND2_X1 U13511 ( .A1(n13297), .A2(n13300), .ZN(n13505) );
  AND2_X1 U13512 ( .A1(n13506), .A2(n13507), .ZN(n13504) );
  OR2_X1 U13513 ( .A1(n13300), .A2(n13297), .ZN(n13507) );
  OR2_X1 U13514 ( .A1(n7954), .A2(n8779), .ZN(n13297) );
  OR3_X1 U13515 ( .A1(n8779), .A2(n8775), .A3(n9796), .ZN(n13300) );
  INV_X1 U13516 ( .A(n13299), .ZN(n13506) );
  OR2_X1 U13517 ( .A1(n13508), .A2(n13509), .ZN(n13299) );
  AND2_X1 U13518 ( .A1(b_12_), .A2(n13510), .ZN(n13509) );
  OR2_X1 U13519 ( .A1(n13511), .A2(n9801), .ZN(n13510) );
  AND2_X1 U13520 ( .A1(a_30_), .A2(n8771), .ZN(n13511) );
  AND2_X1 U13521 ( .A1(b_11_), .A2(n13512), .ZN(n13508) );
  OR2_X1 U13522 ( .A1(n13513), .A2(n7920), .ZN(n13512) );
  AND2_X1 U13523 ( .A1(a_31_), .A2(n8775), .ZN(n13513) );
  XNOR2_X1 U13524 ( .A(n13514), .B(n13515), .ZN(n13301) );
  XOR2_X1 U13525 ( .A(n13516), .B(n13517), .Z(n13515) );
  XOR2_X1 U13526 ( .A(n13518), .B(n13519), .Z(n13305) );
  XOR2_X1 U13527 ( .A(n13520), .B(n13521), .Z(n13519) );
  XOR2_X1 U13528 ( .A(n13522), .B(n13523), .Z(n13309) );
  XOR2_X1 U13529 ( .A(n13524), .B(n13525), .Z(n13523) );
  XOR2_X1 U13530 ( .A(n13526), .B(n13527), .Z(n13313) );
  XOR2_X1 U13531 ( .A(n13528), .B(n13529), .Z(n13527) );
  XOR2_X1 U13532 ( .A(n13530), .B(n13531), .Z(n13317) );
  XOR2_X1 U13533 ( .A(n13532), .B(n13533), .Z(n13531) );
  XOR2_X1 U13534 ( .A(n13534), .B(n13535), .Z(n13321) );
  XOR2_X1 U13535 ( .A(n13536), .B(n13537), .Z(n13535) );
  XOR2_X1 U13536 ( .A(n13538), .B(n13539), .Z(n13325) );
  XOR2_X1 U13537 ( .A(n13540), .B(n13541), .Z(n13539) );
  XOR2_X1 U13538 ( .A(n13542), .B(n13543), .Z(n13329) );
  XOR2_X1 U13539 ( .A(n13544), .B(n13545), .Z(n13543) );
  XOR2_X1 U13540 ( .A(n13546), .B(n13547), .Z(n13333) );
  XOR2_X1 U13541 ( .A(n13548), .B(n13549), .Z(n13547) );
  XOR2_X1 U13542 ( .A(n13550), .B(n13551), .Z(n13337) );
  XOR2_X1 U13543 ( .A(n13552), .B(n13553), .Z(n13551) );
  XOR2_X1 U13544 ( .A(n13554), .B(n13555), .Z(n13341) );
  XOR2_X1 U13545 ( .A(n13556), .B(n13557), .Z(n13555) );
  XOR2_X1 U13546 ( .A(n13558), .B(n13559), .Z(n13345) );
  XOR2_X1 U13547 ( .A(n13560), .B(n13561), .Z(n13559) );
  XOR2_X1 U13548 ( .A(n13562), .B(n13563), .Z(n13349) );
  XOR2_X1 U13549 ( .A(n13564), .B(n13565), .Z(n13563) );
  XOR2_X1 U13550 ( .A(n13566), .B(n13567), .Z(n13353) );
  XOR2_X1 U13551 ( .A(n13568), .B(n13569), .Z(n13567) );
  XOR2_X1 U13552 ( .A(n13570), .B(n13571), .Z(n13357) );
  XOR2_X1 U13553 ( .A(n13572), .B(n13573), .Z(n13571) );
  XOR2_X1 U13554 ( .A(n13574), .B(n13575), .Z(n13361) );
  XOR2_X1 U13555 ( .A(n13576), .B(n13577), .Z(n13575) );
  XOR2_X1 U13556 ( .A(n13578), .B(n13579), .Z(n13364) );
  XOR2_X1 U13557 ( .A(n13580), .B(n13581), .Z(n13579) );
  XOR2_X1 U13558 ( .A(n13582), .B(n13583), .Z(n13368) );
  XOR2_X1 U13559 ( .A(n13584), .B(n8400), .Z(n13583) );
  XOR2_X1 U13560 ( .A(n13585), .B(n13586), .Z(n13372) );
  XOR2_X1 U13561 ( .A(n13587), .B(n13588), .Z(n13586) );
  XOR2_X1 U13562 ( .A(n13589), .B(n13590), .Z(n13376) );
  XOR2_X1 U13563 ( .A(n13591), .B(n13592), .Z(n13590) );
  XOR2_X1 U13564 ( .A(n13593), .B(n13594), .Z(n13380) );
  XOR2_X1 U13565 ( .A(n13595), .B(n13596), .Z(n13594) );
  XOR2_X1 U13566 ( .A(n13597), .B(n13598), .Z(n13384) );
  XOR2_X1 U13567 ( .A(n13599), .B(n13600), .Z(n13598) );
  XOR2_X1 U13568 ( .A(n13601), .B(n13602), .Z(n13388) );
  XOR2_X1 U13569 ( .A(n13603), .B(n13604), .Z(n13602) );
  XOR2_X1 U13570 ( .A(n13605), .B(n13606), .Z(n13392) );
  XOR2_X1 U13571 ( .A(n13607), .B(n13608), .Z(n13606) );
  XOR2_X1 U13572 ( .A(n13609), .B(n13610), .Z(n13396) );
  XOR2_X1 U13573 ( .A(n13611), .B(n13612), .Z(n13610) );
  XOR2_X1 U13574 ( .A(n13613), .B(n13614), .Z(n13400) );
  XOR2_X1 U13575 ( .A(n13615), .B(n13616), .Z(n13614) );
  XOR2_X1 U13576 ( .A(n13617), .B(n13618), .Z(n13404) );
  XOR2_X1 U13577 ( .A(n13619), .B(n13620), .Z(n13618) );
  XOR2_X1 U13578 ( .A(n13621), .B(n13622), .Z(n13408) );
  XOR2_X1 U13579 ( .A(n13623), .B(n13624), .Z(n13622) );
  XOR2_X1 U13580 ( .A(n13625), .B(n13626), .Z(n13412) );
  XOR2_X1 U13581 ( .A(n13627), .B(n13628), .Z(n13626) );
  XNOR2_X1 U13582 ( .A(n13629), .B(n13630), .ZN(n9006) );
  XOR2_X1 U13583 ( .A(n13631), .B(n13632), .Z(n13630) );
  XOR2_X1 U13584 ( .A(n9017), .B(n9016), .Z(n9004) );
  INV_X1 U13585 ( .A(n13633), .ZN(n9016) );
  OR2_X1 U13586 ( .A1(n13634), .A2(n13635), .ZN(n13633) );
  AND2_X1 U13587 ( .A1(n13632), .A2(n13631), .ZN(n13635) );
  AND2_X1 U13588 ( .A1(n13629), .A2(n13636), .ZN(n13634) );
  OR2_X1 U13589 ( .A1(n13631), .A2(n13632), .ZN(n13636) );
  OR2_X1 U13590 ( .A1(n9248), .A2(n8775), .ZN(n13632) );
  OR2_X1 U13591 ( .A1(n13637), .A2(n13638), .ZN(n13631) );
  AND2_X1 U13592 ( .A1(n13628), .A2(n13627), .ZN(n13638) );
  AND2_X1 U13593 ( .A1(n13625), .A2(n13639), .ZN(n13637) );
  OR2_X1 U13594 ( .A1(n13627), .A2(n13628), .ZN(n13639) );
  OR2_X1 U13595 ( .A1(n8730), .A2(n8775), .ZN(n13628) );
  OR2_X1 U13596 ( .A1(n13640), .A2(n13641), .ZN(n13627) );
  AND2_X1 U13597 ( .A1(n13624), .A2(n13623), .ZN(n13641) );
  AND2_X1 U13598 ( .A1(n13621), .A2(n13642), .ZN(n13640) );
  OR2_X1 U13599 ( .A1(n13623), .A2(n13624), .ZN(n13642) );
  OR2_X1 U13600 ( .A1(n8734), .A2(n8775), .ZN(n13624) );
  OR2_X1 U13601 ( .A1(n13643), .A2(n13644), .ZN(n13623) );
  AND2_X1 U13602 ( .A1(n13620), .A2(n13619), .ZN(n13644) );
  AND2_X1 U13603 ( .A1(n13617), .A2(n13645), .ZN(n13643) );
  OR2_X1 U13604 ( .A1(n13619), .A2(n13620), .ZN(n13645) );
  OR2_X1 U13605 ( .A1(n8738), .A2(n8775), .ZN(n13620) );
  OR2_X1 U13606 ( .A1(n13646), .A2(n13647), .ZN(n13619) );
  AND2_X1 U13607 ( .A1(n13616), .A2(n13615), .ZN(n13647) );
  AND2_X1 U13608 ( .A1(n13613), .A2(n13648), .ZN(n13646) );
  OR2_X1 U13609 ( .A1(n13615), .A2(n13616), .ZN(n13648) );
  OR2_X1 U13610 ( .A1(n8742), .A2(n8775), .ZN(n13616) );
  OR2_X1 U13611 ( .A1(n13649), .A2(n13650), .ZN(n13615) );
  AND2_X1 U13612 ( .A1(n13612), .A2(n13611), .ZN(n13650) );
  AND2_X1 U13613 ( .A1(n13609), .A2(n13651), .ZN(n13649) );
  OR2_X1 U13614 ( .A1(n13611), .A2(n13612), .ZN(n13651) );
  OR2_X1 U13615 ( .A1(n8746), .A2(n8775), .ZN(n13612) );
  OR2_X1 U13616 ( .A1(n13652), .A2(n13653), .ZN(n13611) );
  AND2_X1 U13617 ( .A1(n13608), .A2(n13607), .ZN(n13653) );
  AND2_X1 U13618 ( .A1(n13605), .A2(n13654), .ZN(n13652) );
  OR2_X1 U13619 ( .A1(n13607), .A2(n13608), .ZN(n13654) );
  OR2_X1 U13620 ( .A1(n8750), .A2(n8775), .ZN(n13608) );
  OR2_X1 U13621 ( .A1(n13655), .A2(n13656), .ZN(n13607) );
  AND2_X1 U13622 ( .A1(n13604), .A2(n13603), .ZN(n13656) );
  AND2_X1 U13623 ( .A1(n13601), .A2(n13657), .ZN(n13655) );
  OR2_X1 U13624 ( .A1(n13603), .A2(n13604), .ZN(n13657) );
  OR2_X1 U13625 ( .A1(n8754), .A2(n8775), .ZN(n13604) );
  OR2_X1 U13626 ( .A1(n13658), .A2(n13659), .ZN(n13603) );
  AND2_X1 U13627 ( .A1(n13600), .A2(n13599), .ZN(n13659) );
  AND2_X1 U13628 ( .A1(n13597), .A2(n13660), .ZN(n13658) );
  OR2_X1 U13629 ( .A1(n13599), .A2(n13600), .ZN(n13660) );
  OR2_X1 U13630 ( .A1(n8758), .A2(n8775), .ZN(n13600) );
  OR2_X1 U13631 ( .A1(n13661), .A2(n13662), .ZN(n13599) );
  AND2_X1 U13632 ( .A1(n13596), .A2(n13595), .ZN(n13662) );
  AND2_X1 U13633 ( .A1(n13593), .A2(n13663), .ZN(n13661) );
  OR2_X1 U13634 ( .A1(n13595), .A2(n13596), .ZN(n13663) );
  OR2_X1 U13635 ( .A1(n8762), .A2(n8775), .ZN(n13596) );
  OR2_X1 U13636 ( .A1(n13664), .A2(n13665), .ZN(n13595) );
  AND2_X1 U13637 ( .A1(n13592), .A2(n13591), .ZN(n13665) );
  AND2_X1 U13638 ( .A1(n13589), .A2(n13666), .ZN(n13664) );
  OR2_X1 U13639 ( .A1(n13591), .A2(n13592), .ZN(n13666) );
  OR2_X1 U13640 ( .A1(n8766), .A2(n8775), .ZN(n13592) );
  OR2_X1 U13641 ( .A1(n13667), .A2(n13668), .ZN(n13591) );
  AND2_X1 U13642 ( .A1(n13588), .A2(n13587), .ZN(n13668) );
  AND2_X1 U13643 ( .A1(n13585), .A2(n13669), .ZN(n13667) );
  OR2_X1 U13644 ( .A1(n13587), .A2(n13588), .ZN(n13669) );
  OR2_X1 U13645 ( .A1(n8770), .A2(n8775), .ZN(n13588) );
  OR2_X1 U13646 ( .A1(n13670), .A2(n13671), .ZN(n13587) );
  AND2_X1 U13647 ( .A1(n8400), .A2(n13584), .ZN(n13671) );
  AND2_X1 U13648 ( .A1(n13582), .A2(n13672), .ZN(n13670) );
  OR2_X1 U13649 ( .A1(n13584), .A2(n8400), .ZN(n13672) );
  OR2_X1 U13650 ( .A1(n8774), .A2(n8775), .ZN(n8400) );
  OR2_X1 U13651 ( .A1(n13673), .A2(n13674), .ZN(n13584) );
  AND2_X1 U13652 ( .A1(n13581), .A2(n13580), .ZN(n13674) );
  AND2_X1 U13653 ( .A1(n13578), .A2(n13675), .ZN(n13673) );
  OR2_X1 U13654 ( .A1(n13580), .A2(n13581), .ZN(n13675) );
  OR2_X1 U13655 ( .A1(n8778), .A2(n8775), .ZN(n13581) );
  OR2_X1 U13656 ( .A1(n13676), .A2(n13677), .ZN(n13580) );
  AND2_X1 U13657 ( .A1(n13577), .A2(n13576), .ZN(n13677) );
  AND2_X1 U13658 ( .A1(n13574), .A2(n13678), .ZN(n13676) );
  OR2_X1 U13659 ( .A1(n13576), .A2(n13577), .ZN(n13678) );
  OR2_X1 U13660 ( .A1(n8782), .A2(n8775), .ZN(n13577) );
  OR2_X1 U13661 ( .A1(n13679), .A2(n13680), .ZN(n13576) );
  AND2_X1 U13662 ( .A1(n13573), .A2(n13572), .ZN(n13680) );
  AND2_X1 U13663 ( .A1(n13570), .A2(n13681), .ZN(n13679) );
  OR2_X1 U13664 ( .A1(n13572), .A2(n13573), .ZN(n13681) );
  OR2_X1 U13665 ( .A1(n8786), .A2(n8775), .ZN(n13573) );
  OR2_X1 U13666 ( .A1(n13682), .A2(n13683), .ZN(n13572) );
  AND2_X1 U13667 ( .A1(n13569), .A2(n13568), .ZN(n13683) );
  AND2_X1 U13668 ( .A1(n13566), .A2(n13684), .ZN(n13682) );
  OR2_X1 U13669 ( .A1(n13568), .A2(n13569), .ZN(n13684) );
  OR2_X1 U13670 ( .A1(n8790), .A2(n8775), .ZN(n13569) );
  OR2_X1 U13671 ( .A1(n13685), .A2(n13686), .ZN(n13568) );
  AND2_X1 U13672 ( .A1(n13565), .A2(n13564), .ZN(n13686) );
  AND2_X1 U13673 ( .A1(n13562), .A2(n13687), .ZN(n13685) );
  OR2_X1 U13674 ( .A1(n13564), .A2(n13565), .ZN(n13687) );
  OR2_X1 U13675 ( .A1(n8794), .A2(n8775), .ZN(n13565) );
  OR2_X1 U13676 ( .A1(n13688), .A2(n13689), .ZN(n13564) );
  AND2_X1 U13677 ( .A1(n13561), .A2(n13560), .ZN(n13689) );
  AND2_X1 U13678 ( .A1(n13558), .A2(n13690), .ZN(n13688) );
  OR2_X1 U13679 ( .A1(n13560), .A2(n13561), .ZN(n13690) );
  OR2_X1 U13680 ( .A1(n8798), .A2(n8775), .ZN(n13561) );
  OR2_X1 U13681 ( .A1(n13691), .A2(n13692), .ZN(n13560) );
  AND2_X1 U13682 ( .A1(n13557), .A2(n13556), .ZN(n13692) );
  AND2_X1 U13683 ( .A1(n13554), .A2(n13693), .ZN(n13691) );
  OR2_X1 U13684 ( .A1(n13556), .A2(n13557), .ZN(n13693) );
  OR2_X1 U13685 ( .A1(n8802), .A2(n8775), .ZN(n13557) );
  OR2_X1 U13686 ( .A1(n13694), .A2(n13695), .ZN(n13556) );
  AND2_X1 U13687 ( .A1(n13553), .A2(n13552), .ZN(n13695) );
  AND2_X1 U13688 ( .A1(n13550), .A2(n13696), .ZN(n13694) );
  OR2_X1 U13689 ( .A1(n13552), .A2(n13553), .ZN(n13696) );
  OR2_X1 U13690 ( .A1(n8806), .A2(n8775), .ZN(n13553) );
  OR2_X1 U13691 ( .A1(n13697), .A2(n13698), .ZN(n13552) );
  AND2_X1 U13692 ( .A1(n13549), .A2(n13548), .ZN(n13698) );
  AND2_X1 U13693 ( .A1(n13546), .A2(n13699), .ZN(n13697) );
  OR2_X1 U13694 ( .A1(n13548), .A2(n13549), .ZN(n13699) );
  OR2_X1 U13695 ( .A1(n8810), .A2(n8775), .ZN(n13549) );
  OR2_X1 U13696 ( .A1(n13700), .A2(n13701), .ZN(n13548) );
  AND2_X1 U13697 ( .A1(n13545), .A2(n13544), .ZN(n13701) );
  AND2_X1 U13698 ( .A1(n13542), .A2(n13702), .ZN(n13700) );
  OR2_X1 U13699 ( .A1(n13544), .A2(n13545), .ZN(n13702) );
  OR2_X1 U13700 ( .A1(n8140), .A2(n8775), .ZN(n13545) );
  OR2_X1 U13701 ( .A1(n13703), .A2(n13704), .ZN(n13544) );
  AND2_X1 U13702 ( .A1(n13541), .A2(n13540), .ZN(n13704) );
  AND2_X1 U13703 ( .A1(n13538), .A2(n13705), .ZN(n13703) );
  OR2_X1 U13704 ( .A1(n13540), .A2(n13541), .ZN(n13705) );
  OR2_X1 U13705 ( .A1(n8115), .A2(n8775), .ZN(n13541) );
  OR2_X1 U13706 ( .A1(n13706), .A2(n13707), .ZN(n13540) );
  AND2_X1 U13707 ( .A1(n13537), .A2(n13536), .ZN(n13707) );
  AND2_X1 U13708 ( .A1(n13534), .A2(n13708), .ZN(n13706) );
  OR2_X1 U13709 ( .A1(n13536), .A2(n13537), .ZN(n13708) );
  OR2_X1 U13710 ( .A1(n8090), .A2(n8775), .ZN(n13537) );
  OR2_X1 U13711 ( .A1(n13709), .A2(n13710), .ZN(n13536) );
  AND2_X1 U13712 ( .A1(n13533), .A2(n13532), .ZN(n13710) );
  AND2_X1 U13713 ( .A1(n13530), .A2(n13711), .ZN(n13709) );
  OR2_X1 U13714 ( .A1(n13532), .A2(n13533), .ZN(n13711) );
  OR2_X1 U13715 ( .A1(n8065), .A2(n8775), .ZN(n13533) );
  OR2_X1 U13716 ( .A1(n13712), .A2(n13713), .ZN(n13532) );
  AND2_X1 U13717 ( .A1(n13529), .A2(n13528), .ZN(n13713) );
  AND2_X1 U13718 ( .A1(n13526), .A2(n13714), .ZN(n13712) );
  OR2_X1 U13719 ( .A1(n13528), .A2(n13529), .ZN(n13714) );
  OR2_X1 U13720 ( .A1(n8040), .A2(n8775), .ZN(n13529) );
  OR2_X1 U13721 ( .A1(n13715), .A2(n13716), .ZN(n13528) );
  AND2_X1 U13722 ( .A1(n13525), .A2(n13524), .ZN(n13716) );
  AND2_X1 U13723 ( .A1(n13522), .A2(n13717), .ZN(n13715) );
  OR2_X1 U13724 ( .A1(n13524), .A2(n13525), .ZN(n13717) );
  OR2_X1 U13725 ( .A1(n8015), .A2(n8775), .ZN(n13525) );
  OR2_X1 U13726 ( .A1(n13718), .A2(n13719), .ZN(n13524) );
  AND2_X1 U13727 ( .A1(n13521), .A2(n13520), .ZN(n13719) );
  AND2_X1 U13728 ( .A1(n13518), .A2(n13720), .ZN(n13718) );
  OR2_X1 U13729 ( .A1(n13520), .A2(n13521), .ZN(n13720) );
  OR2_X1 U13730 ( .A1(n7979), .A2(n8775), .ZN(n13521) );
  OR2_X1 U13731 ( .A1(n13721), .A2(n13722), .ZN(n13520) );
  AND2_X1 U13732 ( .A1(n13514), .A2(n13517), .ZN(n13722) );
  AND2_X1 U13733 ( .A1(n13723), .A2(n13724), .ZN(n13721) );
  OR2_X1 U13734 ( .A1(n13517), .A2(n13514), .ZN(n13724) );
  OR2_X1 U13735 ( .A1(n7954), .A2(n8775), .ZN(n13514) );
  OR3_X1 U13736 ( .A1(n8775), .A2(n8771), .A3(n9796), .ZN(n13517) );
  INV_X1 U13737 ( .A(n13516), .ZN(n13723) );
  OR2_X1 U13738 ( .A1(n13725), .A2(n13726), .ZN(n13516) );
  AND2_X1 U13739 ( .A1(b_11_), .A2(n13727), .ZN(n13726) );
  OR2_X1 U13740 ( .A1(n13728), .A2(n9801), .ZN(n13727) );
  AND2_X1 U13741 ( .A1(a_30_), .A2(n8767), .ZN(n13728) );
  AND2_X1 U13742 ( .A1(b_10_), .A2(n13729), .ZN(n13725) );
  OR2_X1 U13743 ( .A1(n13730), .A2(n7920), .ZN(n13729) );
  AND2_X1 U13744 ( .A1(a_31_), .A2(n8771), .ZN(n13730) );
  XNOR2_X1 U13745 ( .A(n13731), .B(n13732), .ZN(n13518) );
  XOR2_X1 U13746 ( .A(n13733), .B(n13734), .Z(n13732) );
  XOR2_X1 U13747 ( .A(n13735), .B(n13736), .Z(n13522) );
  XOR2_X1 U13748 ( .A(n13737), .B(n13738), .Z(n13736) );
  XOR2_X1 U13749 ( .A(n13739), .B(n13740), .Z(n13526) );
  XOR2_X1 U13750 ( .A(n13741), .B(n13742), .Z(n13740) );
  XOR2_X1 U13751 ( .A(n13743), .B(n13744), .Z(n13530) );
  XOR2_X1 U13752 ( .A(n13745), .B(n13746), .Z(n13744) );
  XOR2_X1 U13753 ( .A(n13747), .B(n13748), .Z(n13534) );
  XOR2_X1 U13754 ( .A(n13749), .B(n13750), .Z(n13748) );
  XOR2_X1 U13755 ( .A(n13751), .B(n13752), .Z(n13538) );
  XOR2_X1 U13756 ( .A(n13753), .B(n13754), .Z(n13752) );
  XOR2_X1 U13757 ( .A(n13755), .B(n13756), .Z(n13542) );
  XOR2_X1 U13758 ( .A(n13757), .B(n13758), .Z(n13756) );
  XOR2_X1 U13759 ( .A(n13759), .B(n13760), .Z(n13546) );
  XOR2_X1 U13760 ( .A(n13761), .B(n13762), .Z(n13760) );
  XOR2_X1 U13761 ( .A(n13763), .B(n13764), .Z(n13550) );
  XOR2_X1 U13762 ( .A(n13765), .B(n13766), .Z(n13764) );
  XOR2_X1 U13763 ( .A(n13767), .B(n13768), .Z(n13554) );
  XOR2_X1 U13764 ( .A(n13769), .B(n13770), .Z(n13768) );
  XOR2_X1 U13765 ( .A(n13771), .B(n13772), .Z(n13558) );
  XOR2_X1 U13766 ( .A(n13773), .B(n13774), .Z(n13772) );
  XOR2_X1 U13767 ( .A(n13775), .B(n13776), .Z(n13562) );
  XOR2_X1 U13768 ( .A(n13777), .B(n13778), .Z(n13776) );
  XOR2_X1 U13769 ( .A(n13779), .B(n13780), .Z(n13566) );
  XOR2_X1 U13770 ( .A(n13781), .B(n13782), .Z(n13780) );
  XOR2_X1 U13771 ( .A(n13783), .B(n13784), .Z(n13570) );
  XOR2_X1 U13772 ( .A(n13785), .B(n13786), .Z(n13784) );
  XOR2_X1 U13773 ( .A(n13787), .B(n13788), .Z(n13574) );
  XOR2_X1 U13774 ( .A(n13789), .B(n13790), .Z(n13788) );
  XOR2_X1 U13775 ( .A(n13791), .B(n13792), .Z(n13578) );
  XOR2_X1 U13776 ( .A(n13793), .B(n13794), .Z(n13792) );
  XOR2_X1 U13777 ( .A(n13795), .B(n13796), .Z(n13582) );
  XOR2_X1 U13778 ( .A(n13797), .B(n13798), .Z(n13796) );
  XOR2_X1 U13779 ( .A(n13799), .B(n13800), .Z(n13585) );
  XOR2_X1 U13780 ( .A(n13801), .B(n13802), .Z(n13800) );
  XOR2_X1 U13781 ( .A(n13803), .B(n13804), .Z(n13589) );
  XOR2_X1 U13782 ( .A(n13805), .B(n8426), .Z(n13804) );
  XOR2_X1 U13783 ( .A(n13806), .B(n13807), .Z(n13593) );
  XOR2_X1 U13784 ( .A(n13808), .B(n13809), .Z(n13807) );
  XOR2_X1 U13785 ( .A(n13810), .B(n13811), .Z(n13597) );
  XOR2_X1 U13786 ( .A(n13812), .B(n13813), .Z(n13811) );
  XOR2_X1 U13787 ( .A(n13814), .B(n13815), .Z(n13601) );
  XOR2_X1 U13788 ( .A(n13816), .B(n13817), .Z(n13815) );
  XOR2_X1 U13789 ( .A(n13818), .B(n13819), .Z(n13605) );
  XOR2_X1 U13790 ( .A(n13820), .B(n13821), .Z(n13819) );
  XOR2_X1 U13791 ( .A(n13822), .B(n13823), .Z(n13609) );
  XOR2_X1 U13792 ( .A(n13824), .B(n13825), .Z(n13823) );
  XOR2_X1 U13793 ( .A(n13826), .B(n13827), .Z(n13613) );
  XOR2_X1 U13794 ( .A(n13828), .B(n13829), .Z(n13827) );
  XOR2_X1 U13795 ( .A(n13830), .B(n13831), .Z(n13617) );
  XOR2_X1 U13796 ( .A(n13832), .B(n13833), .Z(n13831) );
  XOR2_X1 U13797 ( .A(n13834), .B(n13835), .Z(n13621) );
  XOR2_X1 U13798 ( .A(n13836), .B(n13837), .Z(n13835) );
  XOR2_X1 U13799 ( .A(n13838), .B(n13839), .Z(n13625) );
  XOR2_X1 U13800 ( .A(n13840), .B(n13841), .Z(n13839) );
  XOR2_X1 U13801 ( .A(n13842), .B(n13843), .Z(n13629) );
  XOR2_X1 U13802 ( .A(n13844), .B(n13845), .Z(n13843) );
  XNOR2_X1 U13803 ( .A(n13846), .B(n13847), .ZN(n9017) );
  XOR2_X1 U13804 ( .A(n13848), .B(n13849), .Z(n13847) );
  XOR2_X1 U13805 ( .A(n9028), .B(n9027), .Z(n9015) );
  INV_X1 U13806 ( .A(n13850), .ZN(n9027) );
  OR2_X1 U13807 ( .A1(n13851), .A2(n13852), .ZN(n13850) );
  AND2_X1 U13808 ( .A1(n13849), .A2(n13848), .ZN(n13852) );
  AND2_X1 U13809 ( .A1(n13846), .A2(n13853), .ZN(n13851) );
  OR2_X1 U13810 ( .A1(n13848), .A2(n13849), .ZN(n13853) );
  OR2_X1 U13811 ( .A1(n9248), .A2(n8771), .ZN(n13849) );
  OR2_X1 U13812 ( .A1(n13854), .A2(n13855), .ZN(n13848) );
  AND2_X1 U13813 ( .A1(n13845), .A2(n13844), .ZN(n13855) );
  AND2_X1 U13814 ( .A1(n13842), .A2(n13856), .ZN(n13854) );
  OR2_X1 U13815 ( .A1(n13844), .A2(n13845), .ZN(n13856) );
  OR2_X1 U13816 ( .A1(n8730), .A2(n8771), .ZN(n13845) );
  OR2_X1 U13817 ( .A1(n13857), .A2(n13858), .ZN(n13844) );
  AND2_X1 U13818 ( .A1(n13841), .A2(n13840), .ZN(n13858) );
  AND2_X1 U13819 ( .A1(n13838), .A2(n13859), .ZN(n13857) );
  OR2_X1 U13820 ( .A1(n13840), .A2(n13841), .ZN(n13859) );
  OR2_X1 U13821 ( .A1(n8734), .A2(n8771), .ZN(n13841) );
  OR2_X1 U13822 ( .A1(n13860), .A2(n13861), .ZN(n13840) );
  AND2_X1 U13823 ( .A1(n13837), .A2(n13836), .ZN(n13861) );
  AND2_X1 U13824 ( .A1(n13834), .A2(n13862), .ZN(n13860) );
  OR2_X1 U13825 ( .A1(n13836), .A2(n13837), .ZN(n13862) );
  OR2_X1 U13826 ( .A1(n8738), .A2(n8771), .ZN(n13837) );
  OR2_X1 U13827 ( .A1(n13863), .A2(n13864), .ZN(n13836) );
  AND2_X1 U13828 ( .A1(n13833), .A2(n13832), .ZN(n13864) );
  AND2_X1 U13829 ( .A1(n13830), .A2(n13865), .ZN(n13863) );
  OR2_X1 U13830 ( .A1(n13832), .A2(n13833), .ZN(n13865) );
  OR2_X1 U13831 ( .A1(n8742), .A2(n8771), .ZN(n13833) );
  OR2_X1 U13832 ( .A1(n13866), .A2(n13867), .ZN(n13832) );
  AND2_X1 U13833 ( .A1(n13829), .A2(n13828), .ZN(n13867) );
  AND2_X1 U13834 ( .A1(n13826), .A2(n13868), .ZN(n13866) );
  OR2_X1 U13835 ( .A1(n13828), .A2(n13829), .ZN(n13868) );
  OR2_X1 U13836 ( .A1(n8746), .A2(n8771), .ZN(n13829) );
  OR2_X1 U13837 ( .A1(n13869), .A2(n13870), .ZN(n13828) );
  AND2_X1 U13838 ( .A1(n13825), .A2(n13824), .ZN(n13870) );
  AND2_X1 U13839 ( .A1(n13822), .A2(n13871), .ZN(n13869) );
  OR2_X1 U13840 ( .A1(n13824), .A2(n13825), .ZN(n13871) );
  OR2_X1 U13841 ( .A1(n8750), .A2(n8771), .ZN(n13825) );
  OR2_X1 U13842 ( .A1(n13872), .A2(n13873), .ZN(n13824) );
  AND2_X1 U13843 ( .A1(n13821), .A2(n13820), .ZN(n13873) );
  AND2_X1 U13844 ( .A1(n13818), .A2(n13874), .ZN(n13872) );
  OR2_X1 U13845 ( .A1(n13820), .A2(n13821), .ZN(n13874) );
  OR2_X1 U13846 ( .A1(n8754), .A2(n8771), .ZN(n13821) );
  OR2_X1 U13847 ( .A1(n13875), .A2(n13876), .ZN(n13820) );
  AND2_X1 U13848 ( .A1(n13817), .A2(n13816), .ZN(n13876) );
  AND2_X1 U13849 ( .A1(n13814), .A2(n13877), .ZN(n13875) );
  OR2_X1 U13850 ( .A1(n13816), .A2(n13817), .ZN(n13877) );
  OR2_X1 U13851 ( .A1(n8758), .A2(n8771), .ZN(n13817) );
  OR2_X1 U13852 ( .A1(n13878), .A2(n13879), .ZN(n13816) );
  AND2_X1 U13853 ( .A1(n13813), .A2(n13812), .ZN(n13879) );
  AND2_X1 U13854 ( .A1(n13810), .A2(n13880), .ZN(n13878) );
  OR2_X1 U13855 ( .A1(n13812), .A2(n13813), .ZN(n13880) );
  OR2_X1 U13856 ( .A1(n8762), .A2(n8771), .ZN(n13813) );
  OR2_X1 U13857 ( .A1(n13881), .A2(n13882), .ZN(n13812) );
  AND2_X1 U13858 ( .A1(n13809), .A2(n13808), .ZN(n13882) );
  AND2_X1 U13859 ( .A1(n13806), .A2(n13883), .ZN(n13881) );
  OR2_X1 U13860 ( .A1(n13808), .A2(n13809), .ZN(n13883) );
  OR2_X1 U13861 ( .A1(n8766), .A2(n8771), .ZN(n13809) );
  OR2_X1 U13862 ( .A1(n13884), .A2(n13885), .ZN(n13808) );
  AND2_X1 U13863 ( .A1(n8426), .A2(n13805), .ZN(n13885) );
  AND2_X1 U13864 ( .A1(n13803), .A2(n13886), .ZN(n13884) );
  OR2_X1 U13865 ( .A1(n13805), .A2(n8426), .ZN(n13886) );
  OR2_X1 U13866 ( .A1(n8770), .A2(n8771), .ZN(n8426) );
  OR2_X1 U13867 ( .A1(n13887), .A2(n13888), .ZN(n13805) );
  AND2_X1 U13868 ( .A1(n13802), .A2(n13801), .ZN(n13888) );
  AND2_X1 U13869 ( .A1(n13799), .A2(n13889), .ZN(n13887) );
  OR2_X1 U13870 ( .A1(n13801), .A2(n13802), .ZN(n13889) );
  OR2_X1 U13871 ( .A1(n8774), .A2(n8771), .ZN(n13802) );
  OR2_X1 U13872 ( .A1(n13890), .A2(n13891), .ZN(n13801) );
  AND2_X1 U13873 ( .A1(n13798), .A2(n13797), .ZN(n13891) );
  AND2_X1 U13874 ( .A1(n13795), .A2(n13892), .ZN(n13890) );
  OR2_X1 U13875 ( .A1(n13797), .A2(n13798), .ZN(n13892) );
  OR2_X1 U13876 ( .A1(n8778), .A2(n8771), .ZN(n13798) );
  OR2_X1 U13877 ( .A1(n13893), .A2(n13894), .ZN(n13797) );
  AND2_X1 U13878 ( .A1(n13794), .A2(n13793), .ZN(n13894) );
  AND2_X1 U13879 ( .A1(n13791), .A2(n13895), .ZN(n13893) );
  OR2_X1 U13880 ( .A1(n13793), .A2(n13794), .ZN(n13895) );
  OR2_X1 U13881 ( .A1(n8782), .A2(n8771), .ZN(n13794) );
  OR2_X1 U13882 ( .A1(n13896), .A2(n13897), .ZN(n13793) );
  AND2_X1 U13883 ( .A1(n13790), .A2(n13789), .ZN(n13897) );
  AND2_X1 U13884 ( .A1(n13787), .A2(n13898), .ZN(n13896) );
  OR2_X1 U13885 ( .A1(n13789), .A2(n13790), .ZN(n13898) );
  OR2_X1 U13886 ( .A1(n8786), .A2(n8771), .ZN(n13790) );
  OR2_X1 U13887 ( .A1(n13899), .A2(n13900), .ZN(n13789) );
  AND2_X1 U13888 ( .A1(n13786), .A2(n13785), .ZN(n13900) );
  AND2_X1 U13889 ( .A1(n13783), .A2(n13901), .ZN(n13899) );
  OR2_X1 U13890 ( .A1(n13785), .A2(n13786), .ZN(n13901) );
  OR2_X1 U13891 ( .A1(n8790), .A2(n8771), .ZN(n13786) );
  OR2_X1 U13892 ( .A1(n13902), .A2(n13903), .ZN(n13785) );
  AND2_X1 U13893 ( .A1(n13782), .A2(n13781), .ZN(n13903) );
  AND2_X1 U13894 ( .A1(n13779), .A2(n13904), .ZN(n13902) );
  OR2_X1 U13895 ( .A1(n13781), .A2(n13782), .ZN(n13904) );
  OR2_X1 U13896 ( .A1(n8794), .A2(n8771), .ZN(n13782) );
  OR2_X1 U13897 ( .A1(n13905), .A2(n13906), .ZN(n13781) );
  AND2_X1 U13898 ( .A1(n13778), .A2(n13777), .ZN(n13906) );
  AND2_X1 U13899 ( .A1(n13775), .A2(n13907), .ZN(n13905) );
  OR2_X1 U13900 ( .A1(n13777), .A2(n13778), .ZN(n13907) );
  OR2_X1 U13901 ( .A1(n8798), .A2(n8771), .ZN(n13778) );
  OR2_X1 U13902 ( .A1(n13908), .A2(n13909), .ZN(n13777) );
  AND2_X1 U13903 ( .A1(n13774), .A2(n13773), .ZN(n13909) );
  AND2_X1 U13904 ( .A1(n13771), .A2(n13910), .ZN(n13908) );
  OR2_X1 U13905 ( .A1(n13773), .A2(n13774), .ZN(n13910) );
  OR2_X1 U13906 ( .A1(n8802), .A2(n8771), .ZN(n13774) );
  OR2_X1 U13907 ( .A1(n13911), .A2(n13912), .ZN(n13773) );
  AND2_X1 U13908 ( .A1(n13770), .A2(n13769), .ZN(n13912) );
  AND2_X1 U13909 ( .A1(n13767), .A2(n13913), .ZN(n13911) );
  OR2_X1 U13910 ( .A1(n13769), .A2(n13770), .ZN(n13913) );
  OR2_X1 U13911 ( .A1(n8806), .A2(n8771), .ZN(n13770) );
  OR2_X1 U13912 ( .A1(n13914), .A2(n13915), .ZN(n13769) );
  AND2_X1 U13913 ( .A1(n13766), .A2(n13765), .ZN(n13915) );
  AND2_X1 U13914 ( .A1(n13763), .A2(n13916), .ZN(n13914) );
  OR2_X1 U13915 ( .A1(n13765), .A2(n13766), .ZN(n13916) );
  OR2_X1 U13916 ( .A1(n8810), .A2(n8771), .ZN(n13766) );
  OR2_X1 U13917 ( .A1(n13917), .A2(n13918), .ZN(n13765) );
  AND2_X1 U13918 ( .A1(n13762), .A2(n13761), .ZN(n13918) );
  AND2_X1 U13919 ( .A1(n13759), .A2(n13919), .ZN(n13917) );
  OR2_X1 U13920 ( .A1(n13761), .A2(n13762), .ZN(n13919) );
  OR2_X1 U13921 ( .A1(n8140), .A2(n8771), .ZN(n13762) );
  OR2_X1 U13922 ( .A1(n13920), .A2(n13921), .ZN(n13761) );
  AND2_X1 U13923 ( .A1(n13758), .A2(n13757), .ZN(n13921) );
  AND2_X1 U13924 ( .A1(n13755), .A2(n13922), .ZN(n13920) );
  OR2_X1 U13925 ( .A1(n13757), .A2(n13758), .ZN(n13922) );
  OR2_X1 U13926 ( .A1(n8115), .A2(n8771), .ZN(n13758) );
  OR2_X1 U13927 ( .A1(n13923), .A2(n13924), .ZN(n13757) );
  AND2_X1 U13928 ( .A1(n13754), .A2(n13753), .ZN(n13924) );
  AND2_X1 U13929 ( .A1(n13751), .A2(n13925), .ZN(n13923) );
  OR2_X1 U13930 ( .A1(n13753), .A2(n13754), .ZN(n13925) );
  OR2_X1 U13931 ( .A1(n8090), .A2(n8771), .ZN(n13754) );
  OR2_X1 U13932 ( .A1(n13926), .A2(n13927), .ZN(n13753) );
  AND2_X1 U13933 ( .A1(n13750), .A2(n13749), .ZN(n13927) );
  AND2_X1 U13934 ( .A1(n13747), .A2(n13928), .ZN(n13926) );
  OR2_X1 U13935 ( .A1(n13749), .A2(n13750), .ZN(n13928) );
  OR2_X1 U13936 ( .A1(n8065), .A2(n8771), .ZN(n13750) );
  OR2_X1 U13937 ( .A1(n13929), .A2(n13930), .ZN(n13749) );
  AND2_X1 U13938 ( .A1(n13746), .A2(n13745), .ZN(n13930) );
  AND2_X1 U13939 ( .A1(n13743), .A2(n13931), .ZN(n13929) );
  OR2_X1 U13940 ( .A1(n13745), .A2(n13746), .ZN(n13931) );
  OR2_X1 U13941 ( .A1(n8040), .A2(n8771), .ZN(n13746) );
  OR2_X1 U13942 ( .A1(n13932), .A2(n13933), .ZN(n13745) );
  AND2_X1 U13943 ( .A1(n13742), .A2(n13741), .ZN(n13933) );
  AND2_X1 U13944 ( .A1(n13739), .A2(n13934), .ZN(n13932) );
  OR2_X1 U13945 ( .A1(n13741), .A2(n13742), .ZN(n13934) );
  OR2_X1 U13946 ( .A1(n8015), .A2(n8771), .ZN(n13742) );
  OR2_X1 U13947 ( .A1(n13935), .A2(n13936), .ZN(n13741) );
  AND2_X1 U13948 ( .A1(n13738), .A2(n13737), .ZN(n13936) );
  AND2_X1 U13949 ( .A1(n13735), .A2(n13937), .ZN(n13935) );
  OR2_X1 U13950 ( .A1(n13737), .A2(n13738), .ZN(n13937) );
  OR2_X1 U13951 ( .A1(n7979), .A2(n8771), .ZN(n13738) );
  OR2_X1 U13952 ( .A1(n13938), .A2(n13939), .ZN(n13737) );
  AND2_X1 U13953 ( .A1(n13731), .A2(n13734), .ZN(n13939) );
  AND2_X1 U13954 ( .A1(n13940), .A2(n13941), .ZN(n13938) );
  OR2_X1 U13955 ( .A1(n13734), .A2(n13731), .ZN(n13941) );
  OR2_X1 U13956 ( .A1(n7954), .A2(n8771), .ZN(n13731) );
  OR3_X1 U13957 ( .A1(n8771), .A2(n8767), .A3(n9796), .ZN(n13734) );
  INV_X1 U13958 ( .A(n13733), .ZN(n13940) );
  OR2_X1 U13959 ( .A1(n13942), .A2(n13943), .ZN(n13733) );
  AND2_X1 U13960 ( .A1(b_9_), .A2(n13944), .ZN(n13943) );
  OR2_X1 U13961 ( .A1(n13945), .A2(n7920), .ZN(n13944) );
  AND2_X1 U13962 ( .A1(a_31_), .A2(n8767), .ZN(n13945) );
  AND2_X1 U13963 ( .A1(b_10_), .A2(n13946), .ZN(n13942) );
  OR2_X1 U13964 ( .A1(n13947), .A2(n9801), .ZN(n13946) );
  AND2_X1 U13965 ( .A1(a_30_), .A2(n8763), .ZN(n13947) );
  XNOR2_X1 U13966 ( .A(n13948), .B(n13949), .ZN(n13735) );
  XOR2_X1 U13967 ( .A(n13950), .B(n13951), .Z(n13949) );
  XOR2_X1 U13968 ( .A(n13952), .B(n13953), .Z(n13739) );
  XOR2_X1 U13969 ( .A(n13954), .B(n13955), .Z(n13953) );
  XOR2_X1 U13970 ( .A(n13956), .B(n13957), .Z(n13743) );
  XOR2_X1 U13971 ( .A(n13958), .B(n13959), .Z(n13957) );
  XOR2_X1 U13972 ( .A(n13960), .B(n13961), .Z(n13747) );
  XOR2_X1 U13973 ( .A(n13962), .B(n13963), .Z(n13961) );
  XOR2_X1 U13974 ( .A(n13964), .B(n13965), .Z(n13751) );
  XOR2_X1 U13975 ( .A(n13966), .B(n13967), .Z(n13965) );
  XOR2_X1 U13976 ( .A(n13968), .B(n13969), .Z(n13755) );
  XOR2_X1 U13977 ( .A(n13970), .B(n13971), .Z(n13969) );
  XOR2_X1 U13978 ( .A(n13972), .B(n13973), .Z(n13759) );
  XOR2_X1 U13979 ( .A(n13974), .B(n13975), .Z(n13973) );
  XOR2_X1 U13980 ( .A(n13976), .B(n13977), .Z(n13763) );
  XOR2_X1 U13981 ( .A(n13978), .B(n13979), .Z(n13977) );
  XOR2_X1 U13982 ( .A(n13980), .B(n13981), .Z(n13767) );
  XOR2_X1 U13983 ( .A(n13982), .B(n13983), .Z(n13981) );
  XOR2_X1 U13984 ( .A(n13984), .B(n13985), .Z(n13771) );
  XOR2_X1 U13985 ( .A(n13986), .B(n13987), .Z(n13985) );
  XOR2_X1 U13986 ( .A(n13988), .B(n13989), .Z(n13775) );
  XOR2_X1 U13987 ( .A(n13990), .B(n13991), .Z(n13989) );
  XOR2_X1 U13988 ( .A(n13992), .B(n13993), .Z(n13779) );
  XOR2_X1 U13989 ( .A(n13994), .B(n13995), .Z(n13993) );
  XOR2_X1 U13990 ( .A(n13996), .B(n13997), .Z(n13783) );
  XOR2_X1 U13991 ( .A(n13998), .B(n13999), .Z(n13997) );
  XOR2_X1 U13992 ( .A(n14000), .B(n14001), .Z(n13787) );
  XOR2_X1 U13993 ( .A(n14002), .B(n14003), .Z(n14001) );
  XOR2_X1 U13994 ( .A(n14004), .B(n14005), .Z(n13791) );
  XOR2_X1 U13995 ( .A(n14006), .B(n14007), .Z(n14005) );
  XOR2_X1 U13996 ( .A(n14008), .B(n14009), .Z(n13795) );
  XOR2_X1 U13997 ( .A(n14010), .B(n14011), .Z(n14009) );
  XOR2_X1 U13998 ( .A(n14012), .B(n14013), .Z(n13799) );
  XOR2_X1 U13999 ( .A(n14014), .B(n14015), .Z(n14013) );
  XOR2_X1 U14000 ( .A(n14016), .B(n14017), .Z(n13803) );
  XOR2_X1 U14001 ( .A(n14018), .B(n14019), .Z(n14017) );
  XOR2_X1 U14002 ( .A(n14020), .B(n14021), .Z(n13806) );
  XOR2_X1 U14003 ( .A(n14022), .B(n14023), .Z(n14021) );
  XOR2_X1 U14004 ( .A(n14024), .B(n14025), .Z(n13810) );
  XOR2_X1 U14005 ( .A(n14026), .B(n8452), .Z(n14025) );
  XOR2_X1 U14006 ( .A(n14027), .B(n14028), .Z(n13814) );
  XOR2_X1 U14007 ( .A(n14029), .B(n14030), .Z(n14028) );
  XOR2_X1 U14008 ( .A(n14031), .B(n14032), .Z(n13818) );
  XOR2_X1 U14009 ( .A(n14033), .B(n14034), .Z(n14032) );
  XOR2_X1 U14010 ( .A(n14035), .B(n14036), .Z(n13822) );
  XOR2_X1 U14011 ( .A(n14037), .B(n14038), .Z(n14036) );
  XOR2_X1 U14012 ( .A(n14039), .B(n14040), .Z(n13826) );
  XOR2_X1 U14013 ( .A(n14041), .B(n14042), .Z(n14040) );
  XOR2_X1 U14014 ( .A(n14043), .B(n14044), .Z(n13830) );
  XOR2_X1 U14015 ( .A(n14045), .B(n14046), .Z(n14044) );
  XOR2_X1 U14016 ( .A(n14047), .B(n14048), .Z(n13834) );
  XOR2_X1 U14017 ( .A(n14049), .B(n14050), .Z(n14048) );
  XOR2_X1 U14018 ( .A(n14051), .B(n14052), .Z(n13838) );
  XOR2_X1 U14019 ( .A(n14053), .B(n14054), .Z(n14052) );
  XOR2_X1 U14020 ( .A(n14055), .B(n14056), .Z(n13842) );
  XOR2_X1 U14021 ( .A(n14057), .B(n14058), .Z(n14056) );
  XOR2_X1 U14022 ( .A(n14059), .B(n14060), .Z(n13846) );
  XOR2_X1 U14023 ( .A(n14061), .B(n14062), .Z(n14060) );
  XNOR2_X1 U14024 ( .A(n14063), .B(n14064), .ZN(n9028) );
  XOR2_X1 U14025 ( .A(n14065), .B(n14066), .Z(n14064) );
  XOR2_X1 U14026 ( .A(n7872), .B(n7871), .Z(n9026) );
  INV_X1 U14027 ( .A(n14067), .ZN(n7871) );
  OR2_X1 U14028 ( .A1(n14068), .A2(n14069), .ZN(n14067) );
  AND2_X1 U14029 ( .A1(n14066), .A2(n14065), .ZN(n14069) );
  AND2_X1 U14030 ( .A1(n14063), .A2(n14070), .ZN(n14068) );
  OR2_X1 U14031 ( .A1(n14065), .A2(n14066), .ZN(n14070) );
  OR2_X1 U14032 ( .A1(n9248), .A2(n8767), .ZN(n14066) );
  OR2_X1 U14033 ( .A1(n14071), .A2(n14072), .ZN(n14065) );
  AND2_X1 U14034 ( .A1(n14062), .A2(n14061), .ZN(n14072) );
  AND2_X1 U14035 ( .A1(n14059), .A2(n14073), .ZN(n14071) );
  OR2_X1 U14036 ( .A1(n14061), .A2(n14062), .ZN(n14073) );
  OR2_X1 U14037 ( .A1(n8730), .A2(n8767), .ZN(n14062) );
  OR2_X1 U14038 ( .A1(n14074), .A2(n14075), .ZN(n14061) );
  AND2_X1 U14039 ( .A1(n14058), .A2(n14057), .ZN(n14075) );
  AND2_X1 U14040 ( .A1(n14055), .A2(n14076), .ZN(n14074) );
  OR2_X1 U14041 ( .A1(n14057), .A2(n14058), .ZN(n14076) );
  OR2_X1 U14042 ( .A1(n8734), .A2(n8767), .ZN(n14058) );
  OR2_X1 U14043 ( .A1(n14077), .A2(n14078), .ZN(n14057) );
  AND2_X1 U14044 ( .A1(n14054), .A2(n14053), .ZN(n14078) );
  AND2_X1 U14045 ( .A1(n14051), .A2(n14079), .ZN(n14077) );
  OR2_X1 U14046 ( .A1(n14053), .A2(n14054), .ZN(n14079) );
  OR2_X1 U14047 ( .A1(n8738), .A2(n8767), .ZN(n14054) );
  OR2_X1 U14048 ( .A1(n14080), .A2(n14081), .ZN(n14053) );
  AND2_X1 U14049 ( .A1(n14050), .A2(n14049), .ZN(n14081) );
  AND2_X1 U14050 ( .A1(n14047), .A2(n14082), .ZN(n14080) );
  OR2_X1 U14051 ( .A1(n14049), .A2(n14050), .ZN(n14082) );
  OR2_X1 U14052 ( .A1(n8742), .A2(n8767), .ZN(n14050) );
  OR2_X1 U14053 ( .A1(n14083), .A2(n14084), .ZN(n14049) );
  AND2_X1 U14054 ( .A1(n14046), .A2(n14045), .ZN(n14084) );
  AND2_X1 U14055 ( .A1(n14043), .A2(n14085), .ZN(n14083) );
  OR2_X1 U14056 ( .A1(n14045), .A2(n14046), .ZN(n14085) );
  OR2_X1 U14057 ( .A1(n8746), .A2(n8767), .ZN(n14046) );
  OR2_X1 U14058 ( .A1(n14086), .A2(n14087), .ZN(n14045) );
  AND2_X1 U14059 ( .A1(n14042), .A2(n14041), .ZN(n14087) );
  AND2_X1 U14060 ( .A1(n14039), .A2(n14088), .ZN(n14086) );
  OR2_X1 U14061 ( .A1(n14041), .A2(n14042), .ZN(n14088) );
  OR2_X1 U14062 ( .A1(n8750), .A2(n8767), .ZN(n14042) );
  OR2_X1 U14063 ( .A1(n14089), .A2(n14090), .ZN(n14041) );
  AND2_X1 U14064 ( .A1(n14038), .A2(n14037), .ZN(n14090) );
  AND2_X1 U14065 ( .A1(n14035), .A2(n14091), .ZN(n14089) );
  OR2_X1 U14066 ( .A1(n14037), .A2(n14038), .ZN(n14091) );
  OR2_X1 U14067 ( .A1(n8754), .A2(n8767), .ZN(n14038) );
  OR2_X1 U14068 ( .A1(n14092), .A2(n14093), .ZN(n14037) );
  AND2_X1 U14069 ( .A1(n14034), .A2(n14033), .ZN(n14093) );
  AND2_X1 U14070 ( .A1(n14031), .A2(n14094), .ZN(n14092) );
  OR2_X1 U14071 ( .A1(n14033), .A2(n14034), .ZN(n14094) );
  OR2_X1 U14072 ( .A1(n8758), .A2(n8767), .ZN(n14034) );
  OR2_X1 U14073 ( .A1(n14095), .A2(n14096), .ZN(n14033) );
  AND2_X1 U14074 ( .A1(n14030), .A2(n14029), .ZN(n14096) );
  AND2_X1 U14075 ( .A1(n14027), .A2(n14097), .ZN(n14095) );
  OR2_X1 U14076 ( .A1(n14029), .A2(n14030), .ZN(n14097) );
  OR2_X1 U14077 ( .A1(n8762), .A2(n8767), .ZN(n14030) );
  OR2_X1 U14078 ( .A1(n14098), .A2(n14099), .ZN(n14029) );
  AND2_X1 U14079 ( .A1(n8452), .A2(n14026), .ZN(n14099) );
  AND2_X1 U14080 ( .A1(n14024), .A2(n14100), .ZN(n14098) );
  OR2_X1 U14081 ( .A1(n14026), .A2(n8452), .ZN(n14100) );
  OR2_X1 U14082 ( .A1(n8766), .A2(n8767), .ZN(n8452) );
  OR2_X1 U14083 ( .A1(n14101), .A2(n14102), .ZN(n14026) );
  AND2_X1 U14084 ( .A1(n14023), .A2(n14022), .ZN(n14102) );
  AND2_X1 U14085 ( .A1(n14020), .A2(n14103), .ZN(n14101) );
  OR2_X1 U14086 ( .A1(n14022), .A2(n14023), .ZN(n14103) );
  OR2_X1 U14087 ( .A1(n8770), .A2(n8767), .ZN(n14023) );
  OR2_X1 U14088 ( .A1(n14104), .A2(n14105), .ZN(n14022) );
  AND2_X1 U14089 ( .A1(n14019), .A2(n14018), .ZN(n14105) );
  AND2_X1 U14090 ( .A1(n14016), .A2(n14106), .ZN(n14104) );
  OR2_X1 U14091 ( .A1(n14018), .A2(n14019), .ZN(n14106) );
  OR2_X1 U14092 ( .A1(n8774), .A2(n8767), .ZN(n14019) );
  OR2_X1 U14093 ( .A1(n14107), .A2(n14108), .ZN(n14018) );
  AND2_X1 U14094 ( .A1(n14015), .A2(n14014), .ZN(n14108) );
  AND2_X1 U14095 ( .A1(n14012), .A2(n14109), .ZN(n14107) );
  OR2_X1 U14096 ( .A1(n14014), .A2(n14015), .ZN(n14109) );
  OR2_X1 U14097 ( .A1(n8778), .A2(n8767), .ZN(n14015) );
  OR2_X1 U14098 ( .A1(n14110), .A2(n14111), .ZN(n14014) );
  AND2_X1 U14099 ( .A1(n14011), .A2(n14010), .ZN(n14111) );
  AND2_X1 U14100 ( .A1(n14008), .A2(n14112), .ZN(n14110) );
  OR2_X1 U14101 ( .A1(n14010), .A2(n14011), .ZN(n14112) );
  OR2_X1 U14102 ( .A1(n8782), .A2(n8767), .ZN(n14011) );
  OR2_X1 U14103 ( .A1(n14113), .A2(n14114), .ZN(n14010) );
  AND2_X1 U14104 ( .A1(n14007), .A2(n14006), .ZN(n14114) );
  AND2_X1 U14105 ( .A1(n14004), .A2(n14115), .ZN(n14113) );
  OR2_X1 U14106 ( .A1(n14006), .A2(n14007), .ZN(n14115) );
  OR2_X1 U14107 ( .A1(n8786), .A2(n8767), .ZN(n14007) );
  OR2_X1 U14108 ( .A1(n14116), .A2(n14117), .ZN(n14006) );
  AND2_X1 U14109 ( .A1(n14003), .A2(n14002), .ZN(n14117) );
  AND2_X1 U14110 ( .A1(n14000), .A2(n14118), .ZN(n14116) );
  OR2_X1 U14111 ( .A1(n14002), .A2(n14003), .ZN(n14118) );
  OR2_X1 U14112 ( .A1(n8790), .A2(n8767), .ZN(n14003) );
  OR2_X1 U14113 ( .A1(n14119), .A2(n14120), .ZN(n14002) );
  AND2_X1 U14114 ( .A1(n13999), .A2(n13998), .ZN(n14120) );
  AND2_X1 U14115 ( .A1(n13996), .A2(n14121), .ZN(n14119) );
  OR2_X1 U14116 ( .A1(n13998), .A2(n13999), .ZN(n14121) );
  OR2_X1 U14117 ( .A1(n8794), .A2(n8767), .ZN(n13999) );
  OR2_X1 U14118 ( .A1(n14122), .A2(n14123), .ZN(n13998) );
  AND2_X1 U14119 ( .A1(n13995), .A2(n13994), .ZN(n14123) );
  AND2_X1 U14120 ( .A1(n13992), .A2(n14124), .ZN(n14122) );
  OR2_X1 U14121 ( .A1(n13994), .A2(n13995), .ZN(n14124) );
  OR2_X1 U14122 ( .A1(n8798), .A2(n8767), .ZN(n13995) );
  OR2_X1 U14123 ( .A1(n14125), .A2(n14126), .ZN(n13994) );
  AND2_X1 U14124 ( .A1(n13988), .A2(n13991), .ZN(n14126) );
  AND2_X1 U14125 ( .A1(n14127), .A2(n13990), .ZN(n14125) );
  OR2_X1 U14126 ( .A1(n14128), .A2(n14129), .ZN(n13990) );
  AND2_X1 U14127 ( .A1(n13987), .A2(n13986), .ZN(n14129) );
  AND2_X1 U14128 ( .A1(n13984), .A2(n14130), .ZN(n14128) );
  OR2_X1 U14129 ( .A1(n13986), .A2(n13987), .ZN(n14130) );
  OR2_X1 U14130 ( .A1(n8806), .A2(n8767), .ZN(n13987) );
  OR2_X1 U14131 ( .A1(n14131), .A2(n14132), .ZN(n13986) );
  AND2_X1 U14132 ( .A1(n13980), .A2(n13983), .ZN(n14132) );
  AND2_X1 U14133 ( .A1(n14133), .A2(n13982), .ZN(n14131) );
  OR2_X1 U14134 ( .A1(n14134), .A2(n14135), .ZN(n13982) );
  AND2_X1 U14135 ( .A1(n13976), .A2(n13979), .ZN(n14135) );
  AND2_X1 U14136 ( .A1(n14136), .A2(n13978), .ZN(n14134) );
  OR2_X1 U14137 ( .A1(n14137), .A2(n14138), .ZN(n13978) );
  AND2_X1 U14138 ( .A1(n13972), .A2(n13975), .ZN(n14138) );
  AND2_X1 U14139 ( .A1(n14139), .A2(n13974), .ZN(n14137) );
  OR2_X1 U14140 ( .A1(n14140), .A2(n14141), .ZN(n13974) );
  AND2_X1 U14141 ( .A1(n13968), .A2(n13971), .ZN(n14141) );
  AND2_X1 U14142 ( .A1(n14142), .A2(n13970), .ZN(n14140) );
  OR2_X1 U14143 ( .A1(n14143), .A2(n14144), .ZN(n13970) );
  AND2_X1 U14144 ( .A1(n13964), .A2(n13967), .ZN(n14144) );
  AND2_X1 U14145 ( .A1(n14145), .A2(n13966), .ZN(n14143) );
  OR2_X1 U14146 ( .A1(n14146), .A2(n14147), .ZN(n13966) );
  AND2_X1 U14147 ( .A1(n13960), .A2(n13963), .ZN(n14147) );
  AND2_X1 U14148 ( .A1(n14148), .A2(n13962), .ZN(n14146) );
  OR2_X1 U14149 ( .A1(n14149), .A2(n14150), .ZN(n13962) );
  AND2_X1 U14150 ( .A1(n13956), .A2(n13959), .ZN(n14150) );
  AND2_X1 U14151 ( .A1(n14151), .A2(n13958), .ZN(n14149) );
  OR2_X1 U14152 ( .A1(n14152), .A2(n14153), .ZN(n13958) );
  AND2_X1 U14153 ( .A1(n13952), .A2(n13955), .ZN(n14153) );
  AND2_X1 U14154 ( .A1(n14154), .A2(n13954), .ZN(n14152) );
  OR2_X1 U14155 ( .A1(n14155), .A2(n14156), .ZN(n13954) );
  AND2_X1 U14156 ( .A1(n13948), .A2(n13951), .ZN(n14156) );
  AND2_X1 U14157 ( .A1(n14157), .A2(n14158), .ZN(n14155) );
  OR2_X1 U14158 ( .A1(n13951), .A2(n13948), .ZN(n14158) );
  OR2_X1 U14159 ( .A1(n7954), .A2(n8767), .ZN(n13948) );
  OR3_X1 U14160 ( .A1(n8767), .A2(n8763), .A3(n9796), .ZN(n13951) );
  INV_X1 U14161 ( .A(n13950), .ZN(n14157) );
  OR2_X1 U14162 ( .A1(n14159), .A2(n14160), .ZN(n13950) );
  AND2_X1 U14163 ( .A1(b_9_), .A2(n14161), .ZN(n14160) );
  OR2_X1 U14164 ( .A1(n14162), .A2(n9801), .ZN(n14161) );
  AND2_X1 U14165 ( .A1(a_30_), .A2(n8759), .ZN(n14162) );
  AND2_X1 U14166 ( .A1(b_8_), .A2(n14163), .ZN(n14159) );
  OR2_X1 U14167 ( .A1(n14164), .A2(n7920), .ZN(n14163) );
  AND2_X1 U14168 ( .A1(a_31_), .A2(n8763), .ZN(n14164) );
  OR2_X1 U14169 ( .A1(n13955), .A2(n13952), .ZN(n14154) );
  XNOR2_X1 U14170 ( .A(n14165), .B(n14166), .ZN(n13952) );
  XOR2_X1 U14171 ( .A(n14167), .B(n14168), .Z(n14166) );
  OR2_X1 U14172 ( .A1(n7979), .A2(n8767), .ZN(n13955) );
  OR2_X1 U14173 ( .A1(n13959), .A2(n13956), .ZN(n14151) );
  XOR2_X1 U14174 ( .A(n14169), .B(n14170), .Z(n13956) );
  XOR2_X1 U14175 ( .A(n14171), .B(n14172), .Z(n14170) );
  OR2_X1 U14176 ( .A1(n8015), .A2(n8767), .ZN(n13959) );
  OR2_X1 U14177 ( .A1(n13963), .A2(n13960), .ZN(n14148) );
  XOR2_X1 U14178 ( .A(n14173), .B(n14174), .Z(n13960) );
  XOR2_X1 U14179 ( .A(n14175), .B(n14176), .Z(n14174) );
  OR2_X1 U14180 ( .A1(n8040), .A2(n8767), .ZN(n13963) );
  OR2_X1 U14181 ( .A1(n13967), .A2(n13964), .ZN(n14145) );
  XOR2_X1 U14182 ( .A(n14177), .B(n14178), .Z(n13964) );
  XOR2_X1 U14183 ( .A(n14179), .B(n14180), .Z(n14178) );
  OR2_X1 U14184 ( .A1(n8065), .A2(n8767), .ZN(n13967) );
  OR2_X1 U14185 ( .A1(n13971), .A2(n13968), .ZN(n14142) );
  XOR2_X1 U14186 ( .A(n14181), .B(n14182), .Z(n13968) );
  XOR2_X1 U14187 ( .A(n14183), .B(n14184), .Z(n14182) );
  OR2_X1 U14188 ( .A1(n8090), .A2(n8767), .ZN(n13971) );
  OR2_X1 U14189 ( .A1(n13975), .A2(n13972), .ZN(n14139) );
  XOR2_X1 U14190 ( .A(n14185), .B(n14186), .Z(n13972) );
  XOR2_X1 U14191 ( .A(n14187), .B(n14188), .Z(n14186) );
  OR2_X1 U14192 ( .A1(n8115), .A2(n8767), .ZN(n13975) );
  OR2_X1 U14193 ( .A1(n13979), .A2(n13976), .ZN(n14136) );
  XOR2_X1 U14194 ( .A(n14189), .B(n14190), .Z(n13976) );
  XOR2_X1 U14195 ( .A(n14191), .B(n14192), .Z(n14190) );
  OR2_X1 U14196 ( .A1(n8140), .A2(n8767), .ZN(n13979) );
  OR2_X1 U14197 ( .A1(n13983), .A2(n13980), .ZN(n14133) );
  XOR2_X1 U14198 ( .A(n14193), .B(n14194), .Z(n13980) );
  XOR2_X1 U14199 ( .A(n14195), .B(n14196), .Z(n14194) );
  OR2_X1 U14200 ( .A1(n8810), .A2(n8767), .ZN(n13983) );
  XOR2_X1 U14201 ( .A(n14197), .B(n14198), .Z(n13984) );
  XOR2_X1 U14202 ( .A(n14199), .B(n14200), .Z(n14198) );
  OR2_X1 U14203 ( .A1(n13991), .A2(n13988), .ZN(n14127) );
  XOR2_X1 U14204 ( .A(n14201), .B(n14202), .Z(n13988) );
  XOR2_X1 U14205 ( .A(n14203), .B(n14204), .Z(n14202) );
  OR2_X1 U14206 ( .A1(n8802), .A2(n8767), .ZN(n13991) );
  XOR2_X1 U14207 ( .A(n14205), .B(n14206), .Z(n13992) );
  XOR2_X1 U14208 ( .A(n14207), .B(n14208), .Z(n14206) );
  XOR2_X1 U14209 ( .A(n14209), .B(n14210), .Z(n13996) );
  XOR2_X1 U14210 ( .A(n14211), .B(n14212), .Z(n14210) );
  XOR2_X1 U14211 ( .A(n14213), .B(n14214), .Z(n14000) );
  XOR2_X1 U14212 ( .A(n14215), .B(n14216), .Z(n14214) );
  XOR2_X1 U14213 ( .A(n14217), .B(n14218), .Z(n14004) );
  XOR2_X1 U14214 ( .A(n14219), .B(n14220), .Z(n14218) );
  XOR2_X1 U14215 ( .A(n14221), .B(n14222), .Z(n14008) );
  XOR2_X1 U14216 ( .A(n14223), .B(n14224), .Z(n14222) );
  XOR2_X1 U14217 ( .A(n14225), .B(n14226), .Z(n14012) );
  XOR2_X1 U14218 ( .A(n14227), .B(n14228), .Z(n14226) );
  XOR2_X1 U14219 ( .A(n14229), .B(n14230), .Z(n14016) );
  XOR2_X1 U14220 ( .A(n14231), .B(n14232), .Z(n14230) );
  XOR2_X1 U14221 ( .A(n14233), .B(n14234), .Z(n14020) );
  XOR2_X1 U14222 ( .A(n14235), .B(n14236), .Z(n14234) );
  XOR2_X1 U14223 ( .A(n14237), .B(n14238), .Z(n14024) );
  XOR2_X1 U14224 ( .A(n14239), .B(n14240), .Z(n14238) );
  XOR2_X1 U14225 ( .A(n14241), .B(n14242), .Z(n14027) );
  XOR2_X1 U14226 ( .A(n14243), .B(n14244), .Z(n14242) );
  XOR2_X1 U14227 ( .A(n14245), .B(n14246), .Z(n14031) );
  XOR2_X1 U14228 ( .A(n14247), .B(n8478), .Z(n14246) );
  XOR2_X1 U14229 ( .A(n14248), .B(n14249), .Z(n14035) );
  XOR2_X1 U14230 ( .A(n14250), .B(n14251), .Z(n14249) );
  XOR2_X1 U14231 ( .A(n14252), .B(n14253), .Z(n14039) );
  XOR2_X1 U14232 ( .A(n14254), .B(n14255), .Z(n14253) );
  XOR2_X1 U14233 ( .A(n14256), .B(n14257), .Z(n14043) );
  XOR2_X1 U14234 ( .A(n14258), .B(n14259), .Z(n14257) );
  XOR2_X1 U14235 ( .A(n14260), .B(n14261), .Z(n14047) );
  XOR2_X1 U14236 ( .A(n14262), .B(n14263), .Z(n14261) );
  XOR2_X1 U14237 ( .A(n14264), .B(n14265), .Z(n14051) );
  XOR2_X1 U14238 ( .A(n14266), .B(n14267), .Z(n14265) );
  XOR2_X1 U14239 ( .A(n14268), .B(n14269), .Z(n14055) );
  XOR2_X1 U14240 ( .A(n14270), .B(n14271), .Z(n14269) );
  XOR2_X1 U14241 ( .A(n14272), .B(n14273), .Z(n14059) );
  XOR2_X1 U14242 ( .A(n14274), .B(n14275), .Z(n14273) );
  XOR2_X1 U14243 ( .A(n14276), .B(n14277), .Z(n14063) );
  XOR2_X1 U14244 ( .A(n14278), .B(n14279), .Z(n14277) );
  XNOR2_X1 U14245 ( .A(n14280), .B(n14281), .ZN(n7872) );
  XOR2_X1 U14246 ( .A(n14282), .B(n14283), .Z(n14281) );
  AND2_X1 U14247 ( .A1(n14284), .A2(n9414), .ZN(n7869) );
  OR2_X1 U14248 ( .A1(n14285), .A2(n14286), .ZN(n9414) );
  INV_X1 U14249 ( .A(n14287), .ZN(n14284) );
  AND2_X1 U14250 ( .A1(n14285), .A2(n14286), .ZN(n14287) );
  OR2_X1 U14251 ( .A1(n14288), .A2(n14289), .ZN(n14286) );
  AND2_X1 U14252 ( .A1(n14283), .A2(n14282), .ZN(n14289) );
  AND2_X1 U14253 ( .A1(n14280), .A2(n14290), .ZN(n14288) );
  OR2_X1 U14254 ( .A1(n14282), .A2(n14283), .ZN(n14290) );
  OR2_X1 U14255 ( .A1(n9248), .A2(n8763), .ZN(n14283) );
  OR2_X1 U14256 ( .A1(n14291), .A2(n14292), .ZN(n14282) );
  AND2_X1 U14257 ( .A1(n14279), .A2(n14278), .ZN(n14292) );
  AND2_X1 U14258 ( .A1(n14276), .A2(n14293), .ZN(n14291) );
  OR2_X1 U14259 ( .A1(n14278), .A2(n14279), .ZN(n14293) );
  OR2_X1 U14260 ( .A1(n8730), .A2(n8763), .ZN(n14279) );
  OR2_X1 U14261 ( .A1(n14294), .A2(n14295), .ZN(n14278) );
  AND2_X1 U14262 ( .A1(n14275), .A2(n14274), .ZN(n14295) );
  AND2_X1 U14263 ( .A1(n14272), .A2(n14296), .ZN(n14294) );
  OR2_X1 U14264 ( .A1(n14274), .A2(n14275), .ZN(n14296) );
  OR2_X1 U14265 ( .A1(n8734), .A2(n8763), .ZN(n14275) );
  OR2_X1 U14266 ( .A1(n14297), .A2(n14298), .ZN(n14274) );
  AND2_X1 U14267 ( .A1(n14271), .A2(n14270), .ZN(n14298) );
  AND2_X1 U14268 ( .A1(n14268), .A2(n14299), .ZN(n14297) );
  OR2_X1 U14269 ( .A1(n14270), .A2(n14271), .ZN(n14299) );
  OR2_X1 U14270 ( .A1(n8738), .A2(n8763), .ZN(n14271) );
  OR2_X1 U14271 ( .A1(n14300), .A2(n14301), .ZN(n14270) );
  AND2_X1 U14272 ( .A1(n14267), .A2(n14266), .ZN(n14301) );
  AND2_X1 U14273 ( .A1(n14264), .A2(n14302), .ZN(n14300) );
  OR2_X1 U14274 ( .A1(n14266), .A2(n14267), .ZN(n14302) );
  OR2_X1 U14275 ( .A1(n8742), .A2(n8763), .ZN(n14267) );
  OR2_X1 U14276 ( .A1(n14303), .A2(n14304), .ZN(n14266) );
  AND2_X1 U14277 ( .A1(n14263), .A2(n14262), .ZN(n14304) );
  AND2_X1 U14278 ( .A1(n14260), .A2(n14305), .ZN(n14303) );
  OR2_X1 U14279 ( .A1(n14262), .A2(n14263), .ZN(n14305) );
  OR2_X1 U14280 ( .A1(n8746), .A2(n8763), .ZN(n14263) );
  OR2_X1 U14281 ( .A1(n14306), .A2(n14307), .ZN(n14262) );
  AND2_X1 U14282 ( .A1(n14259), .A2(n14258), .ZN(n14307) );
  AND2_X1 U14283 ( .A1(n14256), .A2(n14308), .ZN(n14306) );
  OR2_X1 U14284 ( .A1(n14258), .A2(n14259), .ZN(n14308) );
  OR2_X1 U14285 ( .A1(n8750), .A2(n8763), .ZN(n14259) );
  OR2_X1 U14286 ( .A1(n14309), .A2(n14310), .ZN(n14258) );
  AND2_X1 U14287 ( .A1(n14255), .A2(n14254), .ZN(n14310) );
  AND2_X1 U14288 ( .A1(n14252), .A2(n14311), .ZN(n14309) );
  OR2_X1 U14289 ( .A1(n14254), .A2(n14255), .ZN(n14311) );
  OR2_X1 U14290 ( .A1(n8754), .A2(n8763), .ZN(n14255) );
  OR2_X1 U14291 ( .A1(n14312), .A2(n14313), .ZN(n14254) );
  AND2_X1 U14292 ( .A1(n14251), .A2(n14250), .ZN(n14313) );
  AND2_X1 U14293 ( .A1(n14248), .A2(n14314), .ZN(n14312) );
  OR2_X1 U14294 ( .A1(n14250), .A2(n14251), .ZN(n14314) );
  OR2_X1 U14295 ( .A1(n8758), .A2(n8763), .ZN(n14251) );
  OR2_X1 U14296 ( .A1(n14315), .A2(n14316), .ZN(n14250) );
  AND2_X1 U14297 ( .A1(n8478), .A2(n14247), .ZN(n14316) );
  AND2_X1 U14298 ( .A1(n14245), .A2(n14317), .ZN(n14315) );
  OR2_X1 U14299 ( .A1(n14247), .A2(n8478), .ZN(n14317) );
  OR2_X1 U14300 ( .A1(n8762), .A2(n8763), .ZN(n8478) );
  OR2_X1 U14301 ( .A1(n14318), .A2(n14319), .ZN(n14247) );
  AND2_X1 U14302 ( .A1(n14244), .A2(n14243), .ZN(n14319) );
  AND2_X1 U14303 ( .A1(n14241), .A2(n14320), .ZN(n14318) );
  OR2_X1 U14304 ( .A1(n14243), .A2(n14244), .ZN(n14320) );
  OR2_X1 U14305 ( .A1(n8766), .A2(n8763), .ZN(n14244) );
  OR2_X1 U14306 ( .A1(n14321), .A2(n14322), .ZN(n14243) );
  AND2_X1 U14307 ( .A1(n14240), .A2(n14239), .ZN(n14322) );
  AND2_X1 U14308 ( .A1(n14237), .A2(n14323), .ZN(n14321) );
  OR2_X1 U14309 ( .A1(n14239), .A2(n14240), .ZN(n14323) );
  OR2_X1 U14310 ( .A1(n8770), .A2(n8763), .ZN(n14240) );
  OR2_X1 U14311 ( .A1(n14324), .A2(n14325), .ZN(n14239) );
  AND2_X1 U14312 ( .A1(n14236), .A2(n14235), .ZN(n14325) );
  AND2_X1 U14313 ( .A1(n14233), .A2(n14326), .ZN(n14324) );
  OR2_X1 U14314 ( .A1(n14235), .A2(n14236), .ZN(n14326) );
  OR2_X1 U14315 ( .A1(n8774), .A2(n8763), .ZN(n14236) );
  OR2_X1 U14316 ( .A1(n14327), .A2(n14328), .ZN(n14235) );
  AND2_X1 U14317 ( .A1(n14232), .A2(n14231), .ZN(n14328) );
  AND2_X1 U14318 ( .A1(n14229), .A2(n14329), .ZN(n14327) );
  OR2_X1 U14319 ( .A1(n14231), .A2(n14232), .ZN(n14329) );
  OR2_X1 U14320 ( .A1(n8778), .A2(n8763), .ZN(n14232) );
  OR2_X1 U14321 ( .A1(n14330), .A2(n14331), .ZN(n14231) );
  AND2_X1 U14322 ( .A1(n14228), .A2(n14227), .ZN(n14331) );
  AND2_X1 U14323 ( .A1(n14225), .A2(n14332), .ZN(n14330) );
  OR2_X1 U14324 ( .A1(n14227), .A2(n14228), .ZN(n14332) );
  OR2_X1 U14325 ( .A1(n8782), .A2(n8763), .ZN(n14228) );
  OR2_X1 U14326 ( .A1(n14333), .A2(n14334), .ZN(n14227) );
  AND2_X1 U14327 ( .A1(n14224), .A2(n14223), .ZN(n14334) );
  AND2_X1 U14328 ( .A1(n14221), .A2(n14335), .ZN(n14333) );
  OR2_X1 U14329 ( .A1(n14223), .A2(n14224), .ZN(n14335) );
  OR2_X1 U14330 ( .A1(n8786), .A2(n8763), .ZN(n14224) );
  OR2_X1 U14331 ( .A1(n14336), .A2(n14337), .ZN(n14223) );
  AND2_X1 U14332 ( .A1(n14220), .A2(n14219), .ZN(n14337) );
  AND2_X1 U14333 ( .A1(n14217), .A2(n14338), .ZN(n14336) );
  OR2_X1 U14334 ( .A1(n14219), .A2(n14220), .ZN(n14338) );
  OR2_X1 U14335 ( .A1(n8790), .A2(n8763), .ZN(n14220) );
  OR2_X1 U14336 ( .A1(n14339), .A2(n14340), .ZN(n14219) );
  AND2_X1 U14337 ( .A1(n14216), .A2(n14215), .ZN(n14340) );
  AND2_X1 U14338 ( .A1(n14213), .A2(n14341), .ZN(n14339) );
  OR2_X1 U14339 ( .A1(n14215), .A2(n14216), .ZN(n14341) );
  OR2_X1 U14340 ( .A1(n8794), .A2(n8763), .ZN(n14216) );
  OR2_X1 U14341 ( .A1(n14342), .A2(n14343), .ZN(n14215) );
  AND2_X1 U14342 ( .A1(n14212), .A2(n14211), .ZN(n14343) );
  AND2_X1 U14343 ( .A1(n14209), .A2(n14344), .ZN(n14342) );
  OR2_X1 U14344 ( .A1(n14211), .A2(n14212), .ZN(n14344) );
  OR2_X1 U14345 ( .A1(n8798), .A2(n8763), .ZN(n14212) );
  OR2_X1 U14346 ( .A1(n14345), .A2(n14346), .ZN(n14211) );
  AND2_X1 U14347 ( .A1(n14208), .A2(n14207), .ZN(n14346) );
  AND2_X1 U14348 ( .A1(n14205), .A2(n14347), .ZN(n14345) );
  OR2_X1 U14349 ( .A1(n14207), .A2(n14208), .ZN(n14347) );
  OR2_X1 U14350 ( .A1(n8802), .A2(n8763), .ZN(n14208) );
  OR2_X1 U14351 ( .A1(n14348), .A2(n14349), .ZN(n14207) );
  AND2_X1 U14352 ( .A1(n14201), .A2(n14204), .ZN(n14349) );
  AND2_X1 U14353 ( .A1(n14350), .A2(n14203), .ZN(n14348) );
  OR2_X1 U14354 ( .A1(n14351), .A2(n14352), .ZN(n14203) );
  AND2_X1 U14355 ( .A1(n14200), .A2(n14199), .ZN(n14352) );
  AND2_X1 U14356 ( .A1(n14197), .A2(n14353), .ZN(n14351) );
  OR2_X1 U14357 ( .A1(n14199), .A2(n14200), .ZN(n14353) );
  OR2_X1 U14358 ( .A1(n8810), .A2(n8763), .ZN(n14200) );
  OR2_X1 U14359 ( .A1(n14354), .A2(n14355), .ZN(n14199) );
  AND2_X1 U14360 ( .A1(n14193), .A2(n14196), .ZN(n14355) );
  AND2_X1 U14361 ( .A1(n14356), .A2(n14195), .ZN(n14354) );
  OR2_X1 U14362 ( .A1(n14357), .A2(n14358), .ZN(n14195) );
  AND2_X1 U14363 ( .A1(n14189), .A2(n14192), .ZN(n14358) );
  AND2_X1 U14364 ( .A1(n14359), .A2(n14191), .ZN(n14357) );
  OR2_X1 U14365 ( .A1(n14360), .A2(n14361), .ZN(n14191) );
  AND2_X1 U14366 ( .A1(n14185), .A2(n14188), .ZN(n14361) );
  AND2_X1 U14367 ( .A1(n14362), .A2(n14187), .ZN(n14360) );
  OR2_X1 U14368 ( .A1(n14363), .A2(n14364), .ZN(n14187) );
  AND2_X1 U14369 ( .A1(n14181), .A2(n14184), .ZN(n14364) );
  AND2_X1 U14370 ( .A1(n14365), .A2(n14183), .ZN(n14363) );
  OR2_X1 U14371 ( .A1(n14366), .A2(n14367), .ZN(n14183) );
  AND2_X1 U14372 ( .A1(n14177), .A2(n14180), .ZN(n14367) );
  AND2_X1 U14373 ( .A1(n14368), .A2(n14179), .ZN(n14366) );
  OR2_X1 U14374 ( .A1(n14369), .A2(n14370), .ZN(n14179) );
  AND2_X1 U14375 ( .A1(n14173), .A2(n14176), .ZN(n14370) );
  AND2_X1 U14376 ( .A1(n14371), .A2(n14175), .ZN(n14369) );
  OR2_X1 U14377 ( .A1(n14372), .A2(n14373), .ZN(n14175) );
  AND2_X1 U14378 ( .A1(n14169), .A2(n14172), .ZN(n14373) );
  AND2_X1 U14379 ( .A1(n14374), .A2(n14171), .ZN(n14372) );
  OR2_X1 U14380 ( .A1(n14375), .A2(n14376), .ZN(n14171) );
  AND2_X1 U14381 ( .A1(n14165), .A2(n14168), .ZN(n14376) );
  AND2_X1 U14382 ( .A1(n14377), .A2(n14378), .ZN(n14375) );
  OR2_X1 U14383 ( .A1(n14168), .A2(n14165), .ZN(n14378) );
  OR2_X1 U14384 ( .A1(n7954), .A2(n8763), .ZN(n14165) );
  OR3_X1 U14385 ( .A1(n8763), .A2(n8759), .A3(n9796), .ZN(n14168) );
  INV_X1 U14386 ( .A(n14167), .ZN(n14377) );
  OR2_X1 U14387 ( .A1(n14379), .A2(n14380), .ZN(n14167) );
  AND2_X1 U14388 ( .A1(b_8_), .A2(n14381), .ZN(n14380) );
  OR2_X1 U14389 ( .A1(n14382), .A2(n9801), .ZN(n14381) );
  AND2_X1 U14390 ( .A1(a_30_), .A2(n8755), .ZN(n14382) );
  AND2_X1 U14391 ( .A1(b_7_), .A2(n14383), .ZN(n14379) );
  OR2_X1 U14392 ( .A1(n14384), .A2(n7920), .ZN(n14383) );
  AND2_X1 U14393 ( .A1(a_31_), .A2(n8759), .ZN(n14384) );
  OR2_X1 U14394 ( .A1(n14172), .A2(n14169), .ZN(n14374) );
  XNOR2_X1 U14395 ( .A(n14385), .B(n14386), .ZN(n14169) );
  XOR2_X1 U14396 ( .A(n14387), .B(n14388), .Z(n14386) );
  OR2_X1 U14397 ( .A1(n7979), .A2(n8763), .ZN(n14172) );
  OR2_X1 U14398 ( .A1(n14176), .A2(n14173), .ZN(n14371) );
  XOR2_X1 U14399 ( .A(n14389), .B(n14390), .Z(n14173) );
  XOR2_X1 U14400 ( .A(n14391), .B(n14392), .Z(n14390) );
  OR2_X1 U14401 ( .A1(n8015), .A2(n8763), .ZN(n14176) );
  OR2_X1 U14402 ( .A1(n14180), .A2(n14177), .ZN(n14368) );
  XOR2_X1 U14403 ( .A(n14393), .B(n14394), .Z(n14177) );
  XOR2_X1 U14404 ( .A(n14395), .B(n14396), .Z(n14394) );
  OR2_X1 U14405 ( .A1(n8040), .A2(n8763), .ZN(n14180) );
  OR2_X1 U14406 ( .A1(n14184), .A2(n14181), .ZN(n14365) );
  XOR2_X1 U14407 ( .A(n14397), .B(n14398), .Z(n14181) );
  XOR2_X1 U14408 ( .A(n14399), .B(n14400), .Z(n14398) );
  OR2_X1 U14409 ( .A1(n8065), .A2(n8763), .ZN(n14184) );
  OR2_X1 U14410 ( .A1(n14188), .A2(n14185), .ZN(n14362) );
  XOR2_X1 U14411 ( .A(n14401), .B(n14402), .Z(n14185) );
  XOR2_X1 U14412 ( .A(n14403), .B(n14404), .Z(n14402) );
  OR2_X1 U14413 ( .A1(n8090), .A2(n8763), .ZN(n14188) );
  OR2_X1 U14414 ( .A1(n14192), .A2(n14189), .ZN(n14359) );
  XOR2_X1 U14415 ( .A(n14405), .B(n14406), .Z(n14189) );
  XOR2_X1 U14416 ( .A(n14407), .B(n14408), .Z(n14406) );
  OR2_X1 U14417 ( .A1(n8115), .A2(n8763), .ZN(n14192) );
  OR2_X1 U14418 ( .A1(n14196), .A2(n14193), .ZN(n14356) );
  XOR2_X1 U14419 ( .A(n14409), .B(n14410), .Z(n14193) );
  XOR2_X1 U14420 ( .A(n14411), .B(n14412), .Z(n14410) );
  OR2_X1 U14421 ( .A1(n8140), .A2(n8763), .ZN(n14196) );
  XOR2_X1 U14422 ( .A(n14413), .B(n14414), .Z(n14197) );
  XOR2_X1 U14423 ( .A(n14415), .B(n14416), .Z(n14414) );
  OR2_X1 U14424 ( .A1(n14204), .A2(n14201), .ZN(n14350) );
  XOR2_X1 U14425 ( .A(n14417), .B(n14418), .Z(n14201) );
  XOR2_X1 U14426 ( .A(n14419), .B(n14420), .Z(n14418) );
  OR2_X1 U14427 ( .A1(n8806), .A2(n8763), .ZN(n14204) );
  XOR2_X1 U14428 ( .A(n14421), .B(n14422), .Z(n14205) );
  XOR2_X1 U14429 ( .A(n14423), .B(n14424), .Z(n14422) );
  XOR2_X1 U14430 ( .A(n14425), .B(n14426), .Z(n14209) );
  XOR2_X1 U14431 ( .A(n14427), .B(n14428), .Z(n14426) );
  XOR2_X1 U14432 ( .A(n14429), .B(n14430), .Z(n14213) );
  XOR2_X1 U14433 ( .A(n14431), .B(n14432), .Z(n14430) );
  XOR2_X1 U14434 ( .A(n14433), .B(n14434), .Z(n14217) );
  XOR2_X1 U14435 ( .A(n14435), .B(n14436), .Z(n14434) );
  XOR2_X1 U14436 ( .A(n14437), .B(n14438), .Z(n14221) );
  XOR2_X1 U14437 ( .A(n14439), .B(n14440), .Z(n14438) );
  XOR2_X1 U14438 ( .A(n14441), .B(n14442), .Z(n14225) );
  XOR2_X1 U14439 ( .A(n14443), .B(n14444), .Z(n14442) );
  XOR2_X1 U14440 ( .A(n14445), .B(n14446), .Z(n14229) );
  XOR2_X1 U14441 ( .A(n14447), .B(n14448), .Z(n14446) );
  XOR2_X1 U14442 ( .A(n14449), .B(n14450), .Z(n14233) );
  XOR2_X1 U14443 ( .A(n14451), .B(n14452), .Z(n14450) );
  XOR2_X1 U14444 ( .A(n14453), .B(n14454), .Z(n14237) );
  XOR2_X1 U14445 ( .A(n14455), .B(n14456), .Z(n14454) );
  XOR2_X1 U14446 ( .A(n14457), .B(n14458), .Z(n14241) );
  XOR2_X1 U14447 ( .A(n14459), .B(n14460), .Z(n14458) );
  XOR2_X1 U14448 ( .A(n14461), .B(n14462), .Z(n14245) );
  XOR2_X1 U14449 ( .A(n14463), .B(n14464), .Z(n14462) );
  XOR2_X1 U14450 ( .A(n14465), .B(n14466), .Z(n14248) );
  XOR2_X1 U14451 ( .A(n14467), .B(n14468), .Z(n14466) );
  XOR2_X1 U14452 ( .A(n14469), .B(n14470), .Z(n14252) );
  XOR2_X1 U14453 ( .A(n14471), .B(n8504), .Z(n14470) );
  XOR2_X1 U14454 ( .A(n14472), .B(n14473), .Z(n14256) );
  XOR2_X1 U14455 ( .A(n14474), .B(n14475), .Z(n14473) );
  XOR2_X1 U14456 ( .A(n14476), .B(n14477), .Z(n14260) );
  XOR2_X1 U14457 ( .A(n14478), .B(n14479), .Z(n14477) );
  XOR2_X1 U14458 ( .A(n14480), .B(n14481), .Z(n14264) );
  XOR2_X1 U14459 ( .A(n14482), .B(n14483), .Z(n14481) );
  XOR2_X1 U14460 ( .A(n14484), .B(n14485), .Z(n14268) );
  XOR2_X1 U14461 ( .A(n14486), .B(n14487), .Z(n14485) );
  XOR2_X1 U14462 ( .A(n14488), .B(n14489), .Z(n14272) );
  XOR2_X1 U14463 ( .A(n14490), .B(n14491), .Z(n14489) );
  XOR2_X1 U14464 ( .A(n14492), .B(n14493), .Z(n14276) );
  XOR2_X1 U14465 ( .A(n14494), .B(n14495), .Z(n14493) );
  XOR2_X1 U14466 ( .A(n14496), .B(n14497), .Z(n14280) );
  XOR2_X1 U14467 ( .A(n14498), .B(n14499), .Z(n14497) );
  XOR2_X1 U14468 ( .A(n9372), .B(n14500), .Z(n14285) );
  XOR2_X1 U14469 ( .A(n9371), .B(n9370), .Z(n14500) );
  OR2_X1 U14470 ( .A1(n9248), .A2(n8759), .ZN(n9370) );
  OR2_X1 U14471 ( .A1(n14501), .A2(n14502), .ZN(n9371) );
  AND2_X1 U14472 ( .A1(n14499), .A2(n14498), .ZN(n14502) );
  AND2_X1 U14473 ( .A1(n14496), .A2(n14503), .ZN(n14501) );
  OR2_X1 U14474 ( .A1(n14498), .A2(n14499), .ZN(n14503) );
  OR2_X1 U14475 ( .A1(n8730), .A2(n8759), .ZN(n14499) );
  OR2_X1 U14476 ( .A1(n14504), .A2(n14505), .ZN(n14498) );
  AND2_X1 U14477 ( .A1(n14495), .A2(n14494), .ZN(n14505) );
  AND2_X1 U14478 ( .A1(n14492), .A2(n14506), .ZN(n14504) );
  OR2_X1 U14479 ( .A1(n14494), .A2(n14495), .ZN(n14506) );
  OR2_X1 U14480 ( .A1(n8734), .A2(n8759), .ZN(n14495) );
  OR2_X1 U14481 ( .A1(n14507), .A2(n14508), .ZN(n14494) );
  AND2_X1 U14482 ( .A1(n14491), .A2(n14490), .ZN(n14508) );
  AND2_X1 U14483 ( .A1(n14488), .A2(n14509), .ZN(n14507) );
  OR2_X1 U14484 ( .A1(n14490), .A2(n14491), .ZN(n14509) );
  OR2_X1 U14485 ( .A1(n8738), .A2(n8759), .ZN(n14491) );
  OR2_X1 U14486 ( .A1(n14510), .A2(n14511), .ZN(n14490) );
  AND2_X1 U14487 ( .A1(n14487), .A2(n14486), .ZN(n14511) );
  AND2_X1 U14488 ( .A1(n14484), .A2(n14512), .ZN(n14510) );
  OR2_X1 U14489 ( .A1(n14486), .A2(n14487), .ZN(n14512) );
  OR2_X1 U14490 ( .A1(n8742), .A2(n8759), .ZN(n14487) );
  OR2_X1 U14491 ( .A1(n14513), .A2(n14514), .ZN(n14486) );
  AND2_X1 U14492 ( .A1(n14483), .A2(n14482), .ZN(n14514) );
  AND2_X1 U14493 ( .A1(n14480), .A2(n14515), .ZN(n14513) );
  OR2_X1 U14494 ( .A1(n14482), .A2(n14483), .ZN(n14515) );
  OR2_X1 U14495 ( .A1(n8746), .A2(n8759), .ZN(n14483) );
  OR2_X1 U14496 ( .A1(n14516), .A2(n14517), .ZN(n14482) );
  AND2_X1 U14497 ( .A1(n14479), .A2(n14478), .ZN(n14517) );
  AND2_X1 U14498 ( .A1(n14476), .A2(n14518), .ZN(n14516) );
  OR2_X1 U14499 ( .A1(n14478), .A2(n14479), .ZN(n14518) );
  OR2_X1 U14500 ( .A1(n8750), .A2(n8759), .ZN(n14479) );
  OR2_X1 U14501 ( .A1(n14519), .A2(n14520), .ZN(n14478) );
  AND2_X1 U14502 ( .A1(n14475), .A2(n14474), .ZN(n14520) );
  AND2_X1 U14503 ( .A1(n14472), .A2(n14521), .ZN(n14519) );
  OR2_X1 U14504 ( .A1(n14474), .A2(n14475), .ZN(n14521) );
  OR2_X1 U14505 ( .A1(n8754), .A2(n8759), .ZN(n14475) );
  OR2_X1 U14506 ( .A1(n14522), .A2(n14523), .ZN(n14474) );
  AND2_X1 U14507 ( .A1(n8504), .A2(n14471), .ZN(n14523) );
  AND2_X1 U14508 ( .A1(n14469), .A2(n14524), .ZN(n14522) );
  OR2_X1 U14509 ( .A1(n14471), .A2(n8504), .ZN(n14524) );
  OR2_X1 U14510 ( .A1(n8758), .A2(n8759), .ZN(n8504) );
  OR2_X1 U14511 ( .A1(n14525), .A2(n14526), .ZN(n14471) );
  AND2_X1 U14512 ( .A1(n14468), .A2(n14467), .ZN(n14526) );
  AND2_X1 U14513 ( .A1(n14465), .A2(n14527), .ZN(n14525) );
  OR2_X1 U14514 ( .A1(n14467), .A2(n14468), .ZN(n14527) );
  OR2_X1 U14515 ( .A1(n8762), .A2(n8759), .ZN(n14468) );
  OR2_X1 U14516 ( .A1(n14528), .A2(n14529), .ZN(n14467) );
  AND2_X1 U14517 ( .A1(n14464), .A2(n14463), .ZN(n14529) );
  AND2_X1 U14518 ( .A1(n14461), .A2(n14530), .ZN(n14528) );
  OR2_X1 U14519 ( .A1(n14463), .A2(n14464), .ZN(n14530) );
  OR2_X1 U14520 ( .A1(n8766), .A2(n8759), .ZN(n14464) );
  OR2_X1 U14521 ( .A1(n14531), .A2(n14532), .ZN(n14463) );
  AND2_X1 U14522 ( .A1(n14460), .A2(n14459), .ZN(n14532) );
  AND2_X1 U14523 ( .A1(n14457), .A2(n14533), .ZN(n14531) );
  OR2_X1 U14524 ( .A1(n14459), .A2(n14460), .ZN(n14533) );
  OR2_X1 U14525 ( .A1(n8770), .A2(n8759), .ZN(n14460) );
  OR2_X1 U14526 ( .A1(n14534), .A2(n14535), .ZN(n14459) );
  AND2_X1 U14527 ( .A1(n14456), .A2(n14455), .ZN(n14535) );
  AND2_X1 U14528 ( .A1(n14453), .A2(n14536), .ZN(n14534) );
  OR2_X1 U14529 ( .A1(n14455), .A2(n14456), .ZN(n14536) );
  OR2_X1 U14530 ( .A1(n8774), .A2(n8759), .ZN(n14456) );
  OR2_X1 U14531 ( .A1(n14537), .A2(n14538), .ZN(n14455) );
  AND2_X1 U14532 ( .A1(n14452), .A2(n14451), .ZN(n14538) );
  AND2_X1 U14533 ( .A1(n14449), .A2(n14539), .ZN(n14537) );
  OR2_X1 U14534 ( .A1(n14451), .A2(n14452), .ZN(n14539) );
  OR2_X1 U14535 ( .A1(n8778), .A2(n8759), .ZN(n14452) );
  OR2_X1 U14536 ( .A1(n14540), .A2(n14541), .ZN(n14451) );
  AND2_X1 U14537 ( .A1(n14448), .A2(n14447), .ZN(n14541) );
  AND2_X1 U14538 ( .A1(n14445), .A2(n14542), .ZN(n14540) );
  OR2_X1 U14539 ( .A1(n14447), .A2(n14448), .ZN(n14542) );
  OR2_X1 U14540 ( .A1(n8782), .A2(n8759), .ZN(n14448) );
  OR2_X1 U14541 ( .A1(n14543), .A2(n14544), .ZN(n14447) );
  AND2_X1 U14542 ( .A1(n14444), .A2(n14443), .ZN(n14544) );
  AND2_X1 U14543 ( .A1(n14441), .A2(n14545), .ZN(n14543) );
  OR2_X1 U14544 ( .A1(n14443), .A2(n14444), .ZN(n14545) );
  OR2_X1 U14545 ( .A1(n8786), .A2(n8759), .ZN(n14444) );
  OR2_X1 U14546 ( .A1(n14546), .A2(n14547), .ZN(n14443) );
  AND2_X1 U14547 ( .A1(n14440), .A2(n14439), .ZN(n14547) );
  AND2_X1 U14548 ( .A1(n14437), .A2(n14548), .ZN(n14546) );
  OR2_X1 U14549 ( .A1(n14439), .A2(n14440), .ZN(n14548) );
  OR2_X1 U14550 ( .A1(n8790), .A2(n8759), .ZN(n14440) );
  OR2_X1 U14551 ( .A1(n14549), .A2(n14550), .ZN(n14439) );
  AND2_X1 U14552 ( .A1(n14436), .A2(n14435), .ZN(n14550) );
  AND2_X1 U14553 ( .A1(n14433), .A2(n14551), .ZN(n14549) );
  OR2_X1 U14554 ( .A1(n14435), .A2(n14436), .ZN(n14551) );
  OR2_X1 U14555 ( .A1(n8794), .A2(n8759), .ZN(n14436) );
  OR2_X1 U14556 ( .A1(n14552), .A2(n14553), .ZN(n14435) );
  AND2_X1 U14557 ( .A1(n14432), .A2(n14431), .ZN(n14553) );
  AND2_X1 U14558 ( .A1(n14429), .A2(n14554), .ZN(n14552) );
  OR2_X1 U14559 ( .A1(n14431), .A2(n14432), .ZN(n14554) );
  OR2_X1 U14560 ( .A1(n8798), .A2(n8759), .ZN(n14432) );
  OR2_X1 U14561 ( .A1(n14555), .A2(n14556), .ZN(n14431) );
  AND2_X1 U14562 ( .A1(n14428), .A2(n14427), .ZN(n14556) );
  AND2_X1 U14563 ( .A1(n14425), .A2(n14557), .ZN(n14555) );
  OR2_X1 U14564 ( .A1(n14427), .A2(n14428), .ZN(n14557) );
  OR2_X1 U14565 ( .A1(n8802), .A2(n8759), .ZN(n14428) );
  OR2_X1 U14566 ( .A1(n14558), .A2(n14559), .ZN(n14427) );
  AND2_X1 U14567 ( .A1(n14424), .A2(n14423), .ZN(n14559) );
  AND2_X1 U14568 ( .A1(n14421), .A2(n14560), .ZN(n14558) );
  OR2_X1 U14569 ( .A1(n14423), .A2(n14424), .ZN(n14560) );
  OR2_X1 U14570 ( .A1(n8806), .A2(n8759), .ZN(n14424) );
  OR2_X1 U14571 ( .A1(n14561), .A2(n14562), .ZN(n14423) );
  AND2_X1 U14572 ( .A1(n14417), .A2(n14420), .ZN(n14562) );
  AND2_X1 U14573 ( .A1(n14563), .A2(n14419), .ZN(n14561) );
  OR2_X1 U14574 ( .A1(n14564), .A2(n14565), .ZN(n14419) );
  AND2_X1 U14575 ( .A1(n14416), .A2(n14415), .ZN(n14565) );
  AND2_X1 U14576 ( .A1(n14413), .A2(n14566), .ZN(n14564) );
  OR2_X1 U14577 ( .A1(n14415), .A2(n14416), .ZN(n14566) );
  OR2_X1 U14578 ( .A1(n8140), .A2(n8759), .ZN(n14416) );
  OR2_X1 U14579 ( .A1(n14567), .A2(n14568), .ZN(n14415) );
  AND2_X1 U14580 ( .A1(n14409), .A2(n14412), .ZN(n14568) );
  AND2_X1 U14581 ( .A1(n14569), .A2(n14411), .ZN(n14567) );
  OR2_X1 U14582 ( .A1(n14570), .A2(n14571), .ZN(n14411) );
  AND2_X1 U14583 ( .A1(n14405), .A2(n14408), .ZN(n14571) );
  AND2_X1 U14584 ( .A1(n14572), .A2(n14407), .ZN(n14570) );
  OR2_X1 U14585 ( .A1(n14573), .A2(n14574), .ZN(n14407) );
  AND2_X1 U14586 ( .A1(n14401), .A2(n14404), .ZN(n14574) );
  AND2_X1 U14587 ( .A1(n14575), .A2(n14403), .ZN(n14573) );
  OR2_X1 U14588 ( .A1(n14576), .A2(n14577), .ZN(n14403) );
  AND2_X1 U14589 ( .A1(n14397), .A2(n14400), .ZN(n14577) );
  AND2_X1 U14590 ( .A1(n14578), .A2(n14399), .ZN(n14576) );
  OR2_X1 U14591 ( .A1(n14579), .A2(n14580), .ZN(n14399) );
  AND2_X1 U14592 ( .A1(n14393), .A2(n14396), .ZN(n14580) );
  AND2_X1 U14593 ( .A1(n14581), .A2(n14395), .ZN(n14579) );
  OR2_X1 U14594 ( .A1(n14582), .A2(n14583), .ZN(n14395) );
  AND2_X1 U14595 ( .A1(n14389), .A2(n14392), .ZN(n14583) );
  AND2_X1 U14596 ( .A1(n14584), .A2(n14391), .ZN(n14582) );
  OR2_X1 U14597 ( .A1(n14585), .A2(n14586), .ZN(n14391) );
  AND2_X1 U14598 ( .A1(n14385), .A2(n14388), .ZN(n14586) );
  AND2_X1 U14599 ( .A1(n14587), .A2(n14588), .ZN(n14585) );
  OR2_X1 U14600 ( .A1(n14388), .A2(n14385), .ZN(n14588) );
  OR2_X1 U14601 ( .A1(n7954), .A2(n8759), .ZN(n14385) );
  OR3_X1 U14602 ( .A1(n8759), .A2(n8755), .A3(n9796), .ZN(n14388) );
  INV_X1 U14603 ( .A(n14387), .ZN(n14587) );
  OR2_X1 U14604 ( .A1(n14589), .A2(n14590), .ZN(n14387) );
  AND2_X1 U14605 ( .A1(b_7_), .A2(n14591), .ZN(n14590) );
  OR2_X1 U14606 ( .A1(n14592), .A2(n9801), .ZN(n14591) );
  AND2_X1 U14607 ( .A1(a_30_), .A2(n8751), .ZN(n14592) );
  AND2_X1 U14608 ( .A1(b_6_), .A2(n14593), .ZN(n14589) );
  OR2_X1 U14609 ( .A1(n14594), .A2(n7920), .ZN(n14593) );
  AND2_X1 U14610 ( .A1(a_31_), .A2(n8755), .ZN(n14594) );
  OR2_X1 U14611 ( .A1(n14392), .A2(n14389), .ZN(n14584) );
  XNOR2_X1 U14612 ( .A(n14595), .B(n14596), .ZN(n14389) );
  XOR2_X1 U14613 ( .A(n14597), .B(n14598), .Z(n14596) );
  OR2_X1 U14614 ( .A1(n7979), .A2(n8759), .ZN(n14392) );
  OR2_X1 U14615 ( .A1(n14396), .A2(n14393), .ZN(n14581) );
  XOR2_X1 U14616 ( .A(n14599), .B(n14600), .Z(n14393) );
  XOR2_X1 U14617 ( .A(n14601), .B(n14602), .Z(n14600) );
  OR2_X1 U14618 ( .A1(n8015), .A2(n8759), .ZN(n14396) );
  OR2_X1 U14619 ( .A1(n14400), .A2(n14397), .ZN(n14578) );
  XOR2_X1 U14620 ( .A(n14603), .B(n14604), .Z(n14397) );
  XOR2_X1 U14621 ( .A(n14605), .B(n14606), .Z(n14604) );
  OR2_X1 U14622 ( .A1(n8040), .A2(n8759), .ZN(n14400) );
  OR2_X1 U14623 ( .A1(n14404), .A2(n14401), .ZN(n14575) );
  XOR2_X1 U14624 ( .A(n14607), .B(n14608), .Z(n14401) );
  XOR2_X1 U14625 ( .A(n14609), .B(n14610), .Z(n14608) );
  OR2_X1 U14626 ( .A1(n8065), .A2(n8759), .ZN(n14404) );
  OR2_X1 U14627 ( .A1(n14408), .A2(n14405), .ZN(n14572) );
  XOR2_X1 U14628 ( .A(n14611), .B(n14612), .Z(n14405) );
  XOR2_X1 U14629 ( .A(n14613), .B(n14614), .Z(n14612) );
  OR2_X1 U14630 ( .A1(n8090), .A2(n8759), .ZN(n14408) );
  OR2_X1 U14631 ( .A1(n14412), .A2(n14409), .ZN(n14569) );
  XOR2_X1 U14632 ( .A(n14615), .B(n14616), .Z(n14409) );
  XOR2_X1 U14633 ( .A(n14617), .B(n14618), .Z(n14616) );
  OR2_X1 U14634 ( .A1(n8115), .A2(n8759), .ZN(n14412) );
  XOR2_X1 U14635 ( .A(n14619), .B(n14620), .Z(n14413) );
  XOR2_X1 U14636 ( .A(n14621), .B(n14622), .Z(n14620) );
  OR2_X1 U14637 ( .A1(n14420), .A2(n14417), .ZN(n14563) );
  XOR2_X1 U14638 ( .A(n14623), .B(n14624), .Z(n14417) );
  XOR2_X1 U14639 ( .A(n14625), .B(n14626), .Z(n14624) );
  OR2_X1 U14640 ( .A1(n8810), .A2(n8759), .ZN(n14420) );
  XOR2_X1 U14641 ( .A(n14627), .B(n14628), .Z(n14421) );
  XOR2_X1 U14642 ( .A(n14629), .B(n14630), .Z(n14628) );
  XOR2_X1 U14643 ( .A(n14631), .B(n14632), .Z(n14425) );
  XOR2_X1 U14644 ( .A(n14633), .B(n14634), .Z(n14632) );
  XOR2_X1 U14645 ( .A(n14635), .B(n14636), .Z(n14429) );
  XOR2_X1 U14646 ( .A(n14637), .B(n14638), .Z(n14636) );
  XOR2_X1 U14647 ( .A(n14639), .B(n14640), .Z(n14433) );
  XOR2_X1 U14648 ( .A(n14641), .B(n14642), .Z(n14640) );
  XOR2_X1 U14649 ( .A(n14643), .B(n14644), .Z(n14437) );
  XOR2_X1 U14650 ( .A(n14645), .B(n14646), .Z(n14644) );
  XOR2_X1 U14651 ( .A(n14647), .B(n14648), .Z(n14441) );
  XOR2_X1 U14652 ( .A(n14649), .B(n14650), .Z(n14648) );
  XOR2_X1 U14653 ( .A(n14651), .B(n14652), .Z(n14445) );
  XOR2_X1 U14654 ( .A(n14653), .B(n14654), .Z(n14652) );
  XOR2_X1 U14655 ( .A(n14655), .B(n14656), .Z(n14449) );
  XOR2_X1 U14656 ( .A(n14657), .B(n14658), .Z(n14656) );
  XOR2_X1 U14657 ( .A(n14659), .B(n14660), .Z(n14453) );
  XOR2_X1 U14658 ( .A(n14661), .B(n14662), .Z(n14660) );
  XOR2_X1 U14659 ( .A(n14663), .B(n14664), .Z(n14457) );
  XOR2_X1 U14660 ( .A(n14665), .B(n14666), .Z(n14664) );
  XOR2_X1 U14661 ( .A(n14667), .B(n14668), .Z(n14461) );
  XOR2_X1 U14662 ( .A(n14669), .B(n14670), .Z(n14668) );
  XOR2_X1 U14663 ( .A(n14671), .B(n14672), .Z(n14465) );
  XOR2_X1 U14664 ( .A(n14673), .B(n14674), .Z(n14672) );
  XOR2_X1 U14665 ( .A(n14675), .B(n14676), .Z(n14469) );
  XOR2_X1 U14666 ( .A(n14677), .B(n14678), .Z(n14676) );
  XOR2_X1 U14667 ( .A(n14679), .B(n14680), .Z(n14472) );
  XOR2_X1 U14668 ( .A(n14681), .B(n14682), .Z(n14680) );
  XOR2_X1 U14669 ( .A(n14683), .B(n14684), .Z(n14476) );
  XOR2_X1 U14670 ( .A(n14685), .B(n8541), .Z(n14684) );
  XOR2_X1 U14671 ( .A(n14686), .B(n14687), .Z(n14480) );
  XOR2_X1 U14672 ( .A(n14688), .B(n14689), .Z(n14687) );
  XOR2_X1 U14673 ( .A(n14690), .B(n14691), .Z(n14484) );
  XOR2_X1 U14674 ( .A(n14692), .B(n14693), .Z(n14691) );
  XOR2_X1 U14675 ( .A(n14694), .B(n14695), .Z(n14488) );
  XOR2_X1 U14676 ( .A(n14696), .B(n14697), .Z(n14695) );
  XOR2_X1 U14677 ( .A(n14698), .B(n14699), .Z(n14492) );
  XOR2_X1 U14678 ( .A(n14700), .B(n14701), .Z(n14699) );
  XOR2_X1 U14679 ( .A(n14702), .B(n14703), .Z(n14496) );
  XOR2_X1 U14680 ( .A(n14704), .B(n14705), .Z(n14703) );
  XOR2_X1 U14681 ( .A(n9379), .B(n14706), .Z(n9372) );
  XOR2_X1 U14682 ( .A(n9378), .B(n9377), .Z(n14706) );
  OR2_X1 U14683 ( .A1(n8730), .A2(n8755), .ZN(n9377) );
  OR2_X1 U14684 ( .A1(n14707), .A2(n14708), .ZN(n9378) );
  AND2_X1 U14685 ( .A1(n14705), .A2(n14704), .ZN(n14708) );
  AND2_X1 U14686 ( .A1(n14702), .A2(n14709), .ZN(n14707) );
  OR2_X1 U14687 ( .A1(n14704), .A2(n14705), .ZN(n14709) );
  OR2_X1 U14688 ( .A1(n8734), .A2(n8755), .ZN(n14705) );
  OR2_X1 U14689 ( .A1(n14710), .A2(n14711), .ZN(n14704) );
  AND2_X1 U14690 ( .A1(n14701), .A2(n14700), .ZN(n14711) );
  AND2_X1 U14691 ( .A1(n14698), .A2(n14712), .ZN(n14710) );
  OR2_X1 U14692 ( .A1(n14700), .A2(n14701), .ZN(n14712) );
  OR2_X1 U14693 ( .A1(n8738), .A2(n8755), .ZN(n14701) );
  OR2_X1 U14694 ( .A1(n14713), .A2(n14714), .ZN(n14700) );
  AND2_X1 U14695 ( .A1(n14697), .A2(n14696), .ZN(n14714) );
  AND2_X1 U14696 ( .A1(n14694), .A2(n14715), .ZN(n14713) );
  OR2_X1 U14697 ( .A1(n14696), .A2(n14697), .ZN(n14715) );
  OR2_X1 U14698 ( .A1(n8742), .A2(n8755), .ZN(n14697) );
  OR2_X1 U14699 ( .A1(n14716), .A2(n14717), .ZN(n14696) );
  AND2_X1 U14700 ( .A1(n14693), .A2(n14692), .ZN(n14717) );
  AND2_X1 U14701 ( .A1(n14690), .A2(n14718), .ZN(n14716) );
  OR2_X1 U14702 ( .A1(n14692), .A2(n14693), .ZN(n14718) );
  OR2_X1 U14703 ( .A1(n8746), .A2(n8755), .ZN(n14693) );
  OR2_X1 U14704 ( .A1(n14719), .A2(n14720), .ZN(n14692) );
  AND2_X1 U14705 ( .A1(n14689), .A2(n14688), .ZN(n14720) );
  AND2_X1 U14706 ( .A1(n14686), .A2(n14721), .ZN(n14719) );
  OR2_X1 U14707 ( .A1(n14688), .A2(n14689), .ZN(n14721) );
  OR2_X1 U14708 ( .A1(n8750), .A2(n8755), .ZN(n14689) );
  OR2_X1 U14709 ( .A1(n14722), .A2(n14723), .ZN(n14688) );
  AND2_X1 U14710 ( .A1(n8541), .A2(n14685), .ZN(n14723) );
  AND2_X1 U14711 ( .A1(n14683), .A2(n14724), .ZN(n14722) );
  OR2_X1 U14712 ( .A1(n14685), .A2(n8541), .ZN(n14724) );
  OR2_X1 U14713 ( .A1(n8754), .A2(n8755), .ZN(n8541) );
  OR2_X1 U14714 ( .A1(n14725), .A2(n14726), .ZN(n14685) );
  AND2_X1 U14715 ( .A1(n14682), .A2(n14681), .ZN(n14726) );
  AND2_X1 U14716 ( .A1(n14679), .A2(n14727), .ZN(n14725) );
  OR2_X1 U14717 ( .A1(n14681), .A2(n14682), .ZN(n14727) );
  OR2_X1 U14718 ( .A1(n8758), .A2(n8755), .ZN(n14682) );
  OR2_X1 U14719 ( .A1(n14728), .A2(n14729), .ZN(n14681) );
  AND2_X1 U14720 ( .A1(n14678), .A2(n14677), .ZN(n14729) );
  AND2_X1 U14721 ( .A1(n14675), .A2(n14730), .ZN(n14728) );
  OR2_X1 U14722 ( .A1(n14677), .A2(n14678), .ZN(n14730) );
  OR2_X1 U14723 ( .A1(n8762), .A2(n8755), .ZN(n14678) );
  OR2_X1 U14724 ( .A1(n14731), .A2(n14732), .ZN(n14677) );
  AND2_X1 U14725 ( .A1(n14674), .A2(n14673), .ZN(n14732) );
  AND2_X1 U14726 ( .A1(n14671), .A2(n14733), .ZN(n14731) );
  OR2_X1 U14727 ( .A1(n14673), .A2(n14674), .ZN(n14733) );
  OR2_X1 U14728 ( .A1(n8766), .A2(n8755), .ZN(n14674) );
  OR2_X1 U14729 ( .A1(n14734), .A2(n14735), .ZN(n14673) );
  AND2_X1 U14730 ( .A1(n14670), .A2(n14669), .ZN(n14735) );
  AND2_X1 U14731 ( .A1(n14667), .A2(n14736), .ZN(n14734) );
  OR2_X1 U14732 ( .A1(n14669), .A2(n14670), .ZN(n14736) );
  OR2_X1 U14733 ( .A1(n8770), .A2(n8755), .ZN(n14670) );
  OR2_X1 U14734 ( .A1(n14737), .A2(n14738), .ZN(n14669) );
  AND2_X1 U14735 ( .A1(n14666), .A2(n14665), .ZN(n14738) );
  AND2_X1 U14736 ( .A1(n14663), .A2(n14739), .ZN(n14737) );
  OR2_X1 U14737 ( .A1(n14665), .A2(n14666), .ZN(n14739) );
  OR2_X1 U14738 ( .A1(n8774), .A2(n8755), .ZN(n14666) );
  OR2_X1 U14739 ( .A1(n14740), .A2(n14741), .ZN(n14665) );
  AND2_X1 U14740 ( .A1(n14662), .A2(n14661), .ZN(n14741) );
  AND2_X1 U14741 ( .A1(n14659), .A2(n14742), .ZN(n14740) );
  OR2_X1 U14742 ( .A1(n14661), .A2(n14662), .ZN(n14742) );
  OR2_X1 U14743 ( .A1(n8778), .A2(n8755), .ZN(n14662) );
  OR2_X1 U14744 ( .A1(n14743), .A2(n14744), .ZN(n14661) );
  AND2_X1 U14745 ( .A1(n14658), .A2(n14657), .ZN(n14744) );
  AND2_X1 U14746 ( .A1(n14655), .A2(n14745), .ZN(n14743) );
  OR2_X1 U14747 ( .A1(n14657), .A2(n14658), .ZN(n14745) );
  OR2_X1 U14748 ( .A1(n8782), .A2(n8755), .ZN(n14658) );
  OR2_X1 U14749 ( .A1(n14746), .A2(n14747), .ZN(n14657) );
  AND2_X1 U14750 ( .A1(n14654), .A2(n14653), .ZN(n14747) );
  AND2_X1 U14751 ( .A1(n14651), .A2(n14748), .ZN(n14746) );
  OR2_X1 U14752 ( .A1(n14653), .A2(n14654), .ZN(n14748) );
  OR2_X1 U14753 ( .A1(n8786), .A2(n8755), .ZN(n14654) );
  OR2_X1 U14754 ( .A1(n14749), .A2(n14750), .ZN(n14653) );
  AND2_X1 U14755 ( .A1(n14650), .A2(n14649), .ZN(n14750) );
  AND2_X1 U14756 ( .A1(n14647), .A2(n14751), .ZN(n14749) );
  OR2_X1 U14757 ( .A1(n14649), .A2(n14650), .ZN(n14751) );
  OR2_X1 U14758 ( .A1(n8790), .A2(n8755), .ZN(n14650) );
  OR2_X1 U14759 ( .A1(n14752), .A2(n14753), .ZN(n14649) );
  AND2_X1 U14760 ( .A1(n14646), .A2(n14645), .ZN(n14753) );
  AND2_X1 U14761 ( .A1(n14643), .A2(n14754), .ZN(n14752) );
  OR2_X1 U14762 ( .A1(n14645), .A2(n14646), .ZN(n14754) );
  OR2_X1 U14763 ( .A1(n8794), .A2(n8755), .ZN(n14646) );
  OR2_X1 U14764 ( .A1(n14755), .A2(n14756), .ZN(n14645) );
  AND2_X1 U14765 ( .A1(n14642), .A2(n14641), .ZN(n14756) );
  AND2_X1 U14766 ( .A1(n14639), .A2(n14757), .ZN(n14755) );
  OR2_X1 U14767 ( .A1(n14641), .A2(n14642), .ZN(n14757) );
  OR2_X1 U14768 ( .A1(n8798), .A2(n8755), .ZN(n14642) );
  OR2_X1 U14769 ( .A1(n14758), .A2(n14759), .ZN(n14641) );
  AND2_X1 U14770 ( .A1(n14638), .A2(n14637), .ZN(n14759) );
  AND2_X1 U14771 ( .A1(n14635), .A2(n14760), .ZN(n14758) );
  OR2_X1 U14772 ( .A1(n14637), .A2(n14638), .ZN(n14760) );
  OR2_X1 U14773 ( .A1(n8802), .A2(n8755), .ZN(n14638) );
  OR2_X1 U14774 ( .A1(n14761), .A2(n14762), .ZN(n14637) );
  AND2_X1 U14775 ( .A1(n14634), .A2(n14633), .ZN(n14762) );
  AND2_X1 U14776 ( .A1(n14631), .A2(n14763), .ZN(n14761) );
  OR2_X1 U14777 ( .A1(n14633), .A2(n14634), .ZN(n14763) );
  OR2_X1 U14778 ( .A1(n8806), .A2(n8755), .ZN(n14634) );
  OR2_X1 U14779 ( .A1(n14764), .A2(n14765), .ZN(n14633) );
  AND2_X1 U14780 ( .A1(n14630), .A2(n14629), .ZN(n14765) );
  AND2_X1 U14781 ( .A1(n14627), .A2(n14766), .ZN(n14764) );
  OR2_X1 U14782 ( .A1(n14629), .A2(n14630), .ZN(n14766) );
  OR2_X1 U14783 ( .A1(n8810), .A2(n8755), .ZN(n14630) );
  OR2_X1 U14784 ( .A1(n14767), .A2(n14768), .ZN(n14629) );
  AND2_X1 U14785 ( .A1(n14623), .A2(n14626), .ZN(n14768) );
  AND2_X1 U14786 ( .A1(n14769), .A2(n14625), .ZN(n14767) );
  OR2_X1 U14787 ( .A1(n14770), .A2(n14771), .ZN(n14625) );
  AND2_X1 U14788 ( .A1(n14622), .A2(n14621), .ZN(n14771) );
  AND2_X1 U14789 ( .A1(n14619), .A2(n14772), .ZN(n14770) );
  OR2_X1 U14790 ( .A1(n14621), .A2(n14622), .ZN(n14772) );
  OR2_X1 U14791 ( .A1(n8115), .A2(n8755), .ZN(n14622) );
  OR2_X1 U14792 ( .A1(n14773), .A2(n14774), .ZN(n14621) );
  AND2_X1 U14793 ( .A1(n14615), .A2(n14618), .ZN(n14774) );
  AND2_X1 U14794 ( .A1(n14775), .A2(n14617), .ZN(n14773) );
  OR2_X1 U14795 ( .A1(n14776), .A2(n14777), .ZN(n14617) );
  AND2_X1 U14796 ( .A1(n14611), .A2(n14614), .ZN(n14777) );
  AND2_X1 U14797 ( .A1(n14778), .A2(n14613), .ZN(n14776) );
  OR2_X1 U14798 ( .A1(n14779), .A2(n14780), .ZN(n14613) );
  AND2_X1 U14799 ( .A1(n14607), .A2(n14610), .ZN(n14780) );
  AND2_X1 U14800 ( .A1(n14781), .A2(n14609), .ZN(n14779) );
  OR2_X1 U14801 ( .A1(n14782), .A2(n14783), .ZN(n14609) );
  AND2_X1 U14802 ( .A1(n14603), .A2(n14606), .ZN(n14783) );
  AND2_X1 U14803 ( .A1(n14784), .A2(n14605), .ZN(n14782) );
  OR2_X1 U14804 ( .A1(n14785), .A2(n14786), .ZN(n14605) );
  AND2_X1 U14805 ( .A1(n14599), .A2(n14602), .ZN(n14786) );
  AND2_X1 U14806 ( .A1(n14787), .A2(n14601), .ZN(n14785) );
  OR2_X1 U14807 ( .A1(n14788), .A2(n14789), .ZN(n14601) );
  AND2_X1 U14808 ( .A1(n14595), .A2(n14598), .ZN(n14789) );
  AND2_X1 U14809 ( .A1(n14790), .A2(n14791), .ZN(n14788) );
  OR2_X1 U14810 ( .A1(n14598), .A2(n14595), .ZN(n14791) );
  OR2_X1 U14811 ( .A1(n7954), .A2(n8755), .ZN(n14595) );
  OR3_X1 U14812 ( .A1(n8755), .A2(n8751), .A3(n9796), .ZN(n14598) );
  INV_X1 U14813 ( .A(n14597), .ZN(n14790) );
  OR2_X1 U14814 ( .A1(n14792), .A2(n14793), .ZN(n14597) );
  AND2_X1 U14815 ( .A1(b_6_), .A2(n14794), .ZN(n14793) );
  OR2_X1 U14816 ( .A1(n14795), .A2(n9801), .ZN(n14794) );
  AND2_X1 U14817 ( .A1(a_30_), .A2(n8747), .ZN(n14795) );
  AND2_X1 U14818 ( .A1(b_5_), .A2(n14796), .ZN(n14792) );
  OR2_X1 U14819 ( .A1(n14797), .A2(n7920), .ZN(n14796) );
  AND2_X1 U14820 ( .A1(a_31_), .A2(n8751), .ZN(n14797) );
  OR2_X1 U14821 ( .A1(n14602), .A2(n14599), .ZN(n14787) );
  XNOR2_X1 U14822 ( .A(n14798), .B(n14799), .ZN(n14599) );
  XOR2_X1 U14823 ( .A(n14800), .B(n14801), .Z(n14799) );
  OR2_X1 U14824 ( .A1(n7979), .A2(n8755), .ZN(n14602) );
  OR2_X1 U14825 ( .A1(n14606), .A2(n14603), .ZN(n14784) );
  XOR2_X1 U14826 ( .A(n14802), .B(n14803), .Z(n14603) );
  XOR2_X1 U14827 ( .A(n14804), .B(n14805), .Z(n14803) );
  OR2_X1 U14828 ( .A1(n8015), .A2(n8755), .ZN(n14606) );
  OR2_X1 U14829 ( .A1(n14610), .A2(n14607), .ZN(n14781) );
  XOR2_X1 U14830 ( .A(n14806), .B(n14807), .Z(n14607) );
  XOR2_X1 U14831 ( .A(n14808), .B(n14809), .Z(n14807) );
  OR2_X1 U14832 ( .A1(n8040), .A2(n8755), .ZN(n14610) );
  OR2_X1 U14833 ( .A1(n14614), .A2(n14611), .ZN(n14778) );
  XOR2_X1 U14834 ( .A(n14810), .B(n14811), .Z(n14611) );
  XOR2_X1 U14835 ( .A(n14812), .B(n14813), .Z(n14811) );
  OR2_X1 U14836 ( .A1(n8065), .A2(n8755), .ZN(n14614) );
  OR2_X1 U14837 ( .A1(n14618), .A2(n14615), .ZN(n14775) );
  XOR2_X1 U14838 ( .A(n14814), .B(n14815), .Z(n14615) );
  XOR2_X1 U14839 ( .A(n14816), .B(n14817), .Z(n14815) );
  OR2_X1 U14840 ( .A1(n8090), .A2(n8755), .ZN(n14618) );
  XOR2_X1 U14841 ( .A(n14818), .B(n14819), .Z(n14619) );
  XOR2_X1 U14842 ( .A(n14820), .B(n14821), .Z(n14819) );
  OR2_X1 U14843 ( .A1(n14626), .A2(n14623), .ZN(n14769) );
  XOR2_X1 U14844 ( .A(n14822), .B(n14823), .Z(n14623) );
  XOR2_X1 U14845 ( .A(n14824), .B(n14825), .Z(n14823) );
  OR2_X1 U14846 ( .A1(n8140), .A2(n8755), .ZN(n14626) );
  XOR2_X1 U14847 ( .A(n14826), .B(n14827), .Z(n14627) );
  XOR2_X1 U14848 ( .A(n14828), .B(n14829), .Z(n14827) );
  XOR2_X1 U14849 ( .A(n14830), .B(n14831), .Z(n14631) );
  XOR2_X1 U14850 ( .A(n14832), .B(n14833), .Z(n14831) );
  XOR2_X1 U14851 ( .A(n14834), .B(n14835), .Z(n14635) );
  XOR2_X1 U14852 ( .A(n14836), .B(n14837), .Z(n14835) );
  XOR2_X1 U14853 ( .A(n14838), .B(n14839), .Z(n14639) );
  XOR2_X1 U14854 ( .A(n14840), .B(n14841), .Z(n14839) );
  XOR2_X1 U14855 ( .A(n14842), .B(n14843), .Z(n14643) );
  XOR2_X1 U14856 ( .A(n14844), .B(n14845), .Z(n14843) );
  XOR2_X1 U14857 ( .A(n14846), .B(n14847), .Z(n14647) );
  XOR2_X1 U14858 ( .A(n14848), .B(n14849), .Z(n14847) );
  XOR2_X1 U14859 ( .A(n14850), .B(n14851), .Z(n14651) );
  XOR2_X1 U14860 ( .A(n14852), .B(n14853), .Z(n14851) );
  XOR2_X1 U14861 ( .A(n14854), .B(n14855), .Z(n14655) );
  XOR2_X1 U14862 ( .A(n14856), .B(n14857), .Z(n14855) );
  XOR2_X1 U14863 ( .A(n14858), .B(n14859), .Z(n14659) );
  XOR2_X1 U14864 ( .A(n14860), .B(n14861), .Z(n14859) );
  XOR2_X1 U14865 ( .A(n14862), .B(n14863), .Z(n14663) );
  XOR2_X1 U14866 ( .A(n14864), .B(n14865), .Z(n14863) );
  XOR2_X1 U14867 ( .A(n14866), .B(n14867), .Z(n14667) );
  XOR2_X1 U14868 ( .A(n14868), .B(n14869), .Z(n14867) );
  XOR2_X1 U14869 ( .A(n14870), .B(n14871), .Z(n14671) );
  XOR2_X1 U14870 ( .A(n14872), .B(n14873), .Z(n14871) );
  XOR2_X1 U14871 ( .A(n14874), .B(n14875), .Z(n14675) );
  XOR2_X1 U14872 ( .A(n14876), .B(n14877), .Z(n14875) );
  XOR2_X1 U14873 ( .A(n14878), .B(n14879), .Z(n14679) );
  XOR2_X1 U14874 ( .A(n14880), .B(n14881), .Z(n14879) );
  XOR2_X1 U14875 ( .A(n14882), .B(n14883), .Z(n14683) );
  XOR2_X1 U14876 ( .A(n14884), .B(n14885), .Z(n14883) );
  XOR2_X1 U14877 ( .A(n14886), .B(n14887), .Z(n14686) );
  XOR2_X1 U14878 ( .A(n14888), .B(n14889), .Z(n14887) );
  XOR2_X1 U14879 ( .A(n14890), .B(n14891), .Z(n14690) );
  XOR2_X1 U14880 ( .A(n14892), .B(n8567), .Z(n14891) );
  XOR2_X1 U14881 ( .A(n14893), .B(n14894), .Z(n14694) );
  XOR2_X1 U14882 ( .A(n14895), .B(n14896), .Z(n14894) );
  XOR2_X1 U14883 ( .A(n14897), .B(n14898), .Z(n14698) );
  XOR2_X1 U14884 ( .A(n14899), .B(n14900), .Z(n14898) );
  XOR2_X1 U14885 ( .A(n14901), .B(n14902), .Z(n14702) );
  XOR2_X1 U14886 ( .A(n14903), .B(n14904), .Z(n14902) );
  XOR2_X1 U14887 ( .A(n9386), .B(n14905), .Z(n9379) );
  XOR2_X1 U14888 ( .A(n9385), .B(n9384), .Z(n14905) );
  OR2_X1 U14889 ( .A1(n8734), .A2(n8751), .ZN(n9384) );
  OR2_X1 U14890 ( .A1(n14906), .A2(n14907), .ZN(n9385) );
  AND2_X1 U14891 ( .A1(n14904), .A2(n14903), .ZN(n14907) );
  AND2_X1 U14892 ( .A1(n14901), .A2(n14908), .ZN(n14906) );
  OR2_X1 U14893 ( .A1(n14903), .A2(n14904), .ZN(n14908) );
  OR2_X1 U14894 ( .A1(n8738), .A2(n8751), .ZN(n14904) );
  OR2_X1 U14895 ( .A1(n14909), .A2(n14910), .ZN(n14903) );
  AND2_X1 U14896 ( .A1(n14900), .A2(n14899), .ZN(n14910) );
  AND2_X1 U14897 ( .A1(n14897), .A2(n14911), .ZN(n14909) );
  OR2_X1 U14898 ( .A1(n14899), .A2(n14900), .ZN(n14911) );
  OR2_X1 U14899 ( .A1(n8742), .A2(n8751), .ZN(n14900) );
  OR2_X1 U14900 ( .A1(n14912), .A2(n14913), .ZN(n14899) );
  AND2_X1 U14901 ( .A1(n14896), .A2(n14895), .ZN(n14913) );
  AND2_X1 U14902 ( .A1(n14893), .A2(n14914), .ZN(n14912) );
  OR2_X1 U14903 ( .A1(n14895), .A2(n14896), .ZN(n14914) );
  OR2_X1 U14904 ( .A1(n8746), .A2(n8751), .ZN(n14896) );
  OR2_X1 U14905 ( .A1(n14915), .A2(n14916), .ZN(n14895) );
  AND2_X1 U14906 ( .A1(n8567), .A2(n14892), .ZN(n14916) );
  AND2_X1 U14907 ( .A1(n14890), .A2(n14917), .ZN(n14915) );
  OR2_X1 U14908 ( .A1(n14892), .A2(n8567), .ZN(n14917) );
  OR2_X1 U14909 ( .A1(n8750), .A2(n8751), .ZN(n8567) );
  OR2_X1 U14910 ( .A1(n14918), .A2(n14919), .ZN(n14892) );
  AND2_X1 U14911 ( .A1(n14889), .A2(n14888), .ZN(n14919) );
  AND2_X1 U14912 ( .A1(n14886), .A2(n14920), .ZN(n14918) );
  OR2_X1 U14913 ( .A1(n14888), .A2(n14889), .ZN(n14920) );
  OR2_X1 U14914 ( .A1(n8754), .A2(n8751), .ZN(n14889) );
  OR2_X1 U14915 ( .A1(n14921), .A2(n14922), .ZN(n14888) );
  AND2_X1 U14916 ( .A1(n14885), .A2(n14884), .ZN(n14922) );
  AND2_X1 U14917 ( .A1(n14882), .A2(n14923), .ZN(n14921) );
  OR2_X1 U14918 ( .A1(n14884), .A2(n14885), .ZN(n14923) );
  OR2_X1 U14919 ( .A1(n8758), .A2(n8751), .ZN(n14885) );
  OR2_X1 U14920 ( .A1(n14924), .A2(n14925), .ZN(n14884) );
  AND2_X1 U14921 ( .A1(n14881), .A2(n14880), .ZN(n14925) );
  AND2_X1 U14922 ( .A1(n14878), .A2(n14926), .ZN(n14924) );
  OR2_X1 U14923 ( .A1(n14880), .A2(n14881), .ZN(n14926) );
  OR2_X1 U14924 ( .A1(n8762), .A2(n8751), .ZN(n14881) );
  OR2_X1 U14925 ( .A1(n14927), .A2(n14928), .ZN(n14880) );
  AND2_X1 U14926 ( .A1(n14877), .A2(n14876), .ZN(n14928) );
  AND2_X1 U14927 ( .A1(n14874), .A2(n14929), .ZN(n14927) );
  OR2_X1 U14928 ( .A1(n14876), .A2(n14877), .ZN(n14929) );
  OR2_X1 U14929 ( .A1(n8766), .A2(n8751), .ZN(n14877) );
  OR2_X1 U14930 ( .A1(n14930), .A2(n14931), .ZN(n14876) );
  AND2_X1 U14931 ( .A1(n14873), .A2(n14872), .ZN(n14931) );
  AND2_X1 U14932 ( .A1(n14870), .A2(n14932), .ZN(n14930) );
  OR2_X1 U14933 ( .A1(n14872), .A2(n14873), .ZN(n14932) );
  OR2_X1 U14934 ( .A1(n8770), .A2(n8751), .ZN(n14873) );
  OR2_X1 U14935 ( .A1(n14933), .A2(n14934), .ZN(n14872) );
  AND2_X1 U14936 ( .A1(n14869), .A2(n14868), .ZN(n14934) );
  AND2_X1 U14937 ( .A1(n14866), .A2(n14935), .ZN(n14933) );
  OR2_X1 U14938 ( .A1(n14868), .A2(n14869), .ZN(n14935) );
  OR2_X1 U14939 ( .A1(n8774), .A2(n8751), .ZN(n14869) );
  OR2_X1 U14940 ( .A1(n14936), .A2(n14937), .ZN(n14868) );
  AND2_X1 U14941 ( .A1(n14865), .A2(n14864), .ZN(n14937) );
  AND2_X1 U14942 ( .A1(n14862), .A2(n14938), .ZN(n14936) );
  OR2_X1 U14943 ( .A1(n14864), .A2(n14865), .ZN(n14938) );
  OR2_X1 U14944 ( .A1(n8778), .A2(n8751), .ZN(n14865) );
  OR2_X1 U14945 ( .A1(n14939), .A2(n14940), .ZN(n14864) );
  AND2_X1 U14946 ( .A1(n14861), .A2(n14860), .ZN(n14940) );
  AND2_X1 U14947 ( .A1(n14858), .A2(n14941), .ZN(n14939) );
  OR2_X1 U14948 ( .A1(n14860), .A2(n14861), .ZN(n14941) );
  OR2_X1 U14949 ( .A1(n8782), .A2(n8751), .ZN(n14861) );
  OR2_X1 U14950 ( .A1(n14942), .A2(n14943), .ZN(n14860) );
  AND2_X1 U14951 ( .A1(n14857), .A2(n14856), .ZN(n14943) );
  AND2_X1 U14952 ( .A1(n14854), .A2(n14944), .ZN(n14942) );
  OR2_X1 U14953 ( .A1(n14856), .A2(n14857), .ZN(n14944) );
  OR2_X1 U14954 ( .A1(n8786), .A2(n8751), .ZN(n14857) );
  OR2_X1 U14955 ( .A1(n14945), .A2(n14946), .ZN(n14856) );
  AND2_X1 U14956 ( .A1(n14853), .A2(n14852), .ZN(n14946) );
  AND2_X1 U14957 ( .A1(n14850), .A2(n14947), .ZN(n14945) );
  OR2_X1 U14958 ( .A1(n14852), .A2(n14853), .ZN(n14947) );
  OR2_X1 U14959 ( .A1(n8790), .A2(n8751), .ZN(n14853) );
  OR2_X1 U14960 ( .A1(n14948), .A2(n14949), .ZN(n14852) );
  AND2_X1 U14961 ( .A1(n14849), .A2(n14848), .ZN(n14949) );
  AND2_X1 U14962 ( .A1(n14846), .A2(n14950), .ZN(n14948) );
  OR2_X1 U14963 ( .A1(n14848), .A2(n14849), .ZN(n14950) );
  OR2_X1 U14964 ( .A1(n8794), .A2(n8751), .ZN(n14849) );
  OR2_X1 U14965 ( .A1(n14951), .A2(n14952), .ZN(n14848) );
  AND2_X1 U14966 ( .A1(n14845), .A2(n14844), .ZN(n14952) );
  AND2_X1 U14967 ( .A1(n14842), .A2(n14953), .ZN(n14951) );
  OR2_X1 U14968 ( .A1(n14844), .A2(n14845), .ZN(n14953) );
  OR2_X1 U14969 ( .A1(n8798), .A2(n8751), .ZN(n14845) );
  OR2_X1 U14970 ( .A1(n14954), .A2(n14955), .ZN(n14844) );
  AND2_X1 U14971 ( .A1(n14841), .A2(n14840), .ZN(n14955) );
  AND2_X1 U14972 ( .A1(n14838), .A2(n14956), .ZN(n14954) );
  OR2_X1 U14973 ( .A1(n14840), .A2(n14841), .ZN(n14956) );
  OR2_X1 U14974 ( .A1(n8802), .A2(n8751), .ZN(n14841) );
  OR2_X1 U14975 ( .A1(n14957), .A2(n14958), .ZN(n14840) );
  AND2_X1 U14976 ( .A1(n14837), .A2(n14836), .ZN(n14958) );
  AND2_X1 U14977 ( .A1(n14834), .A2(n14959), .ZN(n14957) );
  OR2_X1 U14978 ( .A1(n14836), .A2(n14837), .ZN(n14959) );
  OR2_X1 U14979 ( .A1(n8806), .A2(n8751), .ZN(n14837) );
  OR2_X1 U14980 ( .A1(n14960), .A2(n14961), .ZN(n14836) );
  AND2_X1 U14981 ( .A1(n14833), .A2(n14832), .ZN(n14961) );
  AND2_X1 U14982 ( .A1(n14830), .A2(n14962), .ZN(n14960) );
  OR2_X1 U14983 ( .A1(n14832), .A2(n14833), .ZN(n14962) );
  OR2_X1 U14984 ( .A1(n8810), .A2(n8751), .ZN(n14833) );
  OR2_X1 U14985 ( .A1(n14963), .A2(n14964), .ZN(n14832) );
  AND2_X1 U14986 ( .A1(n14829), .A2(n14828), .ZN(n14964) );
  AND2_X1 U14987 ( .A1(n14826), .A2(n14965), .ZN(n14963) );
  OR2_X1 U14988 ( .A1(n14828), .A2(n14829), .ZN(n14965) );
  OR2_X1 U14989 ( .A1(n8140), .A2(n8751), .ZN(n14829) );
  OR2_X1 U14990 ( .A1(n14966), .A2(n14967), .ZN(n14828) );
  AND2_X1 U14991 ( .A1(n14822), .A2(n14825), .ZN(n14967) );
  AND2_X1 U14992 ( .A1(n14968), .A2(n14824), .ZN(n14966) );
  OR2_X1 U14993 ( .A1(n14969), .A2(n14970), .ZN(n14824) );
  AND2_X1 U14994 ( .A1(n14821), .A2(n14820), .ZN(n14970) );
  AND2_X1 U14995 ( .A1(n14818), .A2(n14971), .ZN(n14969) );
  OR2_X1 U14996 ( .A1(n14820), .A2(n14821), .ZN(n14971) );
  OR2_X1 U14997 ( .A1(n8090), .A2(n8751), .ZN(n14821) );
  OR2_X1 U14998 ( .A1(n14972), .A2(n14973), .ZN(n14820) );
  AND2_X1 U14999 ( .A1(n14814), .A2(n14817), .ZN(n14973) );
  AND2_X1 U15000 ( .A1(n14974), .A2(n14816), .ZN(n14972) );
  OR2_X1 U15001 ( .A1(n14975), .A2(n14976), .ZN(n14816) );
  AND2_X1 U15002 ( .A1(n14810), .A2(n14813), .ZN(n14976) );
  AND2_X1 U15003 ( .A1(n14977), .A2(n14812), .ZN(n14975) );
  OR2_X1 U15004 ( .A1(n14978), .A2(n14979), .ZN(n14812) );
  AND2_X1 U15005 ( .A1(n14806), .A2(n14809), .ZN(n14979) );
  AND2_X1 U15006 ( .A1(n14980), .A2(n14808), .ZN(n14978) );
  OR2_X1 U15007 ( .A1(n14981), .A2(n14982), .ZN(n14808) );
  AND2_X1 U15008 ( .A1(n14802), .A2(n14805), .ZN(n14982) );
  AND2_X1 U15009 ( .A1(n14983), .A2(n14804), .ZN(n14981) );
  OR2_X1 U15010 ( .A1(n14984), .A2(n14985), .ZN(n14804) );
  AND2_X1 U15011 ( .A1(n14798), .A2(n14801), .ZN(n14985) );
  AND2_X1 U15012 ( .A1(n14986), .A2(n14987), .ZN(n14984) );
  OR2_X1 U15013 ( .A1(n14801), .A2(n14798), .ZN(n14987) );
  OR2_X1 U15014 ( .A1(n7954), .A2(n8751), .ZN(n14798) );
  OR3_X1 U15015 ( .A1(n8751), .A2(n8747), .A3(n9796), .ZN(n14801) );
  INV_X1 U15016 ( .A(n14800), .ZN(n14986) );
  OR2_X1 U15017 ( .A1(n14988), .A2(n14989), .ZN(n14800) );
  AND2_X1 U15018 ( .A1(b_5_), .A2(n14990), .ZN(n14989) );
  OR2_X1 U15019 ( .A1(n14991), .A2(n9801), .ZN(n14990) );
  AND2_X1 U15020 ( .A1(a_30_), .A2(n8743), .ZN(n14991) );
  AND2_X1 U15021 ( .A1(b_4_), .A2(n14992), .ZN(n14988) );
  OR2_X1 U15022 ( .A1(n14993), .A2(n7920), .ZN(n14992) );
  AND2_X1 U15023 ( .A1(a_31_), .A2(n8747), .ZN(n14993) );
  OR2_X1 U15024 ( .A1(n14805), .A2(n14802), .ZN(n14983) );
  XNOR2_X1 U15025 ( .A(n14994), .B(n14995), .ZN(n14802) );
  XOR2_X1 U15026 ( .A(n14996), .B(n14997), .Z(n14995) );
  OR2_X1 U15027 ( .A1(n7979), .A2(n8751), .ZN(n14805) );
  OR2_X1 U15028 ( .A1(n14809), .A2(n14806), .ZN(n14980) );
  XOR2_X1 U15029 ( .A(n14998), .B(n14999), .Z(n14806) );
  XOR2_X1 U15030 ( .A(n15000), .B(n15001), .Z(n14999) );
  OR2_X1 U15031 ( .A1(n8015), .A2(n8751), .ZN(n14809) );
  OR2_X1 U15032 ( .A1(n14813), .A2(n14810), .ZN(n14977) );
  XOR2_X1 U15033 ( .A(n15002), .B(n15003), .Z(n14810) );
  XOR2_X1 U15034 ( .A(n15004), .B(n15005), .Z(n15003) );
  OR2_X1 U15035 ( .A1(n8040), .A2(n8751), .ZN(n14813) );
  OR2_X1 U15036 ( .A1(n14817), .A2(n14814), .ZN(n14974) );
  XOR2_X1 U15037 ( .A(n15006), .B(n15007), .Z(n14814) );
  XOR2_X1 U15038 ( .A(n15008), .B(n15009), .Z(n15007) );
  OR2_X1 U15039 ( .A1(n8065), .A2(n8751), .ZN(n14817) );
  XOR2_X1 U15040 ( .A(n15010), .B(n15011), .Z(n14818) );
  XOR2_X1 U15041 ( .A(n15012), .B(n15013), .Z(n15011) );
  OR2_X1 U15042 ( .A1(n14825), .A2(n14822), .ZN(n14968) );
  XOR2_X1 U15043 ( .A(n15014), .B(n15015), .Z(n14822) );
  XOR2_X1 U15044 ( .A(n15016), .B(n15017), .Z(n15015) );
  OR2_X1 U15045 ( .A1(n8115), .A2(n8751), .ZN(n14825) );
  XOR2_X1 U15046 ( .A(n15018), .B(n15019), .Z(n14826) );
  XOR2_X1 U15047 ( .A(n15020), .B(n15021), .Z(n15019) );
  XOR2_X1 U15048 ( .A(n15022), .B(n15023), .Z(n14830) );
  XOR2_X1 U15049 ( .A(n15024), .B(n15025), .Z(n15023) );
  XOR2_X1 U15050 ( .A(n15026), .B(n15027), .Z(n14834) );
  XOR2_X1 U15051 ( .A(n15028), .B(n15029), .Z(n15027) );
  XOR2_X1 U15052 ( .A(n15030), .B(n15031), .Z(n14838) );
  XOR2_X1 U15053 ( .A(n15032), .B(n15033), .Z(n15031) );
  XOR2_X1 U15054 ( .A(n15034), .B(n15035), .Z(n14842) );
  XOR2_X1 U15055 ( .A(n15036), .B(n15037), .Z(n15035) );
  XOR2_X1 U15056 ( .A(n15038), .B(n15039), .Z(n14846) );
  XOR2_X1 U15057 ( .A(n15040), .B(n15041), .Z(n15039) );
  XOR2_X1 U15058 ( .A(n15042), .B(n15043), .Z(n14850) );
  XOR2_X1 U15059 ( .A(n15044), .B(n15045), .Z(n15043) );
  XOR2_X1 U15060 ( .A(n15046), .B(n15047), .Z(n14854) );
  XOR2_X1 U15061 ( .A(n15048), .B(n15049), .Z(n15047) );
  XOR2_X1 U15062 ( .A(n15050), .B(n15051), .Z(n14858) );
  XOR2_X1 U15063 ( .A(n15052), .B(n15053), .Z(n15051) );
  XOR2_X1 U15064 ( .A(n15054), .B(n15055), .Z(n14862) );
  XOR2_X1 U15065 ( .A(n15056), .B(n15057), .Z(n15055) );
  XOR2_X1 U15066 ( .A(n15058), .B(n15059), .Z(n14866) );
  XOR2_X1 U15067 ( .A(n15060), .B(n15061), .Z(n15059) );
  XOR2_X1 U15068 ( .A(n15062), .B(n15063), .Z(n14870) );
  XOR2_X1 U15069 ( .A(n15064), .B(n15065), .Z(n15063) );
  XOR2_X1 U15070 ( .A(n15066), .B(n15067), .Z(n14874) );
  XOR2_X1 U15071 ( .A(n15068), .B(n15069), .Z(n15067) );
  XOR2_X1 U15072 ( .A(n15070), .B(n15071), .Z(n14878) );
  XOR2_X1 U15073 ( .A(n15072), .B(n15073), .Z(n15071) );
  XOR2_X1 U15074 ( .A(n15074), .B(n15075), .Z(n14882) );
  XOR2_X1 U15075 ( .A(n15076), .B(n15077), .Z(n15075) );
  XOR2_X1 U15076 ( .A(n15078), .B(n15079), .Z(n14886) );
  XOR2_X1 U15077 ( .A(n15080), .B(n15081), .Z(n15079) );
  XOR2_X1 U15078 ( .A(n15082), .B(n15083), .Z(n14890) );
  XOR2_X1 U15079 ( .A(n15084), .B(n15085), .Z(n15083) );
  XOR2_X1 U15080 ( .A(n15086), .B(n15087), .Z(n14893) );
  XOR2_X1 U15081 ( .A(n15088), .B(n15089), .Z(n15087) );
  XOR2_X1 U15082 ( .A(n15090), .B(n15091), .Z(n14897) );
  XOR2_X1 U15083 ( .A(n15092), .B(n8593), .Z(n15091) );
  XOR2_X1 U15084 ( .A(n15093), .B(n15094), .Z(n14901) );
  XOR2_X1 U15085 ( .A(n15095), .B(n15096), .Z(n15094) );
  XOR2_X1 U15086 ( .A(n9393), .B(n15097), .Z(n9386) );
  XOR2_X1 U15087 ( .A(n9392), .B(n9391), .Z(n15097) );
  OR2_X1 U15088 ( .A1(n8738), .A2(n8747), .ZN(n9391) );
  OR2_X1 U15089 ( .A1(n15098), .A2(n15099), .ZN(n9392) );
  AND2_X1 U15090 ( .A1(n15096), .A2(n15095), .ZN(n15099) );
  AND2_X1 U15091 ( .A1(n15093), .A2(n15100), .ZN(n15098) );
  OR2_X1 U15092 ( .A1(n15095), .A2(n15096), .ZN(n15100) );
  OR2_X1 U15093 ( .A1(n8742), .A2(n8747), .ZN(n15096) );
  OR2_X1 U15094 ( .A1(n15101), .A2(n15102), .ZN(n15095) );
  AND2_X1 U15095 ( .A1(n8593), .A2(n15092), .ZN(n15102) );
  AND2_X1 U15096 ( .A1(n15090), .A2(n15103), .ZN(n15101) );
  OR2_X1 U15097 ( .A1(n15092), .A2(n8593), .ZN(n15103) );
  OR2_X1 U15098 ( .A1(n8746), .A2(n8747), .ZN(n8593) );
  OR2_X1 U15099 ( .A1(n15104), .A2(n15105), .ZN(n15092) );
  AND2_X1 U15100 ( .A1(n15089), .A2(n15088), .ZN(n15105) );
  AND2_X1 U15101 ( .A1(n15086), .A2(n15106), .ZN(n15104) );
  OR2_X1 U15102 ( .A1(n15088), .A2(n15089), .ZN(n15106) );
  OR2_X1 U15103 ( .A1(n8750), .A2(n8747), .ZN(n15089) );
  OR2_X1 U15104 ( .A1(n15107), .A2(n15108), .ZN(n15088) );
  AND2_X1 U15105 ( .A1(n15085), .A2(n15084), .ZN(n15108) );
  AND2_X1 U15106 ( .A1(n15082), .A2(n15109), .ZN(n15107) );
  OR2_X1 U15107 ( .A1(n15084), .A2(n15085), .ZN(n15109) );
  OR2_X1 U15108 ( .A1(n8754), .A2(n8747), .ZN(n15085) );
  OR2_X1 U15109 ( .A1(n15110), .A2(n15111), .ZN(n15084) );
  AND2_X1 U15110 ( .A1(n15081), .A2(n15080), .ZN(n15111) );
  AND2_X1 U15111 ( .A1(n15078), .A2(n15112), .ZN(n15110) );
  OR2_X1 U15112 ( .A1(n15080), .A2(n15081), .ZN(n15112) );
  OR2_X1 U15113 ( .A1(n8758), .A2(n8747), .ZN(n15081) );
  OR2_X1 U15114 ( .A1(n15113), .A2(n15114), .ZN(n15080) );
  AND2_X1 U15115 ( .A1(n15077), .A2(n15076), .ZN(n15114) );
  AND2_X1 U15116 ( .A1(n15074), .A2(n15115), .ZN(n15113) );
  OR2_X1 U15117 ( .A1(n15076), .A2(n15077), .ZN(n15115) );
  OR2_X1 U15118 ( .A1(n8762), .A2(n8747), .ZN(n15077) );
  OR2_X1 U15119 ( .A1(n15116), .A2(n15117), .ZN(n15076) );
  AND2_X1 U15120 ( .A1(n15073), .A2(n15072), .ZN(n15117) );
  AND2_X1 U15121 ( .A1(n15070), .A2(n15118), .ZN(n15116) );
  OR2_X1 U15122 ( .A1(n15072), .A2(n15073), .ZN(n15118) );
  OR2_X1 U15123 ( .A1(n8766), .A2(n8747), .ZN(n15073) );
  OR2_X1 U15124 ( .A1(n15119), .A2(n15120), .ZN(n15072) );
  AND2_X1 U15125 ( .A1(n15069), .A2(n15068), .ZN(n15120) );
  AND2_X1 U15126 ( .A1(n15066), .A2(n15121), .ZN(n15119) );
  OR2_X1 U15127 ( .A1(n15068), .A2(n15069), .ZN(n15121) );
  OR2_X1 U15128 ( .A1(n8770), .A2(n8747), .ZN(n15069) );
  OR2_X1 U15129 ( .A1(n15122), .A2(n15123), .ZN(n15068) );
  AND2_X1 U15130 ( .A1(n15065), .A2(n15064), .ZN(n15123) );
  AND2_X1 U15131 ( .A1(n15062), .A2(n15124), .ZN(n15122) );
  OR2_X1 U15132 ( .A1(n15064), .A2(n15065), .ZN(n15124) );
  OR2_X1 U15133 ( .A1(n8774), .A2(n8747), .ZN(n15065) );
  OR2_X1 U15134 ( .A1(n15125), .A2(n15126), .ZN(n15064) );
  AND2_X1 U15135 ( .A1(n15061), .A2(n15060), .ZN(n15126) );
  AND2_X1 U15136 ( .A1(n15058), .A2(n15127), .ZN(n15125) );
  OR2_X1 U15137 ( .A1(n15060), .A2(n15061), .ZN(n15127) );
  OR2_X1 U15138 ( .A1(n8778), .A2(n8747), .ZN(n15061) );
  OR2_X1 U15139 ( .A1(n15128), .A2(n15129), .ZN(n15060) );
  AND2_X1 U15140 ( .A1(n15057), .A2(n15056), .ZN(n15129) );
  AND2_X1 U15141 ( .A1(n15054), .A2(n15130), .ZN(n15128) );
  OR2_X1 U15142 ( .A1(n15056), .A2(n15057), .ZN(n15130) );
  OR2_X1 U15143 ( .A1(n8782), .A2(n8747), .ZN(n15057) );
  OR2_X1 U15144 ( .A1(n15131), .A2(n15132), .ZN(n15056) );
  AND2_X1 U15145 ( .A1(n15053), .A2(n15052), .ZN(n15132) );
  AND2_X1 U15146 ( .A1(n15050), .A2(n15133), .ZN(n15131) );
  OR2_X1 U15147 ( .A1(n15052), .A2(n15053), .ZN(n15133) );
  OR2_X1 U15148 ( .A1(n8786), .A2(n8747), .ZN(n15053) );
  OR2_X1 U15149 ( .A1(n15134), .A2(n15135), .ZN(n15052) );
  AND2_X1 U15150 ( .A1(n15049), .A2(n15048), .ZN(n15135) );
  AND2_X1 U15151 ( .A1(n15046), .A2(n15136), .ZN(n15134) );
  OR2_X1 U15152 ( .A1(n15048), .A2(n15049), .ZN(n15136) );
  OR2_X1 U15153 ( .A1(n8790), .A2(n8747), .ZN(n15049) );
  OR2_X1 U15154 ( .A1(n15137), .A2(n15138), .ZN(n15048) );
  AND2_X1 U15155 ( .A1(n15045), .A2(n15044), .ZN(n15138) );
  AND2_X1 U15156 ( .A1(n15042), .A2(n15139), .ZN(n15137) );
  OR2_X1 U15157 ( .A1(n15044), .A2(n15045), .ZN(n15139) );
  OR2_X1 U15158 ( .A1(n8794), .A2(n8747), .ZN(n15045) );
  OR2_X1 U15159 ( .A1(n15140), .A2(n15141), .ZN(n15044) );
  AND2_X1 U15160 ( .A1(n15041), .A2(n15040), .ZN(n15141) );
  AND2_X1 U15161 ( .A1(n15038), .A2(n15142), .ZN(n15140) );
  OR2_X1 U15162 ( .A1(n15040), .A2(n15041), .ZN(n15142) );
  OR2_X1 U15163 ( .A1(n8798), .A2(n8747), .ZN(n15041) );
  OR2_X1 U15164 ( .A1(n15143), .A2(n15144), .ZN(n15040) );
  AND2_X1 U15165 ( .A1(n15037), .A2(n15036), .ZN(n15144) );
  AND2_X1 U15166 ( .A1(n15034), .A2(n15145), .ZN(n15143) );
  OR2_X1 U15167 ( .A1(n15036), .A2(n15037), .ZN(n15145) );
  OR2_X1 U15168 ( .A1(n8802), .A2(n8747), .ZN(n15037) );
  OR2_X1 U15169 ( .A1(n15146), .A2(n15147), .ZN(n15036) );
  AND2_X1 U15170 ( .A1(n15033), .A2(n15032), .ZN(n15147) );
  AND2_X1 U15171 ( .A1(n15030), .A2(n15148), .ZN(n15146) );
  OR2_X1 U15172 ( .A1(n15032), .A2(n15033), .ZN(n15148) );
  OR2_X1 U15173 ( .A1(n8806), .A2(n8747), .ZN(n15033) );
  OR2_X1 U15174 ( .A1(n15149), .A2(n15150), .ZN(n15032) );
  AND2_X1 U15175 ( .A1(n15029), .A2(n15028), .ZN(n15150) );
  AND2_X1 U15176 ( .A1(n15026), .A2(n15151), .ZN(n15149) );
  OR2_X1 U15177 ( .A1(n15028), .A2(n15029), .ZN(n15151) );
  OR2_X1 U15178 ( .A1(n8810), .A2(n8747), .ZN(n15029) );
  OR2_X1 U15179 ( .A1(n15152), .A2(n15153), .ZN(n15028) );
  AND2_X1 U15180 ( .A1(n15025), .A2(n15024), .ZN(n15153) );
  AND2_X1 U15181 ( .A1(n15022), .A2(n15154), .ZN(n15152) );
  OR2_X1 U15182 ( .A1(n15024), .A2(n15025), .ZN(n15154) );
  OR2_X1 U15183 ( .A1(n8140), .A2(n8747), .ZN(n15025) );
  OR2_X1 U15184 ( .A1(n15155), .A2(n15156), .ZN(n15024) );
  AND2_X1 U15185 ( .A1(n15021), .A2(n15020), .ZN(n15156) );
  AND2_X1 U15186 ( .A1(n15018), .A2(n15157), .ZN(n15155) );
  OR2_X1 U15187 ( .A1(n15020), .A2(n15021), .ZN(n15157) );
  OR2_X1 U15188 ( .A1(n8115), .A2(n8747), .ZN(n15021) );
  OR2_X1 U15189 ( .A1(n15158), .A2(n15159), .ZN(n15020) );
  AND2_X1 U15190 ( .A1(n15014), .A2(n15017), .ZN(n15159) );
  AND2_X1 U15191 ( .A1(n15160), .A2(n15016), .ZN(n15158) );
  OR2_X1 U15192 ( .A1(n15161), .A2(n15162), .ZN(n15016) );
  AND2_X1 U15193 ( .A1(n15013), .A2(n15012), .ZN(n15162) );
  AND2_X1 U15194 ( .A1(n15010), .A2(n15163), .ZN(n15161) );
  OR2_X1 U15195 ( .A1(n15012), .A2(n15013), .ZN(n15163) );
  OR2_X1 U15196 ( .A1(n8065), .A2(n8747), .ZN(n15013) );
  OR2_X1 U15197 ( .A1(n15164), .A2(n15165), .ZN(n15012) );
  AND2_X1 U15198 ( .A1(n15006), .A2(n15009), .ZN(n15165) );
  AND2_X1 U15199 ( .A1(n15166), .A2(n15008), .ZN(n15164) );
  OR2_X1 U15200 ( .A1(n15167), .A2(n15168), .ZN(n15008) );
  AND2_X1 U15201 ( .A1(n15002), .A2(n15005), .ZN(n15168) );
  AND2_X1 U15202 ( .A1(n15169), .A2(n15004), .ZN(n15167) );
  OR2_X1 U15203 ( .A1(n15170), .A2(n15171), .ZN(n15004) );
  AND2_X1 U15204 ( .A1(n14998), .A2(n15001), .ZN(n15171) );
  AND2_X1 U15205 ( .A1(n15172), .A2(n15000), .ZN(n15170) );
  OR2_X1 U15206 ( .A1(n15173), .A2(n15174), .ZN(n15000) );
  AND2_X1 U15207 ( .A1(n14994), .A2(n14997), .ZN(n15174) );
  AND2_X1 U15208 ( .A1(n15175), .A2(n15176), .ZN(n15173) );
  OR2_X1 U15209 ( .A1(n14997), .A2(n14994), .ZN(n15176) );
  OR2_X1 U15210 ( .A1(n7954), .A2(n8747), .ZN(n14994) );
  OR3_X1 U15211 ( .A1(n8747), .A2(n8743), .A3(n9796), .ZN(n14997) );
  INV_X1 U15212 ( .A(n14996), .ZN(n15175) );
  OR2_X1 U15213 ( .A1(n15177), .A2(n15178), .ZN(n14996) );
  AND2_X1 U15214 ( .A1(b_4_), .A2(n15179), .ZN(n15178) );
  OR2_X1 U15215 ( .A1(n15180), .A2(n9801), .ZN(n15179) );
  AND2_X1 U15216 ( .A1(a_30_), .A2(n8739), .ZN(n15180) );
  AND2_X1 U15217 ( .A1(b_3_), .A2(n15181), .ZN(n15177) );
  OR2_X1 U15218 ( .A1(n15182), .A2(n7920), .ZN(n15181) );
  AND2_X1 U15219 ( .A1(a_31_), .A2(n8743), .ZN(n15182) );
  OR2_X1 U15220 ( .A1(n15001), .A2(n14998), .ZN(n15172) );
  XNOR2_X1 U15221 ( .A(n15183), .B(n15184), .ZN(n14998) );
  XOR2_X1 U15222 ( .A(n15185), .B(n15186), .Z(n15184) );
  OR2_X1 U15223 ( .A1(n7979), .A2(n8747), .ZN(n15001) );
  OR2_X1 U15224 ( .A1(n15005), .A2(n15002), .ZN(n15169) );
  XOR2_X1 U15225 ( .A(n15187), .B(n15188), .Z(n15002) );
  XOR2_X1 U15226 ( .A(n15189), .B(n15190), .Z(n15188) );
  OR2_X1 U15227 ( .A1(n8015), .A2(n8747), .ZN(n15005) );
  OR2_X1 U15228 ( .A1(n15009), .A2(n15006), .ZN(n15166) );
  XOR2_X1 U15229 ( .A(n15191), .B(n15192), .Z(n15006) );
  XOR2_X1 U15230 ( .A(n15193), .B(n15194), .Z(n15192) );
  OR2_X1 U15231 ( .A1(n8040), .A2(n8747), .ZN(n15009) );
  XOR2_X1 U15232 ( .A(n15195), .B(n15196), .Z(n15010) );
  XOR2_X1 U15233 ( .A(n15197), .B(n15198), .Z(n15196) );
  OR2_X1 U15234 ( .A1(n15017), .A2(n15014), .ZN(n15160) );
  XOR2_X1 U15235 ( .A(n15199), .B(n15200), .Z(n15014) );
  XOR2_X1 U15236 ( .A(n15201), .B(n15202), .Z(n15200) );
  OR2_X1 U15237 ( .A1(n8090), .A2(n8747), .ZN(n15017) );
  XOR2_X1 U15238 ( .A(n15203), .B(n15204), .Z(n15018) );
  XOR2_X1 U15239 ( .A(n15205), .B(n15206), .Z(n15204) );
  XOR2_X1 U15240 ( .A(n15207), .B(n15208), .Z(n15022) );
  XOR2_X1 U15241 ( .A(n15209), .B(n15210), .Z(n15208) );
  XOR2_X1 U15242 ( .A(n15211), .B(n15212), .Z(n15026) );
  XOR2_X1 U15243 ( .A(n15213), .B(n15214), .Z(n15212) );
  XOR2_X1 U15244 ( .A(n15215), .B(n15216), .Z(n15030) );
  XOR2_X1 U15245 ( .A(n15217), .B(n15218), .Z(n15216) );
  XOR2_X1 U15246 ( .A(n15219), .B(n15220), .Z(n15034) );
  XOR2_X1 U15247 ( .A(n15221), .B(n15222), .Z(n15220) );
  XOR2_X1 U15248 ( .A(n15223), .B(n15224), .Z(n15038) );
  XOR2_X1 U15249 ( .A(n15225), .B(n15226), .Z(n15224) );
  XOR2_X1 U15250 ( .A(n15227), .B(n15228), .Z(n15042) );
  XOR2_X1 U15251 ( .A(n15229), .B(n15230), .Z(n15228) );
  XOR2_X1 U15252 ( .A(n15231), .B(n15232), .Z(n15046) );
  XOR2_X1 U15253 ( .A(n15233), .B(n15234), .Z(n15232) );
  XOR2_X1 U15254 ( .A(n15235), .B(n15236), .Z(n15050) );
  XOR2_X1 U15255 ( .A(n15237), .B(n15238), .Z(n15236) );
  XOR2_X1 U15256 ( .A(n15239), .B(n15240), .Z(n15054) );
  XOR2_X1 U15257 ( .A(n15241), .B(n15242), .Z(n15240) );
  XOR2_X1 U15258 ( .A(n15243), .B(n15244), .Z(n15058) );
  XOR2_X1 U15259 ( .A(n15245), .B(n15246), .Z(n15244) );
  XOR2_X1 U15260 ( .A(n15247), .B(n15248), .Z(n15062) );
  XOR2_X1 U15261 ( .A(n15249), .B(n15250), .Z(n15248) );
  XOR2_X1 U15262 ( .A(n15251), .B(n15252), .Z(n15066) );
  XOR2_X1 U15263 ( .A(n15253), .B(n15254), .Z(n15252) );
  XOR2_X1 U15264 ( .A(n15255), .B(n15256), .Z(n15070) );
  XOR2_X1 U15265 ( .A(n15257), .B(n15258), .Z(n15256) );
  XOR2_X1 U15266 ( .A(n15259), .B(n15260), .Z(n15074) );
  XOR2_X1 U15267 ( .A(n15261), .B(n15262), .Z(n15260) );
  XOR2_X1 U15268 ( .A(n15263), .B(n15264), .Z(n15078) );
  XOR2_X1 U15269 ( .A(n15265), .B(n15266), .Z(n15264) );
  XOR2_X1 U15270 ( .A(n15267), .B(n15268), .Z(n15082) );
  XOR2_X1 U15271 ( .A(n15269), .B(n15270), .Z(n15268) );
  XOR2_X1 U15272 ( .A(n15271), .B(n15272), .Z(n15086) );
  XOR2_X1 U15273 ( .A(n15273), .B(n15274), .Z(n15272) );
  XOR2_X1 U15274 ( .A(n15275), .B(n15276), .Z(n15090) );
  XOR2_X1 U15275 ( .A(n15277), .B(n15278), .Z(n15276) );
  XOR2_X1 U15276 ( .A(n15279), .B(n15280), .Z(n15093) );
  XOR2_X1 U15277 ( .A(n15281), .B(n15282), .Z(n15280) );
  XOR2_X1 U15278 ( .A(n9399), .B(n15283), .Z(n9393) );
  XOR2_X1 U15279 ( .A(n9398), .B(n8619), .Z(n15283) );
  OR2_X1 U15280 ( .A1(n8742), .A2(n8743), .ZN(n8619) );
  OR2_X1 U15281 ( .A1(n15284), .A2(n15285), .ZN(n9398) );
  AND2_X1 U15282 ( .A1(n15282), .A2(n15281), .ZN(n15285) );
  AND2_X1 U15283 ( .A1(n15279), .A2(n15286), .ZN(n15284) );
  OR2_X1 U15284 ( .A1(n15281), .A2(n15282), .ZN(n15286) );
  OR2_X1 U15285 ( .A1(n8746), .A2(n8743), .ZN(n15282) );
  OR2_X1 U15286 ( .A1(n15287), .A2(n15288), .ZN(n15281) );
  AND2_X1 U15287 ( .A1(n15278), .A2(n15277), .ZN(n15288) );
  AND2_X1 U15288 ( .A1(n15275), .A2(n15289), .ZN(n15287) );
  OR2_X1 U15289 ( .A1(n15277), .A2(n15278), .ZN(n15289) );
  OR2_X1 U15290 ( .A1(n8750), .A2(n8743), .ZN(n15278) );
  OR2_X1 U15291 ( .A1(n15290), .A2(n15291), .ZN(n15277) );
  AND2_X1 U15292 ( .A1(n15274), .A2(n15273), .ZN(n15291) );
  AND2_X1 U15293 ( .A1(n15271), .A2(n15292), .ZN(n15290) );
  OR2_X1 U15294 ( .A1(n15273), .A2(n15274), .ZN(n15292) );
  OR2_X1 U15295 ( .A1(n8754), .A2(n8743), .ZN(n15274) );
  OR2_X1 U15296 ( .A1(n15293), .A2(n15294), .ZN(n15273) );
  AND2_X1 U15297 ( .A1(n15270), .A2(n15269), .ZN(n15294) );
  AND2_X1 U15298 ( .A1(n15267), .A2(n15295), .ZN(n15293) );
  OR2_X1 U15299 ( .A1(n15269), .A2(n15270), .ZN(n15295) );
  OR2_X1 U15300 ( .A1(n8758), .A2(n8743), .ZN(n15270) );
  OR2_X1 U15301 ( .A1(n15296), .A2(n15297), .ZN(n15269) );
  AND2_X1 U15302 ( .A1(n15266), .A2(n15265), .ZN(n15297) );
  AND2_X1 U15303 ( .A1(n15263), .A2(n15298), .ZN(n15296) );
  OR2_X1 U15304 ( .A1(n15265), .A2(n15266), .ZN(n15298) );
  OR2_X1 U15305 ( .A1(n8762), .A2(n8743), .ZN(n15266) );
  OR2_X1 U15306 ( .A1(n15299), .A2(n15300), .ZN(n15265) );
  AND2_X1 U15307 ( .A1(n15262), .A2(n15261), .ZN(n15300) );
  AND2_X1 U15308 ( .A1(n15259), .A2(n15301), .ZN(n15299) );
  OR2_X1 U15309 ( .A1(n15261), .A2(n15262), .ZN(n15301) );
  OR2_X1 U15310 ( .A1(n8766), .A2(n8743), .ZN(n15262) );
  OR2_X1 U15311 ( .A1(n15302), .A2(n15303), .ZN(n15261) );
  AND2_X1 U15312 ( .A1(n15258), .A2(n15257), .ZN(n15303) );
  AND2_X1 U15313 ( .A1(n15255), .A2(n15304), .ZN(n15302) );
  OR2_X1 U15314 ( .A1(n15257), .A2(n15258), .ZN(n15304) );
  OR2_X1 U15315 ( .A1(n8770), .A2(n8743), .ZN(n15258) );
  OR2_X1 U15316 ( .A1(n15305), .A2(n15306), .ZN(n15257) );
  AND2_X1 U15317 ( .A1(n15254), .A2(n15253), .ZN(n15306) );
  AND2_X1 U15318 ( .A1(n15251), .A2(n15307), .ZN(n15305) );
  OR2_X1 U15319 ( .A1(n15253), .A2(n15254), .ZN(n15307) );
  OR2_X1 U15320 ( .A1(n8774), .A2(n8743), .ZN(n15254) );
  OR2_X1 U15321 ( .A1(n15308), .A2(n15309), .ZN(n15253) );
  AND2_X1 U15322 ( .A1(n15250), .A2(n15249), .ZN(n15309) );
  AND2_X1 U15323 ( .A1(n15247), .A2(n15310), .ZN(n15308) );
  OR2_X1 U15324 ( .A1(n15249), .A2(n15250), .ZN(n15310) );
  OR2_X1 U15325 ( .A1(n8778), .A2(n8743), .ZN(n15250) );
  OR2_X1 U15326 ( .A1(n15311), .A2(n15312), .ZN(n15249) );
  AND2_X1 U15327 ( .A1(n15246), .A2(n15245), .ZN(n15312) );
  AND2_X1 U15328 ( .A1(n15243), .A2(n15313), .ZN(n15311) );
  OR2_X1 U15329 ( .A1(n15245), .A2(n15246), .ZN(n15313) );
  OR2_X1 U15330 ( .A1(n8782), .A2(n8743), .ZN(n15246) );
  OR2_X1 U15331 ( .A1(n15314), .A2(n15315), .ZN(n15245) );
  AND2_X1 U15332 ( .A1(n15242), .A2(n15241), .ZN(n15315) );
  AND2_X1 U15333 ( .A1(n15239), .A2(n15316), .ZN(n15314) );
  OR2_X1 U15334 ( .A1(n15241), .A2(n15242), .ZN(n15316) );
  OR2_X1 U15335 ( .A1(n8786), .A2(n8743), .ZN(n15242) );
  OR2_X1 U15336 ( .A1(n15317), .A2(n15318), .ZN(n15241) );
  AND2_X1 U15337 ( .A1(n15238), .A2(n15237), .ZN(n15318) );
  AND2_X1 U15338 ( .A1(n15235), .A2(n15319), .ZN(n15317) );
  OR2_X1 U15339 ( .A1(n15237), .A2(n15238), .ZN(n15319) );
  OR2_X1 U15340 ( .A1(n8790), .A2(n8743), .ZN(n15238) );
  OR2_X1 U15341 ( .A1(n15320), .A2(n15321), .ZN(n15237) );
  AND2_X1 U15342 ( .A1(n15234), .A2(n15233), .ZN(n15321) );
  AND2_X1 U15343 ( .A1(n15231), .A2(n15322), .ZN(n15320) );
  OR2_X1 U15344 ( .A1(n15233), .A2(n15234), .ZN(n15322) );
  OR2_X1 U15345 ( .A1(n8794), .A2(n8743), .ZN(n15234) );
  OR2_X1 U15346 ( .A1(n15323), .A2(n15324), .ZN(n15233) );
  AND2_X1 U15347 ( .A1(n15230), .A2(n15229), .ZN(n15324) );
  AND2_X1 U15348 ( .A1(n15227), .A2(n15325), .ZN(n15323) );
  OR2_X1 U15349 ( .A1(n15229), .A2(n15230), .ZN(n15325) );
  OR2_X1 U15350 ( .A1(n8798), .A2(n8743), .ZN(n15230) );
  OR2_X1 U15351 ( .A1(n15326), .A2(n15327), .ZN(n15229) );
  AND2_X1 U15352 ( .A1(n15226), .A2(n15225), .ZN(n15327) );
  AND2_X1 U15353 ( .A1(n15223), .A2(n15328), .ZN(n15326) );
  OR2_X1 U15354 ( .A1(n15225), .A2(n15226), .ZN(n15328) );
  OR2_X1 U15355 ( .A1(n8802), .A2(n8743), .ZN(n15226) );
  OR2_X1 U15356 ( .A1(n15329), .A2(n15330), .ZN(n15225) );
  AND2_X1 U15357 ( .A1(n15222), .A2(n15221), .ZN(n15330) );
  AND2_X1 U15358 ( .A1(n15219), .A2(n15331), .ZN(n15329) );
  OR2_X1 U15359 ( .A1(n15221), .A2(n15222), .ZN(n15331) );
  OR2_X1 U15360 ( .A1(n8806), .A2(n8743), .ZN(n15222) );
  OR2_X1 U15361 ( .A1(n15332), .A2(n15333), .ZN(n15221) );
  AND2_X1 U15362 ( .A1(n15218), .A2(n15217), .ZN(n15333) );
  AND2_X1 U15363 ( .A1(n15215), .A2(n15334), .ZN(n15332) );
  OR2_X1 U15364 ( .A1(n15217), .A2(n15218), .ZN(n15334) );
  OR2_X1 U15365 ( .A1(n8810), .A2(n8743), .ZN(n15218) );
  OR2_X1 U15366 ( .A1(n15335), .A2(n15336), .ZN(n15217) );
  AND2_X1 U15367 ( .A1(n15214), .A2(n15213), .ZN(n15336) );
  AND2_X1 U15368 ( .A1(n15211), .A2(n15337), .ZN(n15335) );
  OR2_X1 U15369 ( .A1(n15213), .A2(n15214), .ZN(n15337) );
  OR2_X1 U15370 ( .A1(n8140), .A2(n8743), .ZN(n15214) );
  OR2_X1 U15371 ( .A1(n15338), .A2(n15339), .ZN(n15213) );
  AND2_X1 U15372 ( .A1(n15210), .A2(n15209), .ZN(n15339) );
  AND2_X1 U15373 ( .A1(n15207), .A2(n15340), .ZN(n15338) );
  OR2_X1 U15374 ( .A1(n15209), .A2(n15210), .ZN(n15340) );
  OR2_X1 U15375 ( .A1(n8115), .A2(n8743), .ZN(n15210) );
  OR2_X1 U15376 ( .A1(n15341), .A2(n15342), .ZN(n15209) );
  AND2_X1 U15377 ( .A1(n15206), .A2(n15205), .ZN(n15342) );
  AND2_X1 U15378 ( .A1(n15203), .A2(n15343), .ZN(n15341) );
  OR2_X1 U15379 ( .A1(n15205), .A2(n15206), .ZN(n15343) );
  OR2_X1 U15380 ( .A1(n8090), .A2(n8743), .ZN(n15206) );
  OR2_X1 U15381 ( .A1(n15344), .A2(n15345), .ZN(n15205) );
  AND2_X1 U15382 ( .A1(n15199), .A2(n15202), .ZN(n15345) );
  AND2_X1 U15383 ( .A1(n15346), .A2(n15201), .ZN(n15344) );
  OR2_X1 U15384 ( .A1(n15347), .A2(n15348), .ZN(n15201) );
  AND2_X1 U15385 ( .A1(n15198), .A2(n15197), .ZN(n15348) );
  AND2_X1 U15386 ( .A1(n15195), .A2(n15349), .ZN(n15347) );
  OR2_X1 U15387 ( .A1(n15197), .A2(n15198), .ZN(n15349) );
  OR2_X1 U15388 ( .A1(n8040), .A2(n8743), .ZN(n15198) );
  OR2_X1 U15389 ( .A1(n15350), .A2(n15351), .ZN(n15197) );
  AND2_X1 U15390 ( .A1(n15191), .A2(n15194), .ZN(n15351) );
  AND2_X1 U15391 ( .A1(n15352), .A2(n15193), .ZN(n15350) );
  OR2_X1 U15392 ( .A1(n15353), .A2(n15354), .ZN(n15193) );
  AND2_X1 U15393 ( .A1(n15187), .A2(n15190), .ZN(n15354) );
  AND2_X1 U15394 ( .A1(n15355), .A2(n15189), .ZN(n15353) );
  OR2_X1 U15395 ( .A1(n15356), .A2(n15357), .ZN(n15189) );
  AND2_X1 U15396 ( .A1(n15183), .A2(n15186), .ZN(n15357) );
  AND2_X1 U15397 ( .A1(n15358), .A2(n15359), .ZN(n15356) );
  OR2_X1 U15398 ( .A1(n15186), .A2(n15183), .ZN(n15359) );
  OR2_X1 U15399 ( .A1(n7954), .A2(n8743), .ZN(n15183) );
  OR3_X1 U15400 ( .A1(n8743), .A2(n8739), .A3(n9796), .ZN(n15186) );
  INV_X1 U15401 ( .A(n15185), .ZN(n15358) );
  OR2_X1 U15402 ( .A1(n15360), .A2(n15361), .ZN(n15185) );
  AND2_X1 U15403 ( .A1(b_3_), .A2(n15362), .ZN(n15361) );
  OR2_X1 U15404 ( .A1(n15363), .A2(n9801), .ZN(n15362) );
  AND2_X1 U15405 ( .A1(a_30_), .A2(n8735), .ZN(n15363) );
  AND2_X1 U15406 ( .A1(b_2_), .A2(n15364), .ZN(n15360) );
  OR2_X1 U15407 ( .A1(n15365), .A2(n7920), .ZN(n15364) );
  AND2_X1 U15408 ( .A1(a_31_), .A2(n8739), .ZN(n15365) );
  OR2_X1 U15409 ( .A1(n15190), .A2(n15187), .ZN(n15355) );
  XNOR2_X1 U15410 ( .A(n15366), .B(n15367), .ZN(n15187) );
  XOR2_X1 U15411 ( .A(n15368), .B(n15369), .Z(n15367) );
  OR2_X1 U15412 ( .A1(n7979), .A2(n8743), .ZN(n15190) );
  OR2_X1 U15413 ( .A1(n15194), .A2(n15191), .ZN(n15352) );
  XOR2_X1 U15414 ( .A(n15370), .B(n15371), .Z(n15191) );
  XOR2_X1 U15415 ( .A(n15372), .B(n15373), .Z(n15371) );
  OR2_X1 U15416 ( .A1(n8015), .A2(n8743), .ZN(n15194) );
  XOR2_X1 U15417 ( .A(n15374), .B(n15375), .Z(n15195) );
  XOR2_X1 U15418 ( .A(n15376), .B(n15377), .Z(n15375) );
  OR2_X1 U15419 ( .A1(n15202), .A2(n15199), .ZN(n15346) );
  XOR2_X1 U15420 ( .A(n15378), .B(n15379), .Z(n15199) );
  XOR2_X1 U15421 ( .A(n15380), .B(n15381), .Z(n15379) );
  OR2_X1 U15422 ( .A1(n8065), .A2(n8743), .ZN(n15202) );
  XOR2_X1 U15423 ( .A(n15382), .B(n15383), .Z(n15203) );
  XOR2_X1 U15424 ( .A(n15384), .B(n15385), .Z(n15383) );
  XOR2_X1 U15425 ( .A(n15386), .B(n15387), .Z(n15207) );
  XOR2_X1 U15426 ( .A(n15388), .B(n15389), .Z(n15387) );
  XOR2_X1 U15427 ( .A(n15390), .B(n15391), .Z(n15211) );
  XOR2_X1 U15428 ( .A(n15392), .B(n15393), .Z(n15391) );
  XOR2_X1 U15429 ( .A(n15394), .B(n15395), .Z(n15215) );
  XOR2_X1 U15430 ( .A(n15396), .B(n15397), .Z(n15395) );
  XOR2_X1 U15431 ( .A(n15398), .B(n15399), .Z(n15219) );
  XOR2_X1 U15432 ( .A(n15400), .B(n15401), .Z(n15399) );
  XOR2_X1 U15433 ( .A(n15402), .B(n15403), .Z(n15223) );
  XOR2_X1 U15434 ( .A(n15404), .B(n15405), .Z(n15403) );
  XOR2_X1 U15435 ( .A(n15406), .B(n15407), .Z(n15227) );
  XOR2_X1 U15436 ( .A(n15408), .B(n15409), .Z(n15407) );
  XOR2_X1 U15437 ( .A(n15410), .B(n15411), .Z(n15231) );
  XOR2_X1 U15438 ( .A(n15412), .B(n15413), .Z(n15411) );
  XOR2_X1 U15439 ( .A(n15414), .B(n15415), .Z(n15235) );
  XOR2_X1 U15440 ( .A(n15416), .B(n15417), .Z(n15415) );
  XOR2_X1 U15441 ( .A(n15418), .B(n15419), .Z(n15239) );
  XOR2_X1 U15442 ( .A(n15420), .B(n15421), .Z(n15419) );
  XOR2_X1 U15443 ( .A(n15422), .B(n15423), .Z(n15243) );
  XOR2_X1 U15444 ( .A(n15424), .B(n15425), .Z(n15423) );
  XOR2_X1 U15445 ( .A(n15426), .B(n15427), .Z(n15247) );
  XOR2_X1 U15446 ( .A(n15428), .B(n15429), .Z(n15427) );
  XOR2_X1 U15447 ( .A(n15430), .B(n15431), .Z(n15251) );
  XOR2_X1 U15448 ( .A(n15432), .B(n15433), .Z(n15431) );
  XOR2_X1 U15449 ( .A(n15434), .B(n15435), .Z(n15255) );
  XOR2_X1 U15450 ( .A(n15436), .B(n15437), .Z(n15435) );
  XOR2_X1 U15451 ( .A(n15438), .B(n15439), .Z(n15259) );
  XOR2_X1 U15452 ( .A(n15440), .B(n15441), .Z(n15439) );
  XOR2_X1 U15453 ( .A(n15442), .B(n15443), .Z(n15263) );
  XOR2_X1 U15454 ( .A(n15444), .B(n15445), .Z(n15443) );
  XOR2_X1 U15455 ( .A(n15446), .B(n15447), .Z(n15267) );
  XOR2_X1 U15456 ( .A(n15448), .B(n15449), .Z(n15447) );
  XOR2_X1 U15457 ( .A(n15450), .B(n15451), .Z(n15271) );
  XOR2_X1 U15458 ( .A(n15452), .B(n15453), .Z(n15451) );
  XOR2_X1 U15459 ( .A(n15454), .B(n15455), .Z(n15275) );
  XOR2_X1 U15460 ( .A(n15456), .B(n15457), .Z(n15455) );
  XOR2_X1 U15461 ( .A(n15458), .B(n15459), .Z(n15279) );
  XOR2_X1 U15462 ( .A(n15460), .B(n15461), .Z(n15459) );
  XOR2_X1 U15463 ( .A(n9406), .B(n15462), .Z(n9399) );
  XOR2_X1 U15464 ( .A(n9405), .B(n9404), .Z(n15462) );
  OR2_X1 U15465 ( .A1(n8746), .A2(n8739), .ZN(n9404) );
  OR2_X1 U15466 ( .A1(n15463), .A2(n15464), .ZN(n9405) );
  AND2_X1 U15467 ( .A1(n15461), .A2(n15460), .ZN(n15464) );
  AND2_X1 U15468 ( .A1(n15458), .A2(n15465), .ZN(n15463) );
  OR2_X1 U15469 ( .A1(n15460), .A2(n15461), .ZN(n15465) );
  OR2_X1 U15470 ( .A1(n8750), .A2(n8739), .ZN(n15461) );
  OR2_X1 U15471 ( .A1(n15466), .A2(n15467), .ZN(n15460) );
  AND2_X1 U15472 ( .A1(n15457), .A2(n15456), .ZN(n15467) );
  AND2_X1 U15473 ( .A1(n15454), .A2(n15468), .ZN(n15466) );
  OR2_X1 U15474 ( .A1(n15456), .A2(n15457), .ZN(n15468) );
  OR2_X1 U15475 ( .A1(n8754), .A2(n8739), .ZN(n15457) );
  OR2_X1 U15476 ( .A1(n15469), .A2(n15470), .ZN(n15456) );
  AND2_X1 U15477 ( .A1(n15453), .A2(n15452), .ZN(n15470) );
  AND2_X1 U15478 ( .A1(n15450), .A2(n15471), .ZN(n15469) );
  OR2_X1 U15479 ( .A1(n15452), .A2(n15453), .ZN(n15471) );
  OR2_X1 U15480 ( .A1(n8758), .A2(n8739), .ZN(n15453) );
  OR2_X1 U15481 ( .A1(n15472), .A2(n15473), .ZN(n15452) );
  AND2_X1 U15482 ( .A1(n15449), .A2(n15448), .ZN(n15473) );
  AND2_X1 U15483 ( .A1(n15446), .A2(n15474), .ZN(n15472) );
  OR2_X1 U15484 ( .A1(n15448), .A2(n15449), .ZN(n15474) );
  OR2_X1 U15485 ( .A1(n8762), .A2(n8739), .ZN(n15449) );
  OR2_X1 U15486 ( .A1(n15475), .A2(n15476), .ZN(n15448) );
  AND2_X1 U15487 ( .A1(n15445), .A2(n15444), .ZN(n15476) );
  AND2_X1 U15488 ( .A1(n15442), .A2(n15477), .ZN(n15475) );
  OR2_X1 U15489 ( .A1(n15444), .A2(n15445), .ZN(n15477) );
  OR2_X1 U15490 ( .A1(n8766), .A2(n8739), .ZN(n15445) );
  OR2_X1 U15491 ( .A1(n15478), .A2(n15479), .ZN(n15444) );
  AND2_X1 U15492 ( .A1(n15441), .A2(n15440), .ZN(n15479) );
  AND2_X1 U15493 ( .A1(n15438), .A2(n15480), .ZN(n15478) );
  OR2_X1 U15494 ( .A1(n15440), .A2(n15441), .ZN(n15480) );
  OR2_X1 U15495 ( .A1(n8770), .A2(n8739), .ZN(n15441) );
  OR2_X1 U15496 ( .A1(n15481), .A2(n15482), .ZN(n15440) );
  AND2_X1 U15497 ( .A1(n15437), .A2(n15436), .ZN(n15482) );
  AND2_X1 U15498 ( .A1(n15434), .A2(n15483), .ZN(n15481) );
  OR2_X1 U15499 ( .A1(n15436), .A2(n15437), .ZN(n15483) );
  OR2_X1 U15500 ( .A1(n8774), .A2(n8739), .ZN(n15437) );
  OR2_X1 U15501 ( .A1(n15484), .A2(n15485), .ZN(n15436) );
  AND2_X1 U15502 ( .A1(n15433), .A2(n15432), .ZN(n15485) );
  AND2_X1 U15503 ( .A1(n15430), .A2(n15486), .ZN(n15484) );
  OR2_X1 U15504 ( .A1(n15432), .A2(n15433), .ZN(n15486) );
  OR2_X1 U15505 ( .A1(n8778), .A2(n8739), .ZN(n15433) );
  OR2_X1 U15506 ( .A1(n15487), .A2(n15488), .ZN(n15432) );
  AND2_X1 U15507 ( .A1(n15429), .A2(n15428), .ZN(n15488) );
  AND2_X1 U15508 ( .A1(n15426), .A2(n15489), .ZN(n15487) );
  OR2_X1 U15509 ( .A1(n15428), .A2(n15429), .ZN(n15489) );
  OR2_X1 U15510 ( .A1(n8782), .A2(n8739), .ZN(n15429) );
  OR2_X1 U15511 ( .A1(n15490), .A2(n15491), .ZN(n15428) );
  AND2_X1 U15512 ( .A1(n15425), .A2(n15424), .ZN(n15491) );
  AND2_X1 U15513 ( .A1(n15422), .A2(n15492), .ZN(n15490) );
  OR2_X1 U15514 ( .A1(n15424), .A2(n15425), .ZN(n15492) );
  OR2_X1 U15515 ( .A1(n8786), .A2(n8739), .ZN(n15425) );
  OR2_X1 U15516 ( .A1(n15493), .A2(n15494), .ZN(n15424) );
  AND2_X1 U15517 ( .A1(n15421), .A2(n15420), .ZN(n15494) );
  AND2_X1 U15518 ( .A1(n15418), .A2(n15495), .ZN(n15493) );
  OR2_X1 U15519 ( .A1(n15420), .A2(n15421), .ZN(n15495) );
  OR2_X1 U15520 ( .A1(n8790), .A2(n8739), .ZN(n15421) );
  OR2_X1 U15521 ( .A1(n15496), .A2(n15497), .ZN(n15420) );
  AND2_X1 U15522 ( .A1(n15417), .A2(n15416), .ZN(n15497) );
  AND2_X1 U15523 ( .A1(n15414), .A2(n15498), .ZN(n15496) );
  OR2_X1 U15524 ( .A1(n15416), .A2(n15417), .ZN(n15498) );
  OR2_X1 U15525 ( .A1(n8794), .A2(n8739), .ZN(n15417) );
  OR2_X1 U15526 ( .A1(n15499), .A2(n15500), .ZN(n15416) );
  AND2_X1 U15527 ( .A1(n15413), .A2(n15412), .ZN(n15500) );
  AND2_X1 U15528 ( .A1(n15410), .A2(n15501), .ZN(n15499) );
  OR2_X1 U15529 ( .A1(n15412), .A2(n15413), .ZN(n15501) );
  OR2_X1 U15530 ( .A1(n8798), .A2(n8739), .ZN(n15413) );
  OR2_X1 U15531 ( .A1(n15502), .A2(n15503), .ZN(n15412) );
  AND2_X1 U15532 ( .A1(n15409), .A2(n15408), .ZN(n15503) );
  AND2_X1 U15533 ( .A1(n15406), .A2(n15504), .ZN(n15502) );
  OR2_X1 U15534 ( .A1(n15408), .A2(n15409), .ZN(n15504) );
  OR2_X1 U15535 ( .A1(n8802), .A2(n8739), .ZN(n15409) );
  OR2_X1 U15536 ( .A1(n15505), .A2(n15506), .ZN(n15408) );
  AND2_X1 U15537 ( .A1(n15405), .A2(n15404), .ZN(n15506) );
  AND2_X1 U15538 ( .A1(n15402), .A2(n15507), .ZN(n15505) );
  OR2_X1 U15539 ( .A1(n15404), .A2(n15405), .ZN(n15507) );
  OR2_X1 U15540 ( .A1(n8806), .A2(n8739), .ZN(n15405) );
  OR2_X1 U15541 ( .A1(n15508), .A2(n15509), .ZN(n15404) );
  AND2_X1 U15542 ( .A1(n15401), .A2(n15400), .ZN(n15509) );
  AND2_X1 U15543 ( .A1(n15398), .A2(n15510), .ZN(n15508) );
  OR2_X1 U15544 ( .A1(n15400), .A2(n15401), .ZN(n15510) );
  OR2_X1 U15545 ( .A1(n8810), .A2(n8739), .ZN(n15401) );
  OR2_X1 U15546 ( .A1(n15511), .A2(n15512), .ZN(n15400) );
  AND2_X1 U15547 ( .A1(n15397), .A2(n15396), .ZN(n15512) );
  AND2_X1 U15548 ( .A1(n15394), .A2(n15513), .ZN(n15511) );
  OR2_X1 U15549 ( .A1(n15396), .A2(n15397), .ZN(n15513) );
  OR2_X1 U15550 ( .A1(n8140), .A2(n8739), .ZN(n15397) );
  OR2_X1 U15551 ( .A1(n15514), .A2(n15515), .ZN(n15396) );
  AND2_X1 U15552 ( .A1(n15393), .A2(n15392), .ZN(n15515) );
  AND2_X1 U15553 ( .A1(n15390), .A2(n15516), .ZN(n15514) );
  OR2_X1 U15554 ( .A1(n15392), .A2(n15393), .ZN(n15516) );
  OR2_X1 U15555 ( .A1(n8115), .A2(n8739), .ZN(n15393) );
  OR2_X1 U15556 ( .A1(n15517), .A2(n15518), .ZN(n15392) );
  AND2_X1 U15557 ( .A1(n15389), .A2(n15388), .ZN(n15518) );
  AND2_X1 U15558 ( .A1(n15386), .A2(n15519), .ZN(n15517) );
  OR2_X1 U15559 ( .A1(n15388), .A2(n15389), .ZN(n15519) );
  OR2_X1 U15560 ( .A1(n8090), .A2(n8739), .ZN(n15389) );
  OR2_X1 U15561 ( .A1(n15520), .A2(n15521), .ZN(n15388) );
  AND2_X1 U15562 ( .A1(n15385), .A2(n15384), .ZN(n15521) );
  AND2_X1 U15563 ( .A1(n15382), .A2(n15522), .ZN(n15520) );
  OR2_X1 U15564 ( .A1(n15384), .A2(n15385), .ZN(n15522) );
  OR2_X1 U15565 ( .A1(n8065), .A2(n8739), .ZN(n15385) );
  OR2_X1 U15566 ( .A1(n15523), .A2(n15524), .ZN(n15384) );
  AND2_X1 U15567 ( .A1(n15378), .A2(n15381), .ZN(n15524) );
  AND2_X1 U15568 ( .A1(n15525), .A2(n15380), .ZN(n15523) );
  OR2_X1 U15569 ( .A1(n15526), .A2(n15527), .ZN(n15380) );
  AND2_X1 U15570 ( .A1(n15377), .A2(n15376), .ZN(n15527) );
  AND2_X1 U15571 ( .A1(n15374), .A2(n15528), .ZN(n15526) );
  OR2_X1 U15572 ( .A1(n15376), .A2(n15377), .ZN(n15528) );
  OR2_X1 U15573 ( .A1(n8015), .A2(n8739), .ZN(n15377) );
  OR2_X1 U15574 ( .A1(n15529), .A2(n15530), .ZN(n15376) );
  AND2_X1 U15575 ( .A1(n15370), .A2(n15373), .ZN(n15530) );
  AND2_X1 U15576 ( .A1(n15531), .A2(n15372), .ZN(n15529) );
  OR2_X1 U15577 ( .A1(n15532), .A2(n15533), .ZN(n15372) );
  AND2_X1 U15578 ( .A1(n15366), .A2(n15369), .ZN(n15533) );
  AND2_X1 U15579 ( .A1(n15534), .A2(n15535), .ZN(n15532) );
  OR2_X1 U15580 ( .A1(n15369), .A2(n15366), .ZN(n15535) );
  OR2_X1 U15581 ( .A1(n7954), .A2(n8739), .ZN(n15366) );
  OR3_X1 U15582 ( .A1(n8739), .A2(n8735), .A3(n9796), .ZN(n15369) );
  INV_X1 U15583 ( .A(n15368), .ZN(n15534) );
  OR2_X1 U15584 ( .A1(n15536), .A2(n15537), .ZN(n15368) );
  AND2_X1 U15585 ( .A1(b_2_), .A2(n15538), .ZN(n15537) );
  OR2_X1 U15586 ( .A1(n15539), .A2(n9801), .ZN(n15538) );
  AND2_X1 U15587 ( .A1(a_30_), .A2(n8731), .ZN(n15539) );
  AND2_X1 U15588 ( .A1(b_1_), .A2(n15540), .ZN(n15536) );
  OR2_X1 U15589 ( .A1(n15541), .A2(n7920), .ZN(n15540) );
  AND2_X1 U15590 ( .A1(a_31_), .A2(n8735), .ZN(n15541) );
  OR2_X1 U15591 ( .A1(n15373), .A2(n15370), .ZN(n15531) );
  XNOR2_X1 U15592 ( .A(n15542), .B(n15543), .ZN(n15370) );
  XOR2_X1 U15593 ( .A(n15544), .B(n15545), .Z(n15543) );
  OR2_X1 U15594 ( .A1(n7979), .A2(n8739), .ZN(n15373) );
  XOR2_X1 U15595 ( .A(n15546), .B(n15547), .Z(n15374) );
  XOR2_X1 U15596 ( .A(n15548), .B(n15549), .Z(n15547) );
  OR2_X1 U15597 ( .A1(n15381), .A2(n15378), .ZN(n15525) );
  XOR2_X1 U15598 ( .A(n15550), .B(n15551), .Z(n15378) );
  XOR2_X1 U15599 ( .A(n15552), .B(n15553), .Z(n15551) );
  OR2_X1 U15600 ( .A1(n8040), .A2(n8739), .ZN(n15381) );
  XOR2_X1 U15601 ( .A(n15554), .B(n15555), .Z(n15382) );
  XOR2_X1 U15602 ( .A(n15556), .B(n15557), .Z(n15555) );
  XOR2_X1 U15603 ( .A(n15558), .B(n15559), .Z(n15386) );
  XOR2_X1 U15604 ( .A(n15560), .B(n15561), .Z(n15559) );
  XOR2_X1 U15605 ( .A(n15562), .B(n15563), .Z(n15390) );
  XOR2_X1 U15606 ( .A(n15564), .B(n15565), .Z(n15563) );
  XOR2_X1 U15607 ( .A(n15566), .B(n15567), .Z(n15394) );
  XOR2_X1 U15608 ( .A(n15568), .B(n15569), .Z(n15567) );
  XOR2_X1 U15609 ( .A(n15570), .B(n15571), .Z(n15398) );
  XOR2_X1 U15610 ( .A(n15572), .B(n15573), .Z(n15571) );
  XOR2_X1 U15611 ( .A(n15574), .B(n15575), .Z(n15402) );
  XOR2_X1 U15612 ( .A(n15576), .B(n15577), .Z(n15575) );
  XOR2_X1 U15613 ( .A(n15578), .B(n15579), .Z(n15406) );
  XOR2_X1 U15614 ( .A(n15580), .B(n15581), .Z(n15579) );
  XOR2_X1 U15615 ( .A(n15582), .B(n15583), .Z(n15410) );
  XOR2_X1 U15616 ( .A(n15584), .B(n15585), .Z(n15583) );
  XOR2_X1 U15617 ( .A(n15586), .B(n15587), .Z(n15414) );
  XOR2_X1 U15618 ( .A(n15588), .B(n15589), .Z(n15587) );
  XOR2_X1 U15619 ( .A(n15590), .B(n15591), .Z(n15418) );
  XOR2_X1 U15620 ( .A(n15592), .B(n15593), .Z(n15591) );
  XOR2_X1 U15621 ( .A(n15594), .B(n15595), .Z(n15422) );
  XOR2_X1 U15622 ( .A(n15596), .B(n15597), .Z(n15595) );
  XOR2_X1 U15623 ( .A(n15598), .B(n15599), .Z(n15426) );
  XOR2_X1 U15624 ( .A(n15600), .B(n15601), .Z(n15599) );
  XOR2_X1 U15625 ( .A(n15602), .B(n15603), .Z(n15430) );
  XOR2_X1 U15626 ( .A(n15604), .B(n15605), .Z(n15603) );
  XOR2_X1 U15627 ( .A(n15606), .B(n15607), .Z(n15434) );
  XOR2_X1 U15628 ( .A(n15608), .B(n15609), .Z(n15607) );
  XOR2_X1 U15629 ( .A(n15610), .B(n15611), .Z(n15438) );
  XOR2_X1 U15630 ( .A(n15612), .B(n15613), .Z(n15611) );
  XOR2_X1 U15631 ( .A(n15614), .B(n15615), .Z(n15442) );
  XOR2_X1 U15632 ( .A(n15616), .B(n15617), .Z(n15615) );
  XOR2_X1 U15633 ( .A(n15618), .B(n15619), .Z(n15446) );
  XOR2_X1 U15634 ( .A(n15620), .B(n15621), .Z(n15619) );
  XOR2_X1 U15635 ( .A(n15622), .B(n15623), .Z(n15450) );
  XOR2_X1 U15636 ( .A(n15624), .B(n15625), .Z(n15623) );
  XOR2_X1 U15637 ( .A(n15626), .B(n15627), .Z(n15454) );
  XOR2_X1 U15638 ( .A(n15628), .B(n15629), .Z(n15627) );
  XOR2_X1 U15639 ( .A(n15630), .B(n15631), .Z(n15458) );
  XOR2_X1 U15640 ( .A(n15632), .B(n15633), .Z(n15631) );
  XOR2_X1 U15641 ( .A(n15634), .B(n15635), .Z(n9406) );
  XOR2_X1 U15642 ( .A(n15636), .B(n15637), .Z(n15635) );
  AND3_X1 U15643 ( .A1(n8942), .A2(n8940), .A3(n8941), .ZN(n8943) );
  INV_X1 U15644 ( .A(n15638), .ZN(n8941) );
  OR2_X1 U15645 ( .A1(n15639), .A2(n15640), .ZN(n15638) );
  AND2_X1 U15646 ( .A1(n9239), .A2(n9238), .ZN(n15640) );
  AND2_X1 U15647 ( .A1(n9236), .A2(n15641), .ZN(n15639) );
  OR2_X1 U15648 ( .A1(n9238), .A2(n9239), .ZN(n15641) );
  OR2_X1 U15649 ( .A1(n9248), .A2(n8735), .ZN(n9239) );
  OR2_X1 U15650 ( .A1(n15642), .A2(n15643), .ZN(n9238) );
  AND2_X1 U15651 ( .A1(n9258), .A2(n9257), .ZN(n15643) );
  AND2_X1 U15652 ( .A1(n9255), .A2(n15644), .ZN(n15642) );
  OR2_X1 U15653 ( .A1(n9257), .A2(n9258), .ZN(n15644) );
  OR2_X1 U15654 ( .A1(n8730), .A2(n8735), .ZN(n9258) );
  OR2_X1 U15655 ( .A1(n15645), .A2(n15646), .ZN(n9257) );
  AND2_X1 U15656 ( .A1(n8671), .A2(n9289), .ZN(n15646) );
  AND2_X1 U15657 ( .A1(n9287), .A2(n15647), .ZN(n15645) );
  OR2_X1 U15658 ( .A1(n9289), .A2(n8671), .ZN(n15647) );
  OR2_X1 U15659 ( .A1(n8734), .A2(n8735), .ZN(n8671) );
  OR2_X1 U15660 ( .A1(n15648), .A2(n15649), .ZN(n9289) );
  AND2_X1 U15661 ( .A1(n9320), .A2(n9319), .ZN(n15649) );
  AND2_X1 U15662 ( .A1(n9317), .A2(n15650), .ZN(n15648) );
  OR2_X1 U15663 ( .A1(n9319), .A2(n9320), .ZN(n15650) );
  OR2_X1 U15664 ( .A1(n8738), .A2(n8735), .ZN(n9320) );
  OR2_X1 U15665 ( .A1(n15651), .A2(n15652), .ZN(n9319) );
  AND2_X1 U15666 ( .A1(n9366), .A2(n9365), .ZN(n15652) );
  AND2_X1 U15667 ( .A1(n9363), .A2(n15653), .ZN(n15651) );
  OR2_X1 U15668 ( .A1(n9365), .A2(n9366), .ZN(n15653) );
  OR2_X1 U15669 ( .A1(n8742), .A2(n8735), .ZN(n9366) );
  OR2_X1 U15670 ( .A1(n15654), .A2(n15655), .ZN(n9365) );
  AND2_X1 U15671 ( .A1(n9411), .A2(n9410), .ZN(n15655) );
  AND2_X1 U15672 ( .A1(n9408), .A2(n15656), .ZN(n15654) );
  OR2_X1 U15673 ( .A1(n9410), .A2(n9411), .ZN(n15656) );
  OR2_X1 U15674 ( .A1(n8746), .A2(n8735), .ZN(n9411) );
  OR2_X1 U15675 ( .A1(n15657), .A2(n15658), .ZN(n9410) );
  AND2_X1 U15676 ( .A1(n15637), .A2(n15636), .ZN(n15658) );
  AND2_X1 U15677 ( .A1(n15634), .A2(n15659), .ZN(n15657) );
  OR2_X1 U15678 ( .A1(n15636), .A2(n15637), .ZN(n15659) );
  OR2_X1 U15679 ( .A1(n8750), .A2(n8735), .ZN(n15637) );
  OR2_X1 U15680 ( .A1(n15660), .A2(n15661), .ZN(n15636) );
  AND2_X1 U15681 ( .A1(n15633), .A2(n15632), .ZN(n15661) );
  AND2_X1 U15682 ( .A1(n15630), .A2(n15662), .ZN(n15660) );
  OR2_X1 U15683 ( .A1(n15632), .A2(n15633), .ZN(n15662) );
  OR2_X1 U15684 ( .A1(n8754), .A2(n8735), .ZN(n15633) );
  OR2_X1 U15685 ( .A1(n15663), .A2(n15664), .ZN(n15632) );
  AND2_X1 U15686 ( .A1(n15629), .A2(n15628), .ZN(n15664) );
  AND2_X1 U15687 ( .A1(n15626), .A2(n15665), .ZN(n15663) );
  OR2_X1 U15688 ( .A1(n15628), .A2(n15629), .ZN(n15665) );
  OR2_X1 U15689 ( .A1(n8758), .A2(n8735), .ZN(n15629) );
  OR2_X1 U15690 ( .A1(n15666), .A2(n15667), .ZN(n15628) );
  AND2_X1 U15691 ( .A1(n15625), .A2(n15624), .ZN(n15667) );
  AND2_X1 U15692 ( .A1(n15622), .A2(n15668), .ZN(n15666) );
  OR2_X1 U15693 ( .A1(n15624), .A2(n15625), .ZN(n15668) );
  OR2_X1 U15694 ( .A1(n8762), .A2(n8735), .ZN(n15625) );
  OR2_X1 U15695 ( .A1(n15669), .A2(n15670), .ZN(n15624) );
  AND2_X1 U15696 ( .A1(n15621), .A2(n15620), .ZN(n15670) );
  AND2_X1 U15697 ( .A1(n15618), .A2(n15671), .ZN(n15669) );
  OR2_X1 U15698 ( .A1(n15620), .A2(n15621), .ZN(n15671) );
  OR2_X1 U15699 ( .A1(n8766), .A2(n8735), .ZN(n15621) );
  OR2_X1 U15700 ( .A1(n15672), .A2(n15673), .ZN(n15620) );
  AND2_X1 U15701 ( .A1(n15617), .A2(n15616), .ZN(n15673) );
  AND2_X1 U15702 ( .A1(n15614), .A2(n15674), .ZN(n15672) );
  OR2_X1 U15703 ( .A1(n15616), .A2(n15617), .ZN(n15674) );
  OR2_X1 U15704 ( .A1(n8770), .A2(n8735), .ZN(n15617) );
  OR2_X1 U15705 ( .A1(n15675), .A2(n15676), .ZN(n15616) );
  AND2_X1 U15706 ( .A1(n15613), .A2(n15612), .ZN(n15676) );
  AND2_X1 U15707 ( .A1(n15610), .A2(n15677), .ZN(n15675) );
  OR2_X1 U15708 ( .A1(n15612), .A2(n15613), .ZN(n15677) );
  OR2_X1 U15709 ( .A1(n8774), .A2(n8735), .ZN(n15613) );
  OR2_X1 U15710 ( .A1(n15678), .A2(n15679), .ZN(n15612) );
  AND2_X1 U15711 ( .A1(n15609), .A2(n15608), .ZN(n15679) );
  AND2_X1 U15712 ( .A1(n15606), .A2(n15680), .ZN(n15678) );
  OR2_X1 U15713 ( .A1(n15608), .A2(n15609), .ZN(n15680) );
  OR2_X1 U15714 ( .A1(n8778), .A2(n8735), .ZN(n15609) );
  OR2_X1 U15715 ( .A1(n15681), .A2(n15682), .ZN(n15608) );
  AND2_X1 U15716 ( .A1(n15605), .A2(n15604), .ZN(n15682) );
  AND2_X1 U15717 ( .A1(n15602), .A2(n15683), .ZN(n15681) );
  OR2_X1 U15718 ( .A1(n15604), .A2(n15605), .ZN(n15683) );
  OR2_X1 U15719 ( .A1(n8782), .A2(n8735), .ZN(n15605) );
  OR2_X1 U15720 ( .A1(n15684), .A2(n15685), .ZN(n15604) );
  AND2_X1 U15721 ( .A1(n15601), .A2(n15600), .ZN(n15685) );
  AND2_X1 U15722 ( .A1(n15598), .A2(n15686), .ZN(n15684) );
  OR2_X1 U15723 ( .A1(n15600), .A2(n15601), .ZN(n15686) );
  OR2_X1 U15724 ( .A1(n8786), .A2(n8735), .ZN(n15601) );
  OR2_X1 U15725 ( .A1(n15687), .A2(n15688), .ZN(n15600) );
  AND2_X1 U15726 ( .A1(n15597), .A2(n15596), .ZN(n15688) );
  AND2_X1 U15727 ( .A1(n15594), .A2(n15689), .ZN(n15687) );
  OR2_X1 U15728 ( .A1(n15596), .A2(n15597), .ZN(n15689) );
  OR2_X1 U15729 ( .A1(n8790), .A2(n8735), .ZN(n15597) );
  OR2_X1 U15730 ( .A1(n15690), .A2(n15691), .ZN(n15596) );
  AND2_X1 U15731 ( .A1(n15593), .A2(n15592), .ZN(n15691) );
  AND2_X1 U15732 ( .A1(n15590), .A2(n15692), .ZN(n15690) );
  OR2_X1 U15733 ( .A1(n15592), .A2(n15593), .ZN(n15692) );
  OR2_X1 U15734 ( .A1(n8794), .A2(n8735), .ZN(n15593) );
  OR2_X1 U15735 ( .A1(n15693), .A2(n15694), .ZN(n15592) );
  AND2_X1 U15736 ( .A1(n15589), .A2(n15588), .ZN(n15694) );
  AND2_X1 U15737 ( .A1(n15586), .A2(n15695), .ZN(n15693) );
  OR2_X1 U15738 ( .A1(n15588), .A2(n15589), .ZN(n15695) );
  OR2_X1 U15739 ( .A1(n8798), .A2(n8735), .ZN(n15589) );
  OR2_X1 U15740 ( .A1(n15696), .A2(n15697), .ZN(n15588) );
  AND2_X1 U15741 ( .A1(n15585), .A2(n15584), .ZN(n15697) );
  AND2_X1 U15742 ( .A1(n15582), .A2(n15698), .ZN(n15696) );
  OR2_X1 U15743 ( .A1(n15584), .A2(n15585), .ZN(n15698) );
  OR2_X1 U15744 ( .A1(n8802), .A2(n8735), .ZN(n15585) );
  OR2_X1 U15745 ( .A1(n15699), .A2(n15700), .ZN(n15584) );
  AND2_X1 U15746 ( .A1(n15581), .A2(n15580), .ZN(n15700) );
  AND2_X1 U15747 ( .A1(n15578), .A2(n15701), .ZN(n15699) );
  OR2_X1 U15748 ( .A1(n15580), .A2(n15581), .ZN(n15701) );
  OR2_X1 U15749 ( .A1(n8806), .A2(n8735), .ZN(n15581) );
  OR2_X1 U15750 ( .A1(n15702), .A2(n15703), .ZN(n15580) );
  AND2_X1 U15751 ( .A1(n15577), .A2(n15576), .ZN(n15703) );
  AND2_X1 U15752 ( .A1(n15574), .A2(n15704), .ZN(n15702) );
  OR2_X1 U15753 ( .A1(n15576), .A2(n15577), .ZN(n15704) );
  OR2_X1 U15754 ( .A1(n8810), .A2(n8735), .ZN(n15577) );
  OR2_X1 U15755 ( .A1(n15705), .A2(n15706), .ZN(n15576) );
  AND2_X1 U15756 ( .A1(n15573), .A2(n15572), .ZN(n15706) );
  AND2_X1 U15757 ( .A1(n15570), .A2(n15707), .ZN(n15705) );
  OR2_X1 U15758 ( .A1(n15572), .A2(n15573), .ZN(n15707) );
  OR2_X1 U15759 ( .A1(n8140), .A2(n8735), .ZN(n15573) );
  OR2_X1 U15760 ( .A1(n15708), .A2(n15709), .ZN(n15572) );
  AND2_X1 U15761 ( .A1(n15569), .A2(n15568), .ZN(n15709) );
  AND2_X1 U15762 ( .A1(n15566), .A2(n15710), .ZN(n15708) );
  OR2_X1 U15763 ( .A1(n15568), .A2(n15569), .ZN(n15710) );
  OR2_X1 U15764 ( .A1(n8115), .A2(n8735), .ZN(n15569) );
  OR2_X1 U15765 ( .A1(n15711), .A2(n15712), .ZN(n15568) );
  AND2_X1 U15766 ( .A1(n15565), .A2(n15564), .ZN(n15712) );
  AND2_X1 U15767 ( .A1(n15562), .A2(n15713), .ZN(n15711) );
  OR2_X1 U15768 ( .A1(n15564), .A2(n15565), .ZN(n15713) );
  OR2_X1 U15769 ( .A1(n8090), .A2(n8735), .ZN(n15565) );
  OR2_X1 U15770 ( .A1(n15714), .A2(n15715), .ZN(n15564) );
  AND2_X1 U15771 ( .A1(n15561), .A2(n15560), .ZN(n15715) );
  AND2_X1 U15772 ( .A1(n15558), .A2(n15716), .ZN(n15714) );
  OR2_X1 U15773 ( .A1(n15560), .A2(n15561), .ZN(n15716) );
  OR2_X1 U15774 ( .A1(n8065), .A2(n8735), .ZN(n15561) );
  OR2_X1 U15775 ( .A1(n15717), .A2(n15718), .ZN(n15560) );
  AND2_X1 U15776 ( .A1(n15557), .A2(n15556), .ZN(n15718) );
  AND2_X1 U15777 ( .A1(n15554), .A2(n15719), .ZN(n15717) );
  OR2_X1 U15778 ( .A1(n15556), .A2(n15557), .ZN(n15719) );
  OR2_X1 U15779 ( .A1(n8040), .A2(n8735), .ZN(n15557) );
  OR2_X1 U15780 ( .A1(n15720), .A2(n15721), .ZN(n15556) );
  AND2_X1 U15781 ( .A1(n15550), .A2(n15553), .ZN(n15721) );
  AND2_X1 U15782 ( .A1(n15722), .A2(n15552), .ZN(n15720) );
  OR2_X1 U15783 ( .A1(n15723), .A2(n15724), .ZN(n15552) );
  AND2_X1 U15784 ( .A1(n15549), .A2(n15548), .ZN(n15724) );
  AND2_X1 U15785 ( .A1(n15546), .A2(n15725), .ZN(n15723) );
  OR2_X1 U15786 ( .A1(n15548), .A2(n15549), .ZN(n15725) );
  OR2_X1 U15787 ( .A1(n7979), .A2(n8735), .ZN(n15549) );
  OR2_X1 U15788 ( .A1(n15726), .A2(n15727), .ZN(n15548) );
  AND2_X1 U15789 ( .A1(n15542), .A2(n15545), .ZN(n15727) );
  AND2_X1 U15790 ( .A1(n15728), .A2(n15729), .ZN(n15726) );
  OR2_X1 U15791 ( .A1(n15545), .A2(n15542), .ZN(n15729) );
  OR2_X1 U15792 ( .A1(n7954), .A2(n8735), .ZN(n15542) );
  OR3_X1 U15793 ( .A1(n8735), .A2(n8731), .A3(n9796), .ZN(n15545) );
  INV_X1 U15794 ( .A(n15544), .ZN(n15728) );
  OR2_X1 U15795 ( .A1(n15730), .A2(n15731), .ZN(n15544) );
  AND2_X1 U15796 ( .A1(b_1_), .A2(n15732), .ZN(n15731) );
  OR2_X1 U15797 ( .A1(n15733), .A2(n9801), .ZN(n15732) );
  AND2_X1 U15798 ( .A1(n8847), .A2(a_30_), .ZN(n9801) );
  AND2_X1 U15799 ( .A1(a_30_), .A2(n9126), .ZN(n15733) );
  AND2_X1 U15800 ( .A1(b_0_), .A2(n15734), .ZN(n15730) );
  OR2_X1 U15801 ( .A1(n15735), .A2(n7920), .ZN(n15734) );
  AND2_X1 U15802 ( .A1(n7914), .A2(a_31_), .ZN(n7920) );
  AND2_X1 U15803 ( .A1(a_31_), .A2(n8731), .ZN(n15735) );
  XNOR2_X1 U15804 ( .A(n15736), .B(n15737), .ZN(n15546) );
  OR2_X1 U15805 ( .A1(n15738), .A2(n15739), .ZN(n15736) );
  INV_X1 U15806 ( .A(n15740), .ZN(n15739) );
  AND2_X1 U15807 ( .A1(n15741), .A2(n15742), .ZN(n15738) );
  OR2_X1 U15808 ( .A1(n9126), .A2(n7914), .ZN(n15741) );
  OR2_X1 U15809 ( .A1(n15553), .A2(n15550), .ZN(n15722) );
  XOR2_X1 U15810 ( .A(n15743), .B(n15744), .Z(n15550) );
  XOR2_X1 U15811 ( .A(n15745), .B(n15746), .Z(n15743) );
  OR2_X1 U15812 ( .A1(n8015), .A2(n8735), .ZN(n15553) );
  XNOR2_X1 U15813 ( .A(n15747), .B(n15748), .ZN(n15554) );
  XNOR2_X1 U15814 ( .A(n15749), .B(n15750), .ZN(n15747) );
  XNOR2_X1 U15815 ( .A(n15751), .B(n15752), .ZN(n15558) );
  XNOR2_X1 U15816 ( .A(n15753), .B(n15754), .ZN(n15751) );
  XNOR2_X1 U15817 ( .A(n15755), .B(n15756), .ZN(n15562) );
  XNOR2_X1 U15818 ( .A(n15757), .B(n15758), .ZN(n15755) );
  XNOR2_X1 U15819 ( .A(n15759), .B(n15760), .ZN(n15566) );
  XNOR2_X1 U15820 ( .A(n15761), .B(n15762), .ZN(n15759) );
  XNOR2_X1 U15821 ( .A(n15763), .B(n15764), .ZN(n15570) );
  XNOR2_X1 U15822 ( .A(n15765), .B(n15766), .ZN(n15763) );
  XNOR2_X1 U15823 ( .A(n15767), .B(n15768), .ZN(n15574) );
  XNOR2_X1 U15824 ( .A(n15769), .B(n15770), .ZN(n15767) );
  XNOR2_X1 U15825 ( .A(n15771), .B(n15772), .ZN(n15578) );
  XNOR2_X1 U15826 ( .A(n15773), .B(n15774), .ZN(n15771) );
  XNOR2_X1 U15827 ( .A(n15775), .B(n15776), .ZN(n15582) );
  XNOR2_X1 U15828 ( .A(n15777), .B(n15778), .ZN(n15775) );
  XNOR2_X1 U15829 ( .A(n15779), .B(n15780), .ZN(n15586) );
  XNOR2_X1 U15830 ( .A(n15781), .B(n15782), .ZN(n15779) );
  XNOR2_X1 U15831 ( .A(n15783), .B(n15784), .ZN(n15590) );
  XNOR2_X1 U15832 ( .A(n15785), .B(n15786), .ZN(n15783) );
  XNOR2_X1 U15833 ( .A(n15787), .B(n15788), .ZN(n15594) );
  XNOR2_X1 U15834 ( .A(n15789), .B(n15790), .ZN(n15787) );
  XNOR2_X1 U15835 ( .A(n15791), .B(n15792), .ZN(n15598) );
  XNOR2_X1 U15836 ( .A(n15793), .B(n15794), .ZN(n15791) );
  XNOR2_X1 U15837 ( .A(n15795), .B(n15796), .ZN(n15602) );
  XNOR2_X1 U15838 ( .A(n15797), .B(n15798), .ZN(n15795) );
  XNOR2_X1 U15839 ( .A(n15799), .B(n15800), .ZN(n15606) );
  XNOR2_X1 U15840 ( .A(n15801), .B(n15802), .ZN(n15799) );
  XNOR2_X1 U15841 ( .A(n15803), .B(n15804), .ZN(n15610) );
  XNOR2_X1 U15842 ( .A(n15805), .B(n15806), .ZN(n15803) );
  XNOR2_X1 U15843 ( .A(n15807), .B(n15808), .ZN(n15614) );
  XNOR2_X1 U15844 ( .A(n15809), .B(n15810), .ZN(n15807) );
  XNOR2_X1 U15845 ( .A(n15811), .B(n15812), .ZN(n15618) );
  XNOR2_X1 U15846 ( .A(n15813), .B(n15814), .ZN(n15811) );
  XNOR2_X1 U15847 ( .A(n15815), .B(n15816), .ZN(n15622) );
  XNOR2_X1 U15848 ( .A(n15817), .B(n15818), .ZN(n15815) );
  XNOR2_X1 U15849 ( .A(n15819), .B(n15820), .ZN(n15626) );
  XNOR2_X1 U15850 ( .A(n15821), .B(n15822), .ZN(n15819) );
  XOR2_X1 U15851 ( .A(n15823), .B(n15824), .Z(n15630) );
  XOR2_X1 U15852 ( .A(n15825), .B(n15826), .Z(n15824) );
  XOR2_X1 U15853 ( .A(n15827), .B(n15828), .Z(n15634) );
  XOR2_X1 U15854 ( .A(n15829), .B(n15830), .Z(n15828) );
  XOR2_X1 U15855 ( .A(n15831), .B(n15832), .Z(n9408) );
  XOR2_X1 U15856 ( .A(n15833), .B(n15834), .Z(n15832) );
  XOR2_X1 U15857 ( .A(n15835), .B(n15836), .Z(n9363) );
  XOR2_X1 U15858 ( .A(n15837), .B(n15838), .Z(n15836) );
  XOR2_X1 U15859 ( .A(n15839), .B(n15840), .Z(n9317) );
  XOR2_X1 U15860 ( .A(n15841), .B(n15842), .Z(n15840) );
  XOR2_X1 U15861 ( .A(n15843), .B(n15844), .Z(n9287) );
  XOR2_X1 U15862 ( .A(n15845), .B(n15846), .Z(n15844) );
  XOR2_X1 U15863 ( .A(n15847), .B(n15848), .Z(n9255) );
  XOR2_X1 U15864 ( .A(n15849), .B(n15850), .Z(n15848) );
  XOR2_X1 U15865 ( .A(n15851), .B(n15852), .Z(n9236) );
  XOR2_X1 U15866 ( .A(n15853), .B(n8697), .Z(n15852) );
  XOR2_X1 U15867 ( .A(n15854), .B(n9221), .Z(n8940) );
  OR2_X1 U15868 ( .A1(n15855), .A2(n15856), .ZN(n9221) );
  AND2_X1 U15869 ( .A1(n15857), .A2(n15858), .ZN(n15856) );
  AND2_X1 U15870 ( .A1(n15859), .A2(n15860), .ZN(n15855) );
  OR2_X1 U15871 ( .A1(n15858), .A2(n15857), .ZN(n15859) );
  OR2_X1 U15872 ( .A1(n9126), .A2(n9248), .ZN(n15854) );
  XOR2_X1 U15873 ( .A(n15861), .B(n15857), .Z(n8942) );
  OR2_X1 U15874 ( .A1(n15862), .A2(n15863), .ZN(n15857) );
  AND2_X1 U15875 ( .A1(n15851), .A2(n15853), .ZN(n15863) );
  AND2_X1 U15876 ( .A1(n15864), .A2(n8697), .ZN(n15862) );
  OR2_X1 U15877 ( .A1(n8730), .A2(n8731), .ZN(n8697) );
  OR2_X1 U15878 ( .A1(n15853), .A2(n15851), .ZN(n15864) );
  OR2_X1 U15879 ( .A1(n9126), .A2(n8734), .ZN(n15851) );
  OR2_X1 U15880 ( .A1(n15865), .A2(n15866), .ZN(n15853) );
  AND2_X1 U15881 ( .A1(n15847), .A2(n15849), .ZN(n15866) );
  AND2_X1 U15882 ( .A1(n15867), .A2(n15850), .ZN(n15865) );
  OR2_X1 U15883 ( .A1(n9126), .A2(n8738), .ZN(n15850) );
  OR2_X1 U15884 ( .A1(n15849), .A2(n15847), .ZN(n15867) );
  OR2_X1 U15885 ( .A1(n8734), .A2(n8731), .ZN(n15847) );
  INV_X1 U15886 ( .A(a_2_), .ZN(n8734) );
  OR2_X1 U15887 ( .A1(n15868), .A2(n15869), .ZN(n15849) );
  AND2_X1 U15888 ( .A1(n15843), .A2(n15845), .ZN(n15869) );
  AND2_X1 U15889 ( .A1(n15870), .A2(n15846), .ZN(n15868) );
  OR2_X1 U15890 ( .A1(n9126), .A2(n8742), .ZN(n15846) );
  OR2_X1 U15891 ( .A1(n15845), .A2(n15843), .ZN(n15870) );
  OR2_X1 U15892 ( .A1(n8738), .A2(n8731), .ZN(n15843) );
  INV_X1 U15893 ( .A(a_3_), .ZN(n8738) );
  OR2_X1 U15894 ( .A1(n15871), .A2(n15872), .ZN(n15845) );
  AND2_X1 U15895 ( .A1(n15839), .A2(n15841), .ZN(n15872) );
  AND2_X1 U15896 ( .A1(n15873), .A2(n15842), .ZN(n15871) );
  OR2_X1 U15897 ( .A1(n9126), .A2(n8746), .ZN(n15842) );
  OR2_X1 U15898 ( .A1(n15841), .A2(n15839), .ZN(n15873) );
  OR2_X1 U15899 ( .A1(n8742), .A2(n8731), .ZN(n15839) );
  INV_X1 U15900 ( .A(a_4_), .ZN(n8742) );
  OR2_X1 U15901 ( .A1(n15874), .A2(n15875), .ZN(n15841) );
  AND2_X1 U15902 ( .A1(n15835), .A2(n15837), .ZN(n15875) );
  AND2_X1 U15903 ( .A1(n15876), .A2(n15838), .ZN(n15874) );
  OR2_X1 U15904 ( .A1(n9126), .A2(n8750), .ZN(n15838) );
  OR2_X1 U15905 ( .A1(n15837), .A2(n15835), .ZN(n15876) );
  OR2_X1 U15906 ( .A1(n8746), .A2(n8731), .ZN(n15835) );
  INV_X1 U15907 ( .A(a_5_), .ZN(n8746) );
  OR2_X1 U15908 ( .A1(n15877), .A2(n15878), .ZN(n15837) );
  AND2_X1 U15909 ( .A1(n15831), .A2(n15833), .ZN(n15878) );
  AND2_X1 U15910 ( .A1(n15879), .A2(n15834), .ZN(n15877) );
  OR2_X1 U15911 ( .A1(n9126), .A2(n8754), .ZN(n15834) );
  OR2_X1 U15912 ( .A1(n15833), .A2(n15831), .ZN(n15879) );
  OR2_X1 U15913 ( .A1(n8750), .A2(n8731), .ZN(n15831) );
  INV_X1 U15914 ( .A(a_6_), .ZN(n8750) );
  OR2_X1 U15915 ( .A1(n15880), .A2(n15881), .ZN(n15833) );
  AND2_X1 U15916 ( .A1(n15827), .A2(n15829), .ZN(n15881) );
  AND2_X1 U15917 ( .A1(n15882), .A2(n15830), .ZN(n15880) );
  OR2_X1 U15918 ( .A1(n9126), .A2(n8758), .ZN(n15830) );
  OR2_X1 U15919 ( .A1(n15829), .A2(n15827), .ZN(n15882) );
  OR2_X1 U15920 ( .A1(n8754), .A2(n8731), .ZN(n15827) );
  INV_X1 U15921 ( .A(a_7_), .ZN(n8754) );
  OR2_X1 U15922 ( .A1(n15883), .A2(n15884), .ZN(n15829) );
  AND2_X1 U15923 ( .A1(n15823), .A2(n15825), .ZN(n15884) );
  AND2_X1 U15924 ( .A1(n15885), .A2(n15826), .ZN(n15883) );
  OR2_X1 U15925 ( .A1(n9126), .A2(n8762), .ZN(n15826) );
  OR2_X1 U15926 ( .A1(n15825), .A2(n15823), .ZN(n15885) );
  OR2_X1 U15927 ( .A1(n8758), .A2(n8731), .ZN(n15823) );
  INV_X1 U15928 ( .A(a_8_), .ZN(n8758) );
  OR2_X1 U15929 ( .A1(n15886), .A2(n15887), .ZN(n15825) );
  AND2_X1 U15930 ( .A1(n15820), .A2(n15822), .ZN(n15887) );
  AND2_X1 U15931 ( .A1(n15888), .A2(n15821), .ZN(n15886) );
  OR2_X1 U15932 ( .A1(n9126), .A2(n8766), .ZN(n15821) );
  OR2_X1 U15933 ( .A1(n15822), .A2(n15820), .ZN(n15888) );
  OR2_X1 U15934 ( .A1(n8762), .A2(n8731), .ZN(n15820) );
  INV_X1 U15935 ( .A(a_9_), .ZN(n8762) );
  OR2_X1 U15936 ( .A1(n15889), .A2(n15890), .ZN(n15822) );
  AND2_X1 U15937 ( .A1(n15816), .A2(n15818), .ZN(n15890) );
  AND2_X1 U15938 ( .A1(n15891), .A2(n15817), .ZN(n15889) );
  OR2_X1 U15939 ( .A1(n9126), .A2(n8770), .ZN(n15817) );
  OR2_X1 U15940 ( .A1(n15818), .A2(n15816), .ZN(n15891) );
  OR2_X1 U15941 ( .A1(n8766), .A2(n8731), .ZN(n15816) );
  INV_X1 U15942 ( .A(a_10_), .ZN(n8766) );
  OR2_X1 U15943 ( .A1(n15892), .A2(n15893), .ZN(n15818) );
  AND2_X1 U15944 ( .A1(n15812), .A2(n15814), .ZN(n15893) );
  AND2_X1 U15945 ( .A1(n15894), .A2(n15813), .ZN(n15892) );
  OR2_X1 U15946 ( .A1(n9126), .A2(n8774), .ZN(n15813) );
  OR2_X1 U15947 ( .A1(n15814), .A2(n15812), .ZN(n15894) );
  OR2_X1 U15948 ( .A1(n8770), .A2(n8731), .ZN(n15812) );
  INV_X1 U15949 ( .A(a_11_), .ZN(n8770) );
  OR2_X1 U15950 ( .A1(n15895), .A2(n15896), .ZN(n15814) );
  AND2_X1 U15951 ( .A1(n15808), .A2(n15810), .ZN(n15896) );
  AND2_X1 U15952 ( .A1(n15897), .A2(n15809), .ZN(n15895) );
  OR2_X1 U15953 ( .A1(n9126), .A2(n8778), .ZN(n15809) );
  OR2_X1 U15954 ( .A1(n15810), .A2(n15808), .ZN(n15897) );
  OR2_X1 U15955 ( .A1(n8774), .A2(n8731), .ZN(n15808) );
  INV_X1 U15956 ( .A(a_12_), .ZN(n8774) );
  OR2_X1 U15957 ( .A1(n15898), .A2(n15899), .ZN(n15810) );
  AND2_X1 U15958 ( .A1(n15804), .A2(n15806), .ZN(n15899) );
  AND2_X1 U15959 ( .A1(n15900), .A2(n15805), .ZN(n15898) );
  OR2_X1 U15960 ( .A1(n9126), .A2(n8782), .ZN(n15805) );
  OR2_X1 U15961 ( .A1(n15806), .A2(n15804), .ZN(n15900) );
  OR2_X1 U15962 ( .A1(n8778), .A2(n8731), .ZN(n15804) );
  INV_X1 U15963 ( .A(a_13_), .ZN(n8778) );
  OR2_X1 U15964 ( .A1(n15901), .A2(n15902), .ZN(n15806) );
  AND2_X1 U15965 ( .A1(n15800), .A2(n15802), .ZN(n15902) );
  AND2_X1 U15966 ( .A1(n15903), .A2(n15801), .ZN(n15901) );
  OR2_X1 U15967 ( .A1(n9126), .A2(n8786), .ZN(n15801) );
  OR2_X1 U15968 ( .A1(n15802), .A2(n15800), .ZN(n15903) );
  OR2_X1 U15969 ( .A1(n8782), .A2(n8731), .ZN(n15800) );
  INV_X1 U15970 ( .A(a_14_), .ZN(n8782) );
  OR2_X1 U15971 ( .A1(n15904), .A2(n15905), .ZN(n15802) );
  AND2_X1 U15972 ( .A1(n15796), .A2(n15798), .ZN(n15905) );
  AND2_X1 U15973 ( .A1(n15906), .A2(n15797), .ZN(n15904) );
  OR2_X1 U15974 ( .A1(n9126), .A2(n8790), .ZN(n15797) );
  OR2_X1 U15975 ( .A1(n15798), .A2(n15796), .ZN(n15906) );
  OR2_X1 U15976 ( .A1(n8786), .A2(n8731), .ZN(n15796) );
  INV_X1 U15977 ( .A(a_15_), .ZN(n8786) );
  OR2_X1 U15978 ( .A1(n15907), .A2(n15908), .ZN(n15798) );
  AND2_X1 U15979 ( .A1(n15792), .A2(n15794), .ZN(n15908) );
  AND2_X1 U15980 ( .A1(n15909), .A2(n15793), .ZN(n15907) );
  OR2_X1 U15981 ( .A1(n9126), .A2(n8794), .ZN(n15793) );
  OR2_X1 U15982 ( .A1(n15794), .A2(n15792), .ZN(n15909) );
  OR2_X1 U15983 ( .A1(n8790), .A2(n8731), .ZN(n15792) );
  INV_X1 U15984 ( .A(a_16_), .ZN(n8790) );
  OR2_X1 U15985 ( .A1(n15910), .A2(n15911), .ZN(n15794) );
  AND2_X1 U15986 ( .A1(n15788), .A2(n15790), .ZN(n15911) );
  AND2_X1 U15987 ( .A1(n15912), .A2(n15789), .ZN(n15910) );
  OR2_X1 U15988 ( .A1(n9126), .A2(n8798), .ZN(n15789) );
  OR2_X1 U15989 ( .A1(n15790), .A2(n15788), .ZN(n15912) );
  OR2_X1 U15990 ( .A1(n8794), .A2(n8731), .ZN(n15788) );
  INV_X1 U15991 ( .A(a_17_), .ZN(n8794) );
  OR2_X1 U15992 ( .A1(n15913), .A2(n15914), .ZN(n15790) );
  AND2_X1 U15993 ( .A1(n15784), .A2(n15786), .ZN(n15914) );
  AND2_X1 U15994 ( .A1(n15915), .A2(n15785), .ZN(n15913) );
  OR2_X1 U15995 ( .A1(n9126), .A2(n8802), .ZN(n15785) );
  OR2_X1 U15996 ( .A1(n15786), .A2(n15784), .ZN(n15915) );
  OR2_X1 U15997 ( .A1(n8798), .A2(n8731), .ZN(n15784) );
  INV_X1 U15998 ( .A(a_18_), .ZN(n8798) );
  OR2_X1 U15999 ( .A1(n15916), .A2(n15917), .ZN(n15786) );
  AND2_X1 U16000 ( .A1(n15780), .A2(n15782), .ZN(n15917) );
  AND2_X1 U16001 ( .A1(n15918), .A2(n15781), .ZN(n15916) );
  OR2_X1 U16002 ( .A1(n9126), .A2(n8806), .ZN(n15781) );
  OR2_X1 U16003 ( .A1(n15782), .A2(n15780), .ZN(n15918) );
  OR2_X1 U16004 ( .A1(n8802), .A2(n8731), .ZN(n15780) );
  INV_X1 U16005 ( .A(a_19_), .ZN(n8802) );
  OR2_X1 U16006 ( .A1(n15919), .A2(n15920), .ZN(n15782) );
  AND2_X1 U16007 ( .A1(n15776), .A2(n15778), .ZN(n15920) );
  AND2_X1 U16008 ( .A1(n15921), .A2(n15777), .ZN(n15919) );
  OR2_X1 U16009 ( .A1(n9126), .A2(n8810), .ZN(n15777) );
  OR2_X1 U16010 ( .A1(n15778), .A2(n15776), .ZN(n15921) );
  OR2_X1 U16011 ( .A1(n8806), .A2(n8731), .ZN(n15776) );
  INV_X1 U16012 ( .A(a_20_), .ZN(n8806) );
  OR2_X1 U16013 ( .A1(n15922), .A2(n15923), .ZN(n15778) );
  AND2_X1 U16014 ( .A1(n15772), .A2(n15774), .ZN(n15923) );
  AND2_X1 U16015 ( .A1(n15924), .A2(n15773), .ZN(n15922) );
  OR2_X1 U16016 ( .A1(n9126), .A2(n8140), .ZN(n15773) );
  OR2_X1 U16017 ( .A1(n15774), .A2(n15772), .ZN(n15924) );
  OR2_X1 U16018 ( .A1(n8810), .A2(n8731), .ZN(n15772) );
  INV_X1 U16019 ( .A(a_21_), .ZN(n8810) );
  OR2_X1 U16020 ( .A1(n15925), .A2(n15926), .ZN(n15774) );
  AND2_X1 U16021 ( .A1(n15768), .A2(n15770), .ZN(n15926) );
  AND2_X1 U16022 ( .A1(n15927), .A2(n15769), .ZN(n15925) );
  OR2_X1 U16023 ( .A1(n9126), .A2(n8115), .ZN(n15769) );
  OR2_X1 U16024 ( .A1(n15770), .A2(n15768), .ZN(n15927) );
  OR2_X1 U16025 ( .A1(n8140), .A2(n8731), .ZN(n15768) );
  OR2_X1 U16026 ( .A1(n15928), .A2(n15929), .ZN(n15770) );
  AND2_X1 U16027 ( .A1(n15764), .A2(n15766), .ZN(n15929) );
  AND2_X1 U16028 ( .A1(n15930), .A2(n15765), .ZN(n15928) );
  OR2_X1 U16029 ( .A1(n9126), .A2(n8090), .ZN(n15765) );
  OR2_X1 U16030 ( .A1(n15766), .A2(n15764), .ZN(n15930) );
  OR2_X1 U16031 ( .A1(n8115), .A2(n8731), .ZN(n15764) );
  OR2_X1 U16032 ( .A1(n15931), .A2(n15932), .ZN(n15766) );
  AND2_X1 U16033 ( .A1(n15760), .A2(n15762), .ZN(n15932) );
  AND2_X1 U16034 ( .A1(n15933), .A2(n15761), .ZN(n15931) );
  OR2_X1 U16035 ( .A1(n9126), .A2(n8065), .ZN(n15761) );
  OR2_X1 U16036 ( .A1(n15762), .A2(n15760), .ZN(n15933) );
  OR2_X1 U16037 ( .A1(n8090), .A2(n8731), .ZN(n15760) );
  OR2_X1 U16038 ( .A1(n15934), .A2(n15935), .ZN(n15762) );
  AND2_X1 U16039 ( .A1(n15756), .A2(n15758), .ZN(n15935) );
  AND2_X1 U16040 ( .A1(n15936), .A2(n15757), .ZN(n15934) );
  OR2_X1 U16041 ( .A1(n9126), .A2(n8040), .ZN(n15757) );
  OR2_X1 U16042 ( .A1(n15758), .A2(n15756), .ZN(n15936) );
  OR2_X1 U16043 ( .A1(n8065), .A2(n8731), .ZN(n15756) );
  OR2_X1 U16044 ( .A1(n15937), .A2(n15938), .ZN(n15758) );
  AND2_X1 U16045 ( .A1(n15752), .A2(n15754), .ZN(n15938) );
  AND2_X1 U16046 ( .A1(n15939), .A2(n15753), .ZN(n15937) );
  OR2_X1 U16047 ( .A1(n9126), .A2(n8015), .ZN(n15753) );
  OR2_X1 U16048 ( .A1(n15754), .A2(n15752), .ZN(n15939) );
  OR2_X1 U16049 ( .A1(n8040), .A2(n8731), .ZN(n15752) );
  OR2_X1 U16050 ( .A1(n15940), .A2(n15941), .ZN(n15754) );
  AND2_X1 U16051 ( .A1(n15748), .A2(n15750), .ZN(n15941) );
  AND2_X1 U16052 ( .A1(n15942), .A2(n15749), .ZN(n15940) );
  OR2_X1 U16053 ( .A1(n9126), .A2(n7979), .ZN(n15749) );
  OR2_X1 U16054 ( .A1(n15750), .A2(n15748), .ZN(n15942) );
  OR2_X1 U16055 ( .A1(n8015), .A2(n8731), .ZN(n15748) );
  OR2_X1 U16056 ( .A1(n15943), .A2(n15944), .ZN(n15750) );
  AND2_X1 U16057 ( .A1(n15744), .A2(n15746), .ZN(n15944) );
  AND2_X1 U16058 ( .A1(n15745), .A2(n15945), .ZN(n15943) );
  OR2_X1 U16059 ( .A1(n15746), .A2(n15744), .ZN(n15945) );
  OR2_X1 U16060 ( .A1(n7979), .A2(n8731), .ZN(n15744) );
  OR2_X1 U16061 ( .A1(n9126), .A2(n7954), .ZN(n15746) );
  AND2_X1 U16062 ( .A1(n15740), .A2(n15737), .ZN(n15745) );
  OR3_X1 U16063 ( .A1(n9126), .A2(n8731), .A3(n9796), .ZN(n15737) );
  OR2_X1 U16064 ( .A1(n8847), .A2(n7914), .ZN(n9796) );
  INV_X1 U16065 ( .A(a_31_), .ZN(n8847) );
  OR3_X1 U16066 ( .A1(n9126), .A2(n7914), .A3(n15742), .ZN(n15740) );
  OR2_X1 U16067 ( .A1(n7954), .A2(n8731), .ZN(n15742) );
  INV_X1 U16068 ( .A(a_30_), .ZN(n7914) );
  XNOR2_X1 U16069 ( .A(n15858), .B(n15860), .ZN(n15861) );
  OR2_X1 U16070 ( .A1(n9248), .A2(n8731), .ZN(n15860) );
  INV_X1 U16071 ( .A(a_0_), .ZN(n9248) );
  OR2_X1 U16072 ( .A1(n9126), .A2(n8730), .ZN(n15858) );
  INV_X1 U16073 ( .A(a_1_), .ZN(n8730) );
endmodule

