module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n859_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n695_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n823_, new_n431_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_26 );
not g001 ( new_n107_, keyIn_0_20 );
not g002 ( new_n108_, N85 );
and g003 ( new_n109_, new_n108_, N81 );
not g004 ( new_n110_, N81 );
and g005 ( new_n111_, new_n110_, N85 );
or g006 ( new_n112_, new_n109_, new_n111_ );
not g007 ( new_n113_, N93 );
and g008 ( new_n114_, new_n113_, N89 );
not g009 ( new_n115_, N89 );
and g010 ( new_n116_, new_n115_, N93 );
or g011 ( new_n117_, new_n114_, new_n116_ );
not g012 ( new_n118_, new_n117_ );
and g013 ( new_n119_, new_n118_, new_n112_ );
not g014 ( new_n120_, new_n119_ );
or g015 ( new_n121_, new_n118_, new_n112_ );
and g016 ( new_n122_, new_n120_, new_n121_ );
not g017 ( new_n123_, N69 );
and g018 ( new_n124_, new_n123_, N65 );
not g019 ( new_n125_, N65 );
and g020 ( new_n126_, new_n125_, N69 );
or g021 ( new_n127_, new_n124_, new_n126_ );
not g022 ( new_n128_, N77 );
and g023 ( new_n129_, new_n128_, N73 );
not g024 ( new_n130_, N73 );
and g025 ( new_n131_, new_n130_, N77 );
or g026 ( new_n132_, new_n129_, new_n131_ );
not g027 ( new_n133_, new_n132_ );
and g028 ( new_n134_, new_n133_, new_n127_ );
not g029 ( new_n135_, new_n134_ );
or g030 ( new_n136_, new_n133_, new_n127_ );
and g031 ( new_n137_, new_n135_, new_n136_ );
not g032 ( new_n138_, new_n137_ );
and g033 ( new_n139_, new_n138_, new_n122_ );
not g034 ( new_n140_, new_n122_ );
and g035 ( new_n141_, new_n140_, new_n137_ );
or g036 ( new_n142_, new_n139_, new_n141_ );
and g037 ( new_n143_, N129, N137 );
not g038 ( new_n144_, new_n143_ );
and g039 ( new_n145_, new_n142_, new_n144_ );
not g040 ( new_n146_, new_n145_ );
or g041 ( new_n147_, new_n142_, new_n144_ );
and g042 ( new_n148_, new_n146_, new_n147_ );
not g043 ( new_n149_, N17 );
and g044 ( new_n150_, new_n149_, N1 );
not g045 ( new_n151_, N1 );
and g046 ( new_n152_, new_n151_, N17 );
or g047 ( new_n153_, new_n150_, new_n152_ );
not g048 ( new_n154_, N49 );
and g049 ( new_n155_, new_n154_, N33 );
not g050 ( new_n156_, N33 );
and g051 ( new_n157_, new_n156_, N49 );
or g052 ( new_n158_, new_n155_, new_n157_ );
not g053 ( new_n159_, new_n158_ );
and g054 ( new_n160_, new_n159_, new_n153_ );
not g055 ( new_n161_, new_n160_ );
or g056 ( new_n162_, new_n159_, new_n153_ );
and g057 ( new_n163_, new_n161_, new_n162_ );
not g058 ( new_n164_, new_n163_ );
and g059 ( new_n165_, new_n148_, new_n164_ );
not g060 ( new_n166_, new_n165_ );
or g061 ( new_n167_, new_n148_, new_n164_ );
and g062 ( new_n168_, new_n166_, new_n167_ );
not g063 ( new_n169_, new_n168_ );
not g064 ( new_n170_, keyIn_0_17 );
not g065 ( new_n171_, N101 );
and g066 ( new_n172_, new_n171_, N97 );
not g067 ( new_n173_, N97 );
and g068 ( new_n174_, new_n173_, N101 );
or g069 ( new_n175_, new_n172_, new_n174_ );
not g070 ( new_n176_, N109 );
and g071 ( new_n177_, new_n176_, N105 );
not g072 ( new_n178_, N105 );
and g073 ( new_n179_, new_n178_, N109 );
or g074 ( new_n180_, new_n177_, new_n179_ );
not g075 ( new_n181_, new_n180_ );
and g076 ( new_n182_, new_n181_, new_n175_ );
not g077 ( new_n183_, new_n182_ );
or g078 ( new_n184_, new_n181_, new_n175_ );
and g079 ( new_n185_, new_n183_, new_n184_ );
and g080 ( new_n186_, new_n138_, new_n185_ );
not g081 ( new_n187_, new_n185_ );
and g082 ( new_n188_, new_n187_, new_n137_ );
or g083 ( new_n189_, new_n186_, new_n188_ );
and g084 ( new_n190_, N131, N137 );
not g085 ( new_n191_, new_n190_ );
and g086 ( new_n192_, new_n189_, new_n191_ );
not g087 ( new_n193_, new_n192_ );
or g088 ( new_n194_, new_n189_, new_n191_ );
and g089 ( new_n195_, new_n193_, new_n194_ );
not g090 ( new_n196_, N25 );
and g091 ( new_n197_, new_n196_, N9 );
not g092 ( new_n198_, N9 );
and g093 ( new_n199_, new_n198_, N25 );
or g094 ( new_n200_, new_n197_, new_n199_ );
not g095 ( new_n201_, N57 );
and g096 ( new_n202_, new_n201_, N41 );
not g097 ( new_n203_, N41 );
and g098 ( new_n204_, new_n203_, N57 );
or g099 ( new_n205_, new_n202_, new_n204_ );
not g100 ( new_n206_, new_n205_ );
and g101 ( new_n207_, new_n206_, new_n200_ );
not g102 ( new_n208_, new_n207_ );
or g103 ( new_n209_, new_n206_, new_n200_ );
and g104 ( new_n210_, new_n208_, new_n209_ );
not g105 ( new_n211_, new_n210_ );
and g106 ( new_n212_, new_n195_, new_n211_ );
not g107 ( new_n213_, new_n212_ );
or g108 ( new_n214_, new_n195_, new_n211_ );
and g109 ( new_n215_, new_n213_, new_n214_ );
not g110 ( new_n216_, N117 );
and g111 ( new_n217_, new_n216_, N113 );
not g112 ( new_n218_, N113 );
and g113 ( new_n219_, new_n218_, N117 );
or g114 ( new_n220_, new_n217_, new_n219_ );
not g115 ( new_n221_, N125 );
and g116 ( new_n222_, new_n221_, N121 );
not g117 ( new_n223_, N121 );
and g118 ( new_n224_, new_n223_, N125 );
or g119 ( new_n225_, new_n222_, new_n224_ );
not g120 ( new_n226_, new_n225_ );
and g121 ( new_n227_, new_n226_, new_n220_ );
not g122 ( new_n228_, new_n227_ );
or g123 ( new_n229_, new_n226_, new_n220_ );
and g124 ( new_n230_, new_n228_, new_n229_ );
and g125 ( new_n231_, new_n187_, new_n230_ );
not g126 ( new_n232_, new_n230_ );
and g127 ( new_n233_, new_n232_, new_n185_ );
or g128 ( new_n234_, new_n231_, new_n233_ );
and g129 ( new_n235_, N130, N137 );
not g130 ( new_n236_, new_n235_ );
and g131 ( new_n237_, new_n234_, new_n236_ );
not g132 ( new_n238_, new_n237_ );
or g133 ( new_n239_, new_n234_, new_n236_ );
and g134 ( new_n240_, new_n238_, new_n239_ );
not g135 ( new_n241_, N21 );
and g136 ( new_n242_, new_n241_, N5 );
not g137 ( new_n243_, N5 );
and g138 ( new_n244_, new_n243_, N21 );
or g139 ( new_n245_, new_n242_, new_n244_ );
not g140 ( new_n246_, N53 );
and g141 ( new_n247_, new_n246_, N37 );
not g142 ( new_n248_, N37 );
and g143 ( new_n249_, new_n248_, N53 );
or g144 ( new_n250_, new_n247_, new_n249_ );
not g145 ( new_n251_, new_n250_ );
and g146 ( new_n252_, new_n251_, new_n245_ );
not g147 ( new_n253_, new_n252_ );
or g148 ( new_n254_, new_n251_, new_n245_ );
and g149 ( new_n255_, new_n253_, new_n254_ );
not g150 ( new_n256_, new_n255_ );
and g151 ( new_n257_, new_n240_, new_n256_ );
not g152 ( new_n258_, new_n257_ );
or g153 ( new_n259_, new_n240_, new_n256_ );
and g154 ( new_n260_, new_n258_, new_n259_ );
not g155 ( new_n261_, new_n260_ );
and g156 ( new_n262_, new_n261_, new_n168_ );
and g157 ( new_n263_, new_n262_, new_n215_ );
and g158 ( new_n264_, new_n169_, new_n260_ );
and g159 ( new_n265_, new_n264_, new_n215_ );
or g160 ( new_n266_, new_n263_, new_n265_ );
and g161 ( new_n267_, new_n140_, new_n230_ );
and g162 ( new_n268_, new_n232_, new_n122_ );
or g163 ( new_n269_, new_n267_, new_n268_ );
and g164 ( new_n270_, N132, N137 );
not g165 ( new_n271_, new_n270_ );
and g166 ( new_n272_, new_n269_, new_n271_ );
not g167 ( new_n273_, new_n272_ );
or g168 ( new_n274_, new_n269_, new_n271_ );
and g169 ( new_n275_, new_n273_, new_n274_ );
not g170 ( new_n276_, N29 );
and g171 ( new_n277_, new_n276_, N13 );
not g172 ( new_n278_, N13 );
and g173 ( new_n279_, new_n278_, N29 );
or g174 ( new_n280_, new_n277_, new_n279_ );
not g175 ( new_n281_, N61 );
and g176 ( new_n282_, new_n281_, N45 );
not g177 ( new_n283_, N45 );
and g178 ( new_n284_, new_n283_, N61 );
or g179 ( new_n285_, new_n282_, new_n284_ );
not g180 ( new_n286_, new_n285_ );
and g181 ( new_n287_, new_n286_, new_n280_ );
not g182 ( new_n288_, new_n287_ );
or g183 ( new_n289_, new_n286_, new_n280_ );
and g184 ( new_n290_, new_n288_, new_n289_ );
not g185 ( new_n291_, new_n290_ );
and g186 ( new_n292_, new_n275_, new_n291_ );
not g187 ( new_n293_, new_n292_ );
or g188 ( new_n294_, new_n275_, new_n291_ );
and g189 ( new_n295_, new_n293_, new_n294_ );
and g190 ( new_n296_, new_n266_, new_n295_ );
not g191 ( new_n297_, new_n295_ );
and g192 ( new_n298_, new_n297_, new_n215_ );
not g193 ( new_n299_, new_n215_ );
and g194 ( new_n300_, new_n299_, new_n295_ );
or g195 ( new_n301_, new_n298_, new_n300_ );
and g196 ( new_n302_, new_n168_, new_n260_ );
and g197 ( new_n303_, new_n301_, new_n302_ );
or g198 ( new_n304_, new_n296_, new_n303_ );
and g199 ( new_n305_, new_n304_, new_n170_ );
not g200 ( new_n306_, new_n305_ );
or g201 ( new_n307_, new_n304_, new_n170_ );
and g202 ( new_n308_, new_n306_, new_n307_ );
not g203 ( new_n309_, new_n308_ );
not g204 ( new_n310_, keyIn_0_14 );
not g205 ( new_n311_, keyIn_0_6 );
not g206 ( new_n312_, keyIn_0_0 );
and g207 ( new_n313_, new_n243_, N1 );
and g208 ( new_n314_, new_n151_, N5 );
or g209 ( new_n315_, new_n313_, new_n314_ );
and g210 ( new_n316_, new_n315_, new_n312_ );
not g211 ( new_n317_, new_n316_ );
or g212 ( new_n318_, new_n315_, new_n312_ );
and g213 ( new_n319_, new_n317_, new_n318_ );
and g214 ( new_n320_, new_n278_, N9 );
and g215 ( new_n321_, new_n198_, N13 );
or g216 ( new_n322_, new_n320_, new_n321_ );
and g217 ( new_n323_, new_n322_, keyIn_0_1 );
not g218 ( new_n324_, new_n323_ );
or g219 ( new_n325_, new_n322_, keyIn_0_1 );
and g220 ( new_n326_, new_n324_, new_n325_ );
or g221 ( new_n327_, new_n319_, new_n326_ );
not g222 ( new_n328_, new_n327_ );
and g223 ( new_n329_, new_n319_, new_n326_ );
or g224 ( new_n330_, new_n328_, new_n329_ );
and g225 ( new_n331_, new_n330_, new_n311_ );
not g226 ( new_n332_, new_n329_ );
and g227 ( new_n333_, new_n332_, new_n327_ );
and g228 ( new_n334_, new_n333_, keyIn_0_6 );
or g229 ( new_n335_, new_n331_, new_n334_ );
not g230 ( new_n336_, keyIn_0_7 );
or g231 ( new_n337_, new_n156_, N37 );
or g232 ( new_n338_, new_n248_, N33 );
and g233 ( new_n339_, new_n337_, new_n338_ );
or g234 ( new_n340_, new_n339_, keyIn_0_2 );
not g235 ( new_n341_, keyIn_0_2 );
and g236 ( new_n342_, new_n248_, N33 );
and g237 ( new_n343_, new_n156_, N37 );
or g238 ( new_n344_, new_n342_, new_n343_ );
or g239 ( new_n345_, new_n344_, new_n341_ );
and g240 ( new_n346_, new_n345_, new_n340_ );
or g241 ( new_n347_, new_n203_, N45 );
or g242 ( new_n348_, new_n283_, N41 );
and g243 ( new_n349_, new_n347_, new_n348_ );
or g244 ( new_n350_, new_n349_, keyIn_0_3 );
not g245 ( new_n351_, keyIn_0_3 );
and g246 ( new_n352_, new_n283_, N41 );
and g247 ( new_n353_, new_n203_, N45 );
or g248 ( new_n354_, new_n352_, new_n353_ );
or g249 ( new_n355_, new_n354_, new_n351_ );
and g250 ( new_n356_, new_n355_, new_n350_ );
or g251 ( new_n357_, new_n346_, new_n356_ );
and g252 ( new_n358_, new_n344_, new_n341_ );
and g253 ( new_n359_, new_n339_, keyIn_0_2 );
or g254 ( new_n360_, new_n358_, new_n359_ );
and g255 ( new_n361_, new_n354_, new_n351_ );
and g256 ( new_n362_, new_n349_, keyIn_0_3 );
or g257 ( new_n363_, new_n361_, new_n362_ );
or g258 ( new_n364_, new_n360_, new_n363_ );
and g259 ( new_n365_, new_n364_, new_n357_ );
or g260 ( new_n366_, new_n365_, new_n336_ );
and g261 ( new_n367_, new_n360_, new_n363_ );
and g262 ( new_n368_, new_n346_, new_n356_ );
or g263 ( new_n369_, new_n367_, new_n368_ );
or g264 ( new_n370_, new_n369_, keyIn_0_7 );
and g265 ( new_n371_, new_n366_, new_n370_ );
or g266 ( new_n372_, new_n335_, new_n371_ );
or g267 ( new_n373_, new_n333_, keyIn_0_6 );
or g268 ( new_n374_, new_n330_, new_n311_ );
and g269 ( new_n375_, new_n374_, new_n373_ );
and g270 ( new_n376_, new_n369_, keyIn_0_7 );
and g271 ( new_n377_, new_n365_, new_n336_ );
or g272 ( new_n378_, new_n376_, new_n377_ );
or g273 ( new_n379_, new_n375_, new_n378_ );
and g274 ( new_n380_, new_n372_, new_n379_ );
or g275 ( new_n381_, new_n380_, keyIn_0_10 );
not g276 ( new_n382_, keyIn_0_10 );
and g277 ( new_n383_, new_n375_, new_n378_ );
and g278 ( new_n384_, new_n335_, new_n371_ );
or g279 ( new_n385_, new_n383_, new_n384_ );
or g280 ( new_n386_, new_n385_, new_n382_ );
and g281 ( new_n387_, new_n386_, new_n381_ );
and g282 ( new_n388_, N135, N137 );
not g283 ( new_n389_, new_n388_ );
or g284 ( new_n390_, new_n387_, new_n389_ );
and g285 ( new_n391_, new_n385_, new_n382_ );
and g286 ( new_n392_, new_n380_, keyIn_0_10 );
or g287 ( new_n393_, new_n391_, new_n392_ );
or g288 ( new_n394_, new_n393_, new_n388_ );
and g289 ( new_n395_, new_n394_, new_n390_ );
or g290 ( new_n396_, new_n395_, keyIn_0_12 );
not g291 ( new_n397_, keyIn_0_12 );
and g292 ( new_n398_, new_n393_, new_n388_ );
and g293 ( new_n399_, new_n387_, new_n389_ );
or g294 ( new_n400_, new_n398_, new_n399_ );
or g295 ( new_n401_, new_n400_, new_n397_ );
and g296 ( new_n402_, new_n401_, new_n396_ );
and g297 ( new_n403_, new_n115_, N73 );
and g298 ( new_n404_, new_n130_, N89 );
or g299 ( new_n405_, new_n403_, new_n404_ );
and g300 ( new_n406_, new_n223_, N105 );
and g301 ( new_n407_, new_n178_, N121 );
or g302 ( new_n408_, new_n406_, new_n407_ );
not g303 ( new_n409_, new_n408_ );
and g304 ( new_n410_, new_n409_, new_n405_ );
not g305 ( new_n411_, new_n410_ );
or g306 ( new_n412_, new_n409_, new_n405_ );
and g307 ( new_n413_, new_n411_, new_n412_ );
not g308 ( new_n414_, new_n413_ );
or g309 ( new_n415_, new_n402_, new_n414_ );
and g310 ( new_n416_, new_n400_, new_n397_ );
and g311 ( new_n417_, new_n395_, keyIn_0_12 );
or g312 ( new_n418_, new_n416_, new_n417_ );
or g313 ( new_n419_, new_n418_, new_n413_ );
and g314 ( new_n420_, new_n419_, new_n415_ );
or g315 ( new_n421_, new_n420_, new_n310_ );
and g316 ( new_n422_, new_n418_, new_n413_ );
and g317 ( new_n423_, new_n402_, new_n414_ );
or g318 ( new_n424_, new_n422_, new_n423_ );
or g319 ( new_n425_, new_n424_, keyIn_0_14 );
and g320 ( new_n426_, new_n425_, new_n421_ );
and g321 ( new_n427_, new_n241_, N17 );
and g322 ( new_n428_, new_n149_, N21 );
or g323 ( new_n429_, new_n427_, new_n428_ );
and g324 ( new_n430_, new_n276_, N25 );
and g325 ( new_n431_, new_n196_, N29 );
or g326 ( new_n432_, new_n430_, new_n431_ );
not g327 ( new_n433_, new_n432_ );
and g328 ( new_n434_, new_n433_, new_n429_ );
not g329 ( new_n435_, new_n434_ );
or g330 ( new_n436_, new_n433_, new_n429_ );
and g331 ( new_n437_, new_n435_, new_n436_ );
not g332 ( new_n438_, new_n437_ );
and g333 ( new_n439_, new_n246_, N49 );
and g334 ( new_n440_, new_n154_, N53 );
or g335 ( new_n441_, new_n439_, new_n440_ );
and g336 ( new_n442_, new_n441_, keyIn_0_4 );
not g337 ( new_n443_, keyIn_0_4 );
or g338 ( new_n444_, new_n154_, N53 );
or g339 ( new_n445_, new_n246_, N49 );
and g340 ( new_n446_, new_n444_, new_n445_ );
and g341 ( new_n447_, new_n446_, new_n443_ );
or g342 ( new_n448_, new_n442_, new_n447_ );
not g343 ( new_n449_, keyIn_0_5 );
and g344 ( new_n450_, new_n281_, N57 );
and g345 ( new_n451_, new_n201_, N61 );
or g346 ( new_n452_, new_n450_, new_n451_ );
and g347 ( new_n453_, new_n452_, new_n449_ );
or g348 ( new_n454_, new_n201_, N61 );
or g349 ( new_n455_, new_n281_, N57 );
and g350 ( new_n456_, new_n454_, new_n455_ );
and g351 ( new_n457_, new_n456_, keyIn_0_5 );
or g352 ( new_n458_, new_n453_, new_n457_ );
and g353 ( new_n459_, new_n448_, new_n458_ );
or g354 ( new_n460_, new_n446_, new_n443_ );
or g355 ( new_n461_, new_n441_, keyIn_0_4 );
and g356 ( new_n462_, new_n461_, new_n460_ );
or g357 ( new_n463_, new_n456_, keyIn_0_5 );
or g358 ( new_n464_, new_n452_, new_n449_ );
and g359 ( new_n465_, new_n464_, new_n463_ );
and g360 ( new_n466_, new_n462_, new_n465_ );
or g361 ( new_n467_, new_n459_, new_n466_ );
and g362 ( new_n468_, new_n467_, keyIn_0_8 );
not g363 ( new_n469_, keyIn_0_8 );
or g364 ( new_n470_, new_n462_, new_n465_ );
or g365 ( new_n471_, new_n448_, new_n458_ );
and g366 ( new_n472_, new_n471_, new_n470_ );
and g367 ( new_n473_, new_n472_, new_n469_ );
or g368 ( new_n474_, new_n468_, new_n473_ );
and g369 ( new_n475_, new_n474_, new_n438_ );
or g370 ( new_n476_, new_n472_, new_n469_ );
or g371 ( new_n477_, new_n467_, keyIn_0_8 );
and g372 ( new_n478_, new_n476_, new_n477_ );
and g373 ( new_n479_, new_n478_, new_n437_ );
or g374 ( new_n480_, new_n475_, new_n479_ );
and g375 ( new_n481_, N136, N137 );
not g376 ( new_n482_, new_n481_ );
and g377 ( new_n483_, new_n480_, new_n482_ );
not g378 ( new_n484_, new_n483_ );
or g379 ( new_n485_, new_n480_, new_n482_ );
and g380 ( new_n486_, new_n484_, new_n485_ );
and g381 ( new_n487_, new_n113_, N77 );
and g382 ( new_n488_, new_n128_, N93 );
or g383 ( new_n489_, new_n487_, new_n488_ );
and g384 ( new_n490_, new_n221_, N109 );
and g385 ( new_n491_, new_n176_, N125 );
or g386 ( new_n492_, new_n490_, new_n491_ );
not g387 ( new_n493_, new_n492_ );
and g388 ( new_n494_, new_n493_, new_n489_ );
not g389 ( new_n495_, new_n494_ );
or g390 ( new_n496_, new_n493_, new_n489_ );
and g391 ( new_n497_, new_n495_, new_n496_ );
not g392 ( new_n498_, new_n497_ );
and g393 ( new_n499_, new_n486_, new_n498_ );
not g394 ( new_n500_, new_n499_ );
or g395 ( new_n501_, new_n486_, new_n498_ );
and g396 ( new_n502_, new_n500_, new_n501_ );
not g397 ( new_n503_, new_n502_ );
or g398 ( new_n504_, new_n426_, new_n503_ );
or g399 ( new_n505_, new_n504_, new_n309_ );
and g400 ( new_n506_, new_n335_, new_n438_ );
and g401 ( new_n507_, new_n375_, new_n437_ );
or g402 ( new_n508_, new_n506_, new_n507_ );
and g403 ( new_n509_, N133, N137 );
not g404 ( new_n510_, new_n509_ );
and g405 ( new_n511_, new_n508_, new_n510_ );
not g406 ( new_n512_, new_n511_ );
or g407 ( new_n513_, new_n508_, new_n510_ );
and g408 ( new_n514_, new_n512_, new_n513_ );
and g409 ( new_n515_, new_n110_, N65 );
and g410 ( new_n516_, new_n125_, N81 );
or g411 ( new_n517_, new_n515_, new_n516_ );
and g412 ( new_n518_, new_n218_, N97 );
and g413 ( new_n519_, new_n173_, N113 );
or g414 ( new_n520_, new_n518_, new_n519_ );
not g415 ( new_n521_, new_n520_ );
and g416 ( new_n522_, new_n521_, new_n517_ );
not g417 ( new_n523_, new_n522_ );
or g418 ( new_n524_, new_n521_, new_n517_ );
and g419 ( new_n525_, new_n523_, new_n524_ );
not g420 ( new_n526_, new_n525_ );
and g421 ( new_n527_, new_n514_, new_n526_ );
not g422 ( new_n528_, new_n527_ );
or g423 ( new_n529_, new_n514_, new_n526_ );
and g424 ( new_n530_, new_n528_, new_n529_ );
or g425 ( new_n531_, new_n378_, new_n478_ );
or g426 ( new_n532_, new_n474_, new_n371_ );
and g427 ( new_n533_, new_n531_, new_n532_ );
or g428 ( new_n534_, new_n533_, keyIn_0_9 );
not g429 ( new_n535_, keyIn_0_9 );
and g430 ( new_n536_, new_n474_, new_n371_ );
and g431 ( new_n537_, new_n378_, new_n478_ );
or g432 ( new_n538_, new_n536_, new_n537_ );
or g433 ( new_n539_, new_n538_, new_n535_ );
and g434 ( new_n540_, new_n539_, new_n534_ );
and g435 ( new_n541_, N134, N137 );
or g436 ( new_n542_, new_n540_, new_n541_ );
and g437 ( new_n543_, new_n538_, new_n535_ );
and g438 ( new_n544_, new_n533_, keyIn_0_9 );
or g439 ( new_n545_, new_n543_, new_n544_ );
not g440 ( new_n546_, new_n541_ );
or g441 ( new_n547_, new_n545_, new_n546_ );
and g442 ( new_n548_, new_n547_, new_n542_ );
or g443 ( new_n549_, new_n548_, keyIn_0_11 );
not g444 ( new_n550_, keyIn_0_11 );
and g445 ( new_n551_, new_n545_, new_n546_ );
and g446 ( new_n552_, new_n540_, new_n541_ );
or g447 ( new_n553_, new_n551_, new_n552_ );
or g448 ( new_n554_, new_n553_, new_n550_ );
and g449 ( new_n555_, new_n554_, new_n549_ );
and g450 ( new_n556_, new_n108_, N69 );
and g451 ( new_n557_, new_n123_, N85 );
or g452 ( new_n558_, new_n556_, new_n557_ );
and g453 ( new_n559_, new_n216_, N101 );
and g454 ( new_n560_, new_n171_, N117 );
or g455 ( new_n561_, new_n559_, new_n560_ );
not g456 ( new_n562_, new_n561_ );
and g457 ( new_n563_, new_n562_, new_n558_ );
not g458 ( new_n564_, new_n563_ );
or g459 ( new_n565_, new_n562_, new_n558_ );
and g460 ( new_n566_, new_n564_, new_n565_ );
not g461 ( new_n567_, new_n566_ );
or g462 ( new_n568_, new_n555_, new_n567_ );
and g463 ( new_n569_, new_n553_, new_n550_ );
and g464 ( new_n570_, new_n548_, keyIn_0_11 );
or g465 ( new_n571_, new_n569_, new_n570_ );
or g466 ( new_n572_, new_n571_, new_n566_ );
and g467 ( new_n573_, new_n572_, new_n568_ );
or g468 ( new_n574_, new_n573_, keyIn_0_13 );
not g469 ( new_n575_, keyIn_0_13 );
and g470 ( new_n576_, new_n571_, new_n566_ );
and g471 ( new_n577_, new_n555_, new_n567_ );
or g472 ( new_n578_, new_n576_, new_n577_ );
or g473 ( new_n579_, new_n578_, new_n575_ );
and g474 ( new_n580_, new_n579_, new_n574_ );
or g475 ( new_n581_, new_n580_, keyIn_0_15 );
not g476 ( new_n582_, keyIn_0_15 );
and g477 ( new_n583_, new_n578_, new_n575_ );
and g478 ( new_n584_, new_n573_, keyIn_0_13 );
or g479 ( new_n585_, new_n583_, new_n584_ );
or g480 ( new_n586_, new_n585_, new_n582_ );
and g481 ( new_n587_, new_n586_, new_n581_ );
or g482 ( new_n588_, new_n587_, new_n530_ );
or g483 ( new_n589_, new_n588_, new_n505_ );
and g484 ( new_n590_, new_n589_, keyIn_0_18 );
not g485 ( new_n591_, keyIn_0_18 );
not g486 ( new_n592_, new_n426_ );
and g487 ( new_n593_, new_n592_, new_n502_ );
and g488 ( new_n594_, new_n593_, new_n308_ );
not g489 ( new_n595_, new_n530_ );
and g490 ( new_n596_, new_n585_, new_n582_ );
and g491 ( new_n597_, new_n580_, keyIn_0_15 );
or g492 ( new_n598_, new_n596_, new_n597_ );
and g493 ( new_n599_, new_n598_, new_n595_ );
and g494 ( new_n600_, new_n594_, new_n599_ );
and g495 ( new_n601_, new_n600_, new_n591_ );
or g496 ( new_n602_, new_n590_, new_n601_ );
and g497 ( new_n603_, new_n602_, new_n169_ );
or g498 ( new_n604_, new_n603_, new_n107_ );
or g499 ( new_n605_, new_n600_, new_n591_ );
or g500 ( new_n606_, new_n589_, keyIn_0_18 );
and g501 ( new_n607_, new_n606_, new_n605_ );
or g502 ( new_n608_, new_n607_, new_n168_ );
or g503 ( new_n609_, new_n608_, keyIn_0_20 );
and g504 ( new_n610_, new_n609_, new_n604_ );
or g505 ( new_n611_, new_n610_, N1 );
and g506 ( new_n612_, new_n608_, keyIn_0_20 );
and g507 ( new_n613_, new_n603_, new_n107_ );
or g508 ( new_n614_, new_n612_, new_n613_ );
or g509 ( new_n615_, new_n614_, new_n151_ );
and g510 ( new_n616_, new_n615_, new_n611_ );
or g511 ( new_n617_, new_n616_, new_n106_ );
and g512 ( new_n618_, new_n614_, new_n151_ );
and g513 ( new_n619_, new_n610_, N1 );
or g514 ( new_n620_, new_n618_, new_n619_ );
or g515 ( new_n621_, new_n620_, keyIn_0_26 );
and g516 ( N724, new_n621_, new_n617_ );
not g517 ( new_n623_, keyIn_0_27 );
not g518 ( new_n624_, keyIn_0_21 );
and g519 ( new_n625_, new_n602_, new_n261_ );
or g520 ( new_n626_, new_n625_, new_n624_ );
or g521 ( new_n627_, new_n607_, new_n260_ );
or g522 ( new_n628_, new_n627_, keyIn_0_21 );
and g523 ( new_n629_, new_n628_, new_n626_ );
or g524 ( new_n630_, new_n629_, new_n243_ );
and g525 ( new_n631_, new_n627_, keyIn_0_21 );
and g526 ( new_n632_, new_n625_, new_n624_ );
or g527 ( new_n633_, new_n631_, new_n632_ );
or g528 ( new_n634_, new_n633_, N5 );
and g529 ( new_n635_, new_n634_, new_n630_ );
or g530 ( new_n636_, new_n635_, new_n623_ );
and g531 ( new_n637_, new_n633_, N5 );
and g532 ( new_n638_, new_n629_, new_n243_ );
or g533 ( new_n639_, new_n637_, new_n638_ );
or g534 ( new_n640_, new_n639_, keyIn_0_27 );
and g535 ( N725, new_n640_, new_n636_ );
not g536 ( new_n642_, keyIn_0_22 );
and g537 ( new_n643_, new_n602_, new_n299_ );
or g538 ( new_n644_, new_n643_, new_n642_ );
or g539 ( new_n645_, new_n607_, new_n215_ );
or g540 ( new_n646_, new_n645_, keyIn_0_22 );
and g541 ( new_n647_, new_n646_, new_n644_ );
or g542 ( new_n648_, new_n647_, N9 );
and g543 ( new_n649_, new_n645_, keyIn_0_22 );
and g544 ( new_n650_, new_n643_, new_n642_ );
or g545 ( new_n651_, new_n649_, new_n650_ );
or g546 ( new_n652_, new_n651_, new_n198_ );
and g547 ( new_n653_, new_n652_, new_n648_ );
or g548 ( new_n654_, new_n653_, keyIn_0_28 );
not g549 ( new_n655_, keyIn_0_28 );
and g550 ( new_n656_, new_n651_, new_n198_ );
and g551 ( new_n657_, new_n647_, N9 );
or g552 ( new_n658_, new_n656_, new_n657_ );
or g553 ( new_n659_, new_n658_, new_n655_ );
and g554 ( N726, new_n659_, new_n654_ );
not g555 ( new_n661_, keyIn_0_29 );
not g556 ( new_n662_, keyIn_0_23 );
and g557 ( new_n663_, new_n602_, new_n297_ );
or g558 ( new_n664_, new_n663_, new_n662_ );
or g559 ( new_n665_, new_n607_, new_n295_ );
or g560 ( new_n666_, new_n665_, keyIn_0_23 );
and g561 ( new_n667_, new_n666_, new_n664_ );
or g562 ( new_n668_, new_n667_, N13 );
and g563 ( new_n669_, new_n665_, keyIn_0_23 );
and g564 ( new_n670_, new_n663_, new_n662_ );
or g565 ( new_n671_, new_n669_, new_n670_ );
or g566 ( new_n672_, new_n671_, new_n278_ );
and g567 ( new_n673_, new_n672_, new_n668_ );
or g568 ( new_n674_, new_n673_, new_n661_ );
and g569 ( new_n675_, new_n671_, new_n278_ );
and g570 ( new_n676_, new_n667_, N13 );
or g571 ( new_n677_, new_n675_, new_n676_ );
or g572 ( new_n678_, new_n677_, keyIn_0_29 );
and g573 ( N727, new_n678_, new_n674_ );
not g574 ( new_n680_, keyIn_0_19 );
and g575 ( new_n681_, new_n585_, new_n595_ );
and g576 ( new_n682_, new_n308_, new_n503_ );
and g577 ( new_n683_, new_n426_, new_n682_ );
and g578 ( new_n684_, new_n683_, new_n681_ );
or g579 ( new_n685_, new_n684_, new_n680_ );
and g580 ( new_n686_, new_n684_, new_n680_ );
not g581 ( new_n687_, new_n686_ );
and g582 ( new_n688_, new_n687_, new_n685_ );
and g583 ( new_n689_, new_n688_, new_n169_ );
not g584 ( new_n690_, new_n689_ );
and g585 ( new_n691_, new_n690_, N17 );
and g586 ( new_n692_, new_n689_, new_n149_ );
or g587 ( N728, new_n691_, new_n692_ );
not g588 ( new_n694_, keyIn_0_30 );
and g589 ( new_n695_, new_n688_, new_n261_ );
or g590 ( new_n696_, new_n695_, keyIn_0_24 );
and g591 ( new_n697_, new_n695_, keyIn_0_24 );
not g592 ( new_n698_, new_n697_ );
and g593 ( new_n699_, new_n698_, new_n696_ );
not g594 ( new_n700_, new_n699_ );
and g595 ( new_n701_, new_n700_, new_n241_ );
and g596 ( new_n702_, new_n699_, N21 );
or g597 ( new_n703_, new_n701_, new_n702_ );
not g598 ( new_n704_, new_n703_ );
or g599 ( new_n705_, new_n704_, new_n694_ );
or g600 ( new_n706_, new_n703_, keyIn_0_30 );
and g601 ( N729, new_n705_, new_n706_ );
and g602 ( new_n708_, new_n688_, new_n299_ );
not g603 ( new_n709_, new_n708_ );
and g604 ( new_n710_, new_n709_, N25 );
and g605 ( new_n711_, new_n708_, new_n196_ );
or g606 ( N730, new_n710_, new_n711_ );
not g607 ( new_n713_, keyIn_0_25 );
and g608 ( new_n714_, new_n688_, new_n297_ );
not g609 ( new_n715_, new_n714_ );
and g610 ( new_n716_, new_n715_, new_n713_ );
and g611 ( new_n717_, new_n714_, keyIn_0_25 );
or g612 ( new_n718_, new_n716_, new_n717_ );
and g613 ( new_n719_, new_n718_, N29 );
not g614 ( new_n720_, new_n719_ );
or g615 ( new_n721_, new_n718_, N29 );
and g616 ( new_n722_, new_n720_, new_n721_ );
not g617 ( new_n723_, new_n722_ );
and g618 ( new_n724_, new_n723_, keyIn_0_31 );
not g619 ( new_n725_, keyIn_0_31 );
and g620 ( new_n726_, new_n722_, new_n725_ );
or g621 ( N731, new_n724_, new_n726_ );
and g622 ( new_n728_, new_n580_, new_n530_ );
and g623 ( new_n729_, new_n594_, new_n728_ );
and g624 ( new_n730_, new_n729_, new_n169_ );
not g625 ( new_n731_, new_n730_ );
and g626 ( new_n732_, new_n731_, N33 );
and g627 ( new_n733_, new_n730_, new_n156_ );
or g628 ( N732, new_n732_, new_n733_ );
and g629 ( new_n735_, new_n729_, new_n261_ );
not g630 ( new_n736_, new_n735_ );
and g631 ( new_n737_, new_n736_, N37 );
and g632 ( new_n738_, new_n735_, new_n248_ );
or g633 ( N733, new_n737_, new_n738_ );
and g634 ( new_n740_, new_n729_, new_n299_ );
not g635 ( new_n741_, new_n740_ );
and g636 ( new_n742_, new_n741_, N41 );
and g637 ( new_n743_, new_n740_, new_n203_ );
or g638 ( N734, new_n742_, new_n743_ );
and g639 ( new_n745_, new_n729_, new_n297_ );
not g640 ( new_n746_, new_n745_ );
and g641 ( new_n747_, new_n746_, N45 );
and g642 ( new_n748_, new_n745_, new_n283_ );
or g643 ( N735, new_n747_, new_n748_ );
and g644 ( new_n750_, new_n728_, new_n426_ );
and g645 ( new_n751_, new_n750_, new_n682_ );
and g646 ( new_n752_, new_n751_, new_n169_ );
not g647 ( new_n753_, new_n752_ );
and g648 ( new_n754_, new_n753_, N49 );
and g649 ( new_n755_, new_n752_, new_n154_ );
or g650 ( N736, new_n754_, new_n755_ );
and g651 ( new_n757_, new_n751_, new_n261_ );
not g652 ( new_n758_, new_n757_ );
and g653 ( new_n759_, new_n758_, N53 );
and g654 ( new_n760_, new_n757_, new_n246_ );
or g655 ( N737, new_n759_, new_n760_ );
and g656 ( new_n762_, new_n751_, new_n299_ );
not g657 ( new_n763_, new_n762_ );
and g658 ( new_n764_, new_n763_, N57 );
and g659 ( new_n765_, new_n762_, new_n201_ );
or g660 ( N738, new_n764_, new_n765_ );
and g661 ( new_n767_, new_n751_, new_n297_ );
not g662 ( new_n768_, new_n767_ );
and g663 ( new_n769_, new_n768_, N61 );
and g664 ( new_n770_, new_n767_, new_n281_ );
or g665 ( N739, new_n769_, new_n770_ );
not g666 ( new_n772_, keyIn_0_16 );
and g667 ( new_n773_, new_n426_, new_n772_ );
not g668 ( new_n774_, new_n773_ );
and g669 ( new_n775_, new_n592_, keyIn_0_16 );
not g670 ( new_n776_, new_n775_ );
and g671 ( new_n777_, new_n776_, new_n681_ );
and g672 ( new_n778_, new_n777_, new_n774_ );
or g673 ( new_n779_, new_n778_, new_n750_ );
and g674 ( new_n780_, new_n779_, new_n502_ );
and g675 ( new_n781_, new_n426_, new_n503_ );
or g676 ( new_n782_, new_n593_, new_n781_ );
and g677 ( new_n783_, new_n585_, new_n530_ );
and g678 ( new_n784_, new_n782_, new_n783_ );
or g679 ( new_n785_, new_n780_, new_n784_ );
and g680 ( new_n786_, new_n264_, new_n300_ );
and g681 ( new_n787_, new_n785_, new_n786_ );
and g682 ( new_n788_, new_n787_, new_n595_ );
not g683 ( new_n789_, new_n788_ );
and g684 ( new_n790_, new_n789_, N65 );
and g685 ( new_n791_, new_n788_, new_n125_ );
or g686 ( N740, new_n790_, new_n791_ );
and g687 ( new_n793_, new_n787_, new_n580_ );
not g688 ( new_n794_, new_n793_ );
and g689 ( new_n795_, new_n794_, N69 );
and g690 ( new_n796_, new_n793_, new_n123_ );
or g691 ( N741, new_n795_, new_n796_ );
and g692 ( new_n798_, new_n787_, new_n592_ );
not g693 ( new_n799_, new_n798_ );
and g694 ( new_n800_, new_n799_, N73 );
and g695 ( new_n801_, new_n798_, new_n130_ );
or g696 ( N742, new_n800_, new_n801_ );
and g697 ( new_n803_, new_n787_, new_n503_ );
not g698 ( new_n804_, new_n803_ );
and g699 ( new_n805_, new_n804_, N77 );
and g700 ( new_n806_, new_n803_, new_n128_ );
or g701 ( N743, new_n805_, new_n806_ );
and g702 ( new_n808_, new_n265_, new_n297_ );
and g703 ( new_n809_, new_n785_, new_n808_ );
and g704 ( new_n810_, new_n809_, new_n595_ );
not g705 ( new_n811_, new_n810_ );
and g706 ( new_n812_, new_n811_, N81 );
and g707 ( new_n813_, new_n810_, new_n110_ );
or g708 ( N744, new_n812_, new_n813_ );
and g709 ( new_n815_, new_n809_, new_n580_ );
not g710 ( new_n816_, new_n815_ );
and g711 ( new_n817_, new_n816_, N85 );
and g712 ( new_n818_, new_n815_, new_n108_ );
or g713 ( N745, new_n817_, new_n818_ );
and g714 ( new_n820_, new_n809_, new_n592_ );
not g715 ( new_n821_, new_n820_ );
and g716 ( new_n822_, new_n821_, N89 );
and g717 ( new_n823_, new_n820_, new_n115_ );
or g718 ( N746, new_n822_, new_n823_ );
and g719 ( new_n825_, new_n809_, new_n503_ );
not g720 ( new_n826_, new_n825_ );
and g721 ( new_n827_, new_n826_, N93 );
and g722 ( new_n828_, new_n825_, new_n113_ );
or g723 ( N747, new_n827_, new_n828_ );
and g724 ( new_n830_, new_n262_, new_n300_ );
and g725 ( new_n831_, new_n785_, new_n830_ );
and g726 ( new_n832_, new_n831_, new_n595_ );
not g727 ( new_n833_, new_n832_ );
and g728 ( new_n834_, new_n833_, N97 );
and g729 ( new_n835_, new_n832_, new_n173_ );
or g730 ( N748, new_n834_, new_n835_ );
and g731 ( new_n837_, new_n831_, new_n580_ );
not g732 ( new_n838_, new_n837_ );
and g733 ( new_n839_, new_n838_, N101 );
and g734 ( new_n840_, new_n837_, new_n171_ );
or g735 ( N749, new_n839_, new_n840_ );
and g736 ( new_n842_, new_n831_, new_n592_ );
not g737 ( new_n843_, new_n842_ );
and g738 ( new_n844_, new_n843_, N105 );
and g739 ( new_n845_, new_n842_, new_n178_ );
or g740 ( N750, new_n844_, new_n845_ );
and g741 ( new_n847_, new_n831_, new_n503_ );
not g742 ( new_n848_, new_n847_ );
and g743 ( new_n849_, new_n848_, N109 );
and g744 ( new_n850_, new_n847_, new_n176_ );
or g745 ( N751, new_n849_, new_n850_ );
and g746 ( new_n852_, new_n263_, new_n297_ );
and g747 ( new_n853_, new_n785_, new_n852_ );
and g748 ( new_n854_, new_n853_, new_n595_ );
not g749 ( new_n855_, new_n854_ );
and g750 ( new_n856_, new_n855_, N113 );
and g751 ( new_n857_, new_n854_, new_n218_ );
or g752 ( N752, new_n856_, new_n857_ );
and g753 ( new_n859_, new_n853_, new_n580_ );
not g754 ( new_n860_, new_n859_ );
and g755 ( new_n861_, new_n860_, N117 );
and g756 ( new_n862_, new_n859_, new_n216_ );
or g757 ( N753, new_n861_, new_n862_ );
and g758 ( new_n864_, new_n853_, new_n592_ );
not g759 ( new_n865_, new_n864_ );
and g760 ( new_n866_, new_n865_, N121 );
and g761 ( new_n867_, new_n864_, new_n223_ );
or g762 ( N754, new_n866_, new_n867_ );
and g763 ( new_n869_, new_n853_, new_n503_ );
not g764 ( new_n870_, new_n869_ );
and g765 ( new_n871_, new_n870_, N125 );
and g766 ( new_n872_, new_n869_, new_n221_ );
or g767 ( N755, new_n871_, new_n872_ );
endmodule