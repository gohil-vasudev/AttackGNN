module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434;

  OR2_X1 U228 ( .A1(n221), .A2(n222), .ZN(Result_6_) );
  AND2_X1 U229 ( .A1(n223), .A2(n224), .ZN(n222) );
  INV_X1 U230 ( .A(n225), .ZN(n221) );
  OR2_X1 U231 ( .A1(n224), .A2(n223), .ZN(n225) );
  AND2_X1 U232 ( .A1(n226), .A2(n227), .ZN(n223) );
  OR2_X1 U233 ( .A1(n228), .A2(n229), .ZN(n224) );
  OR2_X1 U234 ( .A1(n230), .A2(n231), .ZN(Result_5_) );
  AND2_X1 U235 ( .A1(n232), .A2(n233), .ZN(n231) );
  INV_X1 U236 ( .A(n234), .ZN(n230) );
  OR2_X1 U237 ( .A1(n233), .A2(n232), .ZN(n234) );
  OR2_X1 U238 ( .A1(n235), .A2(n236), .ZN(n232) );
  INV_X1 U239 ( .A(n237), .ZN(n236) );
  OR2_X1 U240 ( .A1(n238), .A2(n239), .ZN(n237) );
  AND2_X1 U241 ( .A1(n239), .A2(n238), .ZN(n235) );
  OR2_X1 U242 ( .A1(n240), .A2(n241), .ZN(Result_4_) );
  AND2_X1 U243 ( .A1(n242), .A2(n243), .ZN(n241) );
  INV_X1 U244 ( .A(n244), .ZN(n240) );
  OR2_X1 U245 ( .A1(n243), .A2(n242), .ZN(n244) );
  OR2_X1 U246 ( .A1(n245), .A2(n246), .ZN(n242) );
  AND2_X1 U247 ( .A1(n247), .A2(n248), .ZN(n246) );
  INV_X1 U248 ( .A(n249), .ZN(n245) );
  OR2_X1 U249 ( .A1(n248), .A2(n247), .ZN(n249) );
  INV_X1 U250 ( .A(n250), .ZN(n247) );
  OR2_X1 U251 ( .A1(n251), .A2(n252), .ZN(Result_3_) );
  AND2_X1 U252 ( .A1(n253), .A2(n254), .ZN(n252) );
  AND2_X1 U253 ( .A1(n255), .A2(n256), .ZN(n251) );
  INV_X1 U254 ( .A(n253), .ZN(n255) );
  AND2_X1 U255 ( .A1(n257), .A2(n258), .ZN(Result_2_) );
  OR2_X1 U256 ( .A1(n259), .A2(n260), .ZN(n257) );
  AND2_X1 U257 ( .A1(n256), .A2(n253), .ZN(n259) );
  OR2_X1 U258 ( .A1(n261), .A2(n262), .ZN(Result_1_) );
  AND2_X1 U259 ( .A1(n263), .A2(n258), .ZN(n262) );
  INV_X1 U260 ( .A(n264), .ZN(n258) );
  AND2_X1 U261 ( .A1(n264), .A2(n265), .ZN(n261) );
  OR3_X1 U262 ( .A1(n266), .A2(n267), .A3(n268), .ZN(Result_0_) );
  AND2_X1 U263 ( .A1(n269), .A2(n270), .ZN(n268) );
  AND2_X1 U264 ( .A1(n263), .A2(n264), .ZN(n267) );
  AND3_X1 U265 ( .A1(n253), .A2(n256), .A3(n260), .ZN(n264) );
  AND2_X1 U266 ( .A1(n271), .A2(n272), .ZN(n260) );
  OR2_X1 U267 ( .A1(n273), .A2(n274), .ZN(n272) );
  INV_X1 U268 ( .A(n254), .ZN(n256) );
  OR2_X1 U269 ( .A1(n275), .A2(n276), .ZN(n254) );
  AND2_X1 U270 ( .A1(n250), .A2(n248), .ZN(n276) );
  AND2_X1 U271 ( .A1(n243), .A2(n277), .ZN(n275) );
  OR2_X1 U272 ( .A1(n248), .A2(n250), .ZN(n277) );
  OR2_X1 U273 ( .A1(n278), .A2(n279), .ZN(n250) );
  OR2_X1 U274 ( .A1(n280), .A2(n281), .ZN(n248) );
  AND2_X1 U275 ( .A1(n238), .A2(n282), .ZN(n281) );
  AND2_X1 U276 ( .A1(n233), .A2(n283), .ZN(n280) );
  OR2_X1 U277 ( .A1(n282), .A2(n238), .ZN(n283) );
  OR2_X1 U278 ( .A1(n284), .A2(n278), .ZN(n238) );
  INV_X1 U279 ( .A(n227), .ZN(n278) );
  INV_X1 U280 ( .A(n239), .ZN(n282) );
  AND2_X1 U281 ( .A1(n285), .A2(Result_7_), .ZN(n239) );
  AND2_X1 U282 ( .A1(n227), .A2(n286), .ZN(Result_7_) );
  AND2_X1 U283 ( .A1(n287), .A2(n288), .ZN(n227) );
  OR2_X1 U284 ( .A1(c_3_), .A2(d_3_), .ZN(n287) );
  INV_X1 U285 ( .A(n289), .ZN(n233) );
  OR2_X1 U286 ( .A1(n290), .A2(n291), .ZN(n289) );
  INV_X1 U287 ( .A(n292), .ZN(n291) );
  OR3_X1 U288 ( .A1(n229), .A2(n293), .A3(n285), .ZN(n292) );
  AND2_X1 U289 ( .A1(n285), .A2(n294), .ZN(n290) );
  OR2_X1 U290 ( .A1(n293), .A2(n229), .ZN(n294) );
  INV_X1 U291 ( .A(n295), .ZN(n285) );
  AND2_X1 U292 ( .A1(n296), .A2(n297), .ZN(n243) );
  INV_X1 U293 ( .A(n298), .ZN(n297) );
  AND2_X1 U294 ( .A1(n299), .A2(n300), .ZN(n298) );
  OR2_X1 U295 ( .A1(n300), .A2(n299), .ZN(n296) );
  OR2_X1 U296 ( .A1(n301), .A2(n302), .ZN(n299) );
  AND2_X1 U297 ( .A1(n303), .A2(n304), .ZN(n302) );
  INV_X1 U298 ( .A(n305), .ZN(n301) );
  OR2_X1 U299 ( .A1(n304), .A2(n303), .ZN(n305) );
  INV_X1 U300 ( .A(n306), .ZN(n303) );
  OR2_X1 U301 ( .A1(n307), .A2(n308), .ZN(n253) );
  AND2_X1 U302 ( .A1(n309), .A2(n310), .ZN(n308) );
  INV_X1 U303 ( .A(n311), .ZN(n307) );
  OR2_X1 U304 ( .A1(n310), .A2(n309), .ZN(n311) );
  OR2_X1 U305 ( .A1(n312), .A2(n313), .ZN(n309) );
  AND2_X1 U306 ( .A1(n314), .A2(n315), .ZN(n313) );
  INV_X1 U307 ( .A(n316), .ZN(n314) );
  AND2_X1 U308 ( .A1(n317), .A2(n316), .ZN(n312) );
  INV_X1 U309 ( .A(n315), .ZN(n317) );
  INV_X1 U310 ( .A(n265), .ZN(n263) );
  OR2_X1 U311 ( .A1(n318), .A2(n266), .ZN(n265) );
  AND2_X1 U312 ( .A1(n319), .A2(n271), .ZN(n318) );
  OR2_X1 U313 ( .A1(n320), .A2(n321), .ZN(n271) );
  INV_X1 U314 ( .A(n273), .ZN(n320) );
  INV_X1 U315 ( .A(n322), .ZN(n319) );
  AND3_X1 U316 ( .A1(n322), .A2(n273), .A3(n274), .ZN(n266) );
  INV_X1 U317 ( .A(n321), .ZN(n274) );
  OR2_X1 U318 ( .A1(n323), .A2(n324), .ZN(n321) );
  AND2_X1 U319 ( .A1(n316), .A2(n315), .ZN(n324) );
  AND2_X1 U320 ( .A1(n310), .A2(n325), .ZN(n323) );
  OR2_X1 U321 ( .A1(n315), .A2(n316), .ZN(n325) );
  OR2_X1 U322 ( .A1(n326), .A2(n327), .ZN(n316) );
  AND2_X1 U323 ( .A1(n306), .A2(n304), .ZN(n327) );
  AND2_X1 U324 ( .A1(n300), .A2(n328), .ZN(n326) );
  OR2_X1 U325 ( .A1(n304), .A2(n306), .ZN(n328) );
  OR2_X1 U326 ( .A1(n228), .A2(n284), .ZN(n306) );
  OR3_X1 U327 ( .A1(n293), .A2(n229), .A3(n295), .ZN(n304) );
  OR2_X1 U328 ( .A1(n228), .A2(n329), .ZN(n295) );
  AND2_X1 U329 ( .A1(n330), .A2(n331), .ZN(n300) );
  OR3_X1 U330 ( .A1(n229), .A2(n332), .A3(n333), .ZN(n331) );
  INV_X1 U331 ( .A(n286), .ZN(n229) );
  OR2_X1 U332 ( .A1(n334), .A2(n335), .ZN(n330) );
  AND2_X1 U333 ( .A1(n286), .A2(n336), .ZN(n335) );
  OR2_X1 U334 ( .A1(n228), .A2(n279), .ZN(n315) );
  AND2_X1 U335 ( .A1(n337), .A2(n338), .ZN(n228) );
  INV_X1 U336 ( .A(n339), .ZN(n338) );
  AND2_X1 U337 ( .A1(n340), .A2(n288), .ZN(n339) );
  OR2_X1 U338 ( .A1(n340), .A2(n288), .ZN(n337) );
  OR2_X1 U339 ( .A1(n341), .A2(n342), .ZN(n340) );
  AND2_X1 U340 ( .A1(c_2_), .A2(n343), .ZN(n342) );
  AND2_X1 U341 ( .A1(d_2_), .A2(n344), .ZN(n341) );
  AND2_X1 U342 ( .A1(n345), .A2(n346), .ZN(n310) );
  INV_X1 U343 ( .A(n347), .ZN(n346) );
  AND2_X1 U344 ( .A1(n348), .A2(n349), .ZN(n347) );
  OR2_X1 U345 ( .A1(n349), .A2(n348), .ZN(n345) );
  OR2_X1 U346 ( .A1(n350), .A2(n351), .ZN(n348) );
  INV_X1 U347 ( .A(n352), .ZN(n351) );
  OR2_X1 U348 ( .A1(n353), .A2(n354), .ZN(n352) );
  AND2_X1 U349 ( .A1(n354), .A2(n353), .ZN(n350) );
  OR2_X1 U350 ( .A1(n293), .A2(n284), .ZN(n353) );
  OR2_X1 U351 ( .A1(n329), .A2(n332), .ZN(n349) );
  AND2_X1 U352 ( .A1(n355), .A2(n356), .ZN(n273) );
  INV_X1 U353 ( .A(n357), .ZN(n356) );
  AND2_X1 U354 ( .A1(n358), .A2(n359), .ZN(n357) );
  OR2_X1 U355 ( .A1(n358), .A2(n359), .ZN(n355) );
  OR2_X1 U356 ( .A1(n360), .A2(n361), .ZN(n358) );
  AND2_X1 U357 ( .A1(n362), .A2(n363), .ZN(n361) );
  AND2_X1 U358 ( .A1(n364), .A2(n365), .ZN(n360) );
  OR2_X1 U359 ( .A1(n366), .A2(n367), .ZN(n322) );
  AND3_X1 U360 ( .A1(n336), .A2(n368), .A3(n270), .ZN(n367) );
  INV_X1 U361 ( .A(n279), .ZN(n270) );
  AND2_X1 U362 ( .A1(n279), .A2(n269), .ZN(n366) );
  INV_X1 U363 ( .A(n368), .ZN(n269) );
  OR2_X1 U364 ( .A1(n369), .A2(n370), .ZN(n368) );
  AND2_X1 U365 ( .A1(n359), .A2(n365), .ZN(n370) );
  AND2_X1 U366 ( .A1(n364), .A2(n371), .ZN(n369) );
  OR2_X1 U367 ( .A1(n365), .A2(n359), .ZN(n371) );
  OR2_X1 U368 ( .A1(n293), .A2(n279), .ZN(n359) );
  INV_X1 U369 ( .A(n363), .ZN(n364) );
  OR2_X1 U370 ( .A1(n354), .A2(n372), .ZN(n363) );
  AND2_X1 U371 ( .A1(n362), .A2(n333), .ZN(n372) );
  INV_X1 U372 ( .A(n365), .ZN(n362) );
  OR2_X1 U373 ( .A1(n284), .A2(n332), .ZN(n365) );
  AND2_X1 U374 ( .A1(n373), .A2(n374), .ZN(n284) );
  INV_X1 U375 ( .A(n375), .ZN(n374) );
  AND2_X1 U376 ( .A1(n376), .A2(n377), .ZN(n375) );
  OR2_X1 U377 ( .A1(n376), .A2(n377), .ZN(n373) );
  OR2_X1 U378 ( .A1(n378), .A2(n379), .ZN(n376) );
  INV_X1 U379 ( .A(n380), .ZN(n379) );
  OR2_X1 U380 ( .A1(n381), .A2(b_1_), .ZN(n380) );
  AND2_X1 U381 ( .A1(b_1_), .A2(n381), .ZN(n378) );
  INV_X1 U382 ( .A(a_1_), .ZN(n381) );
  AND3_X1 U383 ( .A1(n286), .A2(n336), .A3(n333), .ZN(n354) );
  INV_X1 U384 ( .A(n334), .ZN(n333) );
  OR2_X1 U385 ( .A1(n329), .A2(n293), .ZN(n334) );
  AND2_X1 U386 ( .A1(n382), .A2(n383), .ZN(n293) );
  INV_X1 U387 ( .A(n384), .ZN(n383) );
  AND2_X1 U388 ( .A1(n385), .A2(n386), .ZN(n384) );
  OR2_X1 U389 ( .A1(n385), .A2(n386), .ZN(n382) );
  OR2_X1 U390 ( .A1(n387), .A2(n388), .ZN(n385) );
  INV_X1 U391 ( .A(n389), .ZN(n388) );
  OR2_X1 U392 ( .A1(n390), .A2(d_1_), .ZN(n389) );
  AND2_X1 U393 ( .A1(d_1_), .A2(n390), .ZN(n387) );
  INV_X1 U394 ( .A(c_1_), .ZN(n390) );
  INV_X1 U395 ( .A(n226), .ZN(n329) );
  OR2_X1 U396 ( .A1(n391), .A2(n392), .ZN(n226) );
  AND2_X1 U397 ( .A1(n393), .A2(n394), .ZN(n392) );
  INV_X1 U398 ( .A(n395), .ZN(n391) );
  OR2_X1 U399 ( .A1(n393), .A2(n394), .ZN(n395) );
  OR2_X1 U400 ( .A1(n396), .A2(n397), .ZN(n393) );
  AND2_X1 U401 ( .A1(a_2_), .A2(n398), .ZN(n397) );
  AND2_X1 U402 ( .A1(b_2_), .A2(n399), .ZN(n396) );
  INV_X1 U403 ( .A(n332), .ZN(n336) );
  OR2_X1 U404 ( .A1(n400), .A2(n401), .ZN(n332) );
  AND2_X1 U405 ( .A1(n402), .A2(n403), .ZN(n401) );
  INV_X1 U406 ( .A(n404), .ZN(n400) );
  OR2_X1 U407 ( .A1(n403), .A2(n402), .ZN(n404) );
  OR2_X1 U408 ( .A1(n405), .A2(n406), .ZN(n402) );
  AND2_X1 U409 ( .A1(c_0_), .A2(n407), .ZN(n406) );
  INV_X1 U410 ( .A(d_0_), .ZN(n407) );
  AND2_X1 U411 ( .A1(d_0_), .A2(n408), .ZN(n405) );
  INV_X1 U412 ( .A(c_0_), .ZN(n408) );
  OR2_X1 U413 ( .A1(n409), .A2(n410), .ZN(n403) );
  AND2_X1 U414 ( .A1(n411), .A2(c_1_), .ZN(n410) );
  AND2_X1 U415 ( .A1(d_1_), .A2(n412), .ZN(n409) );
  OR2_X1 U416 ( .A1(n411), .A2(c_1_), .ZN(n412) );
  INV_X1 U417 ( .A(n386), .ZN(n411) );
  OR2_X1 U418 ( .A1(n413), .A2(n414), .ZN(n386) );
  AND2_X1 U419 ( .A1(n288), .A2(n344), .ZN(n414) );
  AND2_X1 U420 ( .A1(n415), .A2(n343), .ZN(n413) );
  INV_X1 U421 ( .A(d_2_), .ZN(n343) );
  OR2_X1 U422 ( .A1(n344), .A2(n288), .ZN(n415) );
  INV_X1 U423 ( .A(n416), .ZN(n288) );
  AND2_X1 U424 ( .A1(c_3_), .A2(d_3_), .ZN(n416) );
  INV_X1 U425 ( .A(c_2_), .ZN(n344) );
  AND2_X1 U426 ( .A1(n417), .A2(n394), .ZN(n286) );
  OR2_X1 U427 ( .A1(a_3_), .A2(b_3_), .ZN(n417) );
  OR2_X1 U428 ( .A1(n418), .A2(n419), .ZN(n279) );
  AND2_X1 U429 ( .A1(n420), .A2(n421), .ZN(n419) );
  INV_X1 U430 ( .A(n422), .ZN(n418) );
  OR2_X1 U431 ( .A1(n421), .A2(n420), .ZN(n422) );
  OR2_X1 U432 ( .A1(n423), .A2(n424), .ZN(n420) );
  AND2_X1 U433 ( .A1(a_0_), .A2(n425), .ZN(n424) );
  INV_X1 U434 ( .A(b_0_), .ZN(n425) );
  AND2_X1 U435 ( .A1(b_0_), .A2(n426), .ZN(n423) );
  INV_X1 U436 ( .A(a_0_), .ZN(n426) );
  OR2_X1 U437 ( .A1(n427), .A2(n428), .ZN(n421) );
  AND2_X1 U438 ( .A1(n429), .A2(a_1_), .ZN(n428) );
  AND2_X1 U439 ( .A1(b_1_), .A2(n430), .ZN(n427) );
  OR2_X1 U440 ( .A1(n429), .A2(a_1_), .ZN(n430) );
  INV_X1 U441 ( .A(n377), .ZN(n429) );
  OR2_X1 U442 ( .A1(n431), .A2(n432), .ZN(n377) );
  AND2_X1 U443 ( .A1(n394), .A2(n399), .ZN(n432) );
  AND2_X1 U444 ( .A1(n433), .A2(n398), .ZN(n431) );
  INV_X1 U445 ( .A(b_2_), .ZN(n398) );
  OR2_X1 U446 ( .A1(n399), .A2(n394), .ZN(n433) );
  INV_X1 U447 ( .A(n434), .ZN(n394) );
  AND2_X1 U448 ( .A1(a_3_), .A2(b_3_), .ZN(n434) );
  INV_X1 U449 ( .A(a_2_), .ZN(n399) );
endmodule

