module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, n2982, g2124, n2981,
         n2985, g1430, n2984, n2988, g744, n2987, n2991, g56, n2990, n3742,
         n3741, n8104, g16802, n8103, DFF_1_n1, g16823, n8102, g2950, n4423,
         n4274, g2883, n4330, g22026, g2888, g23358, g2896, n4431, g24473,
         g2892, g25201, g2903, n4305, g26037, g2900, n4291, g26798, g2908,
         n4355, n4273, g2912, n4482, g23357, g2917, n4479, g24476, g2924,
         n4349, g25199, g2920, n4280, DFF_15_n1, n4281, n8099, DFF_16_n1,
         n8098, DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938, g2941,
         g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975,
         g2978, g2981, g2874, g18754, g1506, n4288, g18781, g1501, n4565,
         g18803, g1496, n4557, g18821, g1491, n4326, g18835, g1486, n4390,
         g18852, g1481, n4320, g18866, g1476, n4374, g18883, g1471, n4378,
         g21880, g2877, g19154, g813, n4289, g19163, g809, n4567, g19173, g805,
         n4559, g19184, g801, n4327, g20310, g797, n4391, g20343, g793, n4321,
         g20376, g789, n4375, g20417, g785, n4379, g21878, g2873, g19153, g125,
         n4290, g19162, g121, n4569, g19172, g117, n4561, g19144, g113, n4328,
         g19149, g109, n4392, g19157, g105, n4322, g19167, g101, n4376, g19178,
         g97, n4380, g20874, g2857, g18885, g2200, n4287, g18975, g2195, n4563,
         g18968, g2190, n4555, g18942, g2185, n4325, g18906, g2180, n4389,
         g18867, g2175, n4319, g18836, g2170, n4373, g18957, g2165, n4377,
         g21882, g2878, n4598, n4382, n4383, g3109, n4494, g18669, g18719,
         g3211, g18782, g3084, n4445, g17222, g3085, n4340, g17225, g3086,
         n4337, g17234, g3087, n4344, g17224, g3091, g17228, g3092, g17246,
         g3093, g17226, g3094, g17235, g3095, n4439, g17269, g3096, n4336,
         g25450, g3097, n4433, g25451, g3098, n4434, g25452, g3099, n4443,
         g28420, g3100, n4342, g28421, g28425, g3102, n4343, g29936, g3103,
         n4447, g29939, g3104, n4452, g29941, g3105, g30796, g3106, n4438,
         g30798, g3107, n4437, g30801, g3108, n4334, g17229, g3155, g17247,
         g3158, n4436, g17302, g3161, g17236, g3164, n4339, g17270, g3167,
         n4348, g17340, g3170, n4441, g17248, g3173, n4338, g17303, g3176,
         n4450, g17383, g17271, g3182, n4453, g17341, g3185, n4442, g17429,
         g3088, n4341, n8090, n8089, g3197, n8088, g3201, n4406, g3204, g3207,
         n4329, g3188, n4405, g3133, n8087, DFF_140_n1, g3128, n8086, n8084,
         g3124, n8083, DFF_146_n1, n8082, n8081, n8080, g3112, g3110, g3111,
         n8079, n8078, n8077, DFF_155_n1, n8076, DFF_156_n1, g3151, n4424,
         g3142, n4301, g185, n4384, n4318, n4512, g165, n4369, g22100, g130,
         g22122, g131, g22141, g129, g22123, g133, g22142, g134, g22161, g132,
         g22025, g142, g22027, g143, g22030, g141, g22028, g145, g22031, g146,
         g22037, g22032, g148, g22038, g149, g22047, g147, g22039, g151,
         g22048, g152, g22063, g150, g22049, g154, g22064, g155, g22079, g153,
         g22065, g157, g22080, g158, g22101, g156, g22081, g160, g22102, g161,
         g22124, g159, g22103, g22125, g164, g22143, g162, g25204, g169,
         g25206, g170, g25211, g168, g25207, g172, g25212, g173, g25218, g171,
         g25213, g175, g25219, g176, g25228, g174, g25220, g178, g25229, g179,
         g25239, g177, g30261, g186, g30267, g30275, g192, g30637, g231,
         g30640, g234, g30645, g237, g30668, g195, g30674, g198, g30680, g201,
         g30641, g240, g30646, g243, g30653, g246, g30276, g204, g30284, g207,
         g30292, g210, g30254, g249, g30257, g252, g30262, g30245, g213,
         g30246, g216, g30248, g219, g30258, g258, g30263, g261, g30268, g264,
         g30635, g222, g30636, g225, g30639, g228, g30661, g267, g30669, g270,
         g30675, g273, g25027, g92, g25932, g88, g26529, g83, g27120, g27594,
         g74, g28145, g70, g28634, g65, g29109, g61, g29353, g29579, g52, g180,
         g181, n4506, g309, n4388, g27253, g354, g27255, g343, g27258, g27256,
         g369, g27259, g358, g27265, g361, g27260, g384, g27266, g373, g27277,
         g376, g27267, g398, g27278, g388, g27293, g391, g28732, g408, g28735,
         g411, g28744, g414, g29194, g417, g29197, g420, g29201, g423, g28736,
         g28745, g428, g28754, g426, g26803, g429, g26804, g432, g26807, g435,
         g26805, g438, g26808, g441, g26812, g444, g27759, g448, g27760, g449,
         g27762, g447, g29606, g312, g29608, g313, g29611, g314, g30699, g315,
         g30700, g30702, g317, g30455, g318, g30468, g319, g30482, g320,
         g29167, g322, g29169, g323, g29172, g321, g26655, g403, g26659, g404,
         g26664, g402, g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454,
         DFF_303_n1, g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284,
         n8060, DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1,
         g290, n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055,
         DFF_328_n1, g349, g350, g351, g352, g353, g357, g364, g365, g366,
         g367, g368, g372, g379, g380, g381, g383, g387, g394, g395, g396,
         g397, g324, g337, n4298, n4372, g550, n4313, g554, g18678, g557,
         n4360, g18726, g513, g523, g524, g455, g564, g569, g458, g570, g571,
         g461, g572, g573, g465, g574, g565, g566, g567, g471, g568, g489,
         n4461, g485, n4466, g23067, g486, g23093, g487, g23117, g488, g23385,
         g23399, g24174, g24178, g477, g24207, g478, g24216, g479, g23092,
         g480, g23000, g484, g23022, g464, g24206, g24215, g24228, g528, g535,
         g542, g13149, g543, g544, g21851, g548, g13111, g549, g499, n4541,
         g13160, g558, g559, g27261, g576, g27268, g577, g27279, g575, g27269,
         g579, g27280, g27294, g578, g27281, g582, g27295, g583, g27311, g581,
         g27296, g585, g27312, g586, g27327, g584, g24491, g587, g24498, g590,
         g24507, g593, g24499, g596, g24508, g599, g24519, g602, g28345, g614,
         g28349, g617, g28353, g28342, g605, g28344, g608, g28348, g611,
         g26541, g490, g26545, g493, g26553, g496, g506, n4570, g22578, n4571,
         g525, n8047, n8046, DFF_445_n1, n8045, DFF_446_n1, n8044, n8043, g536,
         g537, g24059, g538, n4492, n8040, n4359, g629, n4295, g16654, g630,
         g20314, g659, g20682, g640, n4404, g23136, g633, n4478, g23324, g653,
         n4422, g24426, g646, n4414, g25185, g660, n4403, g26660, g672, n4413,
         g26776, g27672, g679, n4477, g28199, g686, n4396, g28668, g692, n4418,
         g20875, g699, g20879, g700, g20891, g698, g20880, g702, g20892, g703,
         g20901, g701, g20893, g705, g20902, g706, g20921, g704, g20903, g708,
         g20922, g709, g20944, g707, g20923, g20945, g712, g20966, g710,
         g20946, g714, g20967, g715, g20989, g713, g20968, g717, g20990, g718,
         g21009, g716, g20991, g720, g21010, g721, g21031, g719, g21011, g723,
         g21032, g724, g21051, g722, g20876, g726, g20881, g20894, g725,
         g20924, g729, g20947, g730, g20969, g728, g20948, g732, g20970, g733,
         g20992, g731, g25260, g735, g25262, g736, g25266, g734, g22218, g738,
         g22231, g739, g22242, g737, n4323, n4312, g22126, g818, g22145, g819,
         g22162, g817, g22146, g821, g22163, g822, g22177, g820, g22029, g830,
         g22033, g831, g22040, g829, g22034, g833, g22041, g834, g22054, g832,
         g22042, g836, g22055, g837, g22066, g835, g22056, g22067, g840,
         g22087, g838, g22068, g842, g22088, g843, g22104, g841, g22089, g845,
         g22105, g846, g22127, g844, g22106, g848, g22128, g849, g22147, g847,
         g22129, g851, g22148, g852, g22164, g850, g25209, g857, g25214,
         g25221, g856, g25215, g860, g25222, g861, g25230, g859, g25223, g863,
         g25231, g864, g25240, g862, g25232, g866, g25241, g867, g25248, g865,
         g30269, g873, g30277, g876, g30285, g879, g30643, g918, g30648, g921,
         g30654, g30676, g882, g30681, g885, g30687, g888, g30649, g927,
         g30655, g930, g30662, g933, g30286, g891, g30293, g894, g30298, g897,
         g30259, g936, g30264, g939, g30270, g942, g30247, g900, g30249, g903,
         g30251, g906, g30265, g30271, g948, g30278, g951, g30638, g909,
         g30642, g912, g30647, g915, g30670, g954, g30677, g957, g30682, g960,
         g25042, g780, g25935, g776, g26530, g771, g27123, g767, g27603, g762,
         g28146, g758, g28635, g753, g29110, g29354, g29580, g740, g868, g869,
         n4363, n4364, g1088, n4381, g996, n4387, g27257, g1041, g27262, g1030,
         g27270, g1033, g27263, g1056, g27271, g1045, g27282, g1048, g27272,
         g27283, g1060, g27297, g1063, g27284, g1085, g27298, g1075, g27313,
         g1078, g28738, g1095, g28746, g1098, g28758, g1101, g29198, g1104,
         g29204, g1107, g29209, g1110, g28747, g1114, g28759, g1115, g28767,
         g1113, g26806, g1116, g26809, g26813, g1122, g26810, g1125, g26814,
         g1128, g26818, g1131, g27761, g1135, g27763, g1136, g27765, g1134,
         g29609, g999, g29612, g1000, g29616, g1001, g30701, g1002, g30703,
         g1003, g30705, g1004, g30470, g1005, g30485, g1006, g30500, g29170,
         g1009, g29173, g1010, g29179, g1008, g26661, g1090, g26665, g1091,
         g26669, g1089, g1137, n8027, DFF_649_n1, g1139, n8026, DFF_651_n1,
         g1141, n8025, DFF_653_n1, g967, n8024, DFF_655_n1, g969, DFF_657_n1,
         g971, n8021, DFF_659_n1, g973, n8020, DFF_661_n1, g975, n8019,
         DFF_663_n1, g977, n8018, n4486, n4283, g986, n4432, g992, n4277,
         n8017, g1029, g1036, g1037, g1038, g1040, g1044, g1051, g1052, g1053,
         g1054, g1055, g1059, g1066, g1067, g1068, g1069, g1070, g1074, g1081,
         g1083, g1084, g1011, g1024, n4371, n4316, g1236, n4300, g1240, g18707,
         g1243, n4353, g18763, g1196, n4304, g1199, g1209, g1210, g1142, g1255,
         g1145, g1256, g1257, g1148, g1258, g1259, g1152, g1260, g1251, g1155,
         g1252, g1253, g1158, g1254, g1176, n4460, n4459, g1172, n4465, g23081,
         g1173, g23111, g23126, g1175, g23392, g23406, g24179, g24181, g1164,
         g24213, g1165, g24223, g1166, g23110, g1167, g23014, g1171, g23039,
         g1151, g24212, g24222, g24235, g1214, g1221, g13155, g1229, n4549,
         n4361, g13124, g1235, g1186, n4548, g13171, g1244, g1245, g27273,
         g1262, g27285, g1263, g27299, g1261, g27286, g1265, g27300, g1266,
         g27314, g1264, g27301, g1268, g27315, g1269, g27328, g27316, g1271,
         g27329, g1272, g27339, g1270, g24501, g1273, g24510, g1276, g24521,
         g1279, g24511, g1282, g24522, g1285, g24532, g1288, g28351, g1300,
         g28355, g1303, g28360, g1306, g28346, g1291, g28350, g1294, g28354,
         g1297, g26547, g26557, g1180, g26569, g1183, g1192, n4454, g22615,
         n8009, DFF_783_n1, DFF_792_n1, g1211, n8008, n8007, DFF_795_n1, n8006,
         DFF_796_n1, n8005, n8004, n8003, g1222, g1223, g24072, g1224, n4489,
         n4358, g1315, n4294, g16671, g1316, g20333, g1345, g20717, g1326,
         n4402, g21969, g1319, n4476, g23329, g1339, n4421, g24430, g1332,
         n4412, g25189, g1346, n4401, g26666, g1358, n4411, g26781, g1352,
         n4469, g27678, g1365, n4475, g27718, g1372, n4395, g28321, g1378,
         n4417, g20882, g20896, g1386, g20910, g1384, g20897, g1388, g20911,
         g1389, g20925, g1387, g20912, g1391, g20926, g1392, g20949, g1390,
         g20927, g1394, g20950, g1395, g20972, g1393, g20951, g1397, g20973,
         g1398, g20993, g1396, g20974, g1400, g20994, g21015, g1399, g20995,
         g1403, g21016, g1404, g21033, g1402, g21017, g1406, g21034, g1407,
         g21052, g1405, g21035, g1409, g21053, g1410, g21070, g1408, g20883,
         g1412, g20898, g1413, g20913, g1411, g20952, g1415, g20975, g1416,
         g20996, g20976, g1418, g20997, g1419, g21018, g1417, g25263, g1421,
         g25267, g1422, g25270, g1420, g22234, g1424, g22247, g1425, g22263,
         g1423, n4317, n4515, g1547, n4368, g22149, g1512, g22166, g1513,
         g22178, g1511, g22167, g22179, g1516, g22191, g1514, g22035, g1524,
         g22043, g1525, g22057, g1523, g22044, g1527, g22058, g1528, g22073,
         g1526, g22059, g1530, g22074, g1531, g22090, g1529, g22075, g1533,
         g22091, g1534, g22112, g1532, g22092, g1536, g22113, g22130, g1535,
         g22114, g1539, g22131, g1540, g22150, g1538, g22132, g1542, g22151,
         g1543, g22168, g1541, g22152, g1545, g22169, g1546, g22180, g1544,
         g25217, g1551, g25224, g1552, g25233, g1550, g25225, g1554, g25234,
         g1555, g25242, g25235, g1557, g25243, g1558, g25249, g1556, g25244,
         g1560, g25250, g1561, g25255, g1559, g30279, g1567, g30287, g1570,
         g30294, g1573, g30651, g1612, g30657, g1615, g30663, g1618, g30683,
         g1576, g30688, g1579, g30692, g1582, g30658, g30664, g1624, g30671,
         g1627, g30295, g1585, g30299, g1588, g30302, g1591, g30266, g1630,
         g30272, g1633, g30280, g1636, g30250, g1594, g30252, g1597, g30255,
         g1600, g30273, g1639, g30281, g1642, g30288, g1645, g30644, g1603,
         g30650, g30656, g1609, g30678, g1648, g30684, g1651, g30689, g1654,
         g25056, g1466, g25938, g1462, g26531, g1457, g27129, g1453, g27612,
         g1448, g28147, g1444, g28636, g1439, g29111, g1435, g29355, g29581,
         g1426, g1562, g1563, n4518, g1690, n4386, g27264, g1735, g27274,
         g1724, g27287, g1727, g27275, g1750, g27288, g1739, g27302, g1742,
         g27289, g1765, g27303, g1754, g27317, g1757, g27304, g1779, g27318,
         g27330, g1772, g28749, g1789, g28760, g1792, g28771, g1795, g29205,
         g1798, g29212, g1801, g29218, g1804, g28761, g1808, g28772, g1809,
         g28778, g1807, g26811, g1810, g26815, g1813, g26820, g1816, g26816,
         g1819, g26821, g1822, g26824, g27764, g1829, g27766, g1830, g27768,
         g1828, g29613, g1693, g29617, g1694, g29620, g1695, g30704, g1696,
         g30706, g1697, g30708, g1698, g30487, g1699, g30503, g1700, g30338,
         g1701, g29178, g1703, g29181, g1704, g29184, g1702, g26667, g26670,
         g1785, g26675, g1783, g1831, n7988, DFF_999_n1, g1833, n7987,
         DFF_1001_n1, g1835, n7986, DFF_1003_n1, g1661, n7985, DFF_1005_n1,
         g1663, n7984, DFF_1007_n1, g1665, n7983, DFF_1009_n1, g1667,
         DFF_1011_n1, g1669, n7980, DFF_1013_n1, g1671, n7979, n4484, n4284,
         g1680, n4488, g1686, n4276, n7978, g1723, g1730, g1731, g1732, g1733,
         g1734, g1738, g1745, g1747, g1748, g1749, g1753, g1760, g1761, g1762,
         g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1718, n4296,
         n4315, g1930, n4366, g1934, g18743, g1937, n4311, g18794, g1890,
         n4297, g1893, g1903, g1904, g1836, g1944, g1949, g1950, g1951, g1842,
         g1953, g1846, g1954, g1945, g1849, g1946, g1947, g1852, g1948, g1870,
         n4458, n4457, g1866, n4464, g23097, g1867, g23124, g1868, g23137,
         g1869, g23400, g23413, g24182, g24208, g1858, g24219, g1859, g24231,
         g1860, g23123, g1861, g23030, g1865, g23058, g1845, g24218, g24230,
         g24243, g1908, g1915, g1922, g13164, g1923, DFF_1099_n1, n7971,
         DFF_1100_n1, g13135, g1929, g1880, n4545, g13182, g1938, g1939,
         g27290, g1956, g27305, g1957, g27319, g1955, g27306, g1959, g27320,
         g1960, g27331, g1958, g27321, g1962, g27332, g1963, g27340, g1961,
         g27333, g27341, g1966, g27346, g1964, g24513, g1967, g24524, g1970,
         g24534, g1973, g24525, g1976, g24535, g1979, g24545, g1982, g28357,
         g1994, g28362, g1997, g28366, g2000, g28352, g1985, g28356, g1988,
         g28361, g1991, g26559, g26573, g1874, g26592, g1877, g1886, n4493,
         g22651, n7968, DFF_1133_n1, DFF_1142_n1, g1905, n7967, n7966,
         DFF_1145_n1, n7965, DFF_1146_n1, n7964, n7963, n7962, g1916, g1917,
         g24083, n7960, n4357, g2009, n4293, g16692, g2010, g20353, g2039,
         g20752, g2020, n4400, g21972, g2013, n4474, g23339, g2033, n4420,
         g24434, g2026, n4410, g25194, g2040, n4399, g26671, g2052, n4409,
         g26789, g2046, n4468, g27682, g2059, n4473, g27722, g28325, g2072,
         n4416, g20899, g2079, g20915, g2080, g20934, g2078, g20916, g2082,
         g20935, g2083, g20953, g2081, g20936, g2085, g20954, g2086, g20977,
         g2084, g20955, g2088, g20978, g2089, g20999, g2087, g20979, g2091,
         g21000, g21019, g2090, g21001, g2094, g21020, g2095, g21039, g2093,
         g21021, g2097, g21040, g2098, g21054, g2096, g21041, g2100, g21055,
         g2101, g21071, g2099, g21056, g2103, g21072, g2104, g21080, g2102,
         g20900, g2106, g20917, g20937, g2105, g20980, g2109, g21002, g2110,
         g21022, g2108, g21003, g2112, g21023, g2113, g21042, g2111, g25268,
         g2115, g25271, g2116, g25279, g2114, g22249, g2118, g22267, g2119,
         g22280, g2117, n4324, g2241, n4367, g22170, g2206, g22182, g2207,
         g22192, g2205, g22183, g2209, g22193, g2210, g22200, g2208, g22045,
         g2218, g22060, g2219, g22076, g2217, g22061, g2221, g22077, g2222,
         g22097, g2220, g22078, g2224, g22098, g22115, g2223, g22099, g2227,
         g22116, g2228, g22138, g2226, g22117, g2230, g22139, g2231, g22153,
         g2229, g22140, g2233, g22154, g2234, g22171, g2232, g22155, g2236,
         g22172, g2237, g22184, g2235, g22173, g2239, g22185, g22194, g2238,
         g25227, g2245, g25236, g2246, g25245, g2244, g25237, g2248, g25246,
         g2249, g25251, g2247, g25247, g2251, g25252, g2252, g25256, g2250,
         g25253, g2254, g25257, g2255, g25259, g2253, g30289, g2261, g30296,
         g30300, g2267, g30660, g2306, g30666, g2309, g30672, g2312, g30690,
         g2270, g30693, g2273, g30695, g2276, g30667, g2315, g30673, g2318,
         g30679, g2321, g30301, g2279, g30303, g2282, g30304, g2285, g30274,
         g2324, g30282, g30290, g2330, g30253, g2288, g30256, g2291, g30260,
         g2294, g30283, g2333, g30291, g2336, g30297, g2339, g30652, g2297,
         g30659, g2300, g30665, g2303, g30686, g2342, g30691, g2345, g30694,
         g2348, g25067, g2160, g25940, g26532, g2151, g27131, g2147, g27621,
         g2142, g28148, g2138, g28637, g2133, g29112, g2129, g29357, g29582,
         g2120, g2256, g2257, n4516, g27276, g2429, g27291, g2418, g27307,
         g2421, g27292, g2444, g27308, g2433, g27322, g2436, g27309, g2459,
         g27323, g2448, g27334, g2451, g27324, g2473, g27335, g2463, g27342,
         g2466, g28763, g2483, g28773, g2486, g28782, g29213, g2492, g29221,
         g2495, g29226, g2498, g28774, g2502, g28783, g2503, g28788, g2501,
         g26817, g2504, g26822, g2507, g26825, g2510, g26823, g2513, g26826,
         g2516, g26827, g2519, g27767, g2523, g27769, g2524, g27771, g29618,
         g2387, g29621, g2388, g29623, g2389, g30707, g2390, g30709, g2391,
         g30566, g2392, g30505, g2393, g30341, g2394, g30356, g2395, g29182,
         g2397, g29185, g2398, g29187, g2396, g26672, g2478, g26676, g2479,
         g26025, g2525, n7946, DFF_1349_n1, g2527, n7945, DFF_1351_n1, g2529,
         n7944, DFF_1353_n1, g2355, n7943, DFF_1355_n1, g2357, n7942,
         DFF_1357_n1, g2359, n7941, DFF_1359_n1, g2361, n7940, DFF_1361_n1,
         n7938, DFF_1363_n1, g2365, n7937, n4483, n4285, g2374, n4487, g30055,
         g2380, n4275, n7936, DFF_1378_n1, g2417, g2424, g2425, g2426, g2427,
         g2428, g2432, g2439, g2441, g2442, g2443, g2447, g2454, g2455, g2456,
         g2457, g2458, g2462, g2469, g2470, g2471, g2472, g2412, n4314, n4370,
         g2624, n4299, g2628, g18780, g2631, n4352, g18820, g2584, n4303,
         g2587, g2597, g2598, g2530, g2638, g2643, g2533, g2645, g2536, g2646,
         g2647, g2540, g2648, g2639, g2543, g2640, g2641, g2546, g2642, g2564,
         n4456, n4455, g2560, n4463, g23114, g2561, g23133, g2562, g21970,
         g23407, g23418, g24209, g24214, g2552, g24226, g2553, g24238, g2554,
         g23132, g2555, g23047, g2559, g23076, g2539, g24225, g24237, g24250,
         g2602, g2609, g13175, g2617, n7930, g30072, n7929, g13143, g2623,
         g2574, n4543, g13194, g2632, g2633, g27310, g2650, g27325, g2651,
         g27336, g2649, g27326, g2653, g27337, g2654, g27343, g2652, g27338,
         g2656, g27344, g27347, g2655, g27345, g2659, g27348, g2660, g27354,
         g2658, g24527, g2661, g24537, g2664, g24547, g2667, g24538, g2670,
         g24548, g2673, g24557, g2676, g28364, g2688, g28368, g2691, g28371,
         g2694, g28358, g2679, g28363, g28367, g2685, g26575, g2565, g26596,
         g2568, g26616, g2571, g2580, g22687, n7926, g30061, g2599, n7925,
         n7924, DFF_1495_n1, n7923, DFF_1496_n1, n7922, n7921, n7920, g2611,
         g24092, g2612, n4490, n7918, n4356, g2703, n4292, g16718, g2704,
         g20375, g2733, g20789, g2714, n4398, g21974, g2707, n4472, g23348,
         g2727, n4419, g24438, g2720, n4408, g25197, g2734, n4397, g26677,
         g2746, n4407, g26795, g27243, g2753, n4471, g27724, g2760, n4393,
         g28328, g2766, n4415, g20918, g2773, g20939, g2774, g20962, g2772,
         g20940, g2776, g20963, g2777, g20981, g2775, g20964, g2779, g20982,
         g2780, g21004, g2778, g20983, g2782, g21005, g2783, g21025, g21006,
         g2785, g21026, g2786, g21043, g2784, g21027, g2788, g21044, g2789,
         g21060, g2787, g21045, g2791, g21061, g2792, g21073, g2790, g21062,
         g2794, g21074, g2795, g21081, g2793, g21075, g2797, g21082, g2798,
         g21094, g20919, g2800, g20941, g2801, g20965, g2799, g21007, g2803,
         g21028, g2804, g21046, g2802, g21029, g2806, g21047, g2807, g21063,
         g2805, g25272, g2809, g25280, g2810, g25288, g2808, g22269, g2812,
         g22284, g2813, g22299, g20877, n7913, DFF_1561_n1, g20884, n7912,
         DFF_1562_n1, n4263_Tj_Payload, n4269, g3043, n4268, g3044, n4267,
         g3045, n4266, g3046, n4265, g3047, n4272, g3048, n4271, g3049, n4270,
         g3050, n4259, g3051, n4236, g3052, n4239, g3053, n4237, n4234, g3056,
         n4233, g3057, n4238, g3058, n4235, g3059, n4240, g3060, n4232, g3061,
         n4245, g3062, n4248, g3063, n4246, g3064, n4243, g3065, n4242, g3066,
         n4247, g3067, n4244, g3068, n4249, g3069, n4241, n4254, g3071, n4257,
         g3072, n4255, g3073, n4252, g3074, n4251, g3075, n4256, g3076, n4253,
         g3077, n4258, g3078, n4250, g2997, g25265, g2993, g26048, n7909,
         g23330, g3006, g24445, g3002, g25191, g3013, g26031, g26786, g3024,
         n4262, g3018, n4481, g23359, g3028, n4350, g24446, g3036, n4480,
         g25202, g3032, n7907, DFF_1612_n1, g2987, n4365, g16824, g16844,
         g16853, g16860, g16803, g16835, g16851, g16857, g16866, g3083, n4261,
         N995, n4577, g16845, g16854, g16861, g16880, g18755, g18804, g18837,
         g18868, g18907, g2990, N690, n4578, n4260, n4309, n4308, n4307, n4306,
         n4524, n4525, n4511, n4509, n4499, n4520, n3683, n3887, n3686, n3890,
         n3692, n3896, n4513, n3897, n3424, n3427, n3433, n4529, n4530, n4522,
         n4523, n4521, n3171, n3159, n3163, n3893, n3690, n3689, n3431, n3430,
         n3168, n3160, n3164, n3172, n4527, n4528, n4526, n3167, n3894, n3888,
         n3891, n2302, n2289, n2303, n2275, n4066, n4065, n4606, n4618, n4640,
         n2617, n2351, n2792, n2632, n3936, n3252, n3254, n4102, n3038, n3070,
         n3102, n3130, n3036, n3068, n3128, n2800, n2798, n2616, n2594, n3940,
         n3705, n3933, n3939, n3016, n3000, n3008, n3023, n3700, n4123, n4101,
         n4182, n4073, n3749, n3751, n3758, n3788, n4057, n4122, n4263,
         Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6,
         Tj_OUT7, Tj_OUT8, Tj_OUT5678, Tj_Trigger, n18, n37, n73, n145, n278,
         n306, n307, n310, n318, n372, n529, n530, n557, n567, n588, n602,
         n618, n621, n622, n626, n627, n628, n630, n795, n982, n983, n987,
         n1146, n1330, n1333, n1335, n1497, n1658, n1683, n1684, n1689, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9425, n9426, n9427,
         n9429, n9430, n9431, n9432, n9436, n9438, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9452, n9453, n9454, n9456, n9457,
         n9459, n9460, n9461, n9462, n9463, n9464, n9469, n9470, n9472, n9474,
         n9475, n9477, n9478, n9480, n9481, n9482, n9484, n9486, n9488, n9490,
         n9492, n9493, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9512, n9514,
         n9516, n9518, n9519, n9521, n9522, n9523, n9528, n9529, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9556, n9558, n9562, n9564,
         n9567, n9568, n9569, n9570, n9571, n9572, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9585, n9586, n9587, n9588, n9589, n9595, n9599,
         n9600, n9601, n9602, n9603, n9604, n9607, n9609, n9611, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9627, n9629, n9631,
         n9636, n9637, n9638, n9639, n9642, n9643, n9645, n9650, n9651, n9652,
         n9653, n9654, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9671, n9672, n9673, n9674,
         n9678, n9681, n9683, n9684, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9716, n9717, n9719, n9720, n9722, n9724, n9726, n9727,
         n9728, n9729, n9730, n9732, n9733, n9734, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9754, n9756, n9760, n9762, n9764, n9767, n9769,
         n9771, n9773, n9774, n9775, n9777, n9778, n9780, n9781, n9783, n9784,
         n9786, n9787, n9788, n9790, n9791, n9793, n9794, n9796, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9815, n9817, n9818,
         n9820, n9826, n9829, n9832, n9836, n9837, n9838, n9840, n9841, n9842,
         n9843, n9845, n9847, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9858, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9880, n9882,
         n9884, n9887, n9888, n9889, n9891, n9894, n9897, n9900, n9903, n9906,
         n9908, n9911, n9913, n9916, n9919, n9922, n9925, n9928, n9931, n9934,
         n9944, n9947, n9949, n9954, n9956, n9960, n9965, n9967, n9970, n9972,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9984, n9987, n9991,
         n9992, n9995, n9997, n9998, n9999, n10003, n10004, n10005, n10006,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10039, n10040, n10042, n10043,
         n10045, n10046, n10048, n10049, n10051, n10052, n10054, n10056,
         n10057, n10059, n10060, n10062, n10063, n10065, n10066, n10068,
         n10069, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10164, n10165, n10166, n10167, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10178, n10179, n10180,
         n10181, n10184, n10185, n10186, n10187, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10272,
         n10273, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, U3772_n1, U3776_n1, U3777_n1,
         U3778_n1, U3779_n1, U3780_n1, U3781_n1, U3782_n1, U3783_n1, U3784_n1,
         U3785_n1, U3786_n1, U3787_n1, U3901_n1, U3902_n1, U4467_n1, U4904_n1,
         U4930_n1, U5128_n1, U5141_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1,
         U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1,
         U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5882_n1, U5939_n1,
         U5940_n1, U5941_n1, U5942_n1, U6140_n1, U6460_n1, U6470_n1, U6562_n1,
         U6563_n1, U6718_n1, U7116_n1, U7118_n1, U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n10342), .CLK(n10529), .Q(
        n8104), .QN(n18867) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n10342), .CLK(n10529), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n10342), .CLK(n10529), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n10342), .CLK(n10529), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n10343), .CLK(n10530), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n10343), .CLK(n10530), .Q(
        g2888) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n10343), .CLK(n10530), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n10343), .CLK(n10530), .Q(
        g2892), .QN(n10079) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n10343), .CLK(n10530), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n10343), .CLK(n10530), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n10343), .CLK(n10530), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n10343), .CLK(n10530), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n10343), .CLK(n10530), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n10343), .CLK(n10530), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n10343), .CLK(n10530), .Q(
        g2920), .QN(n10026) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n10343), .CLK(n10530), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n10340), .CLK(n10527), 
        .Q(n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n10340), .CLK(n10527), .Q(
        g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n10340), .CLK(n10527), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n10340), .CLK(n10527), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n10340), .CLK(n10527), .Q(
        g2934), .QN(n10292) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n10340), .CLK(n10527), .Q(
        g2935), .QN(n10275) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n10341), .CLK(n10528), .Q(
        g2938), .QN(n10276) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n10341), .CLK(n10528), .Q(
        g2941), .QN(n10273) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n10341), .CLK(n10528), .Q(
        g2944), .QN(n10279) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n10341), .CLK(n10528), .Q(
        g2947), .QN(n10277) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n10341), .CLK(n10528), .Q(
        g2953), .QN(n10278) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n10341), .CLK(n10528), .Q(
        g2956), .QN(n10280) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n10341), .CLK(n10528), .Q(
        g2959) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n10341), .CLK(n10528), .Q(
        g2962), .QN(n10294) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n10341), .CLK(n10528), .Q(
        g2963), .QN(n10283) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n10341), .CLK(n10528), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n10340), .CLK(n10527), 
        .Q(g2969), .QN(n10286) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n10340), .CLK(n10527), .Q(
        g2972), .QN(n10284) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n10340), .CLK(n10527), .Q(
        g2975), .QN(n10285) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n10340), .CLK(n10527), .Q(
        g2978), .QN(n10281) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n10340), .CLK(n10527), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n10340), .CLK(n10527), .Q(
        g2874), .QN(n10282) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n10341), .CLK(n10528), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n10341), .CLK(n10528), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n10342), .CLK(n10529), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n10342), .CLK(n10529), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n10342), .CLK(n10529), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n10342), .CLK(n10529), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n10342), .CLK(n10529), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n10342), .CLK(n10529), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n10351), .CLK(n10538), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n10351), .CLK(n10538), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n10351), .CLK(n10538), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n10351), .CLK(n10538), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n10351), .CLK(n10538), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n10351), .CLK(n10538), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n10352), .CLK(n10539), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n10352), .CLK(n10539), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n10352), .CLK(n10539), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n10352), .CLK(n10539), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n10352), .CLK(n10539), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n10352), .CLK(n10539), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n10352), .CLK(n10539), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n10352), .CLK(n10539), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n10352), .CLK(n10539), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n10352), .CLK(n10539), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n10352), .CLK(n10539), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n10353), .CLK(n10540), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n10353), .CLK(n10540), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n10353), .CLK(n10540), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n10353), .CLK(n10540), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n10353), .CLK(n10540), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n10354), .CLK(n10541), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n10354), .CLK(n10541), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n10354), .CLK(n10541), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n10354), .CLK(n10541), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n10354), .CLK(n10541), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n10354), .CLK(n10541), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n10354), .CLK(n10541), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n10354), .CLK(n10541), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n10354), .CLK(n10541), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n10354), .CLK(n10541), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n10354), .CLK(n10541), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n10354), .CLK(n10541), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n10355), .CLK(n10542), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n10355), .CLK(n10542), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n10355), .CLK(n10542), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n10355), .CLK(n10542), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n10355), .CLK(n10542), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n10355), .CLK(n10542), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n10355), .CLK(n10542), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n10355), .CLK(n10542), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n10355), .CLK(n10542), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n10355), .CLK(n10542), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n10355), .CLK(n10542), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n10458), .CLK(n10645), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n10466), .CLK(n10653), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n10466), .CLK(n10653), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n10466), .CLK(n10653), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n10468), .CLK(n10655), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n10466), .CLK(n10653), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n10466), .CLK(n10653), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n10467), .CLK(n10654), .Q(
        g3085), .QN(n4340) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n10467), .CLK(n10654), .Q(
        g3086), .QN(n4337) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n10467), .CLK(n10654), 
        .Q(g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n10467), .CLK(n10654), 
        .Q(g3091) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n10467), .CLK(n10654), 
        .Q(g3092) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n10467), .CLK(n10654), 
        .Q(g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n10467), .CLK(n10654), 
        .Q(g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n10467), .CLK(n10654), 
        .Q(g3095), .QN(n4439) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n10467), .CLK(n10654), 
        .Q(g3096), .QN(n4336) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n10468), .CLK(n10655), 
        .Q(g3097), .QN(n4433) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n10468), .CLK(n10655), 
        .Q(g3098), .QN(n4434) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n10468), .CLK(n10655), 
        .Q(g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n10468), .CLK(n10655), 
        .Q(g3100), .QN(n4342) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n10468), .CLK(n10655), 
        .Q(test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n10466), .CLK(n10653), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n10468), .CLK(n10655), 
        .Q(g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n10468), .CLK(n10655), 
        .Q(g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n10468), .CLK(n10655), 
        .Q(g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n10468), .CLK(n10655), 
        .Q(g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n10468), .CLK(n10655), 
        .Q(g3107), .QN(n4437) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n10468), .CLK(n10655), 
        .Q(g3108), .QN(n4334) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n10469), .CLK(n10656), 
        .Q(g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n10469), .CLK(n10656), 
        .Q(g3158), .QN(n4436) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n10469), .CLK(n10656), 
        .Q(g3161) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n10469), .CLK(n10656), 
        .Q(g3164), .QN(n4339) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n10469), .CLK(n10656), 
        .Q(g3167), .QN(n4348) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n10469), .CLK(n10656), 
        .Q(g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n10469), .CLK(n10656), 
        .Q(g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n10469), .CLK(n10656), 
        .Q(g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n10469), .CLK(n10656), 
        .Q(test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n10467), .CLK(n10654), 
        .Q(g3182), .QN(n4453) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n10467), .CLK(n10654), 
        .Q(g3185), .QN(n4442) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n10467), .CLK(n10654), 
        .Q(g3088), .QN(n4341) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n10469), .CLK(n10656), 
        .Q(n8090) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n10470), .CLK(n10657), 
        .Q(n8089), .QN(n18863) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n10470), .CLK(n10657), 
        .Q(g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n10470), .CLK(n10657), 
        .Q(n8088) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n10349), .CLK(n10536), 
        .Q(g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n10349), .CLK(n10536), 
        .Q(g3204), .QN(n10296) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n10349), .CLK(n10536), 
        .Q(g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n10349), .CLK(n10536), 
        .Q(g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n73), .SI(g3188), .SE(n10349), .CLK(n10536), .Q(
        g3133), .QN(n9737) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n10349), .CLK(n10536), 
        .Q(n8087), .QN(DFF_140_n1) );
  SDFFX1 DFF_141_Q_reg ( .D(n278), .SI(n8087), .SE(n10349), .CLK(n10536), .Q(
        g3128) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n10349), .CLK(n10536), 
        .Q(n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n10469), .CLK(n10656), 
        .Q(test_so9), .QN(n9636) );
  SDFFX1 DFF_144_Q_reg ( .D(n310), .SI(test_si10), .SE(n10469), .CLK(n10656), 
        .Q(n8084) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n10349), .CLK(n10536), 
        .Q(g3124), .QN(n9638) );
  SDFFX1 DFF_146_Q_reg ( .D(n318), .SI(g3124), .SE(n10349), .CLK(n10536), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n10349), .CLK(n10536), 
        .Q(n8082), .QN(n18868) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n10350), .CLK(n10537), 
        .Q(n8081), .QN(n18869) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n10350), .CLK(n10537), 
        .Q(n8080) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n10350), .CLK(n10537), 
        .Q(g3112), .QN(n9637) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n10350), .CLK(n10537), 
        .Q(g3110), .QN(n9604) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n10350), .CLK(n10537), 
        .Q(g3111), .QN(n9639) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n10350), .CLK(n10537), 
        .Q(n8079), .QN(n18870) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n10350), .CLK(n10537), 
        .Q(n8078), .QN(n18871) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n10350), .CLK(n10537), 
        .Q(n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n10350), .CLK(n10537), 
        .Q(n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n10350), .CLK(n10537), 
        .Q(g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n10350), .CLK(n10537), 
        .Q(g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n10350), .CLK(n10537), 
        .Q(test_so10), .QN(n10329) );
  SDFFX1 DFF_160_Q_reg ( .D(n73), .SI(test_si11), .SE(n10348), .CLK(n10535), 
        .Q(g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n10348), .CLK(n10535), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n10348), .CLK(n10535), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n10349), .CLK(n10536), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n10363), .CLK(n10550), .Q(
        g130) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n10363), .CLK(n10550), .Q(
        g131) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n10363), .CLK(n10550), .Q(
        g129), .QN(n9877) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n10364), .CLK(n10551), .Q(
        g133) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n10364), .CLK(n10551), .Q(
        g134) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n10364), .CLK(n10551), .Q(
        g132), .QN(n9876) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n10364), .CLK(n10551), .Q(
        g142) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n10364), .CLK(n10551), .Q(
        g143) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n10364), .CLK(n10551), .Q(
        g141), .QN(n9875) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n10364), .CLK(n10551), .Q(
        g145) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n10364), .CLK(n10551), .Q(
        g146) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n10364), .CLK(n10551), .Q(
        test_so11) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n10362), .CLK(n10549), 
        .Q(g148) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n10362), .CLK(n10549), .Q(
        g149) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n10362), .CLK(n10549), .Q(
        g147), .QN(n9874) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n10362), .CLK(n10549), .Q(
        g151) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n10363), .CLK(n10550), .Q(
        g152) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n10363), .CLK(n10550), .Q(
        g150), .QN(n9873) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n10363), .CLK(n10550), .Q(
        g154) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n10363), .CLK(n10550), .Q(
        g155) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n10363), .CLK(n10550), .Q(
        g153), .QN(n9872) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n10359), .CLK(n10546), .Q(
        g157) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n10361), .CLK(n10548), .Q(
        g158) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n10361), .CLK(n10548), .Q(
        g156), .QN(n9871) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n10363), .CLK(n10550), .Q(
        g160) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n10363), .CLK(n10550), .Q(
        g161), .QN(n9832) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n10363), .CLK(n10550), .Q(
        g159) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n10363), .CLK(n10550), .Q(
        test_so12) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n10361), .CLK(n10548), 
        .Q(g164), .QN(n9870) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n10361), .CLK(n10548), .Q(
        g162) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n10361), .CLK(n10548), .Q(
        g169) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n10361), .CLK(n10548), .Q(
        g170), .QN(n9934) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n10361), .CLK(n10548), .Q(
        g168) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n10361), .CLK(n10548), .Q(
        g172) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n10362), .CLK(n10549), .Q(
        g173), .QN(n9931) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n10362), .CLK(n10549), .Q(
        g171) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n10362), .CLK(n10549), .Q(
        g175) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n10362), .CLK(n10549), .Q(
        g176), .QN(n9928) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n10362), .CLK(n10549), .Q(
        g174) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n10362), .CLK(n10549), .Q(
        g178) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n10362), .CLK(n10549), .Q(
        g179), .QN(n9925) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n10362), .CLK(n10549), .Q(
        g177) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n10369), .CLK(n10556), .Q(
        g186), .QN(n9523) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n10369), .CLK(n10556), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n10369), .CLK(n10556), 
        .Q(g192), .QN(n9587) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n10369), .CLK(n10556), .Q(
        g231), .QN(n9522) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n10369), .CLK(n10556), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n10369), .CLK(n10556), .Q(
        g237), .QN(n9470) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n10370), .CLK(n10557), .Q(
        g195), .QN(n9521) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n10370), .CLK(n10557), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n10364), .CLK(n10551), .Q(
        g201), .QN(n9586) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n10364), .CLK(n10551), .Q(
        g240), .QN(n9519) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n10364), .CLK(n10551), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n10365), .CLK(n10552), .Q(
        g246), .QN(n9469) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n10365), .CLK(n10552), .Q(
        g204), .QN(n9518) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n10365), .CLK(n10552), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n10365), .CLK(n10552), .Q(
        g210), .QN(n9575) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n10365), .CLK(n10552), .Q(
        g249), .QN(n9516) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n10365), .CLK(n10552), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n10365), .CLK(n10552), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n10365), .CLK(n10552), 
        .Q(g213), .QN(n9514) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n10365), .CLK(n10552), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n10365), .CLK(n10552), .Q(
        g219), .QN(n9585) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n10365), .CLK(n10552), .Q(
        g258), .QN(n9512) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n10365), .CLK(n10552), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n10366), .CLK(n10553), .Q(
        g264), .QN(n9570) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n10366), .CLK(n10553), .Q(
        g222), .QN(n9421) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n10366), .CLK(n10553), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n10366), .CLK(n10553), .Q(
        g228), .QN(n9427) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n10366), .CLK(n10553), .Q(
        g267), .QN(n9456) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n10366), .CLK(n10553), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n10359), .CLK(n10546), .Q(
        g273), .QN(n9457) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n10359), .CLK(n10546), .Q(
        g92), .QN(n10025) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n10359), .CLK(n10546), .Q(
        g88), .QN(n10306) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n10359), .CLK(n10546), .Q(
        g83), .QN(n10024) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n10359), .CLK(n10546), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n10359), .CLK(n10546), 
        .Q(g74), .QN(n10023) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n10359), .CLK(n10546), .Q(
        g70), .QN(n10317) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n10360), .CLK(n10547), .Q(
        g65), .QN(n10022) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n10360), .CLK(n10547), .Q(
        g61), .QN(n10308) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n10360), .CLK(n10547), .Q(
        g56), .QN(n9603) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n10360), .CLK(n10547), .Q(
        g52), .QN(n9432) );
  SDFFX1 DFF_246_Q_reg ( .D(n37), .SI(g52), .SE(n10360), .CLK(n10547), .Q(g180) );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n10360), .CLK(n10547), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n10360), .CLK(n10547), .Q(
        g181), .QN(n10032) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n10360), .CLK(n10547), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n10360), .CLK(n10547), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n10369), .CLK(n10556), .Q(
        g354), .QN(n9976) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n10369), .CLK(n10556), .Q(
        g343) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n10369), .CLK(n10556), .Q(
        test_so16) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n10368), .CLK(n10555), 
        .Q(g369), .QN(n9954) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n10368), .CLK(n10555), .Q(
        g358) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n10368), .CLK(n10555), .Q(
        g361) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n10368), .CLK(n10555), .Q(
        g384), .QN(n9684) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n10369), .CLK(n10556), .Q(
        g373) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n10368), .CLK(n10555), .Q(
        g376) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n10369), .CLK(n10556), .Q(
        g398), .QN(n9965) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n10369), .CLK(n10556), .Q(
        g388) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n10366), .CLK(n10553), .Q(
        g391) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n10366), .CLK(n10553), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n10366), .CLK(n10553), .Q(
        g411), .QN(n9784) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n10367), .CLK(n10554), .Q(
        g414), .QN(n9783) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n10367), .CLK(n10554), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n10367), .CLK(n10554), .Q(
        g420), .QN(n9781) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n10367), .CLK(n10554), .Q(
        g423), .QN(n9780) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n10367), .CLK(n10554), .Q(
        test_so17) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n10367), .CLK(n10554), 
        .Q(g428) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n10367), .CLK(n10554), .Q(
        g426) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n10367), .CLK(n10554), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n10367), .CLK(n10554), .Q(
        g432), .QN(n9778) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n10367), .CLK(n10554), .Q(
        g435), .QN(n9777) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n10368), .CLK(n10555), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n10368), .CLK(n10555), .Q(
        g441), .QN(n9775) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n10368), .CLK(n10555), .Q(
        g444), .QN(n9774) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n10368), .CLK(n10555), .Q(
        g448), .QN(n10006) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n10368), .CLK(n10555), .Q(
        g449), .QN(n10005) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n10367), .CLK(n10554), .Q(
        g447), .QN(n10004) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n10367), .CLK(n10554), .Q(
        g312), .QN(n9567) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n10368), .CLK(n10555), .Q(
        g313) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n10366), .CLK(n10553), .Q(
        g314) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n10366), .CLK(n10553), .Q(
        g315), .QN(n9564) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n10366), .CLK(n10553), .Q(
        test_so18) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n10359), .CLK(n10546), 
        .Q(g317) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n10361), .CLK(n10548), .Q(
        g318), .QN(n9562) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n10361), .CLK(n10548), .Q(
        g319) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n10359), .CLK(n10546), .Q(
        g320) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n10370), .CLK(n10557), .Q(
        g322), .QN(n9599) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n10370), .CLK(n10557), .Q(
        g323) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n10359), .CLK(n10546), .Q(
        g321) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n10360), .CLK(n10547), .Q(
        g403), .QN(n10003) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n10361), .CLK(n10548), .Q(
        g404) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n10361), .CLK(n10548), .Q(
        g402) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n10455), .CLK(n10642), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n10455), .CLK(n10642), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n10455), .CLK(n10642), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n10455), .CLK(n10642), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n10455), .CLK(n10642), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n10455), .CLK(n10642), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n10357), .CLK(n10544), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n10358), .CLK(n10545), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n10358), .CLK(n10545), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n10358), .CLK(n10545), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n10358), .CLK(n10545), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n10358), .CLK(n10545), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n10358), .CLK(n10545), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n10358), .CLK(n10545), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n10358), .CLK(n10545), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n10358), .CLK(n10545), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n10358), .CLK(n10545), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n10358), .CLK(n10545), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n10368), .CLK(n10555), .Q(
        n8056), .QN(n18872) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n10379), .CLK(n10566), 
        .Q(g305), .QN(n9740) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n10370), .CLK(n10557), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n10370), .CLK(n10557), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n10370), .CLK(
        n10557), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n10370), .CLK(n10557), .Q(
        g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n10370), .CLK(n10557), .Q(
        g351), .QN(n9661) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n10370), .CLK(n10557), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n10370), .CLK(n10557), .Q(
        g353), .QN(n9660) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n10370), .CLK(n10557), .Q(
        g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n10371), .CLK(n10558), .Q(
        g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n10371), .CLK(n10558), .Q(
        g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n10371), .CLK(n10558), .Q(
        g366), .QN(n9450) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n10371), .CLK(n10558), .Q(
        g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n10371), .CLK(n10558), .Q(
        g368), .QN(n9449) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n10371), .CLK(n10558), .Q(
        g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n10371), .CLK(n10558), .Q(
        g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n10371), .CLK(n10558), .Q(
        g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n10371), .CLK(n10558), .Q(
        g381), .QN(n9624) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n10371), .CLK(n10558), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n10371), .CLK(
        n10558), .Q(g383), .QN(n9623) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n10371), .CLK(n10558), .Q(
        g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n10372), .CLK(n10559), .Q(
        g394), .QN(n18862) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n10372), .CLK(n10559), .Q(
        g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n10372), .CLK(n10559), .Q(
        g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n10372), .CLK(n10559), .Q(
        g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n10372), .CLK(n10559), .Q(
        g324), .QN(n9673) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n10372), .CLK(n10559), .Q(
        g5629), .QN(n9671) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n10372), .CLK(n10559), .Q(
        g5648), .QN(n9674) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n10372), .CLK(n10559), .Q(
        g337), .QN(n9672) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n10372), .CLK(n10559), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n10372), .CLK(n10559), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n10372), .CLK(n10559), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(n630), .SI(g550), .SE(n10372), .CLK(n10559), .Q(
        g554), .QN(n10267) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n10373), .CLK(n10560), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n10373), .CLK(n10560), .Q(
        test_so22), .QN(n10326) );
  SDFFX1 DFF_362_Q_reg ( .D(n622), .SI(test_si23), .SE(n10373), .CLK(n10560), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n10373), .CLK(n10560), .Q(
        g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n10373), .CLK(n10560), .Q(
        g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n10373), .CLK(n10560), .Q(
        g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n10373), .CLK(n10560), .Q(
        g569), .QN(n9807) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n10373), .CLK(n10560), .Q(
        g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n10373), .CLK(n10560), .Q(
        g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n10373), .CLK(n10560), .Q(
        g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n10373), .CLK(n10560), .Q(
        g573), .QN(n9808) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n10373), .CLK(n10560), .Q(
        g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n10374), .CLK(n10561), .Q(
        g565), .QN(n9805) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n10374), .CLK(n10561), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n10374), .CLK(n10561), .Q(
        g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n10374), .CLK(n10561), .Q(
        g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n10374), .CLK(n10561), .Q(
        g489), .QN(n9806) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n10374), .CLK(n10561), .Q(
        test_so23), .QN(n10328) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n10374), .CLK(
        n10561), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n10374), .CLK(n10561), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n10374), .CLK(n10561), .Q(
        g486), .QN(n10062) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n10374), .CLK(n10561), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n10374), .CLK(n10561), .Q(
        g488), .QN(n10063) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n10375), .CLK(n10562), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n10375), .CLK(n10562), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n10375), .CLK(n10562), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n10375), .CLK(n10562), .Q(
        g477), .QN(n10068) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n10375), .CLK(n10562), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n10375), .CLK(n10562), .Q(
        g479), .QN(n10069) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n10375), .CLK(n10562), .Q(
        g480), .QN(n10065) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n10375), .CLK(n10562), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n10375), .CLK(n10562), .Q(
        g464), .QN(n10066) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n10375), .CLK(n10562), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n10375), .CLK(n10562), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n10374), .CLK(n10561), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n621), .SI(g471), .SE(n10375), .CLK(n10562), .Q(
        g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n10376), .CLK(n10563), .Q(
        g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n10376), .CLK(n10563), .Q(
        g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n10376), .CLK(n10563), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n10376), .CLK(n10563), .Q(
        g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n10376), .CLK(n10563), .Q(
        g548), .QN(n9416) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n10376), .CLK(n10563), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n10376), .CLK(n10563), .Q(
        g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n10376), .CLK(n10563), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n10376), .CLK(n10563), .Q(
        g559) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n10377), .CLK(n10564), .Q(
        g576) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n10377), .CLK(n10564), .Q(
        g577), .QN(n9616) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n10377), .CLK(n10564), .Q(
        g575) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n10377), .CLK(n10564), .Q(
        g579) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n10377), .CLK(n10564), .Q(
        test_so25), .QN(n10333) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n10377), .CLK(n10564), 
        .Q(g578) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n10377), .CLK(n10564), .Q(
        g582) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n10377), .CLK(n10564), .Q(
        g583), .QN(n9442) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n10377), .CLK(n10564), .Q(
        g581) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n10377), .CLK(n10564), .Q(
        g585) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n10377), .CLK(n10564), .Q(
        g586), .QN(n9650) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n10377), .CLK(n10564), .Q(
        g584) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n10378), .CLK(n10565), .Q(
        g587), .QN(n9710) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n10378), .CLK(n10565), .Q(
        g590), .QN(n9712) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n10378), .CLK(n10565), .Q(
        g593), .QN(n9711) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n10378), .CLK(n10565), .Q(
        g596), .QN(n9698) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n10378), .CLK(n10565), .Q(
        g599), .QN(n9700) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n10378), .CLK(n10565), .Q(
        g602), .QN(n9699) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n10378), .CLK(n10565), .Q(
        g614), .QN(n9714) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n10378), .CLK(n10565), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n10376), .CLK(n10563), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n10378), .CLK(n10565), 
        .Q(g605), .QN(n9716) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n10378), .CLK(n10565), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n10378), .CLK(n10565), .Q(
        g611), .QN(n9717) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n10378), .CLK(n10565), .Q(
        g490), .QN(n9787) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n10379), .CLK(n10566), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n10376), .CLK(n10563), .Q(
        g496), .QN(n9791) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n10376), .CLK(n10563), .Q(
        g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n10379), .CLK(n10566), .Q(
        n4571), .QN(n9713) );
  SDFFX1 DFF_442_Q_reg ( .D(n628), .SI(n4571), .SE(n10379), .CLK(n10566), .Q(
        g16297) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n10379), .CLK(n10566), 
        .Q(g525), .QN(n10036) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n10455), .CLK(n10642), 
        .Q(n8047) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n10455), .CLK(n10642), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n10456), .CLK(n10643), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n10456), .CLK(n10643), 
        .Q(n8044) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n10456), .CLK(n10643), 
        .Q(n8043) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n10456), .CLK(n10643), 
        .Q(test_so27) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n10358), .CLK(
        n10545), .Q(g536) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n10359), .CLK(n10546), 
        .Q(g537) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n10379), .CLK(n10566), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n10379), .CLK(n10566), .Q(
        n8040), .QN(n18855) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n10379), .CLK(n10566), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n10379), .CLK(n10566), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n10379), .CLK(n10566), .Q(
        g630), .QN(n10075) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n10379), .CLK(n10566), .Q(
        g659) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n10380), .CLK(n10567), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(n10380), .CLK(n10567), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n10380), .CLK(n10567), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n10380), .CLK(n10567), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n10380), .CLK(n10567), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(n10380), .CLK(n10567), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n10380), .CLK(n10567), .Q(
        test_so28), .QN(n10325) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n10380), .CLK(n10567), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n10380), .CLK(n10567), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n10380), .CLK(n10567), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n10380), .CLK(n10567), .Q(
        g699) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n10380), .CLK(n10567), .Q(
        g700) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n10381), .CLK(n10568), .Q(
        g698), .QN(n10192) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n10381), .CLK(n10568), .Q(
        g702) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n10381), .CLK(n10568), .Q(
        g703) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n10381), .CLK(n10568), .Q(
        g701), .QN(n10191) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n10381), .CLK(n10568), .Q(
        g705) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n10381), .CLK(n10568), .Q(
        g706) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n10381), .CLK(n10568), .Q(
        g704), .QN(n10190) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n10381), .CLK(n10568), .Q(
        g708) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n10381), .CLK(n10568), .Q(
        g709) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n10381), .CLK(n10568), .Q(
        g707), .QN(n10189) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n10381), .CLK(n10568), .Q(
        test_so29), .QN(n10338) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n10381), .CLK(n10568), 
        .Q(g712) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n10382), .CLK(n10569), .Q(
        g710) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n10382), .CLK(n10569), .Q(
        g714) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n10382), .CLK(n10569), .Q(
        g715) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n10382), .CLK(n10569), .Q(
        g713), .QN(n10187) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n10382), .CLK(n10569), .Q(
        g717) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n10383), .CLK(n10570), .Q(
        g718) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n10383), .CLK(n10570), .Q(
        g716), .QN(n10186) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n10383), .CLK(n10570), .Q(
        g720) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n10383), .CLK(n10570), .Q(
        g721) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n10383), .CLK(n10570), .Q(
        g719), .QN(n10185) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n10383), .CLK(n10570), .Q(
        g723) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n10383), .CLK(n10570), .Q(
        g724) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n10383), .CLK(n10570), .Q(
        g722), .QN(n10184) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n10383), .CLK(n10570), .Q(
        g726) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n10383), .CLK(n10570), .Q(
        test_so30) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n10382), .CLK(n10569), 
        .Q(g725) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n10382), .CLK(n10569), .Q(
        g729), .QN(n10297) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n10382), .CLK(n10569), .Q(
        g730) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n10382), .CLK(n10569), .Q(
        g728) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n10382), .CLK(n10569), .Q(
        g732), .QN(n9889) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n10382), .CLK(n10569), .Q(
        g733), .QN(n9884) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n10382), .CLK(n10569), .Q(
        g731) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n10383), .CLK(n10570), .Q(
        g735) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n10383), .CLK(n10570), .Q(
        g736) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n10384), .CLK(n10571), .Q(
        g734) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n10384), .CLK(n10571), .Q(
        g738), .QN(n10196) );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(n10384), .CLK(n10571), .Q(
        g739) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n10384), .CLK(n10571), .Q(
        g737), .QN(n10263) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n10384), .CLK(n10571), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n10384), .CLK(n10571), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n10384), .CLK(n10571), .Q(
        test_so31), .QN(n10321) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n10385), .CLK(n10572), 
        .Q(g818) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n10388), .CLK(n10575), .Q(
        g819) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n10388), .CLK(n10575), .Q(
        g817), .QN(n9868) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n10385), .CLK(n10572), .Q(
        g821) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n10388), .CLK(n10575), .Q(
        g822) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n10388), .CLK(n10575), .Q(
        g820), .QN(n9867) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n10388), .CLK(n10575), .Q(
        g830) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n10388), .CLK(n10575), .Q(
        g831) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n10388), .CLK(n10575), .Q(
        g829), .QN(n9866) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n10389), .CLK(n10576), .Q(
        g833) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n10389), .CLK(n10576), .Q(
        g834) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n10389), .CLK(n10576), .Q(
        g832), .QN(n9865) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n10389), .CLK(n10576), .Q(
        g836) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n10389), .CLK(n10576), .Q(
        g837) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n10389), .CLK(n10576), .Q(
        g835), .QN(n9864) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n10389), .CLK(n10576), .Q(
        test_so32) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n10387), .CLK(n10574), 
        .Q(g840) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n10387), .CLK(n10574), .Q(
        g838), .QN(n9863) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n10387), .CLK(n10574), .Q(
        g842) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n10387), .CLK(n10574), .Q(
        g843) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n10387), .CLK(n10574), .Q(
        g841), .QN(n9862) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n10387), .CLK(n10574), .Q(
        g845) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n10387), .CLK(n10574), .Q(
        g846) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n10387), .CLK(n10574), .Q(
        g844), .QN(n9861) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n10387), .CLK(n10574), .Q(
        g848) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n10387), .CLK(n10574), .Q(
        g849) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n10387), .CLK(n10574), .Q(
        g847), .QN(n9858) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n10388), .CLK(n10575), .Q(
        g851) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n10388), .CLK(n10575), .Q(
        g852) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n10388), .CLK(n10575), .Q(
        g850), .QN(n9855) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n10388), .CLK(n10575), .Q(
        g857) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n10388), .CLK(n10575), .Q(
        test_so33) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n10384), .CLK(n10571), 
        .Q(g856), .QN(n9922) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n10384), .CLK(n10571), .Q(
        g860) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n10384), .CLK(n10571), .Q(
        g861) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n10384), .CLK(n10571), .Q(
        g859), .QN(n9919) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n10384), .CLK(n10571), .Q(
        g863) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n10385), .CLK(n10572), .Q(
        g864) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n10385), .CLK(n10572), .Q(
        g862), .QN(n9916) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n10385), .CLK(n10572), .Q(
        g866) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n10385), .CLK(n10572), .Q(
        g867) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n10385), .CLK(n10572), .Q(
        g865), .QN(n9913) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n10391), .CLK(n10578), .Q(
        g873), .QN(n9510) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n10391), .CLK(n10578), .Q(
        g876), .QN(n9509) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n10391), .CLK(n10578), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n10391), .CLK(n10578), .Q(
        g918), .QN(n9508) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n10391), .CLK(n10578), .Q(
        g921), .QN(n9529) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n10392), .CLK(n10579), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n10389), .CLK(n10576), 
        .Q(g882), .QN(n9507) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n10389), .CLK(n10576), .Q(
        g885), .QN(n9506) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n10389), .CLK(n10576), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n10389), .CLK(n10576), .Q(
        g927), .QN(n9505) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n10389), .CLK(n10576), .Q(
        g930), .QN(n9528) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n10390), .CLK(n10577), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n10390), .CLK(n10577), .Q(
        g891), .QN(n9504) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n10390), .CLK(n10577), .Q(
        g894), .QN(n9503) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n10390), .CLK(n10577), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n10390), .CLK(n10577), .Q(
        g936), .QN(n9502) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n10390), .CLK(n10577), .Q(
        g939), .QN(n9501) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n10390), .CLK(n10577), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n10390), .CLK(n10577), .Q(
        g900), .QN(n9500) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n10390), .CLK(n10577), .Q(
        g903), .QN(n9499) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n10390), .CLK(n10577), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n10394), .CLK(n10581), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n10395), .CLK(n10582), 
        .Q(g948), .QN(n9498) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n10395), .CLK(n10582), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n10395), .CLK(n10582), .Q(
        g909), .QN(n9497) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n10395), .CLK(n10582), .Q(
        g912), .QN(n9533) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n10390), .CLK(n10577), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n10390), .CLK(n10577), .Q(
        g954), .QN(n9496) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n10391), .CLK(n10578), .Q(
        g957), .QN(n9532) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n10385), .CLK(n10572), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n10385), .CLK(n10572), .Q(
        g780), .QN(n10021) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n10385), .CLK(n10572), .Q(
        g776), .QN(n10314) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n10385), .CLK(n10572), .Q(
        g771), .QN(n10020) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n10385), .CLK(n10572), .Q(
        g767), .QN(n10315) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n10386), .CLK(n10573), .Q(
        g762), .QN(n10019) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n10386), .CLK(n10573), .Q(
        g758), .QN(n10316) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n10386), .CLK(n10573), .Q(
        g753), .QN(n10018) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n10386), .CLK(n10573), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n10386), .CLK(n10573), 
        .Q(g744), .QN(n9602) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n10386), .CLK(n10573), .Q(
        g740), .QN(n9431) );
  SDFFX1 DFF_596_Q_reg ( .D(n37), .SI(g740), .SE(n10386), .CLK(n10573), .Q(
        g868) );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n10386), .CLK(n10573), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n10386), .CLK(n10573), .Q(
        g869), .QN(n10031) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n10386), .CLK(n10573), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n10386), .CLK(n10573), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n10386), .CLK(n10573), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n10387), .CLK(n10574), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n10394), .CLK(n10581), .Q(
        g1041) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n10394), .CLK(n10581), 
        .Q(g1030) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n10394), .CLK(n10581), 
        .Q(g1033), .QN(n9972) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n10394), .CLK(n10581), 
        .Q(g1056) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n10394), .CLK(n10581), 
        .Q(g1045) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n10394), .CLK(n10581), 
        .Q(g1048), .QN(n9949) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n10394), .CLK(n10581), 
        .Q(test_so37) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n10394), .CLK(n10581), 
        .Q(g1060) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n10394), .CLK(n10581), 
        .Q(g1063), .QN(n9683) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n10394), .CLK(n10581), 
        .Q(g1085) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n10394), .CLK(n10581), 
        .Q(g1075) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n10392), .CLK(n10579), 
        .Q(g1078), .QN(n9960) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n10392), .CLK(n10579), 
        .Q(g1095), .QN(n9773) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n10393), .CLK(n10580), 
        .Q(g1098), .QN(n9751) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n10393), .CLK(n10580), 
        .Q(g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n10393), .CLK(n10580), 
        .Q(g1104), .QN(n9771) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n10393), .CLK(n10580), 
        .Q(g1107), .QN(n9750) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n10392), .CLK(n10579), 
        .Q(g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n10392), .CLK(n10579), 
        .Q(g1114) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n10392), .CLK(n10579), 
        .Q(g1115) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n10392), .CLK(n10579), 
        .Q(g1113), .QN(n9999) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n10392), .CLK(n10579), 
        .Q(g1116), .QN(n9769) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n10392), .CLK(n10579), 
        .Q(test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n10392), .CLK(n10579), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n10393), .CLK(n10580), 
        .Q(g1125), .QN(n9767) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n10393), .CLK(n10580), 
        .Q(g1128), .QN(n9749) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n10393), .CLK(n10580), 
        .Q(g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n10393), .CLK(n10580), 
        .Q(g1135), .QN(n9998) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n10393), .CLK(n10580), 
        .Q(g1136), .QN(n9984) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n10392), .CLK(n10579), 
        .Q(g1134), .QN(n9997) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n10393), .CLK(n10580), 
        .Q(g999) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n10393), .CLK(n10580), .Q(
        g1000) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n10392), .CLK(n10579), 
        .Q(g1001), .QN(n9558) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n10391), .CLK(n10578), 
        .Q(g1002) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n10391), .CLK(n10578), 
        .Q(g1003) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n10391), .CLK(n10578), 
        .Q(g1004), .QN(n9556) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n10391), .CLK(n10578), 
        .Q(g1005) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n10391), .CLK(n10578), 
        .Q(g1006) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n10391), .CLK(n10578), 
        .Q(test_so39), .QN(n10339) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n10395), .CLK(n10582), 
        .Q(g1009) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n10395), .CLK(n10582), 
        .Q(g1010) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n10395), .CLK(n10582), 
        .Q(g1008), .QN(n9595) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n10395), .CLK(n10582), 
        .Q(g1090) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n10395), .CLK(n10582), 
        .Q(g1091) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n10395), .CLK(n10582), 
        .Q(g1089), .QN(n9995) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n10395), .CLK(n10582), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n10395), .CLK(n10582), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n10396), .CLK(n10583), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n10396), .CLK(n10583), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n10396), .CLK(n10583), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n10396), .CLK(n10583), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n10396), .CLK(n10583), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n10396), .CLK(n10583), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n10396), .CLK(n10583), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n10396), .CLK(n10583), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n10352), .CLK(n10539), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n10353), .CLK(n10540), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n10353), .CLK(n10540), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n10353), .CLK(n10540), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n10353), .CLK(n10540), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n10353), .CLK(n10540), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n10353), .CLK(n10540), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n10353), .CLK(n10540), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n10393), .CLK(n10580), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n529), .SI(g986), .SE(n10396), .CLK(n10583), .Q(
        g992), .QN(n10028) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n10396), .CLK(n10583), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n10396), .CLK(n10583), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n10396), .CLK(n10583), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n10397), .CLK(n10584), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n10397), .CLK(n10584), .Q(
        g1038), .QN(n9659) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n10397), .CLK(n10584), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n10397), .CLK(
        n10584), .Q(g1040), .QN(n9658) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n10397), .CLK(n10584), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n10397), .CLK(n10584), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n10397), .CLK(n10584), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n10397), .CLK(n10584), .Q(
        g1053), .QN(n9448) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n10397), .CLK(n10584), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n10397), .CLK(n10584), .Q(
        g1055), .QN(n9447) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n10397), .CLK(n10584), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n10397), .CLK(n10584), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n10398), .CLK(n10585), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n10398), .CLK(n10585), .Q(
        g1068), .QN(n9622) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n10398), .CLK(n10585), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n10398), .CLK(n10585), .Q(
        g1070), .QN(n9621) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n10398), .CLK(n10585), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n10398), .CLK(n10585), .Q(
        g1081), .QN(n18861) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n10398), .CLK(n10585), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n10398), .CLK(
        n10585), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n10398), .CLK(n10585), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n10398), .CLK(n10585), .Q(
        g1011), .QN(n9668) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n10398), .CLK(n10585), .Q(
        g5657), .QN(n9666) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n10398), .CLK(n10585), .Q(
        g5686), .QN(n9669) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n10399), .CLK(n10586), .Q(
        g1024), .QN(n9667) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n10399), .CLK(n10586), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n10399), .CLK(n10586), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n10399), .CLK(n10586), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(n987), .SI(g1236), .SE(n10399), .CLK(n10586), .Q(
        g1240), .QN(n10266) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n10399), .CLK(n10586), 
        .Q(g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n10399), .CLK(n10586), 
        .Q(g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n982), .SI(g1196), .SE(n10400), .CLK(n10587), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n10400), .CLK(n10587), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n10400), .CLK(n10587), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n10400), .CLK(n10587), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n10400), .CLK(
        n10587), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n10401), .CLK(n10588), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n10401), .CLK(n10588), .Q(
        g1257), .QN(n18865) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n10401), .CLK(n10588), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n10401), .CLK(n10588), .Q(
        g1259), .QN(n9820) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n10401), .CLK(n10588), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n10401), .CLK(n10588), .Q(
        g1251), .QN(n9817) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n10401), .CLK(n10588), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n10401), .CLK(n10588), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n10401), .CLK(n10588), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n10401), .CLK(n10588), .Q(
        g1176), .QN(n9818) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n10401), .CLK(n10588), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n10401), .CLK(n10588), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n10402), .CLK(n10589), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n10402), .CLK(n10589), 
        .Q(g1173), .QN(n10054) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n10402), .CLK(n10589), 
        .Q(test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n10402), .CLK(n10589), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n10402), .CLK(n10589), 
        .Q(g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n10402), .CLK(n10589), 
        .Q(g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n10402), .CLK(n10589), 
        .Q(g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n10402), .CLK(n10589), 
        .Q(g1164), .QN(n10059) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n10402), .CLK(n10589), 
        .Q(g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n10402), .CLK(n10589), 
        .Q(g1166), .QN(n10060) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n10402), .CLK(n10589), 
        .Q(g1167), .QN(n10056) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n10402), .CLK(n10589), 
        .Q(g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n10403), .CLK(n10590), 
        .Q(g1151), .QN(n10057) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n10403), .CLK(n10590), 
        .Q(g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n10403), .CLK(n10590), 
        .Q(g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n10403), .CLK(n10590), 
        .Q(g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n983), .SI(g1158), .SE(n10403), .CLK(n10590), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n10403), .CLK(n10590), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n10403), .CLK(n10590), .Q(
        test_so45), .QN(n9695) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n10403), .CLK(n10590), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n10403), .CLK(n10590), .Q(
        n4549), .QN(n9414) );
  SDFFX1 DFF_750_Q_reg ( .D(n588), .SI(n4549), .SE(n10403), .CLK(n10590), .Q(
        n4361), .QN(n9415) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n10403), .CLK(n10590), 
        .Q(g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n10403), .CLK(n10590), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n10404), .CLK(n10591), 
        .Q(g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n10404), .CLK(n10591), .Q(
        g1245), .QN(n10078) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n10404), .CLK(n10591), 
        .Q(g1262), .QN(n9611) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n10405), .CLK(n10592), 
        .Q(g1263) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n10405), .CLK(n10592), 
        .Q(g1261) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n10405), .CLK(n10592), 
        .Q(g1265), .QN(n9631) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n10405), .CLK(n10592), 
        .Q(g1266) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n10404), .CLK(n10591), 
        .Q(g1264) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n10404), .CLK(n10591), 
        .Q(g1268), .QN(n9438) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n10404), .CLK(n10591), 
        .Q(g1269) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n10404), .CLK(n10591), 
        .Q(test_so46) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n10404), .CLK(n10591), 
        .Q(g1271), .QN(n9645) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n10405), .CLK(n10592), 
        .Q(g1272) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n10405), .CLK(n10592), 
        .Q(g1270) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n10405), .CLK(n10592), 
        .Q(g1273), .QN(n9707) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n10405), .CLK(n10592), 
        .Q(g1276), .QN(n9709) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n10405), .CLK(n10592), 
        .Q(g1279), .QN(n9708) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n10405), .CLK(n10592), 
        .Q(g1282), .QN(n9694) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n10405), .CLK(n10592), 
        .Q(g1285), .QN(n9697) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n10405), .CLK(n10592), 
        .Q(g1288), .QN(n9696) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n10406), .CLK(n10593), 
        .Q(g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n10406), .CLK(n10593), 
        .Q(g1303), .QN(n9727) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n10404), .CLK(n10591), 
        .Q(g1306), .QN(n9726) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n10406), .CLK(n10593), 
        .Q(g1291), .QN(n9733) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n10406), .CLK(n10593), 
        .Q(g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n10406), .CLK(n10593), 
        .Q(g1297), .QN(n9734) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n10406), .CLK(n10593), 
        .Q(test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n10404), .CLK(n10591), 
        .Q(g1180), .QN(n9794) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n10404), .CLK(n10591), 
        .Q(g1183), .QN(n9790) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n10404), .CLK(n10591), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n10406), .CLK(n10593), 
        .Q(n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n627), .SI(n8009), .SE(n10406), .CLK(n10593), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n10406), .CLK(n10593), 
        .Q(g1211), .QN(n10035) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n10407), .CLK(n10594), 
        .Q(n8008) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n10407), .CLK(n10594), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n10407), .CLK(n10594), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n10407), .CLK(n10594), 
        .Q(n8005) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n10407), .CLK(n10594), 
        .Q(n8004) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n10407), .CLK(n10594), 
        .Q(n8003) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n10407), .CLK(n10594), 
        .Q(g1222) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n10407), .CLK(n10594), 
        .Q(g1223) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n10407), .CLK(n10594), 
        .Q(g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n10407), .CLK(n10594), .Q(
        test_so48), .QN(n18858) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n10345), .CLK(n10532), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n10345), .CLK(n10532), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n10399), .CLK(n10586), 
        .Q(g1316), .QN(n10074) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n10399), .CLK(n10586), 
        .Q(g1345) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n10399), .CLK(n10586), 
        .Q(g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(n10399), .CLK(n10586), 
        .Q(g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n10399), .CLK(n10586), 
        .Q(g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n10400), .CLK(n10587), 
        .Q(g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n10400), .CLK(n10587), 
        .Q(g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(n10400), .CLK(n10587), 
        .Q(g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n10400), .CLK(n10587), 
        .Q(g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n10400), .CLK(n10587), 
        .Q(g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n10400), .CLK(n10587), 
        .Q(g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n10400), .CLK(n10587), 
        .Q(g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n10407), .CLK(n10594), 
        .Q(test_so49), .QN(n10337) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n10407), .CLK(n10594), 
        .Q(g1386) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n10408), .CLK(n10595), 
        .Q(g1384) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n10408), .CLK(n10595), 
        .Q(g1388) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n10408), .CLK(n10595), 
        .Q(g1389) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n10408), .CLK(n10595), 
        .Q(g1387), .QN(n10181) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n10408), .CLK(n10595), 
        .Q(g1391) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n10408), .CLK(n10595), 
        .Q(g1392) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n10408), .CLK(n10595), 
        .Q(g1390), .QN(n10180) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n10408), .CLK(n10595), 
        .Q(g1394) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n10408), .CLK(n10595), 
        .Q(g1395) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n10408), .CLK(n10595), 
        .Q(g1393), .QN(n10179) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n10408), .CLK(n10595), 
        .Q(g1397) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n10408), .CLK(n10595), 
        .Q(g1398) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n10409), .CLK(n10596), 
        .Q(g1396), .QN(n10178) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n10409), .CLK(n10596), 
        .Q(g1400) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n10409), .CLK(n10596), 
        .Q(test_so50) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n10409), .CLK(n10596), 
        .Q(g1399) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n10409), .CLK(n10596), 
        .Q(g1403) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n10409), .CLK(n10596), 
        .Q(g1404) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n10409), .CLK(n10596), 
        .Q(g1402), .QN(n10176) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n10409), .CLK(n10596), 
        .Q(g1406) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n10409), .CLK(n10596), 
        .Q(g1407) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n10409), .CLK(n10596), 
        .Q(g1405), .QN(n10175) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n10409), .CLK(n10596), 
        .Q(g1409) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n10409), .CLK(n10596), 
        .Q(g1410) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n10410), .CLK(n10597), 
        .Q(g1408), .QN(n10174) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n10410), .CLK(n10597), 
        .Q(g1412) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n10410), .CLK(n10597), 
        .Q(g1413) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n10410), .CLK(n10597), 
        .Q(g1411), .QN(n10173) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n10410), .CLK(n10597), 
        .Q(g1415), .QN(n10298) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n10410), .CLK(n10597), 
        .Q(g1416) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n10410), .CLK(n10597), 
        .Q(test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n10406), .CLK(n10593), 
        .Q(g1418), .QN(n9888) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n10406), .CLK(n10593), 
        .Q(g1419), .QN(n9882) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n10406), .CLK(n10593), 
        .Q(g1417) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n10410), .CLK(n10597), 
        .Q(g1421) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n10410), .CLK(n10597), 
        .Q(g1422) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n10410), .CLK(n10597), 
        .Q(g1420) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n10410), .CLK(n10597), 
        .Q(g1424), .QN(n10195) );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(n10410), .CLK(n10597), 
        .Q(g1425) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n10411), .CLK(n10598), 
        .Q(g1423), .QN(n10262) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n10411), .CLK(n10598), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n10411), .CLK(n10598), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n10411), .CLK(n10598), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n10411), .CLK(n10598), 
        .Q(g1512) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n10415), .CLK(n10602), 
        .Q(g1513) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n10416), .CLK(n10603), 
        .Q(g1511), .QN(n9854) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n10411), .CLK(n10598), 
        .Q(test_so52) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n10416), .CLK(n10603), 
        .Q(g1516) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n10416), .CLK(n10603), 
        .Q(g1514), .QN(n9853) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n10417), .CLK(n10604), 
        .Q(g1524) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n10417), .CLK(n10604), 
        .Q(g1525) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n10417), .CLK(n10604), 
        .Q(g1523), .QN(n9852) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n10417), .CLK(n10604), 
        .Q(g1527) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n10417), .CLK(n10604), 
        .Q(g1528) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n10417), .CLK(n10604), 
        .Q(g1526), .QN(n9851) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n10417), .CLK(n10604), 
        .Q(g1530) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n10417), .CLK(n10604), 
        .Q(g1531) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n10417), .CLK(n10604), 
        .Q(g1529), .QN(n9850) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n10417), .CLK(n10604), 
        .Q(g1533) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n10417), .CLK(n10604), 
        .Q(g1534) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n10417), .CLK(n10604), 
        .Q(g1532), .QN(n9849) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n10418), .CLK(n10605), 
        .Q(g1536) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n10418), .CLK(n10605), 
        .Q(test_so53) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n10415), .CLK(n10602), 
        .Q(g1535) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n10415), .CLK(n10602), 
        .Q(g1539) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n10415), .CLK(n10602), 
        .Q(g1540) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n10415), .CLK(n10602), 
        .Q(g1538), .QN(n9847) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n10415), .CLK(n10602), 
        .Q(g1542) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n10415), .CLK(n10602), 
        .Q(g1543), .QN(n9829) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n10415), .CLK(n10602), 
        .Q(g1541) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n10416), .CLK(n10603), 
        .Q(g1545) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n10416), .CLK(n10603), 
        .Q(g1546), .QN(n9845) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n10416), .CLK(n10603), 
        .Q(g1544) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n10416), .CLK(n10603), 
        .Q(g1551) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n10416), .CLK(n10603), 
        .Q(g1552), .QN(n9911) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n10416), .CLK(n10603), 
        .Q(g1550) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n10416), .CLK(n10603), 
        .Q(g1554) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n10416), .CLK(n10603), 
        .Q(g1555), .QN(n9908) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n10416), .CLK(n10603), 
        .Q(test_so54) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n10411), .CLK(n10598), 
        .Q(g1557) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n10411), .CLK(n10598), 
        .Q(g1558), .QN(n9906) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n10411), .CLK(n10598), 
        .Q(g1556) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n10411), .CLK(n10598), 
        .Q(g1560) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n10411), .CLK(n10598), 
        .Q(g1561), .QN(n9903) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n10411), .CLK(n10598), 
        .Q(g1559) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n10422), .CLK(n10609), 
        .Q(g1567), .QN(n9495) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n10422), .CLK(n10609), 
        .Q(g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n10422), .CLK(n10609), 
        .Q(g1573), .QN(n9581) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n10422), .CLK(n10609), 
        .Q(g1612), .QN(n9493) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n10422), .CLK(n10609), 
        .Q(g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n10422), .CLK(n10609), 
        .Q(g1618), .QN(n9464) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n10422), .CLK(n10609), 
        .Q(g1576), .QN(n9492) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n10423), .CLK(n10610), 
        .Q(g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n10423), .CLK(n10610), 
        .Q(g1582), .QN(n9580) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n10423), .CLK(n10610), 
        .Q(test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n10423), .CLK(n10610), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n10423), .CLK(n10610), 
        .Q(g1627), .QN(n9463) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n10423), .CLK(n10610), 
        .Q(g1585), .QN(n9490) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n10423), .CLK(n10610), 
        .Q(g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n10418), .CLK(n10605), 
        .Q(g1591), .QN(n9572) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n10418), .CLK(n10605), 
        .Q(g1630), .QN(n9488) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n10418), .CLK(n10605), 
        .Q(g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n10418), .CLK(n10605), 
        .Q(g1636), .QN(n9462) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n10418), .CLK(n10605), 
        .Q(g1594), .QN(n9486) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n10418), .CLK(n10605), 
        .Q(g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n10418), .CLK(n10605), 
        .Q(g1600), .QN(n9579) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n10418), .CLK(n10605), 
        .Q(g1639), .QN(n9484) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n10418), .CLK(n10605), 
        .Q(g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n10418), .CLK(n10605), 
        .Q(g1645), .QN(n9569) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n10419), .CLK(n10606), 
        .Q(g1603), .QN(n9420) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n10419), .CLK(n10606), 
        .Q(test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n10419), .CLK(n10606), 
        .Q(g1609), .QN(n9426) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n10419), .CLK(n10606), 
        .Q(g1648), .QN(n9453) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n10419), .CLK(n10606), 
        .Q(g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n10412), .CLK(n10599), 
        .Q(g1654), .QN(n9454) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n10412), .CLK(n10599), 
        .Q(g1466), .QN(n10017) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n10412), .CLK(n10599), 
        .Q(g1462), .QN(n10307) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n10412), .CLK(n10599), 
        .Q(g1457), .QN(n10016) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n10412), .CLK(n10599), 
        .Q(g1453), .QN(n10312) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n10412), .CLK(n10599), 
        .Q(g1448), .QN(n10015) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n10412), .CLK(n10599), 
        .Q(g1444), .QN(n10318) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n10412), .CLK(n10599), 
        .Q(g1439), .QN(n10014) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n10412), .CLK(n10599), 
        .Q(g1435), .QN(n10309) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n10413), .CLK(n10600), 
        .Q(g1430), .QN(n9601) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n10413), .CLK(n10600), 
        .Q(g1426), .QN(n9430) );
  SDFFX1 DFF_946_Q_reg ( .D(n37), .SI(g1426), .SE(n10413), .CLK(n10600), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n10413), .CLK(n10600), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n10413), .CLK(
        n10600), .Q(g1563), .QN(n10030) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n10413), .CLK(n10600), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n10413), .CLK(n10600), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n10421), .CLK(n10608), 
        .Q(g1735) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n10421), .CLK(n10608), 
        .Q(g1724), .QN(n9970) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n10422), .CLK(n10609), 
        .Q(g1727) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n10422), .CLK(n10609), 
        .Q(g1750) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n10422), .CLK(n10609), 
        .Q(g1739), .QN(n9947) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n10421), .CLK(n10608), 
        .Q(g1742) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n10421), .CLK(n10608), 
        .Q(g1765) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n10421), .CLK(n10608), 
        .Q(g1754), .QN(n9681) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n10421), .CLK(n10608), 
        .Q(g1757) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n10422), .CLK(n10609), 
        .Q(g1779) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n10422), .CLK(n10609), 
        .Q(test_so58), .QN(n10331) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n10419), .CLK(n10606), 
        .Q(g1772) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n10419), .CLK(n10606), 
        .Q(g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n10421), .CLK(n10608), 
        .Q(g1792), .QN(n9748) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n10421), .CLK(n10608), 
        .Q(g1795), .QN(n9764) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n10421), .CLK(n10608), 
        .Q(g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n10421), .CLK(n10608), 
        .Q(g1801), .QN(n9747) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n10419), .CLK(n10606), 
        .Q(g1804), .QN(n9762) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n10419), .CLK(n10606), 
        .Q(g1808) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n10420), .CLK(n10607), 
        .Q(g1809), .QN(n9982) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n10420), .CLK(n10607), 
        .Q(g1807) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n10420), .CLK(n10607), 
        .Q(g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n10420), .CLK(n10607), 
        .Q(g1813), .QN(n9746) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n10420), .CLK(n10607), 
        .Q(g1816), .QN(n9760) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n10420), .CLK(n10607), 
        .Q(g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n10420), .CLK(n10607), 
        .Q(g1822), .QN(n9745) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n10421), .CLK(n10608), 
        .Q(test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n10420), .CLK(n10607), 
        .Q(g1829), .QN(n9992) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n10420), .CLK(n10607), 
        .Q(g1830), .QN(n9981) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n10420), .CLK(n10607), 
        .Q(g1828), .QN(n9991) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n10420), .CLK(n10607), 
        .Q(g1693) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n10420), .CLK(n10607), 
        .Q(g1694), .QN(n9539) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n10419), .CLK(n10606), 
        .Q(g1695) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n10419), .CLK(n10606), 
        .Q(g1696) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n10419), .CLK(n10606), 
        .Q(g1697), .QN(n9538) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n10412), .CLK(n10599), 
        .Q(g1698) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n10413), .CLK(n10600), 
        .Q(g1699) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n10412), .CLK(n10599), 
        .Q(g1700), .QN(n9537) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n10413), .CLK(n10600), 
        .Q(g1701) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n10423), .CLK(n10610), 
        .Q(g1703) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n10423), .CLK(n10610), 
        .Q(g1704), .QN(n9589) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n10412), .CLK(n10599), 
        .Q(g1702) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n10413), .CLK(n10600), 
        .Q(test_so60) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n10414), .CLK(n10601), 
        .Q(g1785), .QN(n9980) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n10414), .CLK(n10601), 
        .Q(g1783) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n10414), .CLK(n10601), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n10414), .CLK(n10601), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n10414), .CLK(n10601), 
        .Q(g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n10414), .CLK(n10601), 
        .Q(n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n10414), .CLK(n10601), 
        .Q(g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n10414), .CLK(n10601), 
        .Q(n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n10414), .CLK(n10601), 
        .Q(g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n10414), .CLK(n10601), 
        .Q(n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n10414), .CLK(n10601), 
        .Q(g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n10414), .CLK(n10601), 
        .Q(n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n10415), .CLK(n10602), 
        .Q(g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n10415), .CLK(n10602), 
        .Q(n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n10415), .CLK(n10602), 
        .Q(g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n10415), .CLK(n10602), 
        .Q(test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n10342), .CLK(n10529), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n10342), .CLK(n10529), 
        .Q(n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n10351), .CLK(n10538), 
        .Q(g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n10351), .CLK(n10538), 
        .Q(n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n10421), .CLK(n10608), 
        .Q(g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n530), .SI(g1680), .SE(n10423), .CLK(n10610), .Q(
        g1686), .QN(n10027) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n10423), .CLK(n10610), 
        .Q(n7978) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n10423), .CLK(n10610), 
        .Q(g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n10424), .CLK(n10611), 
        .Q(g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n10424), .CLK(n10611), 
        .Q(g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n10424), .CLK(n10611), 
        .Q(g1732), .QN(n9657) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n10424), .CLK(n10611), 
        .Q(g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n10424), .CLK(n10611), 
        .Q(g1734), .QN(n9656) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n10424), .CLK(n10611), 
        .Q(g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n10424), .CLK(n10611), 
        .Q(g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n10424), .CLK(n10611), 
        .Q(test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n10424), .CLK(
        n10611), .Q(g1747), .QN(n9446) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n10424), .CLK(n10611), 
        .Q(g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n10424), .CLK(n10611), 
        .Q(g1749), .QN(n9445) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n10424), .CLK(n10611), 
        .Q(g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n10425), .CLK(n10612), 
        .Q(g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n10425), .CLK(n10612), 
        .Q(g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n10425), .CLK(n10612), 
        .Q(g1762), .QN(n9620) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n10425), .CLK(n10612), 
        .Q(g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n10425), .CLK(n10612), 
        .Q(g1764), .QN(n9619) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n10425), .CLK(n10612), 
        .Q(g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n10425), .CLK(n10612), 
        .Q(g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n10425), .CLK(n10612), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n10425), .CLK(n10612), 
        .Q(g1777), .QN(n9665) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n10425), .CLK(n10612), 
        .Q(g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n10425), .CLK(n10612), 
        .Q(g1705), .QN(n9663) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n10425), .CLK(n10612), 
        .Q(test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n10426), .CLK(
        n10613), .Q(g5738), .QN(n9664) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n10426), .CLK(n10613), 
        .Q(g1718), .QN(n9662) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n10426), .CLK(n10613), 
        .Q(g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n10426), .CLK(n10613), 
        .Q(g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n10426), .CLK(n10613), 
        .Q(g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(n1335), .SI(g1930), .SE(n10426), .CLK(n10613), 
        .Q(g1934), .QN(n10265) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n10426), .CLK(n10613), 
        .Q(g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n10426), .CLK(n10613), 
        .Q(g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1333), .SI(g1890), .SE(n10427), .CLK(n10614), 
        .Q(g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n10427), .CLK(n10614), 
        .Q(g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n10427), .CLK(n10614), 
        .Q(g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n10427), .CLK(n10614), 
        .Q(g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n10428), .CLK(n10615), 
        .Q(g1949), .QN(n9815) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n10428), .CLK(n10615), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n10428), .CLK(n10615), 
        .Q(g1951), .QN(n18864) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n10428), .CLK(n10615), 
        .Q(test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n10428), .CLK(
        n10615), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n10428), .CLK(n10615), 
        .Q(g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n10428), .CLK(n10615), 
        .Q(g1945), .QN(n9813) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n10428), .CLK(n10615), 
        .Q(g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n10428), .CLK(n10615), 
        .Q(g1947), .QN(n18866) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n10428), .CLK(n10615), 
        .Q(g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n10428), .CLK(n10615), 
        .Q(g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n10428), .CLK(n10615), 
        .Q(g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n10429), .CLK(n10616), 
        .Q(g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n10429), .CLK(n10616), 
        .Q(g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n10429), .CLK(n10616), 
        .Q(g1867), .QN(n10045) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n10429), .CLK(n10616), 
        .Q(g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n10429), .CLK(n10616), 
        .Q(g1869), .QN(n10046) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n10429), .CLK(n10616), 
        .Q(g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n10429), .CLK(n10616), 
        .Q(test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n10429), .CLK(n10616), .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n10429), .CLK(n10616), 
        .Q(g1858), .QN(n10051) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n10429), .CLK(n10616), 
        .Q(g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n10429), .CLK(n10616), 
        .Q(g1860), .QN(n10052) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n10429), .CLK(n10616), 
        .Q(g1861), .QN(n10048) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n10430), .CLK(n10617), 
        .Q(g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n10430), .CLK(n10617), 
        .Q(g1845), .QN(n10049) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n10430), .CLK(n10617), 
        .Q(g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n10430), .CLK(n10617), 
        .Q(g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n10430), .CLK(n10617), 
        .Q(g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1330), .SI(g1852), .SE(n10430), .CLK(n10617), 
        .Q(g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n10430), .CLK(n10617), 
        .Q(g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n10430), .CLK(n10617), 
        .Q(g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n10430), .CLK(n10617), 
        .Q(g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n10430), .CLK(n10617), 
        .Q(test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n618), .SI(test_si67), .SE(n10430), .CLK(n10617), 
        .Q(n7971), .QN(DFF_1100_n1) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n10430), .CLK(n10617), 
        .Q(g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n10431), .CLK(n10618), 
        .Q(g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n10431), .CLK(n10618), 
        .Q(g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n10431), .CLK(n10618), 
        .Q(g1939), .QN(n10077) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n10432), .CLK(n10619), 
        .Q(g1956) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n10432), .CLK(n10619), 
        .Q(g1957) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n10432), .CLK(n10619), 
        .Q(g1955), .QN(n9609) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n10432), .CLK(n10619), 
        .Q(g1959) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n10432), .CLK(n10619), 
        .Q(g1960) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n10431), .CLK(n10618), 
        .Q(g1958), .QN(n9629) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n10431), .CLK(n10618), 
        .Q(g1962) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n10431), .CLK(n10618), 
        .Q(g1963) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n10431), .CLK(n10618), 
        .Q(g1961), .QN(n9436) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n10431), .CLK(n10618), 
        .Q(test_so67) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n10432), .CLK(n10619), .Q(g1966) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n10432), .CLK(n10619), 
        .Q(g1964), .QN(n9643) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n10432), .CLK(n10619), 
        .Q(g1967), .QN(n9704) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n10432), .CLK(n10619), 
        .Q(g1970), .QN(n9706) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n10432), .CLK(n10619), 
        .Q(g1973), .QN(n9705) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n10432), .CLK(n10619), 
        .Q(g1976), .QN(n9691) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n10432), .CLK(n10619), 
        .Q(g1979), .QN(n9693) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n10433), .CLK(n10620), 
        .Q(g1982), .QN(n9692) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n10433), .CLK(n10620), 
        .Q(g1994), .QN(n9722) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n10433), .CLK(n10620), 
        .Q(g1997), .QN(n9724) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n10431), .CLK(n10618), 
        .Q(g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n10433), .CLK(n10620), 
        .Q(g1985), .QN(n9730) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n10433), .CLK(n10620), 
        .Q(g1988), .QN(n9732) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n10433), .CLK(n10620), 
        .Q(g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n10433), .CLK(n10620), 
        .Q(test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n10431), .CLK(n10618), .Q(g1874), .QN(n9793) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n10431), .CLK(n10618), 
        .Q(g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n10431), .CLK(n10618), 
        .Q(g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n10433), .CLK(n10620), 
        .Q(n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n626), .SI(n7968), .SE(n10433), .CLK(n10620), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n10433), .CLK(n10620), 
        .Q(g1905), .QN(n10034) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n10433), .CLK(n10620), .Q(n7967) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n10433), .CLK(
        n10620), .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n10434), .CLK(
        n10621), .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n10434), .CLK(
        n10621), .Q(n7964) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n10434), .CLK(
        n10621), .Q(n7963) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n10434), .CLK(
        n10621), .Q(n7962) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n10434), .CLK(
        n10621), .Q(g1916) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n10434), .CLK(
        n10621), .Q(g1917) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n10434), .CLK(n10621), 
        .Q(test_so69) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n10351), .CLK(n10538), 
        .Q(n7960), .QN(n18857) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n10351), .CLK(n10538), 
        .Q(g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n10351), .CLK(n10538), 
        .Q(g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n10426), .CLK(n10613), 
        .Q(g2010), .QN(n10073) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n10426), .CLK(n10613), 
        .Q(g2039) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n10426), .CLK(n10613), 
        .Q(g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(n10426), .CLK(n10613), 
        .Q(g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n10427), .CLK(n10614), 
        .Q(g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n10427), .CLK(n10614), 
        .Q(g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n10427), .CLK(n10614), 
        .Q(g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(n10427), .CLK(n10614), 
        .Q(g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n10427), .CLK(n10614), 
        .Q(g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n10427), .CLK(n10614), 
        .Q(g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n10427), .CLK(n10614), 
        .Q(test_so70), .QN(n10323) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n10427), .CLK(n10614), .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n10435), .CLK(n10622), 
        .Q(g2079) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n10435), .CLK(n10622), 
        .Q(g2080) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n10435), .CLK(n10622), 
        .Q(g2078), .QN(n10172) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n10435), .CLK(n10622), 
        .Q(g2082) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n10435), .CLK(n10622), 
        .Q(g2083) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n10435), .CLK(n10622), 
        .Q(g2081), .QN(n10171) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n10435), .CLK(n10622), 
        .Q(g2085) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n10435), .CLK(n10622), 
        .Q(g2086) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n10436), .CLK(n10623), 
        .Q(g2084), .QN(n10170) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n10436), .CLK(n10623), 
        .Q(g2088) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n10436), .CLK(n10623), 
        .Q(g2089) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n10436), .CLK(n10623), 
        .Q(g2087), .QN(n10169) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n10436), .CLK(n10623), 
        .Q(g2091) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n10436), .CLK(n10623), 
        .Q(test_so71) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n10435), .CLK(n10622), .Q(g2090) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n10435), .CLK(n10622), 
        .Q(g2094) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n10436), .CLK(n10623), 
        .Q(g2095) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n10436), .CLK(n10623), 
        .Q(g2093), .QN(n10167) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n10436), .CLK(n10623), 
        .Q(g2097) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n10436), .CLK(n10623), 
        .Q(g2098) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n10436), .CLK(n10623), 
        .Q(g2096), .QN(n10166) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n10436), .CLK(n10623), 
        .Q(g2100) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n10437), .CLK(n10624), 
        .Q(g2101) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n10437), .CLK(n10624), 
        .Q(g2099), .QN(n10165) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n10437), .CLK(n10624), 
        .Q(g2103) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n10437), .CLK(n10624), 
        .Q(g2104) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n10437), .CLK(n10624), 
        .Q(g2102), .QN(n10164) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n10437), .CLK(n10624), 
        .Q(g2106) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n10437), .CLK(n10624), 
        .Q(test_so72), .QN(n10336) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n10434), .CLK(n10621), .Q(g2105) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n10434), .CLK(n10621), 
        .Q(g2109), .QN(n10299) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n10434), .CLK(n10621), 
        .Q(g2110) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n10434), .CLK(n10621), 
        .Q(g2108) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n10434), .CLK(n10621), 
        .Q(g2112), .QN(n9887) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n10435), .CLK(n10622), 
        .Q(g2113), .QN(n9880) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n10435), .CLK(n10622), 
        .Q(g2111) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n10437), .CLK(n10624), 
        .Q(g2115) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n10437), .CLK(n10624), 
        .Q(g2116) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n10437), .CLK(n10624), 
        .Q(g2114) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n10437), .CLK(n10624), 
        .Q(g2118), .QN(n10194) );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(n10437), .CLK(n10624), 
        .Q(g2119) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n10438), .CLK(n10625), 
        .Q(g2117), .QN(n10261) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n10438), .CLK(n10625), 
        .Q(g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n10438), .CLK(n10625), 
        .Q(test_so73), .QN(n10320) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n10438), .CLK(
        n10625), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n10438), .CLK(n10625), 
        .Q(g2206) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n10438), .CLK(n10625), 
        .Q(g2207) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n10439), .CLK(n10626), 
        .Q(g2205), .QN(n9843) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n10344), .CLK(n10531), 
        .Q(g2209) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n10438), .CLK(n10625), 
        .Q(g2210) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n10439), .CLK(n10626), 
        .Q(g2208), .QN(n9842) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n10439), .CLK(n10626), 
        .Q(g2218) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n10439), .CLK(n10626), 
        .Q(g2219) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n10439), .CLK(n10626), 
        .Q(g2217), .QN(n9841) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n10439), .CLK(n10626), 
        .Q(g2221) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n10439), .CLK(n10626), 
        .Q(g2222) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n10440), .CLK(n10627), 
        .Q(g2220), .QN(n9840) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n10440), .CLK(n10627), 
        .Q(g2224) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n10440), .CLK(n10627), 
        .Q(test_so74) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n10438), .CLK(n10625), .Q(g2223) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n10438), .CLK(n10625), 
        .Q(g2227) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n10438), .CLK(n10625), 
        .Q(g2228) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n10438), .CLK(n10625), 
        .Q(g2226), .QN(n9838) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n10438), .CLK(n10625), 
        .Q(g2230) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n10439), .CLK(n10626), 
        .Q(g2231) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n10439), .CLK(n10626), 
        .Q(g2229), .QN(n9837) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n10439), .CLK(n10626), 
        .Q(g2233) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n10439), .CLK(n10626), 
        .Q(g2234) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n10439), .CLK(n10626), 
        .Q(g2232), .QN(n9836) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n10441), .CLK(n10628), 
        .Q(g2236) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n10441), .CLK(n10628), 
        .Q(g2237), .QN(n9826) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n10441), .CLK(n10628), 
        .Q(g2235) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n10441), .CLK(n10628), 
        .Q(g2239) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n10441), .CLK(n10628), 
        .Q(test_so75) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n10440), .CLK(n10627), .Q(g2238) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n10440), .CLK(n10627), 
        .Q(g2245) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n10440), .CLK(n10627), 
        .Q(g2246), .QN(n9900) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n10440), .CLK(n10627), 
        .Q(g2244) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n10440), .CLK(n10627), 
        .Q(g2248) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n10440), .CLK(n10627), 
        .Q(g2249), .QN(n9897) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n10440), .CLK(n10627), 
        .Q(g2247) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n10440), .CLK(n10627), 
        .Q(g2251) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n10440), .CLK(n10627), 
        .Q(g2252), .QN(n9894) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n10441), .CLK(n10628), 
        .Q(g2250) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n10441), .CLK(n10628), 
        .Q(g2254) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n10441), .CLK(n10628), 
        .Q(g2255), .QN(n9891) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n10441), .CLK(n10628), 
        .Q(g2253) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n10452), .CLK(n10639), 
        .Q(g2261), .QN(n9482) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n10452), .CLK(n10639), 
        .Q(test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n10452), .CLK(n10639), .Q(g2267), .QN(n9578) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n10452), .CLK(n10639), 
        .Q(g2306), .QN(n9481) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n10453), .CLK(n10640), 
        .Q(g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n10453), .CLK(n10640), 
        .Q(g2312), .QN(n9461) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n10453), .CLK(n10640), 
        .Q(g2270), .QN(n9480) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n10453), .CLK(n10640), 
        .Q(g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n10453), .CLK(n10640), 
        .Q(g2276), .QN(n9577) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n10453), .CLK(n10640), 
        .Q(g2315), .QN(n9478) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n10453), .CLK(n10640), 
        .Q(g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n10443), .CLK(n10630), 
        .Q(g2321), .QN(n9460) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n10444), .CLK(n10631), 
        .Q(g2279), .QN(n9477) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n10444), .CLK(n10631), 
        .Q(g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n10442), .CLK(n10629), 
        .Q(g2285), .QN(n9571) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n10443), .CLK(n10630), 
        .Q(g2324), .QN(n9475) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n10443), .CLK(n10630), 
        .Q(test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n10443), .CLK(n10630), .Q(g2330), .QN(n9459) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n10443), .CLK(n10630), 
        .Q(g2288), .QN(n9474) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n10443), .CLK(n10630), 
        .Q(g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n10443), .CLK(n10630), 
        .Q(g2294), .QN(n9576) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n10443), .CLK(n10630), 
        .Q(g2333), .QN(n9472) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n10443), .CLK(n10630), 
        .Q(g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n10443), .CLK(n10630), 
        .Q(g2339), .QN(n9568) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n10443), .CLK(n10630), 
        .Q(g2297), .QN(n9419) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n10443), .CLK(n10630), 
        .Q(g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n10441), .CLK(n10628), 
        .Q(g2303), .QN(n9425) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n10441), .CLK(n10628), 
        .Q(g2342), .QN(n9418) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n10441), .CLK(n10628), 
        .Q(g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n10442), .CLK(n10629), 
        .Q(g2348), .QN(n9417) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n10442), .CLK(n10629), 
        .Q(g2160), .QN(n10013) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n10442), .CLK(n10629), 
        .Q(test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n10442), .CLK(n10629), .Q(g2151), .QN(n10012) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n10442), .CLK(n10629), 
        .Q(g2147), .QN(n10313) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n10442), .CLK(n10629), 
        .Q(g2142), .QN(n10011) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n10442), .CLK(n10629), 
        .Q(g2138), .QN(n10319) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n10442), .CLK(n10629), 
        .Q(g2133), .QN(n10010) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n10442), .CLK(n10629), 
        .Q(g2129), .QN(n10310) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n10442), .CLK(n10629), 
        .Q(g2124), .QN(n9600) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n10442), .CLK(n10629), 
        .Q(g2120), .QN(n9429) );
  SDFFX1 DFF_1296_Q_reg ( .D(n37), .SI(g2120), .SE(n10344), .CLK(n10531), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n10344), .CLK(n10531), 
        .Q(g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n10344), .CLK(n10531), 
        .Q(g2257), .QN(n10029) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n10344), .CLK(n10531), 
        .Q(g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n10344), .CLK(n10531), 
        .Q(test_so79), .QN(n10322) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n10452), .CLK(n10639), .Q(g2429) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n10452), .CLK(n10639), 
        .Q(g2418), .QN(n9967) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n10452), .CLK(n10639), 
        .Q(g2421) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n10452), .CLK(n10639), 
        .Q(g2444) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n10452), .CLK(n10639), 
        .Q(g2433), .QN(n9944) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n10451), .CLK(n10638), 
        .Q(g2436) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n10451), .CLK(n10638), 
        .Q(g2459) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n10452), .CLK(n10639), 
        .Q(g2448), .QN(n9678) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n10451), .CLK(n10638), 
        .Q(g2451) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n10452), .CLK(n10639), 
        .Q(g2473) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n10452), .CLK(n10639), 
        .Q(g2463), .QN(n9956) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n10444), .CLK(n10631), 
        .Q(g2466) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n10445), .CLK(n10632), 
        .Q(g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n10446), .CLK(n10633), 
        .Q(g2486), .QN(n9744) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n10446), .CLK(n10633), 
        .Q(test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n10445), .CLK(n10632), .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n10445), .CLK(n10632), 
        .Q(g2495), .QN(n9743) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n10445), .CLK(n10632), 
        .Q(g2498), .QN(n9756) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n10445), .CLK(n10632), 
        .Q(g2502) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n10445), .CLK(n10632), 
        .Q(g2503), .QN(n9979) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n10445), .CLK(n10632), 
        .Q(g2501) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n10445), .CLK(n10632), 
        .Q(g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n10445), .CLK(n10632), 
        .Q(g2507), .QN(n9742) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n10445), .CLK(n10632), 
        .Q(g2510), .QN(n9754) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n10446), .CLK(n10633), 
        .Q(g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n10446), .CLK(n10633), 
        .Q(g2516), .QN(n9741) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n10446), .CLK(n10633), 
        .Q(g2519), .QN(n9752) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n10446), .CLK(n10633), 
        .Q(g2523), .QN(n9987) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n10445), .CLK(n10632), 
        .Q(g2524), .QN(n9978) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n10445), .CLK(n10632), 
        .Q(test_so81) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n10444), .CLK(n10631), .Q(g2387) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n10444), .CLK(n10631), 
        .Q(g2388), .QN(n9536) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n10444), .CLK(n10631), 
        .Q(g2389) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n10444), .CLK(n10631), 
        .Q(g2390) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n10444), .CLK(n10631), 
        .Q(g2391), .QN(n9535) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n10444), .CLK(n10631), 
        .Q(g2392) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n10444), .CLK(n10631), 
        .Q(g2393) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n10444), .CLK(n10631), 
        .Q(g2394), .QN(n9534) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n10444), .CLK(n10631), 
        .Q(g2395) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n10453), .CLK(n10640), 
        .Q(g2397) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n10453), .CLK(n10640), 
        .Q(g2398), .QN(n9588) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n10344), .CLK(n10531), 
        .Q(g2396) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n10344), .CLK(n10531), 
        .Q(g2478) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n10344), .CLK(n10531), 
        .Q(g2479), .QN(n9977) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n10344), .CLK(n10531), 
        .Q(test_so82) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n10355), .CLK(n10542), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n10356), .CLK(n10543), 
        .Q(n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n10356), .CLK(n10543), 
        .Q(g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n10356), .CLK(n10543), 
        .Q(n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n10356), .CLK(n10543), 
        .Q(g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n10356), .CLK(n10543), 
        .Q(n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n10356), .CLK(n10543), 
        .Q(g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n10356), .CLK(n10543), 
        .Q(n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n10356), .CLK(n10543), 
        .Q(g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n10356), .CLK(n10543), 
        .Q(n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n10356), .CLK(n10543), 
        .Q(g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n10356), .CLK(n10543), 
        .Q(n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n10356), .CLK(n10543), 
        .Q(g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n10357), .CLK(n10544), 
        .Q(n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n10357), .CLK(n10544), 
        .Q(test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n10357), .CLK(
        n10544), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n10458), .CLK(n10645), 
        .Q(g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n10458), .CLK(n10645), 
        .Q(n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n10458), .CLK(n10645), 
        .Q(g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n10458), .CLK(n10645), 
        .Q(g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n10459), .CLK(n10646), 
        .Q(n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n10459), .CLK(n10646), 
        .Q(g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n10459), .CLK(n10646), 
        .Q(g2424), .QN(n18859) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n10459), .CLK(n10646), 
        .Q(g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n10459), .CLK(n10646), 
        .Q(g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n10459), .CLK(n10646), 
        .Q(g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n10459), .CLK(n10646), 
        .Q(g2428), .QN(n9653) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n10459), .CLK(n10646), 
        .Q(g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n10459), .CLK(n10646), 
        .Q(g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n10459), .CLK(n10646), 
        .Q(test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n10459), .CLK(
        n10646), .Q(g2441), .QN(n9444) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n10459), .CLK(n10646), 
        .Q(g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n10460), .CLK(n10647), 
        .Q(g2443), .QN(n9443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n10460), .CLK(n10647), 
        .Q(g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n10460), .CLK(n10647), 
        .Q(g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n10460), .CLK(n10647), 
        .Q(g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n10460), .CLK(n10647), 
        .Q(g2456), .QN(n9618) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n10460), .CLK(n10647), 
        .Q(g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n10460), .CLK(n10647), 
        .Q(g2458), .QN(n9617) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n10460), .CLK(n10647), 
        .Q(g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n10460), .CLK(n10647), 
        .Q(g2469), .QN(n18860) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n10460), .CLK(n10647), 
        .Q(g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n10460), .CLK(n10647), 
        .Q(g2471), .QN(n9452) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n10460), .CLK(n10647), 
        .Q(g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n10461), .CLK(n10648), 
        .Q(test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n10345), .CLK(n10532), 
        .Q(g5747), .QN(n9651) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n10345), .CLK(n10532), 
        .Q(g5796), .QN(n9654) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n10345), .CLK(n10532), 
        .Q(g2412), .QN(n9652) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n10345), .CLK(n10532), 
        .Q(g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n10345), .CLK(n10532), 
        .Q(g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n10345), .CLK(n10532), 
        .Q(g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(n1689), .SI(g2624), .SE(n10346), .CLK(n10533), 
        .Q(g2628), .QN(n10264) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n10346), .CLK(n10533), 
        .Q(g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n10346), .CLK(n10533), 
        .Q(g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1684), .SI(g2584), .SE(n10448), .CLK(n10635), 
        .Q(g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n10448), .CLK(n10635), 
        .Q(g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n10448), .CLK(n10635), 
        .Q(g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n10448), .CLK(n10635), 
        .Q(g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n10448), .CLK(n10635), 
        .Q(g2643), .QN(n9811) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n10448), .CLK(n10635), 
        .Q(test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n10448), .CLK(
        n10635), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n10448), .CLK(n10635), 
        .Q(g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n10448), .CLK(n10635), 
        .Q(g2647), .QN(n9812) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n10446), .CLK(n10633), 
        .Q(g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n10446), .CLK(n10633), 
        .Q(g2639), .QN(n9809) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n10447), .CLK(n10634), 
        .Q(g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n10447), .CLK(n10634), 
        .Q(g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n10447), .CLK(n10634), 
        .Q(g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n10447), .CLK(n10634), 
        .Q(g2564), .QN(n9810) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n10447), .CLK(n10634), 
        .Q(g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n10447), .CLK(n10634), 
        .Q(g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n10447), .CLK(n10634), 
        .Q(g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n10447), .CLK(n10634), 
        .Q(g2561), .QN(n10037) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n10447), .CLK(n10634), 
        .Q(g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n10447), .CLK(n10634), 
        .Q(test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n10448), .CLK(n10635), .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n10448), .CLK(n10635), 
        .Q(g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n10448), .CLK(n10635), 
        .Q(g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n10449), .CLK(n10636), 
        .Q(g2552), .QN(n10042) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n10449), .CLK(n10636), 
        .Q(g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n10449), .CLK(n10636), 
        .Q(g2554), .QN(n10043) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n10446), .CLK(n10633), 
        .Q(g2555), .QN(n10039) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n10446), .CLK(n10633), 
        .Q(g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n10446), .CLK(n10633), 
        .Q(g2539), .QN(n10040) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n10446), .CLK(n10633), 
        .Q(g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n10447), .CLK(n10634), 
        .Q(g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n10447), .CLK(n10634), 
        .Q(g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1683), .SI(g2546), .SE(n10449), .CLK(n10636), 
        .Q(g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n10449), .CLK(n10636), 
        .Q(g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n10449), .CLK(n10636), 
        .Q(test_so88), .QN(n9688) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n10449), .CLK(n10636), .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n10449), .CLK(n10636), 
        .Q(n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n10451), .CLK(n10638), 
        .Q(n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n10449), .CLK(n10636), 
        .Q(g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n10449), .CLK(n10636), 
        .Q(g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n10449), .CLK(n10636), 
        .Q(g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n10449), .CLK(n10636), 
        .Q(g2633), .QN(n10076) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n10450), .CLK(n10637), 
        .Q(g2650) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n10451), .CLK(n10638), 
        .Q(g2651), .QN(n9607) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n10451), .CLK(n10638), 
        .Q(g2649) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n10451), .CLK(n10638), 
        .Q(g2653) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n10451), .CLK(n10638), 
        .Q(g2654), .QN(n9627) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n10451), .CLK(n10638), 
        .Q(g2652) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n10451), .CLK(n10638), 
        .Q(g2656) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n10451), .CLK(n10638), 
        .Q(test_so89), .QN(n10332) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n10450), .CLK(n10637), .Q(g2655) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n10450), .CLK(n10637), 
        .Q(g2659) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n10450), .CLK(n10637), 
        .Q(g2660), .QN(n9642) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n10450), .CLK(n10637), 
        .Q(g2658) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n10450), .CLK(n10637), 
        .Q(g2661), .QN(n9701) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n10450), .CLK(n10637), 
        .Q(g2664), .QN(n9703) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n10450), .CLK(n10637), 
        .Q(g2667), .QN(n9702) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n10450), .CLK(n10637), 
        .Q(g2670), .QN(n9687) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n10450), .CLK(n10637), 
        .Q(g2673), .QN(n9690) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n10450), .CLK(n10637), 
        .Q(g2676), .QN(n9689) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n10450), .CLK(n10637), 
        .Q(g2688), .QN(n9719) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n10451), .CLK(n10638), 
        .Q(g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n10346), .CLK(n10533), 
        .Q(g2694), .QN(n9720) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n10461), .CLK(n10648), 
        .Q(g2679), .QN(n9728) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n10461), .CLK(n10648), 
        .Q(test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n10461), .CLK(n10648), .Q(g2685), .QN(n9729) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n10461), .CLK(n10648), 
        .Q(g2565), .QN(n9786) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n10461), .CLK(n10648), 
        .Q(g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n10461), .CLK(n10648), 
        .Q(g2571), .QN(n9788) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n10461), .CLK(n10648), 
        .Q(g2580), .QN(n9796) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n10347), .CLK(n10534), 
        .Q(n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n10347), .CLK(n10534), 
        .Q(g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n10347), .CLK(n10534), 
        .Q(g2599), .QN(n10033) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n10357), .CLK(
        n10544), .Q(n7925) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n10357), .CLK(
        n10544), .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n10357), .CLK(
        n10544), .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n10357), .CLK(
        n10544), .Q(n7922) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n10357), .CLK(
        n10544), .Q(n7921) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n10357), .CLK(
        n10544), .Q(n7920) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n10357), .CLK(
        n10544), .Q(test_so91) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n10357), .CLK(
        n10544), .Q(g2611) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n10461), .CLK(n10648), 
        .Q(g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n10461), .CLK(n10648), 
        .Q(n7918), .QN(n18856) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n10461), .CLK(n10648), 
        .Q(g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n10462), .CLK(n10649), 
        .Q(g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n10462), .CLK(n10649), 
        .Q(g2704), .QN(n10072) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n10462), .CLK(n10649), 
        .Q(g2733) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n10462), .CLK(n10649), 
        .Q(g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(n10462), .CLK(n10649), 
        .Q(g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n10462), .CLK(n10649), 
        .Q(g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n10462), .CLK(n10649), 
        .Q(g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n10462), .CLK(n10649), 
        .Q(g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(n10462), .CLK(n10649), 
        .Q(g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n10462), .CLK(n10649), 
        .Q(test_so92), .QN(n10324) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n10462), .CLK(n10649), .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n10462), .CLK(n10649), 
        .Q(g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n10463), .CLK(n10650), 
        .Q(g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n10463), .CLK(n10650), 
        .Q(g2773) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n10463), .CLK(n10650), 
        .Q(g2774) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n10463), .CLK(n10650), 
        .Q(g2772), .QN(n10162) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n10464), .CLK(n10651), 
        .Q(g2776) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n10464), .CLK(n10651), 
        .Q(g2777) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n10464), .CLK(n10651), 
        .Q(g2775), .QN(n10161) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n10464), .CLK(n10651), 
        .Q(g2779) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n10464), .CLK(n10651), 
        .Q(g2780) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n10464), .CLK(n10651), 
        .Q(g2778), .QN(n10160) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n10464), .CLK(n10651), 
        .Q(g2782) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n10464), .CLK(n10651), 
        .Q(g2783) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n10464), .CLK(n10651), 
        .Q(test_so93), .QN(n10334) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n10464), .CLK(n10651), .Q(g2785) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n10464), .CLK(n10651), 
        .Q(g2786) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n10465), .CLK(n10652), 
        .Q(g2784), .QN(n10159) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n10465), .CLK(n10652), 
        .Q(g2788) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n10465), .CLK(n10652), 
        .Q(g2789) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n10465), .CLK(n10652), 
        .Q(g2787), .QN(n10158) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n10465), .CLK(n10652), 
        .Q(g2791) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n10465), .CLK(n10652), 
        .Q(g2792) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n10465), .CLK(n10652), 
        .Q(g2790), .QN(n10157) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n10465), .CLK(n10652), 
        .Q(g2794) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n10465), .CLK(n10652), 
        .Q(g2795) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n10465), .CLK(n10652), 
        .Q(g2793), .QN(n10156) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n10465), .CLK(n10652), 
        .Q(g2797) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n10465), .CLK(n10652), 
        .Q(g2798) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n10466), .CLK(n10653), 
        .Q(test_so94), .QN(n10335) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n10463), .CLK(n10650), .Q(g2800) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n10463), .CLK(n10650), 
        .Q(g2801) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n10463), .CLK(n10650), 
        .Q(g2799), .QN(n10155) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n10463), .CLK(n10650), 
        .Q(g2803), .QN(n10300) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n10463), .CLK(n10650), 
        .Q(g2804) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n10463), .CLK(n10650), 
        .Q(g2802) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n10463), .CLK(n10650), 
        .Q(g2806) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n10463), .CLK(n10650), 
        .Q(g2807), .QN(n9878) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n10464), .CLK(n10651), 
        .Q(g2805) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n10466), .CLK(n10653), 
        .Q(g2809) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n10466), .CLK(n10653), 
        .Q(g2810) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n10347), .CLK(n10534), 
        .Q(g2808) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n10466), .CLK(n10653), 
        .Q(g2812), .QN(n10193) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n10466), .CLK(n10653), 
        .Q(g2813) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n10466), .CLK(n10653), 
        .Q(test_so95) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n10345), .CLK(n10532), .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n10345), .CLK(n10532), 
        .Q(n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263_Tj_Payload), .SI(n7912), .SE(n10345), .CLK(
        n10532), .Q(n4598), .QN(n10302) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n10455), .CLK(n10642), 
        .Q(g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n10456), .CLK(n10643), 
        .Q(g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n10456), .CLK(n10643), 
        .Q(g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n10456), .CLK(n10643), 
        .Q(g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n10456), .CLK(n10643), 
        .Q(g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n10457), .CLK(n10644), 
        .Q(g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n10457), .CLK(n10644), 
        .Q(g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n10457), .CLK(n10644), 
        .Q(g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n10457), .CLK(n10644), 
        .Q(g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n10457), .CLK(n10644), 
        .Q(g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n10458), .CLK(n10645), 
        .Q(g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n10458), .CLK(n10645), 
        .Q(test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n10453), .CLK(n10640), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n10453), .CLK(n10640), 
        .Q(g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n10453), .CLK(n10640), 
        .Q(g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n10454), .CLK(n10641), 
        .Q(g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n10454), .CLK(n10641), 
        .Q(g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n10454), .CLK(n10641), 
        .Q(g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n10454), .CLK(n10641), 
        .Q(g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n10454), .CLK(n10641), 
        .Q(g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n10454), .CLK(n10641), 
        .Q(g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n10454), .CLK(n10641), 
        .Q(g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n10454), .CLK(n10641), 
        .Q(g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n10454), .CLK(n10641), 
        .Q(g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n10454), .CLK(n10641), 
        .Q(g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n10455), .CLK(n10642), 
        .Q(g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n10455), .CLK(n10642), 
        .Q(test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n10348), .CLK(n10535), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n10348), .CLK(n10535), 
        .Q(g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n10348), .CLK(n10535), 
        .Q(g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n10348), .CLK(n10535), 
        .Q(g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n10348), .CLK(n10535), 
        .Q(g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n10348), .CLK(n10535), 
        .Q(g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n10348), .CLK(n10535), 
        .Q(g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n10346), .CLK(n10533), 
        .Q(g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n10347), .CLK(n10534), 
        .Q(g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n10347), .CLK(n10534), 
        .Q(g2993), .QN(n10303) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n10347), .CLK(n10534), 
        .Q(n7909), .QN(n18873) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(n10347), .CLK(n10534), 
        .Q(g3006), .QN(n10305) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n10347), .CLK(n10534), 
        .Q(g3002), .QN(n10304) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n10347), .CLK(n10534), 
        .Q(g3013), .QN(n10311) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n10347), .CLK(n10534), 
        .Q(test_so98), .QN(n10327) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n10347), .CLK(n10534), .Q(g3024) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n10346), .CLK(n10533), 
        .Q(g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(n10346), .CLK(n10533), 
        .Q(g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n10346), .CLK(n10533), 
        .Q(g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n10346), .CLK(n10533), 
        .Q(g3032), .QN(n9736) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n10346), .CLK(n10533), 
        .Q(g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n10346), .CLK(n10533), 
        .Q(n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n10346), .CLK(n10533), 
        .Q(g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n10455), .CLK(n10642), 
        .Q(g8275), .QN(n10288) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n10456), .CLK(n10643), 
        .Q(g8274), .QN(n10290) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n10456), .CLK(n10643), 
        .Q(g8273), .QN(n18874) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n10456), .CLK(n10643), 
        .Q(g8272), .QN(n18875) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n10456), .CLK(n10643), 
        .Q(g8268), .QN(n18876) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n10457), .CLK(n10644), 
        .Q(g8269), .QN(n10291) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n10457), .CLK(n10644), 
        .Q(test_so99), .QN(n10330) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n10457), .CLK(
        n10644), .Q(g8271), .QN(n10289) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n10457), .CLK(n10644), 
        .Q(g3083), .QN(n10293) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n10457), .CLK(n10644), 
        .Q(g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n10457), .CLK(n10644), .Q(
        n4577), .QN(n9739) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n10457), .CLK(n10644), 
        .Q(g8266), .QN(n18877) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n10458), .CLK(n10645), 
        .Q(g8265), .QN(n18878) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n10458), .CLK(n10645), 
        .Q(g8264) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n10458), .CLK(n10645), 
        .Q(g8262), .QN(n18879) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n10458), .CLK(n10645), 
        .Q(g8263), .QN(n10272) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n10458), .CLK(n10645), 
        .Q(g8260), .QN(n10268) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n10348), .CLK(n10535), 
        .Q(g8261), .QN(n10269) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n10454), .CLK(n10641), 
        .Q(g8259), .QN(n10270) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n10454), .CLK(n10641), 
        .Q(g2990), .QN(n10295) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n10348), .CLK(n10535), .Q(
        n4578), .QN(n9738) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n10470), .CLK(n10657), 
        .Q(test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n10379), .CLK(n10566), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n10345), .CLK(n10532), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n10351), .CLK(n10538), 
        .Q(g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n10461), .CLK(n10648), 
        .Q(g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n10344), .CLK(n10531), 
        .Q(g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n10413), .CLK(n10600), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n10413), .CLK(n10600), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n10344), .CLK(n10531), 
        .Q(n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n10360), .CLK(n10547), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n10360), .CLK(n10547), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n145), .IN2(n3016), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n3023), .IN2(n3000), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n3008), .IN2(n3068), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n3128), .IN2(n3036), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(n3758), .IN2(n3788), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n3751), .IN2(n3749), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n2792), .IN2(n2632), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n2351), .IN2(n567), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(n4263), .Q(n4263_Tj_Payload)
         );
  NBUFFX2 U10157 ( .INP(n10514), .Z(n10341) );
  NBUFFX2 U10158 ( .INP(n10514), .Z(n10340) );
  NBUFFX2 U10159 ( .INP(n10476), .Z(n10454) );
  NBUFFX2 U10160 ( .INP(n10475), .Z(n10457) );
  NBUFFX2 U10161 ( .INP(n10472), .Z(n10465) );
  NBUFFX2 U10162 ( .INP(n10473), .Z(n10464) );
  NBUFFX2 U10163 ( .INP(n10473), .Z(n10463) );
  NBUFFX2 U10164 ( .INP(n10473), .Z(n10462) );
  NBUFFX2 U10165 ( .INP(n10512), .Z(n10347) );
  NBUFFX2 U10166 ( .INP(n10477), .Z(n10450) );
  NBUFFX2 U10167 ( .INP(n10478), .Z(n10449) );
  NBUFFX2 U10168 ( .INP(n10478), .Z(n10447) );
  NBUFFX2 U10169 ( .INP(n10478), .Z(n10448) );
  NBUFFX2 U10170 ( .INP(n10512), .Z(n10346) );
  NBUFFX2 U10171 ( .INP(n10474), .Z(n10461) );
  NBUFFX2 U10172 ( .INP(n10474), .Z(n10460) );
  NBUFFX2 U10173 ( .INP(n10474), .Z(n10459) );
  NBUFFX2 U10174 ( .INP(n10509), .Z(n10356) );
  NBUFFX2 U10175 ( .INP(n10479), .Z(n10446) );
  NBUFFX2 U10176 ( .INP(n10479), .Z(n10445) );
  NBUFFX2 U10177 ( .INP(n10477), .Z(n10451) );
  NBUFFX2 U10178 ( .INP(n10480), .Z(n10442) );
  NBUFFX2 U10179 ( .INP(n10479), .Z(n10444) );
  NBUFFX2 U10180 ( .INP(n10480), .Z(n10443) );
  NBUFFX2 U10181 ( .INP(n10476), .Z(n10453) );
  NBUFFX2 U10182 ( .INP(n10477), .Z(n10452) );
  NBUFFX2 U10183 ( .INP(n10480), .Z(n10441) );
  NBUFFX2 U10184 ( .INP(n10481), .Z(n10440) );
  NBUFFX2 U10185 ( .INP(n10513), .Z(n10344) );
  NBUFFX2 U10186 ( .INP(n10481), .Z(n10439) );
  NBUFFX2 U10187 ( .INP(n10481), .Z(n10438) );
  NBUFFX2 U10188 ( .INP(n10482), .Z(n10437) );
  NBUFFX2 U10189 ( .INP(n10482), .Z(n10436) );
  NBUFFX2 U10190 ( .INP(n10482), .Z(n10435) );
  NBUFFX2 U10191 ( .INP(n10483), .Z(n10434) );
  NBUFFX2 U10192 ( .INP(n10483), .Z(n10433) );
  NBUFFX2 U10193 ( .INP(n10483), .Z(n10432) );
  NBUFFX2 U10194 ( .INP(n10484), .Z(n10431) );
  NBUFFX2 U10195 ( .INP(n10484), .Z(n10430) );
  NBUFFX2 U10196 ( .INP(n10484), .Z(n10429) );
  NBUFFX2 U10197 ( .INP(n10485), .Z(n10428) );
  NBUFFX2 U10198 ( .INP(n10485), .Z(n10427) );
  NBUFFX2 U10199 ( .INP(n10485), .Z(n10426) );
  NBUFFX2 U10200 ( .INP(n10486), .Z(n10425) );
  NBUFFX2 U10201 ( .INP(n10486), .Z(n10424) );
  NBUFFX2 U10202 ( .INP(n10489), .Z(n10414) );
  NBUFFX2 U10203 ( .INP(n10487), .Z(n10420) );
  NBUFFX2 U10204 ( .INP(n10487), .Z(n10421) );
  NBUFFX2 U10205 ( .INP(n10490), .Z(n10413) );
  NBUFFX2 U10206 ( .INP(n10490), .Z(n10412) );
  NBUFFX2 U10207 ( .INP(n10488), .Z(n10419) );
  NBUFFX2 U10208 ( .INP(n10486), .Z(n10423) );
  NBUFFX2 U10209 ( .INP(n10487), .Z(n10422) );
  NBUFFX2 U10210 ( .INP(n10488), .Z(n10418) );
  NBUFFX2 U10211 ( .INP(n10488), .Z(n10417) );
  NBUFFX2 U10212 ( .INP(n10489), .Z(n10416) );
  NBUFFX2 U10213 ( .INP(n10489), .Z(n10415) );
  NBUFFX2 U10214 ( .INP(n10490), .Z(n10411) );
  NBUFFX2 U10215 ( .INP(n10491), .Z(n10410) );
  NBUFFX2 U10216 ( .INP(n10491), .Z(n10409) );
  NBUFFX2 U10217 ( .INP(n10491), .Z(n10408) );
  NBUFFX2 U10218 ( .INP(n10512), .Z(n10345) );
  NBUFFX2 U10219 ( .INP(n10492), .Z(n10407) );
  NBUFFX2 U10220 ( .INP(n10492), .Z(n10406) );
  NBUFFX2 U10221 ( .INP(n10492), .Z(n10405) );
  NBUFFX2 U10222 ( .INP(n10493), .Z(n10404) );
  NBUFFX2 U10223 ( .INP(n10493), .Z(n10403) );
  NBUFFX2 U10224 ( .INP(n10493), .Z(n10402) );
  NBUFFX2 U10225 ( .INP(n10494), .Z(n10401) );
  NBUFFX2 U10226 ( .INP(n10494), .Z(n10400) );
  NBUFFX2 U10227 ( .INP(n10494), .Z(n10399) );
  NBUFFX2 U10228 ( .INP(n10495), .Z(n10398) );
  NBUFFX2 U10229 ( .INP(n10495), .Z(n10397) );
  NBUFFX2 U10230 ( .INP(n10495), .Z(n10396) );
  NBUFFX2 U10231 ( .INP(n10496), .Z(n10393) );
  NBUFFX2 U10232 ( .INP(n10499), .Z(n10386) );
  NBUFFX2 U10233 ( .INP(n10496), .Z(n10395) );
  NBUFFX2 U10234 ( .INP(n10496), .Z(n10394) );
  NBUFFX2 U10235 ( .INP(n10497), .Z(n10390) );
  NBUFFX2 U10236 ( .INP(n10497), .Z(n10392) );
  NBUFFX2 U10237 ( .INP(n10497), .Z(n10391) );
  NBUFFX2 U10238 ( .INP(n10498), .Z(n10387) );
  NBUFFX2 U10239 ( .INP(n10498), .Z(n10389) );
  NBUFFX2 U10240 ( .INP(n10498), .Z(n10388) );
  NBUFFX2 U10241 ( .INP(n10499), .Z(n10385) );
  NBUFFX2 U10242 ( .INP(n10499), .Z(n10384) );
  NBUFFX2 U10243 ( .INP(n10500), .Z(n10383) );
  NBUFFX2 U10244 ( .INP(n10500), .Z(n10382) );
  NBUFFX2 U10245 ( .INP(n10500), .Z(n10381) );
  NBUFFX2 U10246 ( .INP(n10501), .Z(n10380) );
  NBUFFX2 U10247 ( .INP(n10475), .Z(n10456) );
  NBUFFX2 U10248 ( .INP(n10501), .Z(n10378) );
  NBUFFX2 U10249 ( .INP(n10502), .Z(n10377) );
  NBUFFX2 U10250 ( .INP(n10502), .Z(n10376) );
  NBUFFX2 U10251 ( .INP(n10502), .Z(n10375) );
  NBUFFX2 U10252 ( .INP(n10503), .Z(n10374) );
  NBUFFX2 U10253 ( .INP(n10503), .Z(n10373) );
  NBUFFX2 U10254 ( .INP(n10503), .Z(n10372) );
  NBUFFX2 U10255 ( .INP(n10504), .Z(n10371) );
  NBUFFX2 U10256 ( .INP(n10501), .Z(n10379) );
  NBUFFX2 U10257 ( .INP(n10508), .Z(n10358) );
  NBUFFX2 U10258 ( .INP(n10508), .Z(n10357) );
  NBUFFX2 U10259 ( .INP(n10476), .Z(n10455) );
  NBUFFX2 U10260 ( .INP(n10505), .Z(n10367) );
  NBUFFX2 U10261 ( .INP(n10505), .Z(n10368) );
  NBUFFX2 U10262 ( .INP(n10507), .Z(n10360) );
  NBUFFX2 U10263 ( .INP(n10505), .Z(n10366) );
  NBUFFX2 U10264 ( .INP(n10506), .Z(n10365) );
  NBUFFX2 U10265 ( .INP(n10504), .Z(n10370) );
  NBUFFX2 U10266 ( .INP(n10504), .Z(n10369) );
  NBUFFX2 U10267 ( .INP(n10507), .Z(n10361) );
  NBUFFX2 U10268 ( .INP(n10508), .Z(n10359) );
  NBUFFX2 U10269 ( .INP(n10507), .Z(n10362) );
  NBUFFX2 U10270 ( .INP(n10506), .Z(n10364) );
  NBUFFX2 U10271 ( .INP(n10506), .Z(n10363) );
  NBUFFX2 U10272 ( .INP(n10511), .Z(n10348) );
  NBUFFX2 U10273 ( .INP(n10511), .Z(n10350) );
  NBUFFX2 U10274 ( .INP(n10511), .Z(n10349) );
  NBUFFX2 U10275 ( .INP(n10471), .Z(n10469) );
  NBUFFX2 U10276 ( .INP(n10472), .Z(n10467) );
  NBUFFX2 U10277 ( .INP(n10471), .Z(n10468) );
  NBUFFX2 U10278 ( .INP(n10472), .Z(n10466) );
  NBUFFX2 U10279 ( .INP(n10475), .Z(n10458) );
  NBUFFX2 U10280 ( .INP(n10509), .Z(n10355) );
  NBUFFX2 U10281 ( .INP(n10509), .Z(n10354) );
  NBUFFX2 U10282 ( .INP(n10510), .Z(n10353) );
  NBUFFX2 U10283 ( .INP(n10510), .Z(n10352) );
  NBUFFX2 U10284 ( .INP(n10510), .Z(n10351) );
  NBUFFX2 U10285 ( .INP(n10513), .Z(n10343) );
  NBUFFX2 U10286 ( .INP(n10513), .Z(n10342) );
  NBUFFX2 U10287 ( .INP(n10701), .Z(n10528) );
  NBUFFX2 U10288 ( .INP(n10701), .Z(n10527) );
  NBUFFX2 U10289 ( .INP(n10663), .Z(n10641) );
  NBUFFX2 U10290 ( .INP(n10662), .Z(n10644) );
  NBUFFX2 U10291 ( .INP(n10659), .Z(n10652) );
  NBUFFX2 U10292 ( .INP(n10660), .Z(n10651) );
  NBUFFX2 U10293 ( .INP(n10660), .Z(n10650) );
  NBUFFX2 U10294 ( .INP(n10660), .Z(n10649) );
  NBUFFX2 U10295 ( .INP(n10699), .Z(n10534) );
  NBUFFX2 U10296 ( .INP(n10664), .Z(n10637) );
  NBUFFX2 U10297 ( .INP(n10665), .Z(n10636) );
  NBUFFX2 U10298 ( .INP(n10665), .Z(n10634) );
  NBUFFX2 U10299 ( .INP(n10665), .Z(n10635) );
  NBUFFX2 U10300 ( .INP(n10699), .Z(n10533) );
  NBUFFX2 U10301 ( .INP(n10661), .Z(n10648) );
  NBUFFX2 U10302 ( .INP(n10661), .Z(n10647) );
  NBUFFX2 U10303 ( .INP(n10661), .Z(n10646) );
  NBUFFX2 U10304 ( .INP(n10696), .Z(n10543) );
  NBUFFX2 U10305 ( .INP(n10666), .Z(n10633) );
  NBUFFX2 U10306 ( .INP(n10666), .Z(n10632) );
  NBUFFX2 U10307 ( .INP(n10664), .Z(n10638) );
  NBUFFX2 U10308 ( .INP(n10667), .Z(n10629) );
  NBUFFX2 U10309 ( .INP(n10666), .Z(n10631) );
  NBUFFX2 U10310 ( .INP(n10667), .Z(n10630) );
  NBUFFX2 U10311 ( .INP(n10663), .Z(n10640) );
  NBUFFX2 U10312 ( .INP(n10664), .Z(n10639) );
  NBUFFX2 U10313 ( .INP(n10667), .Z(n10628) );
  NBUFFX2 U10314 ( .INP(n10668), .Z(n10627) );
  NBUFFX2 U10315 ( .INP(n10700), .Z(n10531) );
  NBUFFX2 U10316 ( .INP(n10668), .Z(n10626) );
  NBUFFX2 U10317 ( .INP(n10668), .Z(n10625) );
  NBUFFX2 U10318 ( .INP(n10669), .Z(n10624) );
  NBUFFX2 U10319 ( .INP(n10669), .Z(n10623) );
  NBUFFX2 U10320 ( .INP(n10669), .Z(n10622) );
  NBUFFX2 U10321 ( .INP(n10670), .Z(n10621) );
  NBUFFX2 U10322 ( .INP(n10670), .Z(n10620) );
  NBUFFX2 U10323 ( .INP(n10670), .Z(n10619) );
  NBUFFX2 U10324 ( .INP(n10671), .Z(n10618) );
  NBUFFX2 U10325 ( .INP(n10671), .Z(n10617) );
  NBUFFX2 U10326 ( .INP(n10671), .Z(n10616) );
  NBUFFX2 U10327 ( .INP(n10672), .Z(n10615) );
  NBUFFX2 U10328 ( .INP(n10672), .Z(n10614) );
  NBUFFX2 U10329 ( .INP(n10672), .Z(n10613) );
  NBUFFX2 U10330 ( .INP(n10673), .Z(n10612) );
  NBUFFX2 U10331 ( .INP(n10673), .Z(n10611) );
  NBUFFX2 U10332 ( .INP(n10676), .Z(n10601) );
  NBUFFX2 U10333 ( .INP(n10674), .Z(n10607) );
  NBUFFX2 U10334 ( .INP(n10674), .Z(n10608) );
  NBUFFX2 U10335 ( .INP(n10677), .Z(n10600) );
  NBUFFX2 U10336 ( .INP(n10677), .Z(n10599) );
  NBUFFX2 U10337 ( .INP(n10675), .Z(n10606) );
  NBUFFX2 U10338 ( .INP(n10673), .Z(n10610) );
  NBUFFX2 U10339 ( .INP(n10674), .Z(n10609) );
  NBUFFX2 U10340 ( .INP(n10675), .Z(n10605) );
  NBUFFX2 U10341 ( .INP(n10675), .Z(n10604) );
  NBUFFX2 U10342 ( .INP(n10676), .Z(n10603) );
  NBUFFX2 U10343 ( .INP(n10676), .Z(n10602) );
  NBUFFX2 U10344 ( .INP(n10677), .Z(n10598) );
  NBUFFX2 U10345 ( .INP(n10678), .Z(n10597) );
  NBUFFX2 U10346 ( .INP(n10678), .Z(n10596) );
  NBUFFX2 U10347 ( .INP(n10678), .Z(n10595) );
  NBUFFX2 U10348 ( .INP(n10699), .Z(n10532) );
  NBUFFX2 U10349 ( .INP(n10679), .Z(n10594) );
  NBUFFX2 U10350 ( .INP(n10679), .Z(n10593) );
  NBUFFX2 U10351 ( .INP(n10679), .Z(n10592) );
  NBUFFX2 U10352 ( .INP(n10680), .Z(n10591) );
  NBUFFX2 U10353 ( .INP(n10680), .Z(n10590) );
  NBUFFX2 U10354 ( .INP(n10680), .Z(n10589) );
  NBUFFX2 U10355 ( .INP(n10681), .Z(n10588) );
  NBUFFX2 U10356 ( .INP(n10681), .Z(n10587) );
  NBUFFX2 U10357 ( .INP(n10681), .Z(n10586) );
  NBUFFX2 U10358 ( .INP(n10682), .Z(n10585) );
  NBUFFX2 U10359 ( .INP(n10682), .Z(n10584) );
  NBUFFX2 U10360 ( .INP(n10682), .Z(n10583) );
  NBUFFX2 U10361 ( .INP(n10683), .Z(n10580) );
  NBUFFX2 U10362 ( .INP(n10686), .Z(n10573) );
  NBUFFX2 U10363 ( .INP(n10683), .Z(n10582) );
  NBUFFX2 U10364 ( .INP(n10683), .Z(n10581) );
  NBUFFX2 U10365 ( .INP(n10684), .Z(n10577) );
  NBUFFX2 U10366 ( .INP(n10684), .Z(n10579) );
  NBUFFX2 U10367 ( .INP(n10684), .Z(n10578) );
  NBUFFX2 U10368 ( .INP(n10685), .Z(n10574) );
  NBUFFX2 U10369 ( .INP(n10685), .Z(n10576) );
  NBUFFX2 U10370 ( .INP(n10685), .Z(n10575) );
  NBUFFX2 U10371 ( .INP(n10686), .Z(n10572) );
  NBUFFX2 U10372 ( .INP(n10686), .Z(n10571) );
  NBUFFX2 U10373 ( .INP(n10687), .Z(n10570) );
  NBUFFX2 U10374 ( .INP(n10687), .Z(n10569) );
  NBUFFX2 U10375 ( .INP(n10687), .Z(n10568) );
  NBUFFX2 U10376 ( .INP(n10688), .Z(n10567) );
  NBUFFX2 U10377 ( .INP(n10662), .Z(n10643) );
  NBUFFX2 U10378 ( .INP(n10688), .Z(n10565) );
  NBUFFX2 U10379 ( .INP(n10689), .Z(n10564) );
  NBUFFX2 U10380 ( .INP(n10689), .Z(n10563) );
  NBUFFX2 U10381 ( .INP(n10689), .Z(n10562) );
  NBUFFX2 U10382 ( .INP(n10690), .Z(n10561) );
  NBUFFX2 U10383 ( .INP(n10690), .Z(n10560) );
  NBUFFX2 U10384 ( .INP(n10690), .Z(n10559) );
  NBUFFX2 U10385 ( .INP(n10691), .Z(n10558) );
  NBUFFX2 U10386 ( .INP(n10688), .Z(n10566) );
  NBUFFX2 U10387 ( .INP(n10695), .Z(n10545) );
  NBUFFX2 U10388 ( .INP(n10695), .Z(n10544) );
  NBUFFX2 U10389 ( .INP(n10663), .Z(n10642) );
  NBUFFX2 U10390 ( .INP(n10692), .Z(n10554) );
  NBUFFX2 U10391 ( .INP(n10692), .Z(n10555) );
  NBUFFX2 U10392 ( .INP(n10694), .Z(n10547) );
  NBUFFX2 U10393 ( .INP(n10692), .Z(n10553) );
  NBUFFX2 U10394 ( .INP(n10693), .Z(n10552) );
  NBUFFX2 U10395 ( .INP(n10691), .Z(n10557) );
  NBUFFX2 U10396 ( .INP(n10691), .Z(n10556) );
  NBUFFX2 U10397 ( .INP(n10694), .Z(n10548) );
  NBUFFX2 U10398 ( .INP(n10695), .Z(n10546) );
  NBUFFX2 U10399 ( .INP(n10694), .Z(n10549) );
  NBUFFX2 U10400 ( .INP(n10693), .Z(n10551) );
  NBUFFX2 U10401 ( .INP(n10693), .Z(n10550) );
  NBUFFX2 U10402 ( .INP(n10698), .Z(n10535) );
  NBUFFX2 U10403 ( .INP(n10698), .Z(n10537) );
  NBUFFX2 U10404 ( .INP(n10698), .Z(n10536) );
  NBUFFX2 U10405 ( .INP(n10658), .Z(n10656) );
  NBUFFX2 U10406 ( .INP(n10659), .Z(n10654) );
  NBUFFX2 U10407 ( .INP(n10658), .Z(n10655) );
  NBUFFX2 U10408 ( .INP(n10659), .Z(n10653) );
  NBUFFX2 U10409 ( .INP(n10662), .Z(n10645) );
  NBUFFX2 U10410 ( .INP(n10696), .Z(n10542) );
  NBUFFX2 U10411 ( .INP(n10696), .Z(n10541) );
  NBUFFX2 U10412 ( .INP(n10697), .Z(n10540) );
  NBUFFX2 U10413 ( .INP(n10697), .Z(n10539) );
  NBUFFX2 U10414 ( .INP(n10697), .Z(n10538) );
  NBUFFX2 U10415 ( .INP(n10700), .Z(n10530) );
  NBUFFX2 U10416 ( .INP(n10700), .Z(n10529) );
  NBUFFX2 U10417 ( .INP(n10471), .Z(n10470) );
  NBUFFX2 U10418 ( .INP(n10658), .Z(n10657) );
  NBUFFX2 U10419 ( .INP(n10710), .Z(n10660) );
  NBUFFX2 U10420 ( .INP(n10523), .Z(n10473) );
  NBUFFX2 U10421 ( .INP(n10710), .Z(n10661) );
  NBUFFX2 U10422 ( .INP(n10523), .Z(n10474) );
  NBUFFX2 U10423 ( .INP(n10710), .Z(n10658) );
  NBUFFX2 U10424 ( .INP(n10523), .Z(n10471) );
  NBUFFX2 U10425 ( .INP(n10710), .Z(n10659) );
  NBUFFX2 U10426 ( .INP(n10523), .Z(n10472) );
  NBUFFX2 U10427 ( .INP(n10709), .Z(n10665) );
  NBUFFX2 U10428 ( .INP(n10522), .Z(n10478) );
  NBUFFX2 U10429 ( .INP(n10709), .Z(n10666) );
  NBUFFX2 U10430 ( .INP(n10522), .Z(n10479) );
  NBUFFX2 U10431 ( .INP(n10709), .Z(n10664) );
  NBUFFX2 U10432 ( .INP(n10522), .Z(n10477) );
  NBUFFX2 U10433 ( .INP(n10708), .Z(n10667) );
  NBUFFX2 U10434 ( .INP(n10521), .Z(n10480) );
  NBUFFX2 U10435 ( .INP(n10708), .Z(n10668) );
  NBUFFX2 U10436 ( .INP(n10521), .Z(n10481) );
  NBUFFX2 U10437 ( .INP(n10708), .Z(n10669) );
  NBUFFX2 U10438 ( .INP(n10521), .Z(n10482) );
  NBUFFX2 U10439 ( .INP(n10708), .Z(n10670) );
  NBUFFX2 U10440 ( .INP(n10521), .Z(n10483) );
  NBUFFX2 U10441 ( .INP(n10708), .Z(n10671) );
  NBUFFX2 U10442 ( .INP(n10521), .Z(n10484) );
  NBUFFX2 U10443 ( .INP(n10707), .Z(n10672) );
  NBUFFX2 U10444 ( .INP(n10520), .Z(n10485) );
  NBUFFX2 U10445 ( .INP(n10707), .Z(n10673) );
  NBUFFX2 U10446 ( .INP(n10520), .Z(n10486) );
  NBUFFX2 U10447 ( .INP(n10707), .Z(n10674) );
  NBUFFX2 U10448 ( .INP(n10520), .Z(n10487) );
  NBUFFX2 U10449 ( .INP(n10707), .Z(n10675) );
  NBUFFX2 U10450 ( .INP(n10520), .Z(n10488) );
  NBUFFX2 U10451 ( .INP(n10707), .Z(n10676) );
  NBUFFX2 U10452 ( .INP(n10520), .Z(n10489) );
  NBUFFX2 U10453 ( .INP(n10706), .Z(n10677) );
  NBUFFX2 U10454 ( .INP(n10519), .Z(n10490) );
  NBUFFX2 U10455 ( .INP(n10706), .Z(n10678) );
  NBUFFX2 U10456 ( .INP(n10519), .Z(n10491) );
  NBUFFX2 U10457 ( .INP(n10702), .Z(n10699) );
  NBUFFX2 U10458 ( .INP(n10515), .Z(n10512) );
  NBUFFX2 U10459 ( .INP(n10706), .Z(n10679) );
  NBUFFX2 U10460 ( .INP(n10519), .Z(n10492) );
  NBUFFX2 U10461 ( .INP(n10706), .Z(n10680) );
  NBUFFX2 U10462 ( .INP(n10519), .Z(n10493) );
  NBUFFX2 U10463 ( .INP(n10706), .Z(n10681) );
  NBUFFX2 U10464 ( .INP(n10519), .Z(n10494) );
  NBUFFX2 U10465 ( .INP(n10705), .Z(n10682) );
  NBUFFX2 U10466 ( .INP(n10518), .Z(n10495) );
  NBUFFX2 U10467 ( .INP(n10705), .Z(n10683) );
  NBUFFX2 U10468 ( .INP(n10518), .Z(n10496) );
  NBUFFX2 U10469 ( .INP(n10705), .Z(n10684) );
  NBUFFX2 U10470 ( .INP(n10518), .Z(n10497) );
  NBUFFX2 U10471 ( .INP(n10705), .Z(n10685) );
  NBUFFX2 U10472 ( .INP(n10518), .Z(n10498) );
  NBUFFX2 U10473 ( .INP(n10705), .Z(n10686) );
  NBUFFX2 U10474 ( .INP(n10518), .Z(n10499) );
  NBUFFX2 U10475 ( .INP(n10704), .Z(n10687) );
  NBUFFX2 U10476 ( .INP(n10517), .Z(n10500) );
  NBUFFX2 U10477 ( .INP(n10704), .Z(n10689) );
  NBUFFX2 U10478 ( .INP(n10517), .Z(n10502) );
  NBUFFX2 U10479 ( .INP(n10704), .Z(n10690) );
  NBUFFX2 U10480 ( .INP(n10517), .Z(n10503) );
  NBUFFX2 U10481 ( .INP(n10704), .Z(n10688) );
  NBUFFX2 U10482 ( .INP(n10517), .Z(n10501) );
  NBUFFX2 U10483 ( .INP(n10709), .Z(n10663) );
  NBUFFX2 U10484 ( .INP(n10522), .Z(n10476) );
  NBUFFX2 U10485 ( .INP(n10703), .Z(n10692) );
  NBUFFX2 U10486 ( .INP(n10516), .Z(n10505) );
  NBUFFX2 U10487 ( .INP(n10704), .Z(n10691) );
  NBUFFX2 U10488 ( .INP(n10517), .Z(n10504) );
  NBUFFX2 U10489 ( .INP(n10703), .Z(n10695) );
  NBUFFX2 U10490 ( .INP(n10516), .Z(n10508) );
  NBUFFX2 U10491 ( .INP(n10703), .Z(n10694) );
  NBUFFX2 U10492 ( .INP(n10516), .Z(n10507) );
  NBUFFX2 U10493 ( .INP(n10703), .Z(n10693) );
  NBUFFX2 U10494 ( .INP(n10516), .Z(n10506) );
  NBUFFX2 U10495 ( .INP(n10702), .Z(n10698) );
  NBUFFX2 U10496 ( .INP(n10515), .Z(n10511) );
  NBUFFX2 U10497 ( .INP(n10709), .Z(n10662) );
  NBUFFX2 U10498 ( .INP(n10522), .Z(n10475) );
  NBUFFX2 U10499 ( .INP(n10703), .Z(n10696) );
  NBUFFX2 U10500 ( .INP(n10516), .Z(n10509) );
  NBUFFX2 U10501 ( .INP(n10702), .Z(n10697) );
  NBUFFX2 U10502 ( .INP(n10515), .Z(n10510) );
  NBUFFX2 U10503 ( .INP(n10702), .Z(n10700) );
  NBUFFX2 U10504 ( .INP(n10515), .Z(n10513) );
  NBUFFX2 U10505 ( .INP(n10702), .Z(n10701) );
  NBUFFX2 U10506 ( .INP(n10515), .Z(n10514) );
  NBUFFX2 U10507 ( .INP(n10526), .Z(n10515) );
  NBUFFX2 U10508 ( .INP(n10526), .Z(n10516) );
  NBUFFX2 U10509 ( .INP(n10526), .Z(n10517) );
  NBUFFX2 U10510 ( .INP(n10525), .Z(n10518) );
  NBUFFX2 U10511 ( .INP(n10525), .Z(n10519) );
  NBUFFX2 U10512 ( .INP(n10525), .Z(n10520) );
  NBUFFX2 U10513 ( .INP(n10524), .Z(n10521) );
  NBUFFX2 U10514 ( .INP(n10524), .Z(n10522) );
  NBUFFX2 U10515 ( .INP(n10524), .Z(n10523) );
  NBUFFX2 U10516 ( .INP(test_se), .Z(n10524) );
  NBUFFX2 U10517 ( .INP(test_se), .Z(n10525) );
  NBUFFX2 U10518 ( .INP(test_se), .Z(n10526) );
  NBUFFX2 U10519 ( .INP(n10713), .Z(n10702) );
  NBUFFX2 U10520 ( .INP(n10713), .Z(n10703) );
  NBUFFX2 U10521 ( .INP(n10713), .Z(n10704) );
  NBUFFX2 U10522 ( .INP(n10712), .Z(n10705) );
  NBUFFX2 U10523 ( .INP(n10712), .Z(n10706) );
  NBUFFX2 U10524 ( .INP(n10712), .Z(n10707) );
  NBUFFX2 U10525 ( .INP(n10711), .Z(n10708) );
  NBUFFX2 U10526 ( .INP(n10711), .Z(n10709) );
  NBUFFX2 U10527 ( .INP(n10711), .Z(n10710) );
  NBUFFX2 U10528 ( .INP(CK), .Z(n10711) );
  NBUFFX2 U10529 ( .INP(CK), .Z(n10712) );
  NBUFFX2 U10530 ( .INP(CK), .Z(n10713) );
  INVX0 U10531 ( .INP(n10714), .ZN(n987) );
  NOR2X0 U10532 ( .IN1(n10715), .IN2(n10716), .QN(n10714) );
  NOR2X0 U10533 ( .IN1(g1236), .IN2(n10266), .QN(n10716) );
  INVX0 U10534 ( .INP(n10717), .ZN(n983) );
  INVX0 U10535 ( .INP(n10718), .ZN(n795) );
  INVX0 U10536 ( .INP(g27380), .ZN(n73) );
  INVX0 U10537 ( .INP(n10719), .ZN(n630) );
  NOR2X0 U10538 ( .IN1(n10720), .IN2(n10721), .QN(n10719) );
  NOR2X0 U10539 ( .IN1(g550), .IN2(n10267), .QN(n10721) );
  INVX0 U10540 ( .INP(n10722), .ZN(n628) );
  INVX0 U10541 ( .INP(n10723), .ZN(n627) );
  INVX0 U10542 ( .INP(n10724), .ZN(n602) );
  INVX0 U10543 ( .INP(n10725), .ZN(n557) );
  INVX0 U10544 ( .INP(n10726), .ZN(n529) );
  NAND2X0 U10545 ( .IN1(n10727), .IN2(n10728), .QN(n4281) );
  NAND2X0 U10546 ( .IN1(n10294), .IN2(n10729), .QN(n10728) );
  INVX0 U10547 ( .INP(n10730), .ZN(n10727) );
  NOR2X0 U10548 ( .IN1(n10729), .IN2(n10294), .QN(n10730) );
  NAND2X0 U10549 ( .IN1(n10731), .IN2(n10732), .QN(n4280) );
  NAND2X0 U10550 ( .IN1(n10292), .IN2(n10733), .QN(n10732) );
  INVX0 U10551 ( .INP(n10734), .ZN(n10731) );
  NOR2X0 U10552 ( .IN1(n10733), .IN2(n10292), .QN(n10734) );
  NAND2X0 U10553 ( .IN1(g2879), .IN2(n10735), .QN(n4279) );
  NAND2X0 U10554 ( .IN1(DFF_18_n1), .IN2(g8021), .QN(n10735) );
  NOR2X0 U10555 ( .IN1(n10736), .IN2(n10737), .QN(n4278) );
  NOR2X0 U10556 ( .IN1(n10738), .IN2(n10739), .QN(n10737) );
  NOR2X0 U10557 ( .IN1(n10740), .IN2(n10741), .QN(n10736) );
  NAND2X0 U10558 ( .IN1(n10742), .IN2(n10743), .QN(n10741) );
  NOR2X0 U10559 ( .IN1(n10744), .IN2(n10745), .QN(n10743) );
  NAND2X0 U10560 ( .IN1(n10746), .IN2(n10747), .QN(n10745) );
  NOR2X0 U10561 ( .IN1(n10748), .IN2(n10749), .QN(n10747) );
  NOR2X0 U10562 ( .IN1(n10022), .IN2(n10750), .QN(n10749) );
  NOR2X0 U10563 ( .IN1(n10751), .IN2(g65), .QN(n10748) );
  NOR2X0 U10564 ( .IN1(n10752), .IN2(n10753), .QN(n10746) );
  NOR2X0 U10565 ( .IN1(n10306), .IN2(n10754), .QN(n10753) );
  NOR2X0 U10566 ( .IN1(n10755), .IN2(g88), .QN(n10752) );
  NAND2X0 U10567 ( .IN1(n10756), .IN2(n10757), .QN(n10744) );
  NAND2X0 U10568 ( .IN1(n10308), .IN2(n10758), .QN(n10757) );
  NAND2X0 U10569 ( .IN1(n10759), .IN2(g61), .QN(n10756) );
  NOR2X0 U10570 ( .IN1(n10760), .IN2(n10761), .QN(n10742) );
  NAND2X0 U10571 ( .IN1(n10762), .IN2(n10763), .QN(n10761) );
  NOR2X0 U10572 ( .IN1(n10764), .IN2(n10765), .QN(n10763) );
  NOR2X0 U10573 ( .IN1(n10024), .IN2(n10766), .QN(n10765) );
  NOR2X0 U10574 ( .IN1(n10767), .IN2(g83), .QN(n10764) );
  NOR2X0 U10575 ( .IN1(n10768), .IN2(n10769), .QN(n10762) );
  NOR2X0 U10576 ( .IN1(n9603), .IN2(n10770), .QN(n10769) );
  NOR2X0 U10577 ( .IN1(n10771), .IN2(g56), .QN(n10768) );
  NAND2X0 U10578 ( .IN1(n10772), .IN2(n10773), .QN(n10760) );
  NAND2X0 U10579 ( .IN1(n10023), .IN2(n10774), .QN(n10773) );
  NAND2X0 U10580 ( .IN1(n10775), .IN2(g74), .QN(n10772) );
  NAND2X0 U10581 ( .IN1(n10776), .IN2(n10777), .QN(n10740) );
  NOR2X0 U10582 ( .IN1(n10778), .IN2(n10779), .QN(n10777) );
  NAND2X0 U10583 ( .IN1(n10780), .IN2(n10781), .QN(n10779) );
  NOR2X0 U10584 ( .IN1(n10782), .IN2(n10783), .QN(n10778) );
  NOR2X0 U10585 ( .IN1(test_so15), .IN2(n10784), .QN(n10783) );
  INVX0 U10586 ( .INP(n10785), .ZN(n10782) );
  NAND2X0 U10587 ( .IN1(n10784), .IN2(test_so15), .QN(n10785) );
  NOR2X0 U10588 ( .IN1(n10786), .IN2(n10787), .QN(n10776) );
  NAND2X0 U10589 ( .IN1(n10788), .IN2(n10789), .QN(n10787) );
  NOR2X0 U10590 ( .IN1(n10790), .IN2(n10791), .QN(n10789) );
  NOR2X0 U10591 ( .IN1(n9432), .IN2(n10792), .QN(n10791) );
  NOR2X0 U10592 ( .IN1(n10793), .IN2(g52), .QN(n10790) );
  NOR2X0 U10593 ( .IN1(n10794), .IN2(n10795), .QN(n10788) );
  NOR2X0 U10594 ( .IN1(n10025), .IN2(n10796), .QN(n10795) );
  NOR2X0 U10595 ( .IN1(n4513), .IN2(g92), .QN(n10794) );
  NAND2X0 U10596 ( .IN1(n10797), .IN2(n10798), .QN(n10786) );
  NAND2X0 U10597 ( .IN1(n10317), .IN2(n10799), .QN(n10798) );
  NAND2X0 U10598 ( .IN1(n10800), .IN2(g70), .QN(n10797) );
  NOR2X0 U10599 ( .IN1(n10801), .IN2(n10802), .QN(n4277) );
  NOR2X0 U10600 ( .IN1(n10803), .IN2(n10804), .QN(n10802) );
  NOR2X0 U10601 ( .IN1(n10805), .IN2(n10806), .QN(n10801) );
  NAND2X0 U10602 ( .IN1(n10807), .IN2(n10808), .QN(n10806) );
  NOR2X0 U10603 ( .IN1(n10809), .IN2(n10810), .QN(n10808) );
  NAND2X0 U10604 ( .IN1(n10811), .IN2(n10812), .QN(n10810) );
  NOR2X0 U10605 ( .IN1(n10813), .IN2(n10814), .QN(n10812) );
  NOR2X0 U10606 ( .IN1(n10018), .IN2(n10815), .QN(n10814) );
  NOR2X0 U10607 ( .IN1(n10816), .IN2(g753), .QN(n10813) );
  NOR2X0 U10608 ( .IN1(n10817), .IN2(n10818), .QN(n10811) );
  NOR2X0 U10609 ( .IN1(n10316), .IN2(n10819), .QN(n10818) );
  NOR2X0 U10610 ( .IN1(n10820), .IN2(g758), .QN(n10817) );
  NAND2X0 U10611 ( .IN1(n10821), .IN2(n10822), .QN(n10809) );
  NAND2X0 U10612 ( .IN1(n10019), .IN2(n10823), .QN(n10822) );
  NAND2X0 U10613 ( .IN1(n10824), .IN2(g762), .QN(n10821) );
  NOR2X0 U10614 ( .IN1(n10825), .IN2(n10826), .QN(n10807) );
  NAND2X0 U10615 ( .IN1(n10827), .IN2(n10828), .QN(n10826) );
  NOR2X0 U10616 ( .IN1(n10829), .IN2(n10830), .QN(n10828) );
  NOR2X0 U10617 ( .IN1(n10021), .IN2(n10831), .QN(n10830) );
  NOR2X0 U10618 ( .IN1(n10832), .IN2(g780), .QN(n10829) );
  NOR2X0 U10619 ( .IN1(n10833), .IN2(n10834), .QN(n10827) );
  NOR2X0 U10620 ( .IN1(n10314), .IN2(n10835), .QN(n10834) );
  NOR2X0 U10621 ( .IN1(n10836), .IN2(g776), .QN(n10833) );
  NAND2X0 U10622 ( .IN1(n10837), .IN2(n10838), .QN(n10825) );
  NAND2X0 U10623 ( .IN1(n10315), .IN2(n10839), .QN(n10838) );
  NAND2X0 U10624 ( .IN1(n10840), .IN2(g767), .QN(n10837) );
  NAND2X0 U10625 ( .IN1(n10841), .IN2(n10842), .QN(n10805) );
  NOR2X0 U10626 ( .IN1(n10843), .IN2(n10844), .QN(n10842) );
  NAND2X0 U10627 ( .IN1(n10845), .IN2(n10780), .QN(n10844) );
  NOR2X0 U10628 ( .IN1(n10846), .IN2(n10847), .QN(n10843) );
  NOR2X0 U10629 ( .IN1(test_so36), .IN2(n10848), .QN(n10847) );
  INVX0 U10630 ( .INP(n10849), .ZN(n10846) );
  NAND2X0 U10631 ( .IN1(n10848), .IN2(test_so36), .QN(n10849) );
  NOR2X0 U10632 ( .IN1(n10850), .IN2(n10851), .QN(n10841) );
  NAND2X0 U10633 ( .IN1(n10852), .IN2(n10853), .QN(n10851) );
  NOR2X0 U10634 ( .IN1(n10854), .IN2(n10855), .QN(n10853) );
  NOR2X0 U10635 ( .IN1(n9431), .IN2(n10856), .QN(n10855) );
  NOR2X0 U10636 ( .IN1(n10857), .IN2(g740), .QN(n10854) );
  NOR2X0 U10637 ( .IN1(n10858), .IN2(n10859), .QN(n10852) );
  NOR2X0 U10638 ( .IN1(n10020), .IN2(n10860), .QN(n10859) );
  NOR2X0 U10639 ( .IN1(n10861), .IN2(g771), .QN(n10858) );
  NAND2X0 U10640 ( .IN1(n10862), .IN2(n10863), .QN(n10850) );
  NAND2X0 U10641 ( .IN1(n9602), .IN2(n10864), .QN(n10863) );
  NAND2X0 U10642 ( .IN1(n10865), .IN2(g744), .QN(n10862) );
  NOR2X0 U10643 ( .IN1(n10866), .IN2(n10867), .QN(n4276) );
  NOR2X0 U10644 ( .IN1(n10868), .IN2(n10869), .QN(n10867) );
  NOR2X0 U10645 ( .IN1(n10870), .IN2(n10871), .QN(n10866) );
  NAND2X0 U10646 ( .IN1(n10872), .IN2(n10873), .QN(n10871) );
  NOR2X0 U10647 ( .IN1(n10874), .IN2(n10875), .QN(n10873) );
  NAND2X0 U10648 ( .IN1(n10876), .IN2(n10877), .QN(n10875) );
  NOR2X0 U10649 ( .IN1(n10878), .IN2(n10879), .QN(n10877) );
  NOR2X0 U10650 ( .IN1(n10014), .IN2(n10880), .QN(n10879) );
  NOR2X0 U10651 ( .IN1(n10881), .IN2(g1439), .QN(n10878) );
  NOR2X0 U10652 ( .IN1(n10882), .IN2(n10883), .QN(n10876) );
  NOR2X0 U10653 ( .IN1(n10309), .IN2(n10884), .QN(n10883) );
  NOR2X0 U10654 ( .IN1(n10885), .IN2(g1435), .QN(n10882) );
  NAND2X0 U10655 ( .IN1(n10886), .IN2(n10887), .QN(n10874) );
  NAND2X0 U10656 ( .IN1(n10017), .IN2(n10888), .QN(n10887) );
  NAND2X0 U10657 ( .IN1(n10889), .IN2(g1466), .QN(n10886) );
  NOR2X0 U10658 ( .IN1(n10890), .IN2(n10891), .QN(n10872) );
  NAND2X0 U10659 ( .IN1(n10892), .IN2(n10893), .QN(n10891) );
  NOR2X0 U10660 ( .IN1(n10894), .IN2(n10895), .QN(n10893) );
  NOR2X0 U10661 ( .IN1(n10016), .IN2(n10896), .QN(n10895) );
  NOR2X0 U10662 ( .IN1(n10897), .IN2(g1457), .QN(n10894) );
  NOR2X0 U10663 ( .IN1(n10898), .IN2(n10899), .QN(n10892) );
  NOR2X0 U10664 ( .IN1(n9601), .IN2(n10900), .QN(n10899) );
  NOR2X0 U10665 ( .IN1(n10901), .IN2(g1430), .QN(n10898) );
  NAND2X0 U10666 ( .IN1(n10902), .IN2(n10903), .QN(n10890) );
  NAND2X0 U10667 ( .IN1(n10015), .IN2(n10904), .QN(n10903) );
  NAND2X0 U10668 ( .IN1(n10905), .IN2(g1448), .QN(n10902) );
  NAND2X0 U10669 ( .IN1(n10906), .IN2(n10907), .QN(n10870) );
  NOR2X0 U10670 ( .IN1(n10908), .IN2(n10909), .QN(n10907) );
  NAND2X0 U10671 ( .IN1(n10910), .IN2(n10780), .QN(n10909) );
  NAND2X0 U10672 ( .IN1(n10911), .IN2(n10912), .QN(n10908) );
  NAND2X0 U10673 ( .IN1(n10312), .IN2(n10913), .QN(n10912) );
  NAND2X0 U10674 ( .IN1(n10914), .IN2(g1453), .QN(n10911) );
  NOR2X0 U10675 ( .IN1(n10915), .IN2(n10916), .QN(n10906) );
  NAND2X0 U10676 ( .IN1(n10917), .IN2(n10918), .QN(n10916) );
  NOR2X0 U10677 ( .IN1(n10919), .IN2(n10920), .QN(n10918) );
  NOR2X0 U10678 ( .IN1(n10307), .IN2(n10921), .QN(n10920) );
  NOR2X0 U10679 ( .IN1(n10922), .IN2(g1462), .QN(n10919) );
  NOR2X0 U10680 ( .IN1(n10923), .IN2(n10924), .QN(n10917) );
  NOR2X0 U10681 ( .IN1(n10318), .IN2(n10925), .QN(n10924) );
  NOR2X0 U10682 ( .IN1(n10926), .IN2(g1444), .QN(n10923) );
  NAND2X0 U10683 ( .IN1(n10927), .IN2(n10928), .QN(n10915) );
  NAND2X0 U10684 ( .IN1(n9430), .IN2(n10929), .QN(n10928) );
  NAND2X0 U10685 ( .IN1(n10930), .IN2(g1426), .QN(n10927) );
  NOR2X0 U10686 ( .IN1(n10931), .IN2(n10932), .QN(n4275) );
  NOR2X0 U10687 ( .IN1(n10933), .IN2(n10934), .QN(n10932) );
  NOR2X0 U10688 ( .IN1(n10935), .IN2(n10936), .QN(n10931) );
  NAND2X0 U10689 ( .IN1(n10937), .IN2(n10938), .QN(n10936) );
  NOR2X0 U10690 ( .IN1(n10939), .IN2(n10940), .QN(n10938) );
  NAND2X0 U10691 ( .IN1(n10941), .IN2(n10942), .QN(n10940) );
  NOR2X0 U10692 ( .IN1(n10943), .IN2(n10944), .QN(n10942) );
  NOR2X0 U10693 ( .IN1(n10010), .IN2(n10945), .QN(n10944) );
  NOR2X0 U10694 ( .IN1(n10946), .IN2(g2133), .QN(n10943) );
  NOR2X0 U10695 ( .IN1(n10947), .IN2(n10948), .QN(n10941) );
  NOR2X0 U10696 ( .IN1(n10310), .IN2(n10949), .QN(n10948) );
  NOR2X0 U10697 ( .IN1(n10950), .IN2(g2129), .QN(n10947) );
  NAND2X0 U10698 ( .IN1(n10951), .IN2(n10952), .QN(n10939) );
  NAND2X0 U10699 ( .IN1(n10013), .IN2(n10953), .QN(n10952) );
  NAND2X0 U10700 ( .IN1(n10954), .IN2(g2160), .QN(n10951) );
  NOR2X0 U10701 ( .IN1(n10955), .IN2(n10956), .QN(n10937) );
  NAND2X0 U10702 ( .IN1(n10957), .IN2(n10958), .QN(n10956) );
  NOR2X0 U10703 ( .IN1(n10959), .IN2(n10960), .QN(n10958) );
  NOR2X0 U10704 ( .IN1(n10012), .IN2(n10961), .QN(n10960) );
  NOR2X0 U10705 ( .IN1(n10962), .IN2(g2151), .QN(n10959) );
  NOR2X0 U10706 ( .IN1(n10963), .IN2(n10964), .QN(n10957) );
  NOR2X0 U10707 ( .IN1(n9600), .IN2(n10965), .QN(n10964) );
  NOR2X0 U10708 ( .IN1(n10966), .IN2(g2124), .QN(n10963) );
  NAND2X0 U10709 ( .IN1(n10967), .IN2(n10968), .QN(n10955) );
  NAND2X0 U10710 ( .IN1(n10011), .IN2(n10969), .QN(n10968) );
  NAND2X0 U10711 ( .IN1(n10970), .IN2(g2142), .QN(n10967) );
  NAND2X0 U10712 ( .IN1(n10971), .IN2(n10972), .QN(n10935) );
  NOR2X0 U10713 ( .IN1(n10973), .IN2(n10974), .QN(n10972) );
  NAND2X0 U10714 ( .IN1(n10975), .IN2(n10780), .QN(n10974) );
  NOR2X0 U10715 ( .IN1(n10976), .IN2(n10977), .QN(n10973) );
  NOR2X0 U10716 ( .IN1(test_so78), .IN2(n10978), .QN(n10977) );
  INVX0 U10717 ( .INP(n10979), .ZN(n10976) );
  NAND2X0 U10718 ( .IN1(n10978), .IN2(test_so78), .QN(n10979) );
  NOR2X0 U10719 ( .IN1(n10980), .IN2(n10981), .QN(n10971) );
  NAND2X0 U10720 ( .IN1(n10982), .IN2(n10983), .QN(n10981) );
  NOR2X0 U10721 ( .IN1(n10984), .IN2(n10985), .QN(n10983) );
  NOR2X0 U10722 ( .IN1(n9429), .IN2(n10986), .QN(n10985) );
  NOR2X0 U10723 ( .IN1(n10987), .IN2(g2120), .QN(n10984) );
  NOR2X0 U10724 ( .IN1(n10988), .IN2(n10989), .QN(n10982) );
  NOR2X0 U10725 ( .IN1(n10313), .IN2(n10990), .QN(n10989) );
  NOR2X0 U10726 ( .IN1(n10991), .IN2(g2147), .QN(n10988) );
  NAND2X0 U10727 ( .IN1(n10992), .IN2(n10993), .QN(n10980) );
  NAND2X0 U10728 ( .IN1(n10319), .IN2(n10994), .QN(n10993) );
  NAND2X0 U10729 ( .IN1(n10995), .IN2(g2138), .QN(n10992) );
  NAND2X0 U10730 ( .IN1(n10996), .IN2(n10997), .QN(n4274) );
  INVX0 U10731 ( .INP(n10998), .ZN(n10997) );
  NOR2X0 U10732 ( .IN1(n10999), .IN2(n11000), .QN(n10996) );
  NOR2X0 U10733 ( .IN1(n4423), .IN2(g2883), .QN(n11000) );
  NOR2X0 U10734 ( .IN1(n4330), .IN2(g2950), .QN(n10999) );
  NAND2X0 U10735 ( .IN1(n11001), .IN2(n11002), .QN(n4273) );
  NAND2X0 U10736 ( .IN1(n11003), .IN2(n11004), .QN(n11002) );
  NAND2X0 U10737 ( .IN1(n4482), .IN2(n11005), .QN(n11003) );
  NAND2X0 U10738 ( .IN1(n2426), .IN2(n11006), .QN(n4272) );
  NAND2X0 U10739 ( .IN1(n11007), .IN2(n11008), .QN(n11006) );
  NOR2X0 U10740 ( .IN1(n11009), .IN2(n11010), .QN(n11007) );
  NOR2X0 U10741 ( .IN1(test_so27), .IN2(n11011), .QN(n11010) );
  NOR2X0 U10742 ( .IN1(n11012), .IN2(n11013), .QN(n11009) );
  NAND2X0 U10743 ( .IN1(n11014), .IN2(n11015), .QN(n4271) );
  NAND2X0 U10744 ( .IN1(n2446), .IN2(n11016), .QN(n11015) );
  NAND2X0 U10745 ( .IN1(n11017), .IN2(n11008), .QN(n11014) );
  NOR2X0 U10746 ( .IN1(n11018), .IN2(n11019), .QN(n11017) );
  NOR2X0 U10747 ( .IN1(n11011), .IN2(g536), .QN(n11019) );
  NOR2X0 U10748 ( .IN1(n11012), .IN2(n11020), .QN(n11018) );
  NAND2X0 U10749 ( .IN1(n11021), .IN2(n11022), .QN(n4270) );
  NAND2X0 U10750 ( .IN1(n2446), .IN2(n11023), .QN(n11022) );
  NAND2X0 U10751 ( .IN1(n11024), .IN2(n11008), .QN(n11021) );
  NOR2X0 U10752 ( .IN1(n11025), .IN2(n11026), .QN(n11024) );
  NOR2X0 U10753 ( .IN1(n11011), .IN2(g537), .QN(n11026) );
  NOR2X0 U10754 ( .IN1(n11012), .IN2(n11027), .QN(n11025) );
  NAND2X0 U10755 ( .IN1(n11028), .IN2(n11029), .QN(n4269) );
  NAND2X0 U10756 ( .IN1(n11030), .IN2(n11008), .QN(n11029) );
  NOR2X0 U10757 ( .IN1(n11031), .IN2(n11032), .QN(n11030) );
  NOR2X0 U10758 ( .IN1(n11011), .IN2(n8047), .QN(n11032) );
  NOR2X0 U10759 ( .IN1(n11012), .IN2(n11033), .QN(n11031) );
  NAND2X0 U10760 ( .IN1(n11034), .IN2(n2440), .QN(n4268) );
  NOR2X0 U10761 ( .IN1(n11035), .IN2(n11036), .QN(n11034) );
  NOR2X0 U10762 ( .IN1(n11037), .IN2(n11038), .QN(n11035) );
  NAND2X0 U10763 ( .IN1(n11039), .IN2(n11040), .QN(n11038) );
  NAND2X0 U10764 ( .IN1(n11041), .IN2(n11042), .QN(n11040) );
  NAND2X0 U10765 ( .IN1(n11043), .IN2(DFF_445_n1), .QN(n11039) );
  NAND2X0 U10766 ( .IN1(n11044), .IN2(n2440), .QN(n4267) );
  NOR2X0 U10767 ( .IN1(n11045), .IN2(n11036), .QN(n11044) );
  NOR2X0 U10768 ( .IN1(n11037), .IN2(n11046), .QN(n11045) );
  NAND2X0 U10769 ( .IN1(n11047), .IN2(n11048), .QN(n11046) );
  NAND2X0 U10770 ( .IN1(n11049), .IN2(n11042), .QN(n11048) );
  NAND2X0 U10771 ( .IN1(n11043), .IN2(DFF_446_n1), .QN(n11047) );
  NAND2X0 U10772 ( .IN1(n11028), .IN2(n11050), .QN(n4266) );
  NAND2X0 U10773 ( .IN1(n11051), .IN2(n11008), .QN(n11050) );
  NOR2X0 U10774 ( .IN1(n11052), .IN2(n11053), .QN(n11051) );
  NOR2X0 U10775 ( .IN1(n11011), .IN2(n8044), .QN(n11053) );
  NOR2X0 U10776 ( .IN1(n11012), .IN2(n11054), .QN(n11052) );
  NOR2X0 U10777 ( .IN1(n11036), .IN2(n11055), .QN(n11028) );
  INVX0 U10778 ( .INP(n11056), .ZN(n11055) );
  NAND2X0 U10779 ( .IN1(n2446), .IN2(n2445), .QN(n11056) );
  INVX0 U10780 ( .INP(n2426), .ZN(n11036) );
  NAND2X0 U10781 ( .IN1(n2426), .IN2(n11057), .QN(n4265) );
  NAND2X0 U10782 ( .IN1(n11058), .IN2(n11008), .QN(n11057) );
  NOR2X0 U10783 ( .IN1(n11059), .IN2(n11060), .QN(n11058) );
  NOR2X0 U10784 ( .IN1(n11011), .IN2(n8043), .QN(n11060) );
  INVX0 U10785 ( .INP(n11043), .ZN(n11011) );
  NOR2X0 U10786 ( .IN1(n11012), .IN2(n11061), .QN(n11059) );
  INVX0 U10787 ( .INP(n11042), .ZN(n11012) );
  NAND2X0 U10788 ( .IN1(DFF_1562_n1), .IN2(n11062), .QN(n4263) );
  NAND2X0 U10789 ( .IN1(n11063), .IN2(n11064), .QN(n4262) );
  NAND2X0 U10790 ( .IN1(n11065), .IN2(n11066), .QN(n11063) );
  NAND2X0 U10791 ( .IN1(n4481), .IN2(n11067), .QN(n11066) );
  NOR2X0 U10792 ( .IN1(n11068), .IN2(n11069), .QN(n4261) );
  NOR2X0 U10793 ( .IN1(n11070), .IN2(n11071), .QN(n11069) );
  NOR2X0 U10794 ( .IN1(n11072), .IN2(n11073), .QN(n11068) );
  INVX0 U10795 ( .INP(n11071), .ZN(n11072) );
  NAND2X0 U10796 ( .IN1(n11074), .IN2(n11075), .QN(n4260) );
  NAND2X0 U10797 ( .IN1(n11070), .IN2(n11076), .QN(n11075) );
  NAND2X0 U10798 ( .IN1(n11077), .IN2(n11073), .QN(n11074) );
  INVX0 U10799 ( .INP(n11070), .ZN(n11073) );
  NOR2X0 U10800 ( .IN1(g3231), .IN2(n18871), .QN(n11070) );
  INVX0 U10801 ( .INP(n11076), .ZN(n11077) );
  NAND2X0 U10802 ( .IN1(n11078), .IN2(n11079), .QN(n4259) );
  NAND2X0 U10803 ( .IN1(n11080), .IN2(test_so22), .QN(n11079) );
  NOR2X0 U10804 ( .IN1(n11081), .IN2(n11082), .QN(n11080) );
  INVX0 U10805 ( .INP(n11083), .ZN(n11082) );
  NAND2X0 U10806 ( .IN1(n11084), .IN2(n11085), .QN(n11083) );
  NOR2X0 U10807 ( .IN1(n11085), .IN2(n11084), .QN(n11081) );
  NOR2X0 U10808 ( .IN1(n11086), .IN2(n11087), .QN(n11084) );
  NOR2X0 U10809 ( .IN1(n11088), .IN2(n11020), .QN(n11087) );
  INVX0 U10810 ( .INP(n11089), .ZN(n11086) );
  NAND2X0 U10811 ( .IN1(n11088), .IN2(n11020), .QN(n11089) );
  NAND2X0 U10812 ( .IN1(n11090), .IN2(n11091), .QN(n11020) );
  NOR2X0 U10813 ( .IN1(n11092), .IN2(n11093), .QN(n11090) );
  NOR2X0 U10814 ( .IN1(n11094), .IN2(n11095), .QN(n11093) );
  NOR2X0 U10815 ( .IN1(n11096), .IN2(n11097), .QN(n11092) );
  NAND2X0 U10816 ( .IN1(n11098), .IN2(n11099), .QN(n11088) );
  NAND2X0 U10817 ( .IN1(n11049), .IN2(n11100), .QN(n11099) );
  INVX0 U10818 ( .INP(n11101), .ZN(n11098) );
  NOR2X0 U10819 ( .IN1(n11100), .IN2(n11049), .QN(n11101) );
  INVX0 U10820 ( .INP(n11102), .ZN(n11049) );
  NAND2X0 U10821 ( .IN1(n11103), .IN2(n11104), .QN(n11102) );
  NOR2X0 U10822 ( .IN1(n11105), .IN2(n11106), .QN(n11103) );
  NOR2X0 U10823 ( .IN1(n11107), .IN2(n11095), .QN(n11106) );
  NOR2X0 U10824 ( .IN1(n11096), .IN2(n11108), .QN(n11105) );
  NAND2X0 U10825 ( .IN1(n11109), .IN2(n11110), .QN(n11100) );
  NAND2X0 U10826 ( .IN1(n11111), .IN2(n11112), .QN(n11110) );
  NAND2X0 U10827 ( .IN1(n11113), .IN2(n11114), .QN(n11112) );
  NAND2X0 U10828 ( .IN1(n11115), .IN2(n11033), .QN(n11114) );
  NAND2X0 U10829 ( .IN1(n11116), .IN2(n11013), .QN(n11113) );
  NOR2X0 U10830 ( .IN1(n11117), .IN2(n11118), .QN(n11111) );
  NOR2X0 U10831 ( .IN1(n11041), .IN2(n11054), .QN(n11118) );
  NOR2X0 U10832 ( .IN1(n11119), .IN2(n11120), .QN(n11117) );
  NAND2X0 U10833 ( .IN1(n11121), .IN2(n11122), .QN(n11109) );
  NAND2X0 U10834 ( .IN1(n11123), .IN2(n11124), .QN(n11122) );
  NAND2X0 U10835 ( .IN1(n11041), .IN2(n11054), .QN(n11124) );
  INVX0 U10836 ( .INP(n11120), .ZN(n11041) );
  NAND2X0 U10837 ( .IN1(n11119), .IN2(n11120), .QN(n11123) );
  NAND2X0 U10838 ( .IN1(n11125), .IN2(n11104), .QN(n11120) );
  NOR2X0 U10839 ( .IN1(n11126), .IN2(n11127), .QN(n11125) );
  NOR2X0 U10840 ( .IN1(n11128), .IN2(n11129), .QN(n11127) );
  NOR2X0 U10841 ( .IN1(n11130), .IN2(n11131), .QN(n11126) );
  INVX0 U10842 ( .INP(n11054), .ZN(n11119) );
  NAND2X0 U10843 ( .IN1(n11132), .IN2(n11104), .QN(n11054) );
  NOR2X0 U10844 ( .IN1(n11133), .IN2(n11134), .QN(n11132) );
  NOR2X0 U10845 ( .IN1(n11135), .IN2(n11129), .QN(n11134) );
  NOR2X0 U10846 ( .IN1(n11130), .IN2(n11136), .QN(n11133) );
  NOR2X0 U10847 ( .IN1(n11137), .IN2(n11138), .QN(n11121) );
  NOR2X0 U10848 ( .IN1(n11115), .IN2(n11033), .QN(n11138) );
  INVX0 U10849 ( .INP(n11013), .ZN(n11115) );
  NOR2X0 U10850 ( .IN1(n11116), .IN2(n11013), .QN(n11137) );
  NAND2X0 U10851 ( .IN1(n11139), .IN2(n11140), .QN(n11013) );
  NOR2X0 U10852 ( .IN1(n11141), .IN2(n11142), .QN(n11139) );
  NOR2X0 U10853 ( .IN1(n11143), .IN2(n11129), .QN(n11142) );
  NOR2X0 U10854 ( .IN1(n11130), .IN2(n11144), .QN(n11141) );
  INVX0 U10855 ( .INP(n11033), .ZN(n11116) );
  NAND2X0 U10856 ( .IN1(n11145), .IN2(n11104), .QN(n11033) );
  NOR2X0 U10857 ( .IN1(n11146), .IN2(n11147), .QN(n11145) );
  NOR2X0 U10858 ( .IN1(n11148), .IN2(n11095), .QN(n11147) );
  NOR2X0 U10859 ( .IN1(n11096), .IN2(n11149), .QN(n11146) );
  NAND2X0 U10860 ( .IN1(n11150), .IN2(n11151), .QN(n11085) );
  INVX0 U10861 ( .INP(n11152), .ZN(n11151) );
  NOR2X0 U10862 ( .IN1(n11027), .IN2(n11153), .QN(n11152) );
  NAND2X0 U10863 ( .IN1(n11153), .IN2(n11027), .QN(n11150) );
  NAND2X0 U10864 ( .IN1(n11154), .IN2(n11104), .QN(n11027) );
  NOR2X0 U10865 ( .IN1(n11155), .IN2(n11156), .QN(n11154) );
  NOR2X0 U10866 ( .IN1(n11157), .IN2(n11129), .QN(n11156) );
  NOR2X0 U10867 ( .IN1(n11130), .IN2(n11158), .QN(n11155) );
  INVX0 U10868 ( .INP(n11061), .ZN(n11153) );
  NAND2X0 U10869 ( .IN1(n11159), .IN2(n11091), .QN(n11061) );
  NOR2X0 U10870 ( .IN1(n11160), .IN2(n11161), .QN(n11159) );
  NOR2X0 U10871 ( .IN1(n11162), .IN2(n11095), .QN(n11161) );
  NOR2X0 U10872 ( .IN1(n11096), .IN2(n11163), .QN(n11160) );
  NOR2X0 U10873 ( .IN1(n11164), .IN2(n11165), .QN(n11078) );
  NOR2X0 U10874 ( .IN1(n4360), .IN2(n11166), .QN(n11165) );
  NOR2X0 U10875 ( .IN1(n11167), .IN2(n11168), .QN(n11166) );
  NOR2X0 U10876 ( .IN1(n11169), .IN2(n11023), .QN(n11168) );
  INVX0 U10877 ( .INP(n11016), .ZN(n11169) );
  NOR2X0 U10878 ( .IN1(n11170), .IN2(n11016), .QN(n11167) );
  NAND2X0 U10879 ( .IN1(n11171), .IN2(n11091), .QN(n11016) );
  INVX0 U10880 ( .INP(n11172), .ZN(n11091) );
  NAND2X0 U10881 ( .IN1(n11104), .IN2(n567), .QN(n11172) );
  NAND2X0 U10882 ( .IN1(n11173), .IN2(n11174), .QN(n567) );
  NOR2X0 U10883 ( .IN1(n11175), .IN2(n11176), .QN(n11171) );
  NOR2X0 U10884 ( .IN1(n11177), .IN2(n11095), .QN(n11176) );
  NAND2X0 U10885 ( .IN1(n11096), .IN2(n11178), .QN(n11095) );
  NOR2X0 U10886 ( .IN1(n11096), .IN2(n11179), .QN(n11175) );
  INVX0 U10887 ( .INP(n11023), .ZN(n11170) );
  NAND2X0 U10888 ( .IN1(n11180), .IN2(n11140), .QN(n11023) );
  INVX0 U10889 ( .INP(n11181), .ZN(n11140) );
  NAND2X0 U10890 ( .IN1(n11104), .IN2(n11182), .QN(n11181) );
  NAND2X0 U10891 ( .IN1(n11173), .IN2(n11183), .QN(n11182) );
  NOR2X0 U10892 ( .IN1(n10725), .IN2(n4541), .QN(n11104) );
  NOR2X0 U10893 ( .IN1(n11184), .IN2(n11185), .QN(n11180) );
  NOR2X0 U10894 ( .IN1(n11186), .IN2(n11129), .QN(n11185) );
  NAND2X0 U10895 ( .IN1(n11130), .IN2(n11178), .QN(n11129) );
  NOR2X0 U10896 ( .IN1(n11130), .IN2(n11187), .QN(n11184) );
  NOR2X0 U10897 ( .IN1(n11188), .IN2(n11189), .QN(n11164) );
  NAND2X0 U10898 ( .IN1(n11008), .IN2(n11043), .QN(n11189) );
  NOR2X0 U10899 ( .IN1(n11042), .IN2(n10725), .QN(n11043) );
  NAND2X0 U10900 ( .IN1(n11190), .IN2(n11191), .QN(n10725) );
  NOR2X0 U10901 ( .IN1(g563), .IN2(n11192), .QN(n11191) );
  NOR2X0 U10902 ( .IN1(n4298), .IN2(g499), .QN(n11192) );
  NOR2X0 U10903 ( .IN1(g559), .IN2(g21851), .QN(n11190) );
  NAND2X0 U10904 ( .IN1(n11193), .IN2(n11194), .QN(n11188) );
  NAND2X0 U10905 ( .IN1(n18855), .IN2(n11195), .QN(n11194) );
  NAND2X0 U10906 ( .IN1(n4492), .IN2(g3229), .QN(n11193) );
  NAND2X0 U10907 ( .IN1(n11196), .IN2(n11197), .QN(n4258) );
  NAND2X0 U10908 ( .IN1(n2361), .IN2(n11198), .QN(n11197) );
  NAND2X0 U10909 ( .IN1(n11199), .IN2(n11200), .QN(n11196) );
  NOR2X0 U10910 ( .IN1(n11201), .IN2(n11202), .QN(n11199) );
  NOR2X0 U10911 ( .IN1(n11203), .IN2(g2611), .QN(n11202) );
  NOR2X0 U10912 ( .IN1(n11204), .IN2(n11205), .QN(n11201) );
  NAND2X0 U10913 ( .IN1(n11206), .IN2(n2375), .QN(n4257) );
  NOR2X0 U10914 ( .IN1(n11207), .IN2(n11208), .QN(n11206) );
  NOR2X0 U10915 ( .IN1(n11209), .IN2(n11210), .QN(n11208) );
  NAND2X0 U10916 ( .IN1(n11211), .IN2(n11212), .QN(n11210) );
  NAND2X0 U10917 ( .IN1(n11213), .IN2(n11214), .QN(n11212) );
  NAND2X0 U10918 ( .IN1(n11215), .IN2(DFF_1495_n1), .QN(n11211) );
  NAND2X0 U10919 ( .IN1(n11216), .IN2(n11217), .QN(n4256) );
  NAND2X0 U10920 ( .IN1(n11218), .IN2(n11200), .QN(n11217) );
  NOR2X0 U10921 ( .IN1(n11219), .IN2(n11220), .QN(n11218) );
  NOR2X0 U10922 ( .IN1(n11203), .IN2(n7920), .QN(n11220) );
  NOR2X0 U10923 ( .IN1(n11204), .IN2(n11221), .QN(n11219) );
  NAND2X0 U10924 ( .IN1(n11222), .IN2(n2375), .QN(n4255) );
  NOR2X0 U10925 ( .IN1(n11207), .IN2(n11223), .QN(n11222) );
  NOR2X0 U10926 ( .IN1(n11209), .IN2(n11224), .QN(n11223) );
  NAND2X0 U10927 ( .IN1(n11225), .IN2(n11226), .QN(n11224) );
  NAND2X0 U10928 ( .IN1(n11227), .IN2(n11214), .QN(n11226) );
  NAND2X0 U10929 ( .IN1(n11215), .IN2(DFF_1496_n1), .QN(n11225) );
  NAND2X0 U10930 ( .IN1(n11228), .IN2(n11229), .QN(n4254) );
  NAND2X0 U10931 ( .IN1(n11230), .IN2(n11200), .QN(n11229) );
  NOR2X0 U10932 ( .IN1(n11231), .IN2(n11232), .QN(n11230) );
  NOR2X0 U10933 ( .IN1(n11203), .IN2(n7925), .QN(n11232) );
  NOR2X0 U10934 ( .IN1(n11204), .IN2(n11233), .QN(n11231) );
  NAND2X0 U10935 ( .IN1(n11234), .IN2(n11235), .QN(n4253) );
  NAND2X0 U10936 ( .IN1(n2361), .IN2(n11236), .QN(n11235) );
  NAND2X0 U10937 ( .IN1(n11237), .IN2(n11200), .QN(n11234) );
  NOR2X0 U10938 ( .IN1(n11238), .IN2(n11239), .QN(n11237) );
  NOR2X0 U10939 ( .IN1(test_so91), .IN2(n11203), .QN(n11239) );
  NOR2X0 U10940 ( .IN1(n11204), .IN2(n11240), .QN(n11238) );
  NAND2X0 U10941 ( .IN1(n11228), .IN2(n11241), .QN(n4252) );
  NAND2X0 U10942 ( .IN1(n11242), .IN2(n11200), .QN(n11241) );
  NOR2X0 U10943 ( .IN1(n11243), .IN2(n11244), .QN(n11242) );
  NOR2X0 U10944 ( .IN1(n11203), .IN2(n7922), .QN(n11244) );
  NOR2X0 U10945 ( .IN1(n11204), .IN2(n11245), .QN(n11243) );
  NOR2X0 U10946 ( .IN1(n11207), .IN2(n11246), .QN(n11228) );
  INVX0 U10947 ( .INP(n11247), .ZN(n11246) );
  NAND2X0 U10948 ( .IN1(n2361), .IN2(n2374), .QN(n11247) );
  INVX0 U10949 ( .INP(n11216), .ZN(n11207) );
  NAND2X0 U10950 ( .IN1(n11216), .IN2(n11248), .QN(n4251) );
  NAND2X0 U10951 ( .IN1(n11249), .IN2(n11200), .QN(n11248) );
  NOR2X0 U10952 ( .IN1(n11250), .IN2(n11251), .QN(n11249) );
  NOR2X0 U10953 ( .IN1(n11203), .IN2(n7921), .QN(n11251) );
  INVX0 U10954 ( .INP(n11215), .ZN(n11203) );
  NOR2X0 U10955 ( .IN1(n11204), .IN2(n11252), .QN(n11250) );
  INVX0 U10956 ( .INP(n11214), .ZN(n11204) );
  NAND2X0 U10957 ( .IN1(n2361), .IN2(n11253), .QN(n11216) );
  NAND2X0 U10958 ( .IN1(n11254), .IN2(n11255), .QN(n4250) );
  NAND2X0 U10959 ( .IN1(n11256), .IN2(g2631), .QN(n11255) );
  NAND2X0 U10960 ( .IN1(n11257), .IN2(n11258), .QN(n11256) );
  NAND2X0 U10961 ( .IN1(n11259), .IN2(n11236), .QN(n11258) );
  INVX0 U10962 ( .INP(n11198), .ZN(n11259) );
  NAND2X0 U10963 ( .IN1(n11260), .IN2(n11198), .QN(n11257) );
  NAND2X0 U10964 ( .IN1(n11261), .IN2(n11262), .QN(n11198) );
  NOR2X0 U10965 ( .IN1(n11263), .IN2(n11264), .QN(n11261) );
  NOR2X0 U10966 ( .IN1(n11265), .IN2(n11266), .QN(n11264) );
  NOR2X0 U10967 ( .IN1(n11267), .IN2(n11268), .QN(n11263) );
  INVX0 U10968 ( .INP(n11236), .ZN(n11260) );
  NAND2X0 U10969 ( .IN1(n11269), .IN2(n11270), .QN(n11236) );
  NOR2X0 U10970 ( .IN1(n11271), .IN2(n11272), .QN(n11269) );
  NOR2X0 U10971 ( .IN1(n11273), .IN2(n11274), .QN(n11272) );
  NOR2X0 U10972 ( .IN1(n11275), .IN2(n11276), .QN(n11271) );
  NOR2X0 U10973 ( .IN1(n11277), .IN2(n11278), .QN(n11254) );
  NOR2X0 U10974 ( .IN1(n4303), .IN2(n11279), .QN(n11278) );
  NAND2X0 U10975 ( .IN1(n11280), .IN2(n11281), .QN(n11279) );
  INVX0 U10976 ( .INP(n11282), .ZN(n11281) );
  NOR2X0 U10977 ( .IN1(n11283), .IN2(n11284), .QN(n11282) );
  NAND2X0 U10978 ( .IN1(n11284), .IN2(n11283), .QN(n11280) );
  NOR2X0 U10979 ( .IN1(n11285), .IN2(n11286), .QN(n11283) );
  INVX0 U10980 ( .INP(n11287), .ZN(n11286) );
  NAND2X0 U10981 ( .IN1(n11288), .IN2(n11213), .QN(n11287) );
  NOR2X0 U10982 ( .IN1(n11288), .IN2(n11213), .QN(n11285) );
  INVX0 U10983 ( .INP(n11289), .ZN(n11213) );
  NAND2X0 U10984 ( .IN1(n11290), .IN2(n11291), .QN(n11289) );
  NOR2X0 U10985 ( .IN1(n11292), .IN2(n11293), .QN(n11290) );
  NOR2X0 U10986 ( .IN1(n11294), .IN2(n11266), .QN(n11293) );
  NOR2X0 U10987 ( .IN1(n11267), .IN2(n11295), .QN(n11292) );
  NOR2X0 U10988 ( .IN1(n11296), .IN2(n11297), .QN(n11288) );
  NOR2X0 U10989 ( .IN1(n11298), .IN2(n11227), .QN(n11297) );
  INVX0 U10990 ( .INP(n11299), .ZN(n11296) );
  NAND2X0 U10991 ( .IN1(n11227), .IN2(n11298), .QN(n11299) );
  NAND2X0 U10992 ( .IN1(n11300), .IN2(n11301), .QN(n11298) );
  NAND2X0 U10993 ( .IN1(n11302), .IN2(n11303), .QN(n11301) );
  NAND2X0 U10994 ( .IN1(n11304), .IN2(n11305), .QN(n11303) );
  NAND2X0 U10995 ( .IN1(n11306), .IN2(n11252), .QN(n11305) );
  NAND2X0 U10996 ( .IN1(n11307), .IN2(n11233), .QN(n11304) );
  NOR2X0 U10997 ( .IN1(n11308), .IN2(n11309), .QN(n11302) );
  NOR2X0 U10998 ( .IN1(n11310), .IN2(n11240), .QN(n11309) );
  NOR2X0 U10999 ( .IN1(n11311), .IN2(n11205), .QN(n11308) );
  NAND2X0 U11000 ( .IN1(n11312), .IN2(n11313), .QN(n11300) );
  NAND2X0 U11001 ( .IN1(n11314), .IN2(n11315), .QN(n11313) );
  NAND2X0 U11002 ( .IN1(n11310), .IN2(n11240), .QN(n11315) );
  INVX0 U11003 ( .INP(n11205), .ZN(n11310) );
  NAND2X0 U11004 ( .IN1(n11311), .IN2(n11205), .QN(n11314) );
  NAND2X0 U11005 ( .IN1(n11316), .IN2(n11291), .QN(n11205) );
  NOR2X0 U11006 ( .IN1(n11317), .IN2(n11318), .QN(n11316) );
  NOR2X0 U11007 ( .IN1(n11319), .IN2(n11266), .QN(n11318) );
  NOR2X0 U11008 ( .IN1(n11267), .IN2(n11320), .QN(n11317) );
  INVX0 U11009 ( .INP(n11240), .ZN(n11311) );
  NAND2X0 U11010 ( .IN1(n11321), .IN2(n11270), .QN(n11240) );
  NOR2X0 U11011 ( .IN1(n11322), .IN2(n11323), .QN(n11321) );
  NOR2X0 U11012 ( .IN1(n11324), .IN2(n11274), .QN(n11323) );
  NOR2X0 U11013 ( .IN1(n11275), .IN2(n11325), .QN(n11322) );
  NOR2X0 U11014 ( .IN1(n11326), .IN2(n11327), .QN(n11312) );
  NOR2X0 U11015 ( .IN1(n11306), .IN2(n11252), .QN(n11327) );
  INVX0 U11016 ( .INP(n11233), .ZN(n11306) );
  NOR2X0 U11017 ( .IN1(n11307), .IN2(n11233), .QN(n11326) );
  NAND2X0 U11018 ( .IN1(n11328), .IN2(n11291), .QN(n11233) );
  NOR2X0 U11019 ( .IN1(n11329), .IN2(n11330), .QN(n11328) );
  NOR2X0 U11020 ( .IN1(n11331), .IN2(n11274), .QN(n11330) );
  NOR2X0 U11021 ( .IN1(n11275), .IN2(n11332), .QN(n11329) );
  INVX0 U11022 ( .INP(n11252), .ZN(n11307) );
  NAND2X0 U11023 ( .IN1(n11333), .IN2(n11270), .QN(n11252) );
  INVX0 U11024 ( .INP(n11334), .ZN(n11270) );
  NAND2X0 U11025 ( .IN1(n11291), .IN2(n2351), .QN(n11334) );
  NOR2X0 U11026 ( .IN1(n11335), .IN2(n11336), .QN(n11333) );
  NOR2X0 U11027 ( .IN1(n11337), .IN2(n11274), .QN(n11336) );
  NOR2X0 U11028 ( .IN1(n11275), .IN2(n11338), .QN(n11335) );
  INVX0 U11029 ( .INP(n11339), .ZN(n11227) );
  NAND2X0 U11030 ( .IN1(n11340), .IN2(n11291), .QN(n11339) );
  NOR2X0 U11031 ( .IN1(n11341), .IN2(n11342), .QN(n11340) );
  NOR2X0 U11032 ( .IN1(n11343), .IN2(n11274), .QN(n11342) );
  NAND2X0 U11033 ( .IN1(n11275), .IN2(n11344), .QN(n11274) );
  NOR2X0 U11034 ( .IN1(n11275), .IN2(n11345), .QN(n11341) );
  NAND2X0 U11035 ( .IN1(n11346), .IN2(n11347), .QN(n11284) );
  INVX0 U11036 ( .INP(n11348), .ZN(n11347) );
  NOR2X0 U11037 ( .IN1(n11221), .IN2(n11349), .QN(n11348) );
  NAND2X0 U11038 ( .IN1(n11349), .IN2(n11221), .QN(n11346) );
  NAND2X0 U11039 ( .IN1(n11350), .IN2(n11262), .QN(n11221) );
  INVX0 U11040 ( .INP(n11351), .ZN(n11262) );
  NAND2X0 U11041 ( .IN1(n11291), .IN2(n11352), .QN(n11351) );
  NAND2X0 U11042 ( .IN1(n11353), .IN2(n11354), .QN(n11352) );
  NOR2X0 U11043 ( .IN1(n11355), .IN2(n11356), .QN(n11350) );
  NOR2X0 U11044 ( .IN1(n11357), .IN2(n11266), .QN(n11356) );
  NOR2X0 U11045 ( .IN1(n11267), .IN2(n11358), .QN(n11355) );
  INVX0 U11046 ( .INP(n11245), .ZN(n11349) );
  NAND2X0 U11047 ( .IN1(n11359), .IN2(n11291), .QN(n11245) );
  NOR2X0 U11048 ( .IN1(n11253), .IN2(n4543), .QN(n11291) );
  NOR2X0 U11049 ( .IN1(n11360), .IN2(n11361), .QN(n11359) );
  NOR2X0 U11050 ( .IN1(n11362), .IN2(n11266), .QN(n11361) );
  NAND2X0 U11051 ( .IN1(n11267), .IN2(n11344), .QN(n11266) );
  NOR2X0 U11052 ( .IN1(n11267), .IN2(n11363), .QN(n11360) );
  NOR2X0 U11053 ( .IN1(n11364), .IN2(n11365), .QN(n11277) );
  NAND2X0 U11054 ( .IN1(n11200), .IN2(n11215), .QN(n11365) );
  NOR2X0 U11055 ( .IN1(n11253), .IN2(n11214), .QN(n11215) );
  NAND2X0 U11056 ( .IN1(n11366), .IN2(n10076), .QN(n11253) );
  NOR2X0 U11057 ( .IN1(g2637), .IN2(g30072), .QN(n11366) );
  NAND2X0 U11058 ( .IN1(n11367), .IN2(n11368), .QN(n11364) );
  NAND2X0 U11059 ( .IN1(n18856), .IN2(n11195), .QN(n11368) );
  NAND2X0 U11060 ( .IN1(n4490), .IN2(g3229), .QN(n11367) );
  NAND2X0 U11061 ( .IN1(n11369), .IN2(n11370), .QN(n4249) );
  NAND2X0 U11062 ( .IN1(n2289), .IN2(n11371), .QN(n11370) );
  NAND2X0 U11063 ( .IN1(n11372), .IN2(n11373), .QN(n11369) );
  NOR2X0 U11064 ( .IN1(n11374), .IN2(n11375), .QN(n11372) );
  NOR2X0 U11065 ( .IN1(n11376), .IN2(g1917), .QN(n11375) );
  NOR2X0 U11066 ( .IN1(n11377), .IN2(n11378), .QN(n11374) );
  NAND2X0 U11067 ( .IN1(n11379), .IN2(n2303), .QN(n4248) );
  NOR2X0 U11068 ( .IN1(n11380), .IN2(n11381), .QN(n11379) );
  NOR2X0 U11069 ( .IN1(n11382), .IN2(n11383), .QN(n11380) );
  NAND2X0 U11070 ( .IN1(n11384), .IN2(n11385), .QN(n11383) );
  NAND2X0 U11071 ( .IN1(n11386), .IN2(n11387), .QN(n11385) );
  NAND2X0 U11072 ( .IN1(n11388), .IN2(DFF_1145_n1), .QN(n11384) );
  NAND2X0 U11073 ( .IN1(n2275), .IN2(n11389), .QN(n4247) );
  NAND2X0 U11074 ( .IN1(n11390), .IN2(n11373), .QN(n11389) );
  NOR2X0 U11075 ( .IN1(n11391), .IN2(n11392), .QN(n11390) );
  NOR2X0 U11076 ( .IN1(n11376), .IN2(n7962), .QN(n11392) );
  NOR2X0 U11077 ( .IN1(n11377), .IN2(n11393), .QN(n11391) );
  NAND2X0 U11078 ( .IN1(n11394), .IN2(n2303), .QN(n4246) );
  NOR2X0 U11079 ( .IN1(n11395), .IN2(n11381), .QN(n11394) );
  NOR2X0 U11080 ( .IN1(n11382), .IN2(n11396), .QN(n11395) );
  NAND2X0 U11081 ( .IN1(n11397), .IN2(n11398), .QN(n11396) );
  NAND2X0 U11082 ( .IN1(n11399), .IN2(n11387), .QN(n11398) );
  NAND2X0 U11083 ( .IN1(n11388), .IN2(DFF_1146_n1), .QN(n11397) );
  NAND2X0 U11084 ( .IN1(n11400), .IN2(n11401), .QN(n4245) );
  NAND2X0 U11085 ( .IN1(n11402), .IN2(n11373), .QN(n11401) );
  NOR2X0 U11086 ( .IN1(n11403), .IN2(n11404), .QN(n11402) );
  NOR2X0 U11087 ( .IN1(n11376), .IN2(n7967), .QN(n11404) );
  NOR2X0 U11088 ( .IN1(n11377), .IN2(n11405), .QN(n11403) );
  NAND2X0 U11089 ( .IN1(n11406), .IN2(n11407), .QN(n4244) );
  NAND2X0 U11090 ( .IN1(n2289), .IN2(n11408), .QN(n11407) );
  NAND2X0 U11091 ( .IN1(n11409), .IN2(n11373), .QN(n11406) );
  NOR2X0 U11092 ( .IN1(n11410), .IN2(n11411), .QN(n11409) );
  NOR2X0 U11093 ( .IN1(n11376), .IN2(g1916), .QN(n11411) );
  NOR2X0 U11094 ( .IN1(n11377), .IN2(n11412), .QN(n11410) );
  NAND2X0 U11095 ( .IN1(n11400), .IN2(n11413), .QN(n4243) );
  NAND2X0 U11096 ( .IN1(n11414), .IN2(n11373), .QN(n11413) );
  NOR2X0 U11097 ( .IN1(n11415), .IN2(n11416), .QN(n11414) );
  NOR2X0 U11098 ( .IN1(n11376), .IN2(n7964), .QN(n11416) );
  NOR2X0 U11099 ( .IN1(n11377), .IN2(n11417), .QN(n11415) );
  NOR2X0 U11100 ( .IN1(n11381), .IN2(n11418), .QN(n11400) );
  INVX0 U11101 ( .INP(n11419), .ZN(n11418) );
  NAND2X0 U11102 ( .IN1(n2289), .IN2(n2302), .QN(n11419) );
  INVX0 U11103 ( .INP(n2275), .ZN(n11381) );
  NAND2X0 U11104 ( .IN1(n2275), .IN2(n11420), .QN(n4242) );
  NAND2X0 U11105 ( .IN1(n11421), .IN2(n11373), .QN(n11420) );
  NOR2X0 U11106 ( .IN1(n11422), .IN2(n11423), .QN(n11421) );
  NOR2X0 U11107 ( .IN1(n11376), .IN2(n7963), .QN(n11423) );
  INVX0 U11108 ( .INP(n11388), .ZN(n11376) );
  NOR2X0 U11109 ( .IN1(n11377), .IN2(n11424), .QN(n11422) );
  INVX0 U11110 ( .INP(n11387), .ZN(n11377) );
  NAND2X0 U11111 ( .IN1(n11425), .IN2(n11426), .QN(n4241) );
  NAND2X0 U11112 ( .IN1(n11427), .IN2(g1937), .QN(n11426) );
  NAND2X0 U11113 ( .IN1(n11428), .IN2(n11429), .QN(n11427) );
  NAND2X0 U11114 ( .IN1(n11430), .IN2(n11408), .QN(n11429) );
  INVX0 U11115 ( .INP(n11371), .ZN(n11430) );
  NAND2X0 U11116 ( .IN1(n11431), .IN2(n11371), .QN(n11428) );
  NAND2X0 U11117 ( .IN1(n11432), .IN2(n11433), .QN(n11371) );
  NOR2X0 U11118 ( .IN1(n11434), .IN2(n11435), .QN(n11432) );
  NOR2X0 U11119 ( .IN1(n11436), .IN2(n11437), .QN(n11435) );
  NOR2X0 U11120 ( .IN1(n11438), .IN2(n11439), .QN(n11434) );
  INVX0 U11121 ( .INP(n11408), .ZN(n11431) );
  NAND2X0 U11122 ( .IN1(n11440), .IN2(n11441), .QN(n11408) );
  NOR2X0 U11123 ( .IN1(n11442), .IN2(n11443), .QN(n11440) );
  NOR2X0 U11124 ( .IN1(n11444), .IN2(n11445), .QN(n11443) );
  NOR2X0 U11125 ( .IN1(n11446), .IN2(n11447), .QN(n11442) );
  NOR2X0 U11126 ( .IN1(n11448), .IN2(n11449), .QN(n11425) );
  NOR2X0 U11127 ( .IN1(n4297), .IN2(n11450), .QN(n11449) );
  NAND2X0 U11128 ( .IN1(n11451), .IN2(n11452), .QN(n11450) );
  INVX0 U11129 ( .INP(n11453), .ZN(n11452) );
  NOR2X0 U11130 ( .IN1(n11454), .IN2(n11455), .QN(n11453) );
  NAND2X0 U11131 ( .IN1(n11455), .IN2(n11454), .QN(n11451) );
  NOR2X0 U11132 ( .IN1(n11456), .IN2(n11457), .QN(n11454) );
  INVX0 U11133 ( .INP(n11458), .ZN(n11457) );
  NAND2X0 U11134 ( .IN1(n11459), .IN2(n11386), .QN(n11458) );
  NOR2X0 U11135 ( .IN1(n11459), .IN2(n11386), .QN(n11456) );
  INVX0 U11136 ( .INP(n11460), .ZN(n11386) );
  NAND2X0 U11137 ( .IN1(n11461), .IN2(n11462), .QN(n11460) );
  NOR2X0 U11138 ( .IN1(n11463), .IN2(n11464), .QN(n11461) );
  NOR2X0 U11139 ( .IN1(n11465), .IN2(n11437), .QN(n11464) );
  NOR2X0 U11140 ( .IN1(n11438), .IN2(n11466), .QN(n11463) );
  NOR2X0 U11141 ( .IN1(n11467), .IN2(n11468), .QN(n11459) );
  NOR2X0 U11142 ( .IN1(n11469), .IN2(n11399), .QN(n11468) );
  INVX0 U11143 ( .INP(n11470), .ZN(n11467) );
  NAND2X0 U11144 ( .IN1(n11399), .IN2(n11469), .QN(n11470) );
  NAND2X0 U11145 ( .IN1(n11471), .IN2(n11472), .QN(n11469) );
  NAND2X0 U11146 ( .IN1(n11473), .IN2(n11474), .QN(n11472) );
  NAND2X0 U11147 ( .IN1(n11475), .IN2(n11476), .QN(n11474) );
  NAND2X0 U11148 ( .IN1(n11477), .IN2(n11424), .QN(n11476) );
  NAND2X0 U11149 ( .IN1(n11478), .IN2(n11405), .QN(n11475) );
  NOR2X0 U11150 ( .IN1(n11479), .IN2(n11480), .QN(n11473) );
  NOR2X0 U11151 ( .IN1(n11481), .IN2(n11412), .QN(n11480) );
  NOR2X0 U11152 ( .IN1(n11482), .IN2(n11378), .QN(n11479) );
  NAND2X0 U11153 ( .IN1(n11483), .IN2(n11484), .QN(n11471) );
  NAND2X0 U11154 ( .IN1(n11485), .IN2(n11486), .QN(n11484) );
  NAND2X0 U11155 ( .IN1(n11481), .IN2(n11412), .QN(n11486) );
  INVX0 U11156 ( .INP(n11378), .ZN(n11481) );
  NAND2X0 U11157 ( .IN1(n11482), .IN2(n11378), .QN(n11485) );
  NAND2X0 U11158 ( .IN1(n11487), .IN2(n11462), .QN(n11378) );
  NOR2X0 U11159 ( .IN1(n11488), .IN2(n11489), .QN(n11487) );
  NOR2X0 U11160 ( .IN1(n11490), .IN2(n11437), .QN(n11489) );
  NOR2X0 U11161 ( .IN1(n11438), .IN2(n11491), .QN(n11488) );
  INVX0 U11162 ( .INP(n11412), .ZN(n11482) );
  NAND2X0 U11163 ( .IN1(n11492), .IN2(n11441), .QN(n11412) );
  NOR2X0 U11164 ( .IN1(n11493), .IN2(n11494), .QN(n11492) );
  NOR2X0 U11165 ( .IN1(n11495), .IN2(n11445), .QN(n11494) );
  NOR2X0 U11166 ( .IN1(n11446), .IN2(n11496), .QN(n11493) );
  NOR2X0 U11167 ( .IN1(n11497), .IN2(n11498), .QN(n11483) );
  NOR2X0 U11168 ( .IN1(n11477), .IN2(n11424), .QN(n11498) );
  INVX0 U11169 ( .INP(n11405), .ZN(n11477) );
  NOR2X0 U11170 ( .IN1(n11478), .IN2(n11405), .QN(n11497) );
  NAND2X0 U11171 ( .IN1(n11499), .IN2(n11462), .QN(n11405) );
  NOR2X0 U11172 ( .IN1(n11500), .IN2(n11501), .QN(n11499) );
  NOR2X0 U11173 ( .IN1(n11502), .IN2(n11445), .QN(n11501) );
  NOR2X0 U11174 ( .IN1(n11446), .IN2(n11503), .QN(n11500) );
  INVX0 U11175 ( .INP(n11424), .ZN(n11478) );
  NAND2X0 U11176 ( .IN1(n11504), .IN2(n11441), .QN(n11424) );
  INVX0 U11177 ( .INP(n11505), .ZN(n11441) );
  NAND2X0 U11178 ( .IN1(n11462), .IN2(n11506), .QN(n11505) );
  NAND2X0 U11179 ( .IN1(n11507), .IN2(n11508), .QN(n11506) );
  NOR2X0 U11180 ( .IN1(n11509), .IN2(n11510), .QN(n11504) );
  NOR2X0 U11181 ( .IN1(n11511), .IN2(n11445), .QN(n11510) );
  NOR2X0 U11182 ( .IN1(n11446), .IN2(n11512), .QN(n11509) );
  INVX0 U11183 ( .INP(n11513), .ZN(n11399) );
  NAND2X0 U11184 ( .IN1(n11514), .IN2(n11462), .QN(n11513) );
  NOR2X0 U11185 ( .IN1(n11515), .IN2(n11516), .QN(n11514) );
  NOR2X0 U11186 ( .IN1(n11517), .IN2(n11445), .QN(n11516) );
  NAND2X0 U11187 ( .IN1(n11446), .IN2(n11518), .QN(n11445) );
  NOR2X0 U11188 ( .IN1(n11446), .IN2(n11519), .QN(n11515) );
  NAND2X0 U11189 ( .IN1(n11520), .IN2(n11521), .QN(n11455) );
  INVX0 U11190 ( .INP(n11522), .ZN(n11521) );
  NOR2X0 U11191 ( .IN1(n11393), .IN2(n11523), .QN(n11522) );
  NAND2X0 U11192 ( .IN1(n11523), .IN2(n11393), .QN(n11520) );
  NAND2X0 U11193 ( .IN1(n11524), .IN2(n11433), .QN(n11393) );
  INVX0 U11194 ( .INP(n11525), .ZN(n11433) );
  NAND2X0 U11195 ( .IN1(n11462), .IN2(n11526), .QN(n11525) );
  NAND2X0 U11196 ( .IN1(n11507), .IN2(n11527), .QN(n11526) );
  NOR2X0 U11197 ( .IN1(n11528), .IN2(n11529), .QN(n11524) );
  NOR2X0 U11198 ( .IN1(n11530), .IN2(n11437), .QN(n11529) );
  NOR2X0 U11199 ( .IN1(n11438), .IN2(n11531), .QN(n11528) );
  INVX0 U11200 ( .INP(n11417), .ZN(n11523) );
  NAND2X0 U11201 ( .IN1(n11532), .IN2(n11462), .QN(n11417) );
  NOR2X0 U11202 ( .IN1(n10724), .IN2(n4545), .QN(n11462) );
  NOR2X0 U11203 ( .IN1(n11533), .IN2(n11534), .QN(n11532) );
  NOR2X0 U11204 ( .IN1(n11535), .IN2(n11437), .QN(n11534) );
  NAND2X0 U11205 ( .IN1(n11438), .IN2(n11518), .QN(n11437) );
  NOR2X0 U11206 ( .IN1(n11438), .IN2(n11536), .QN(n11533) );
  NOR2X0 U11207 ( .IN1(n11537), .IN2(n11538), .QN(n11448) );
  NAND2X0 U11208 ( .IN1(n11373), .IN2(n11388), .QN(n11538) );
  NOR2X0 U11209 ( .IN1(n10724), .IN2(n11387), .QN(n11388) );
  NAND2X0 U11210 ( .IN1(n11539), .IN2(n10077), .QN(n10724) );
  NOR2X0 U11211 ( .IN1(g1943), .IN2(n618), .QN(n11539) );
  NAND2X0 U11212 ( .IN1(n11540), .IN2(n11541), .QN(n11537) );
  INVX0 U11213 ( .INP(n11542), .ZN(n11541) );
  NOR2X0 U11214 ( .IN1(n11195), .IN2(test_so69), .QN(n11542) );
  NAND2X0 U11215 ( .IN1(n18857), .IN2(n11195), .QN(n11540) );
  NAND2X0 U11216 ( .IN1(n11543), .IN2(n11544), .QN(n4240) );
  NAND2X0 U11217 ( .IN1(n2217), .IN2(n11545), .QN(n11544) );
  NAND2X0 U11218 ( .IN1(n11546), .IN2(n11547), .QN(n11543) );
  NOR2X0 U11219 ( .IN1(n11548), .IN2(n11549), .QN(n11546) );
  NOR2X0 U11220 ( .IN1(n11550), .IN2(g1223), .QN(n11549) );
  NOR2X0 U11221 ( .IN1(n11551), .IN2(n11552), .QN(n11548) );
  NAND2X0 U11222 ( .IN1(n11553), .IN2(n2231), .QN(n4239) );
  NOR2X0 U11223 ( .IN1(n11554), .IN2(n11555), .QN(n11553) );
  NOR2X0 U11224 ( .IN1(n11556), .IN2(n11557), .QN(n11555) );
  NAND2X0 U11225 ( .IN1(n11558), .IN2(n11559), .QN(n11557) );
  NAND2X0 U11226 ( .IN1(n11560), .IN2(n11561), .QN(n11559) );
  NAND2X0 U11227 ( .IN1(n11562), .IN2(DFF_795_n1), .QN(n11558) );
  NAND2X0 U11228 ( .IN1(n11563), .IN2(n11564), .QN(n4238) );
  NAND2X0 U11229 ( .IN1(n11565), .IN2(n11547), .QN(n11564) );
  NOR2X0 U11230 ( .IN1(n11566), .IN2(n11567), .QN(n11565) );
  NOR2X0 U11231 ( .IN1(n11550), .IN2(n8003), .QN(n11567) );
  NOR2X0 U11232 ( .IN1(n11551), .IN2(n11568), .QN(n11566) );
  NAND2X0 U11233 ( .IN1(n11569), .IN2(n2231), .QN(n4237) );
  NOR2X0 U11234 ( .IN1(n11554), .IN2(n11570), .QN(n11569) );
  NOR2X0 U11235 ( .IN1(n11556), .IN2(n11571), .QN(n11570) );
  NAND2X0 U11236 ( .IN1(n11572), .IN2(n11573), .QN(n11571) );
  NAND2X0 U11237 ( .IN1(n11574), .IN2(n11561), .QN(n11573) );
  NAND2X0 U11238 ( .IN1(n11562), .IN2(DFF_796_n1), .QN(n11572) );
  NAND2X0 U11239 ( .IN1(n11575), .IN2(n11576), .QN(n4236) );
  NAND2X0 U11240 ( .IN1(n11577), .IN2(n11547), .QN(n11576) );
  NOR2X0 U11241 ( .IN1(n11578), .IN2(n11579), .QN(n11577) );
  NOR2X0 U11242 ( .IN1(n11550), .IN2(n8008), .QN(n11579) );
  NOR2X0 U11243 ( .IN1(n11551), .IN2(n11580), .QN(n11578) );
  NAND2X0 U11244 ( .IN1(n11581), .IN2(n11582), .QN(n4235) );
  NAND2X0 U11245 ( .IN1(n2217), .IN2(n11583), .QN(n11582) );
  NAND2X0 U11246 ( .IN1(n11584), .IN2(n11547), .QN(n11581) );
  NOR2X0 U11247 ( .IN1(n11585), .IN2(n11586), .QN(n11584) );
  NOR2X0 U11248 ( .IN1(n11550), .IN2(g1222), .QN(n11586) );
  NOR2X0 U11249 ( .IN1(n11551), .IN2(n11587), .QN(n11585) );
  NAND2X0 U11250 ( .IN1(n11575), .IN2(n11588), .QN(n4234) );
  NAND2X0 U11251 ( .IN1(n11589), .IN2(n11547), .QN(n11588) );
  NOR2X0 U11252 ( .IN1(n11590), .IN2(n11591), .QN(n11589) );
  NOR2X0 U11253 ( .IN1(n11550), .IN2(n8005), .QN(n11591) );
  NOR2X0 U11254 ( .IN1(n11551), .IN2(n11592), .QN(n11590) );
  NOR2X0 U11255 ( .IN1(n11554), .IN2(n11593), .QN(n11575) );
  INVX0 U11256 ( .INP(n11594), .ZN(n11593) );
  NAND2X0 U11257 ( .IN1(n2217), .IN2(n2230), .QN(n11594) );
  INVX0 U11258 ( .INP(n11563), .ZN(n11554) );
  NAND2X0 U11259 ( .IN1(n11563), .IN2(n11595), .QN(n4233) );
  NAND2X0 U11260 ( .IN1(n11596), .IN2(n11547), .QN(n11595) );
  NOR2X0 U11261 ( .IN1(n11597), .IN2(n11598), .QN(n11596) );
  NOR2X0 U11262 ( .IN1(n11550), .IN2(n8004), .QN(n11598) );
  INVX0 U11263 ( .INP(n11562), .ZN(n11550) );
  NOR2X0 U11264 ( .IN1(n11551), .IN2(n11599), .QN(n11597) );
  INVX0 U11265 ( .INP(n11561), .ZN(n11551) );
  NAND2X0 U11266 ( .IN1(n2217), .IN2(n11600), .QN(n11563) );
  NAND2X0 U11267 ( .IN1(n11601), .IN2(n11602), .QN(n4232) );
  NAND2X0 U11268 ( .IN1(n11603), .IN2(g1243), .QN(n11602) );
  NAND2X0 U11269 ( .IN1(n11604), .IN2(n11605), .QN(n11603) );
  NAND2X0 U11270 ( .IN1(n11606), .IN2(n11583), .QN(n11605) );
  INVX0 U11271 ( .INP(n11545), .ZN(n11606) );
  NAND2X0 U11272 ( .IN1(n11607), .IN2(n11545), .QN(n11604) );
  NAND2X0 U11273 ( .IN1(n11608), .IN2(n11609), .QN(n11545) );
  NOR2X0 U11274 ( .IN1(n11610), .IN2(n11611), .QN(n11608) );
  NOR2X0 U11275 ( .IN1(n11612), .IN2(n11613), .QN(n11611) );
  NOR2X0 U11276 ( .IN1(n11614), .IN2(n11615), .QN(n11610) );
  INVX0 U11277 ( .INP(n11583), .ZN(n11607) );
  NAND2X0 U11278 ( .IN1(n11616), .IN2(n11617), .QN(n11583) );
  NOR2X0 U11279 ( .IN1(n11618), .IN2(n11619), .QN(n11616) );
  NOR2X0 U11280 ( .IN1(n11620), .IN2(n11621), .QN(n11619) );
  NOR2X0 U11281 ( .IN1(n11622), .IN2(n11623), .QN(n11618) );
  NOR2X0 U11282 ( .IN1(n11624), .IN2(n11625), .QN(n11601) );
  NOR2X0 U11283 ( .IN1(n4304), .IN2(n11626), .QN(n11625) );
  NAND2X0 U11284 ( .IN1(n11627), .IN2(n11628), .QN(n11626) );
  INVX0 U11285 ( .INP(n11629), .ZN(n11628) );
  NOR2X0 U11286 ( .IN1(n11630), .IN2(n11631), .QN(n11629) );
  NAND2X0 U11287 ( .IN1(n11631), .IN2(n11630), .QN(n11627) );
  NOR2X0 U11288 ( .IN1(n11632), .IN2(n11633), .QN(n11630) );
  INVX0 U11289 ( .INP(n11634), .ZN(n11633) );
  NAND2X0 U11290 ( .IN1(n11635), .IN2(n11560), .QN(n11634) );
  NOR2X0 U11291 ( .IN1(n11635), .IN2(n11560), .QN(n11632) );
  INVX0 U11292 ( .INP(n11636), .ZN(n11560) );
  NAND2X0 U11293 ( .IN1(n11637), .IN2(n11638), .QN(n11636) );
  NOR2X0 U11294 ( .IN1(n11639), .IN2(n11640), .QN(n11637) );
  NOR2X0 U11295 ( .IN1(n11641), .IN2(n11613), .QN(n11640) );
  NOR2X0 U11296 ( .IN1(n11614), .IN2(n11642), .QN(n11639) );
  NOR2X0 U11297 ( .IN1(n11643), .IN2(n11644), .QN(n11635) );
  NOR2X0 U11298 ( .IN1(n11645), .IN2(n11574), .QN(n11644) );
  INVX0 U11299 ( .INP(n11646), .ZN(n11643) );
  NAND2X0 U11300 ( .IN1(n11574), .IN2(n11645), .QN(n11646) );
  NAND2X0 U11301 ( .IN1(n11647), .IN2(n11648), .QN(n11645) );
  NAND2X0 U11302 ( .IN1(n11649), .IN2(n11650), .QN(n11648) );
  NAND2X0 U11303 ( .IN1(n11651), .IN2(n11652), .QN(n11650) );
  NAND2X0 U11304 ( .IN1(n11653), .IN2(n11599), .QN(n11652) );
  NAND2X0 U11305 ( .IN1(n11654), .IN2(n11580), .QN(n11651) );
  NOR2X0 U11306 ( .IN1(n11655), .IN2(n11656), .QN(n11649) );
  NOR2X0 U11307 ( .IN1(n11657), .IN2(n11587), .QN(n11656) );
  NOR2X0 U11308 ( .IN1(n11658), .IN2(n11552), .QN(n11655) );
  NAND2X0 U11309 ( .IN1(n11659), .IN2(n11660), .QN(n11647) );
  NAND2X0 U11310 ( .IN1(n11661), .IN2(n11662), .QN(n11660) );
  NAND2X0 U11311 ( .IN1(n11657), .IN2(n11587), .QN(n11662) );
  INVX0 U11312 ( .INP(n11552), .ZN(n11657) );
  NAND2X0 U11313 ( .IN1(n11658), .IN2(n11552), .QN(n11661) );
  NAND2X0 U11314 ( .IN1(n11663), .IN2(n11638), .QN(n11552) );
  NOR2X0 U11315 ( .IN1(n11664), .IN2(n11665), .QN(n11663) );
  NOR2X0 U11316 ( .IN1(n11666), .IN2(n11613), .QN(n11665) );
  NOR2X0 U11317 ( .IN1(n11614), .IN2(n11667), .QN(n11664) );
  INVX0 U11318 ( .INP(n11587), .ZN(n11658) );
  NAND2X0 U11319 ( .IN1(n11668), .IN2(n11617), .QN(n11587) );
  NOR2X0 U11320 ( .IN1(n11669), .IN2(n11670), .QN(n11668) );
  NOR2X0 U11321 ( .IN1(n11671), .IN2(n11621), .QN(n11670) );
  NOR2X0 U11322 ( .IN1(n11622), .IN2(n11672), .QN(n11669) );
  NOR2X0 U11323 ( .IN1(n11673), .IN2(n11674), .QN(n11659) );
  NOR2X0 U11324 ( .IN1(n11653), .IN2(n11599), .QN(n11674) );
  INVX0 U11325 ( .INP(n11580), .ZN(n11653) );
  NOR2X0 U11326 ( .IN1(n11654), .IN2(n11580), .QN(n11673) );
  NAND2X0 U11327 ( .IN1(n11675), .IN2(n11638), .QN(n11580) );
  NOR2X0 U11328 ( .IN1(n11676), .IN2(n11677), .QN(n11675) );
  NOR2X0 U11329 ( .IN1(n11678), .IN2(n11621), .QN(n11677) );
  NOR2X0 U11330 ( .IN1(n11622), .IN2(n11679), .QN(n11676) );
  INVX0 U11331 ( .INP(n11599), .ZN(n11654) );
  NAND2X0 U11332 ( .IN1(n11680), .IN2(n11617), .QN(n11599) );
  INVX0 U11333 ( .INP(n11681), .ZN(n11617) );
  NAND2X0 U11334 ( .IN1(n11638), .IN2(n11682), .QN(n11681) );
  NAND2X0 U11335 ( .IN1(n11683), .IN2(n11684), .QN(n11682) );
  NOR2X0 U11336 ( .IN1(n11685), .IN2(n11686), .QN(n11680) );
  NOR2X0 U11337 ( .IN1(n11687), .IN2(n11621), .QN(n11686) );
  NOR2X0 U11338 ( .IN1(n11622), .IN2(n11688), .QN(n11685) );
  INVX0 U11339 ( .INP(n11689), .ZN(n11574) );
  NAND2X0 U11340 ( .IN1(n11690), .IN2(n11638), .QN(n11689) );
  NOR2X0 U11341 ( .IN1(n11691), .IN2(n11692), .QN(n11690) );
  NOR2X0 U11342 ( .IN1(n11693), .IN2(n11621), .QN(n11692) );
  NAND2X0 U11343 ( .IN1(n11622), .IN2(n11694), .QN(n11621) );
  NOR2X0 U11344 ( .IN1(n11622), .IN2(n11695), .QN(n11691) );
  NAND2X0 U11345 ( .IN1(n11696), .IN2(n11697), .QN(n11631) );
  INVX0 U11346 ( .INP(n11698), .ZN(n11697) );
  NOR2X0 U11347 ( .IN1(n11568), .IN2(n11699), .QN(n11698) );
  NAND2X0 U11348 ( .IN1(n11699), .IN2(n11568), .QN(n11696) );
  NAND2X0 U11349 ( .IN1(n11700), .IN2(n11609), .QN(n11568) );
  INVX0 U11350 ( .INP(n11701), .ZN(n11609) );
  NAND2X0 U11351 ( .IN1(n11638), .IN2(n11702), .QN(n11701) );
  NAND2X0 U11352 ( .IN1(n11683), .IN2(n11703), .QN(n11702) );
  NOR2X0 U11353 ( .IN1(n11704), .IN2(n11705), .QN(n11700) );
  NOR2X0 U11354 ( .IN1(n11706), .IN2(n11613), .QN(n11705) );
  NOR2X0 U11355 ( .IN1(n11614), .IN2(n11707), .QN(n11704) );
  INVX0 U11356 ( .INP(n11592), .ZN(n11699) );
  NAND2X0 U11357 ( .IN1(n11708), .IN2(n11638), .QN(n11592) );
  NOR2X0 U11358 ( .IN1(n11600), .IN2(n4548), .QN(n11638) );
  NOR2X0 U11359 ( .IN1(n11709), .IN2(n11710), .QN(n11708) );
  NOR2X0 U11360 ( .IN1(n11711), .IN2(n11613), .QN(n11710) );
  NAND2X0 U11361 ( .IN1(n11614), .IN2(n11694), .QN(n11613) );
  NOR2X0 U11362 ( .IN1(n11614), .IN2(n11712), .QN(n11709) );
  NOR2X0 U11363 ( .IN1(n11713), .IN2(n11714), .QN(n11624) );
  NAND2X0 U11364 ( .IN1(n11547), .IN2(n11562), .QN(n11714) );
  NOR2X0 U11365 ( .IN1(n11600), .IN2(n11561), .QN(n11562) );
  NAND2X0 U11366 ( .IN1(n11715), .IN2(n10078), .QN(n11600) );
  NOR2X0 U11367 ( .IN1(g1249), .IN2(n588), .QN(n11715) );
  NAND2X0 U11368 ( .IN1(n11716), .IN2(n11717), .QN(n11713) );
  NAND2X0 U11369 ( .IN1(n4489), .IN2(g3229), .QN(n11717) );
  NAND2X0 U11370 ( .IN1(n11195), .IN2(n18858), .QN(n11716) );
  INVX0 U11371 ( .INP(n11718), .ZN(n3788) );
  INVX0 U11372 ( .INP(n11719), .ZN(n3758) );
  INVX0 U11373 ( .INP(n11720), .ZN(n3751) );
  INVX0 U11374 ( .INP(n11721), .ZN(n372) );
  INVX0 U11375 ( .INP(n11722), .ZN(n37) );
  NAND2X0 U11376 ( .IN1(n3896), .IN2(g88), .QN(n4528) );
  NAND2X0 U11377 ( .IN1(n3890), .IN2(g1462), .QN(n4527) );
  NAND2X0 U11378 ( .IN1(n3887), .IN2(test_so78), .QN(n4526) );
  NAND2X0 U11379 ( .IN1(n3692), .IN2(test_so15), .QN(n4521) );
  NAND2X0 U11380 ( .IN1(n3686), .IN2(g1453), .QN(n4523) );
  NAND2X0 U11381 ( .IN1(n3683), .IN2(g2147), .QN(n4522) );
  NAND2X0 U11382 ( .IN1(n11723), .IN2(n11724), .QN(n3254) );
  INVX0 U11383 ( .INP(n11725), .ZN(n11723) );
  NOR2X0 U11384 ( .IN1(n11726), .IN2(n11727), .QN(n11725) );
  INVX0 U11385 ( .INP(g24734), .ZN(n318) );
  INVX0 U11386 ( .INP(g25435), .ZN(n310) );
  INVX0 U11387 ( .INP(n11728), .ZN(n306) );
  NAND2X0 U11388 ( .IN1(n11729), .IN2(n11730), .QN(n3023) );
  NOR2X0 U11389 ( .IN1(n4388), .IN2(n11731), .QN(n11730) );
  NOR2X0 U11390 ( .IN1(n11732), .IN2(n11733), .QN(n11729) );
  NAND2X0 U11391 ( .IN1(n11734), .IN2(n11735), .QN(n3016) );
  NOR2X0 U11392 ( .IN1(n4387), .IN2(n11736), .QN(n11735) );
  NOR2X0 U11393 ( .IN1(n11737), .IN2(n11738), .QN(n11734) );
  NAND2X0 U11394 ( .IN1(n11739), .IN2(n11740), .QN(n3008) );
  NOR2X0 U11395 ( .IN1(n4386), .IN2(n11741), .QN(n11740) );
  NOR2X0 U11396 ( .IN1(n11742), .IN2(n11743), .QN(n11739) );
  NAND2X0 U11397 ( .IN1(n11744), .IN2(n11745), .QN(n3000) );
  NOR2X0 U11398 ( .IN1(n10322), .IN2(n11746), .QN(n11745) );
  NOR2X0 U11399 ( .IN1(n11747), .IN2(n11748), .QN(n11744) );
  NAND2X0 U11400 ( .IN1(n11749), .IN2(n11750), .QN(n2800) );
  INVX0 U11401 ( .INP(n11751), .ZN(n11750) );
  NOR2X0 U11402 ( .IN1(n11752), .IN2(n11753), .QN(n11751) );
  NAND2X0 U11403 ( .IN1(n11752), .IN2(n11753), .QN(n11749) );
  NAND2X0 U11404 ( .IN1(n11754), .IN2(n11755), .QN(n11752) );
  NAND2X0 U11405 ( .IN1(n11756), .IN2(n11757), .QN(n11755) );
  NAND2X0 U11406 ( .IN1(n11758), .IN2(n11759), .QN(n11757) );
  NOR2X0 U11407 ( .IN1(n11760), .IN2(n11761), .QN(n11758) );
  NOR2X0 U11408 ( .IN1(n11762), .IN2(n11763), .QN(n11761) );
  INVX0 U11409 ( .INP(n11764), .ZN(n11763) );
  NOR2X0 U11410 ( .IN1(n11765), .IN2(n4387), .QN(n11764) );
  NOR2X0 U11411 ( .IN1(n11766), .IN2(n11767), .QN(n11760) );
  NAND2X0 U11412 ( .IN1(n11768), .IN2(n11753), .QN(n11754) );
  NOR2X0 U11413 ( .IN1(n11769), .IN2(n11770), .QN(n11768) );
  NAND2X0 U11414 ( .IN1(n11759), .IN2(n11762), .QN(n11769) );
  INVX0 U11415 ( .INP(g26135), .ZN(n278) );
  NAND2X0 U11416 ( .IN1(n11771), .IN2(n11772), .QN(n2719) );
  NAND2X0 U11417 ( .IN1(n10771), .IN2(n11773), .QN(n11772) );
  NAND2X0 U11418 ( .IN1(n11774), .IN2(n10770), .QN(n11771) );
  NAND2X0 U11419 ( .IN1(n11775), .IN2(n11776), .QN(n2686) );
  NAND2X0 U11420 ( .IN1(n10901), .IN2(n11777), .QN(n11776) );
  NAND2X0 U11421 ( .IN1(n4530), .IN2(n10900), .QN(n11775) );
  NAND2X0 U11422 ( .IN1(n11778), .IN2(n11779), .QN(n2671) );
  NAND2X0 U11423 ( .IN1(n10966), .IN2(n11780), .QN(n11779) );
  NAND2X0 U11424 ( .IN1(n4529), .IN2(n10965), .QN(n11778) );
  NAND2X0 U11425 ( .IN1(n11781), .IN2(n11782), .QN(n2616) );
  NAND2X0 U11426 ( .IN1(n11766), .IN2(n11783), .QN(n11782) );
  INVX0 U11427 ( .INP(n11784), .ZN(n11781) );
  NOR2X0 U11428 ( .IN1(n11783), .IN2(n11766), .QN(n11784) );
  NAND2X0 U11429 ( .IN1(n11785), .IN2(n11786), .QN(n11783) );
  NAND2X0 U11430 ( .IN1(n11787), .IN2(n11753), .QN(n11786) );
  NOR2X0 U11431 ( .IN1(n11788), .IN2(n11789), .QN(n11785) );
  NOR2X0 U11432 ( .IN1(n11790), .IN2(n11762), .QN(n11789) );
  NOR2X0 U11433 ( .IN1(n11791), .IN2(n11792), .QN(n11790) );
  NOR2X0 U11434 ( .IN1(n11793), .IN2(n11794), .QN(n11792) );
  NAND2X0 U11435 ( .IN1(n11767), .IN2(n11795), .QN(n11794) );
  NOR2X0 U11436 ( .IN1(n11796), .IN2(n11797), .QN(n11767) );
  NOR2X0 U11437 ( .IN1(n11798), .IN2(n11799), .QN(n11797) );
  NAND2X0 U11438 ( .IN1(n11800), .IN2(n11759), .QN(n11793) );
  NAND2X0 U11439 ( .IN1(n11801), .IN2(n11802), .QN(n11800) );
  INVX0 U11440 ( .INP(n2632), .ZN(n11802) );
  INVX0 U11441 ( .INP(n11803), .ZN(n11791) );
  NAND2X0 U11442 ( .IN1(n2632), .IN2(n11804), .QN(n11803) );
  NOR2X0 U11443 ( .IN1(n11756), .IN2(n11796), .QN(n11804) );
  NOR2X0 U11444 ( .IN1(n11766), .IN2(n11805), .QN(n11788) );
  NOR2X0 U11445 ( .IN1(n11799), .IN2(n11806), .QN(n11805) );
  NAND2X0 U11446 ( .IN1(n11807), .IN2(n11759), .QN(n11806) );
  NAND2X0 U11447 ( .IN1(n11808), .IN2(n11809), .QN(n11807) );
  NAND2X0 U11448 ( .IN1(n11795), .IN2(n11798), .QN(n11809) );
  NOR2X0 U11449 ( .IN1(n11753), .IN2(n11810), .QN(n11795) );
  INVX0 U11450 ( .INP(n11811), .ZN(n11810) );
  INVX0 U11451 ( .INP(n11812), .ZN(n11808) );
  NOR2X0 U11452 ( .IN1(n11042), .IN2(n11008), .QN(n2446) );
  INVX0 U11453 ( .INP(n11037), .ZN(n11008) );
  NAND2X0 U11454 ( .IN1(n4360), .IN2(n11813), .QN(n11037) );
  NAND2X0 U11455 ( .IN1(n10036), .IN2(n10326), .QN(n11813) );
  NAND2X0 U11456 ( .IN1(n10326), .IN2(n11814), .QN(n11042) );
  NAND2X0 U11457 ( .IN1(n4360), .IN2(n10036), .QN(n11814) );
  NAND2X0 U11458 ( .IN1(g499), .IN2(n11815), .QN(n2445) );
  NAND2X0 U11459 ( .IN1(n11816), .IN2(n11817), .QN(n11815) );
  NOR2X0 U11460 ( .IN1(n11173), .IN2(n11818), .QN(n11817) );
  NOR2X0 U11461 ( .IN1(n4295), .IN2(g734), .QN(n11818) );
  INVX0 U11462 ( .INP(n11178), .ZN(n11173) );
  NAND2X0 U11463 ( .IN1(n11819), .IN2(n11820), .QN(n11178) );
  NOR2X0 U11464 ( .IN1(n11821), .IN2(n11822), .QN(n11820) );
  NAND2X0 U11465 ( .IN1(n11823), .IN2(n11144), .QN(n11822) );
  NOR2X0 U11466 ( .IN1(n11177), .IN2(n11094), .QN(n11823) );
  NAND2X0 U11467 ( .IN1(n11824), .IN2(n11187), .QN(n11821) );
  NOR2X0 U11468 ( .IN1(n11825), .IN2(n11162), .QN(n11824) );
  INVX0 U11469 ( .INP(n11826), .ZN(n11825) );
  NOR2X0 U11470 ( .IN1(n11827), .IN2(n11828), .QN(n11819) );
  NAND2X0 U11471 ( .IN1(n11829), .IN2(n11107), .QN(n11828) );
  NOR2X0 U11472 ( .IN1(n11136), .IN2(n11131), .QN(n11829) );
  NAND2X0 U11473 ( .IN1(n11830), .IN2(n11148), .QN(n11827) );
  NOR2X0 U11474 ( .IN1(n11831), .IN2(n11158), .QN(n11830) );
  NOR2X0 U11475 ( .IN1(n11832), .IN2(n11833), .QN(n11831) );
  NAND2X0 U11476 ( .IN1(n11834), .IN2(n11835), .QN(n11833) );
  NAND2X0 U11477 ( .IN1(n10196), .IN2(g6677), .QN(n11835) );
  NAND2X0 U11478 ( .IN1(n10263), .IN2(g629), .QN(n11834) );
  NOR2X0 U11479 ( .IN1(n4359), .IN2(g739), .QN(n11832) );
  NOR2X0 U11480 ( .IN1(n11836), .IN2(n11837), .QN(n11816) );
  NOR2X0 U11481 ( .IN1(n4359), .IN2(g736), .QN(n11837) );
  NOR2X0 U11482 ( .IN1(n4309), .IN2(g735), .QN(n11836) );
  NAND2X0 U11483 ( .IN1(g2574), .IN2(n11838), .QN(n2374) );
  NAND2X0 U11484 ( .IN1(n11839), .IN2(n11840), .QN(n11838) );
  NOR2X0 U11485 ( .IN1(n11353), .IN2(n11841), .QN(n11840) );
  NOR2X0 U11486 ( .IN1(n4292), .IN2(g2808), .QN(n11841) );
  NOR2X0 U11487 ( .IN1(n11842), .IN2(n11843), .QN(n11839) );
  NOR2X0 U11488 ( .IN1(n4356), .IN2(g2810), .QN(n11843) );
  NOR2X0 U11489 ( .IN1(n4306), .IN2(g2809), .QN(n11842) );
  NOR2X0 U11490 ( .IN1(n11214), .IN2(n11200), .QN(n2361) );
  INVX0 U11491 ( .INP(n11209), .ZN(n11200) );
  NAND2X0 U11492 ( .IN1(n4352), .IN2(n11844), .QN(n11209) );
  NAND2X0 U11493 ( .IN1(n4303), .IN2(n10033), .QN(n11844) );
  NAND2X0 U11494 ( .IN1(n4303), .IN2(n11845), .QN(n11214) );
  NAND2X0 U11495 ( .IN1(n4352), .IN2(n10033), .QN(n11845) );
  NAND2X0 U11496 ( .IN1(n11353), .IN2(n11846), .QN(n2351) );
  INVX0 U11497 ( .INP(n11344), .ZN(n11353) );
  NAND2X0 U11498 ( .IN1(n11847), .IN2(n11848), .QN(n11344) );
  NOR2X0 U11499 ( .IN1(n11849), .IN2(n11850), .QN(n11848) );
  NAND2X0 U11500 ( .IN1(n11851), .IN2(n11358), .QN(n11850) );
  NOR2X0 U11501 ( .IN1(n11273), .IN2(n11324), .QN(n11851) );
  NAND2X0 U11502 ( .IN1(n11852), .IN2(n11338), .QN(n11849) );
  NOR2X0 U11503 ( .IN1(n11265), .IN2(n11853), .QN(n11852) );
  INVX0 U11504 ( .INP(n11854), .ZN(n11853) );
  NOR2X0 U11505 ( .IN1(n11855), .IN2(n11856), .QN(n11847) );
  NAND2X0 U11506 ( .IN1(n11857), .IN2(n11343), .QN(n11856) );
  NOR2X0 U11507 ( .IN1(n11363), .IN2(n11295), .QN(n11857) );
  NAND2X0 U11508 ( .IN1(n11858), .IN2(n11331), .QN(n11855) );
  NOR2X0 U11509 ( .IN1(n11859), .IN2(n11320), .QN(n11858) );
  NOR2X0 U11510 ( .IN1(n11860), .IN2(n11861), .QN(n11859) );
  NAND2X0 U11511 ( .IN1(n11862), .IN2(n11863), .QN(n11861) );
  NAND2X0 U11512 ( .IN1(n10193), .IN2(g7425), .QN(n11863) );
  INVX0 U11513 ( .INP(n11864), .ZN(n11862) );
  NOR2X0 U11514 ( .IN1(n4292), .IN2(test_so95), .QN(n11864) );
  NOR2X0 U11515 ( .IN1(n4356), .IN2(g2813), .QN(n11860) );
  NAND2X0 U11516 ( .IN1(g1880), .IN2(n11865), .QN(n2302) );
  NAND2X0 U11517 ( .IN1(n11866), .IN2(n11867), .QN(n11865) );
  NOR2X0 U11518 ( .IN1(n11507), .IN2(n11868), .QN(n11867) );
  NOR2X0 U11519 ( .IN1(n4293), .IN2(g2114), .QN(n11868) );
  INVX0 U11520 ( .INP(n11518), .ZN(n11507) );
  NAND2X0 U11521 ( .IN1(n11869), .IN2(n11870), .QN(n11518) );
  NOR2X0 U11522 ( .IN1(n11871), .IN2(n11872), .QN(n11870) );
  NAND2X0 U11523 ( .IN1(n11873), .IN2(n11531), .QN(n11872) );
  NOR2X0 U11524 ( .IN1(n11444), .IN2(n11495), .QN(n11873) );
  NAND2X0 U11525 ( .IN1(n11874), .IN2(n11512), .QN(n11871) );
  NOR2X0 U11526 ( .IN1(n11436), .IN2(n11875), .QN(n11874) );
  INVX0 U11527 ( .INP(n11876), .ZN(n11875) );
  NOR2X0 U11528 ( .IN1(n11877), .IN2(n11878), .QN(n11869) );
  NAND2X0 U11529 ( .IN1(n11879), .IN2(n11490), .QN(n11878) );
  NOR2X0 U11530 ( .IN1(n11466), .IN2(n11519), .QN(n11879) );
  NAND2X0 U11531 ( .IN1(n11880), .IN2(n11535), .QN(n11877) );
  NOR2X0 U11532 ( .IN1(n11881), .IN2(n11503), .QN(n11880) );
  NOR2X0 U11533 ( .IN1(n11882), .IN2(n11883), .QN(n11881) );
  NAND2X0 U11534 ( .IN1(n11884), .IN2(n11885), .QN(n11883) );
  NAND2X0 U11535 ( .IN1(n10194), .IN2(g7229), .QN(n11885) );
  NAND2X0 U11536 ( .IN1(n10261), .IN2(g2009), .QN(n11884) );
  NOR2X0 U11537 ( .IN1(n4357), .IN2(g2119), .QN(n11882) );
  NOR2X0 U11538 ( .IN1(n11886), .IN2(n11887), .QN(n11866) );
  NOR2X0 U11539 ( .IN1(n4357), .IN2(g2116), .QN(n11887) );
  NOR2X0 U11540 ( .IN1(n4307), .IN2(g2115), .QN(n11886) );
  NOR2X0 U11541 ( .IN1(n11387), .IN2(n11373), .QN(n2289) );
  INVX0 U11542 ( .INP(n11382), .ZN(n11373) );
  NAND2X0 U11543 ( .IN1(n4311), .IN2(n11888), .QN(n11382) );
  NAND2X0 U11544 ( .IN1(n4297), .IN2(n10034), .QN(n11888) );
  NAND2X0 U11545 ( .IN1(n4297), .IN2(n11889), .QN(n11387) );
  NAND2X0 U11546 ( .IN1(n4311), .IN2(n10034), .QN(n11889) );
  NAND2X0 U11547 ( .IN1(g1186), .IN2(n11890), .QN(n2230) );
  NAND2X0 U11548 ( .IN1(n11891), .IN2(n11892), .QN(n11890) );
  NOR2X0 U11549 ( .IN1(n11683), .IN2(n11893), .QN(n11892) );
  NOR2X0 U11550 ( .IN1(n4294), .IN2(g1420), .QN(n11893) );
  INVX0 U11551 ( .INP(n11694), .ZN(n11683) );
  NAND2X0 U11552 ( .IN1(n11894), .IN2(n11895), .QN(n11694) );
  NOR2X0 U11553 ( .IN1(n11896), .IN2(n11897), .QN(n11895) );
  NAND2X0 U11554 ( .IN1(n11898), .IN2(n11707), .QN(n11897) );
  NOR2X0 U11555 ( .IN1(n11620), .IN2(n11671), .QN(n11898) );
  NAND2X0 U11556 ( .IN1(n11899), .IN2(n11688), .QN(n11896) );
  NOR2X0 U11557 ( .IN1(n11612), .IN2(n11900), .QN(n11899) );
  INVX0 U11558 ( .INP(n11901), .ZN(n11900) );
  NOR2X0 U11559 ( .IN1(n11902), .IN2(n11903), .QN(n11894) );
  NAND2X0 U11560 ( .IN1(n11904), .IN2(n11666), .QN(n11903) );
  NOR2X0 U11561 ( .IN1(n11642), .IN2(n11695), .QN(n11904) );
  NAND2X0 U11562 ( .IN1(n11905), .IN2(n11711), .QN(n11902) );
  NOR2X0 U11563 ( .IN1(n11906), .IN2(n11679), .QN(n11905) );
  NOR2X0 U11564 ( .IN1(n11907), .IN2(n11908), .QN(n11906) );
  NAND2X0 U11565 ( .IN1(n11909), .IN2(n11910), .QN(n11908) );
  NAND2X0 U11566 ( .IN1(n10195), .IN2(g6979), .QN(n11910) );
  NAND2X0 U11567 ( .IN1(n10262), .IN2(g1315), .QN(n11909) );
  NOR2X0 U11568 ( .IN1(n4358), .IN2(g1425), .QN(n11907) );
  NOR2X0 U11569 ( .IN1(n11911), .IN2(n11912), .QN(n11891) );
  NOR2X0 U11570 ( .IN1(n4358), .IN2(g1422), .QN(n11912) );
  NOR2X0 U11571 ( .IN1(n4308), .IN2(g1421), .QN(n11911) );
  NOR2X0 U11572 ( .IN1(n11561), .IN2(n11547), .QN(n2217) );
  INVX0 U11573 ( .INP(n11556), .ZN(n11547) );
  NAND2X0 U11574 ( .IN1(n4353), .IN2(n11913), .QN(n11556) );
  NAND2X0 U11575 ( .IN1(n4304), .IN2(n10035), .QN(n11913) );
  NAND2X0 U11576 ( .IN1(n4304), .IN2(n11914), .QN(n11561) );
  NAND2X0 U11577 ( .IN1(n4353), .IN2(n10035), .QN(n11914) );
  INVX0 U11578 ( .INP(n11915), .ZN(n1689) );
  NOR2X0 U11579 ( .IN1(n11916), .IN2(n11917), .QN(n11915) );
  NOR2X0 U11580 ( .IN1(g2624), .IN2(n10264), .QN(n11917) );
  INVX0 U11581 ( .INP(n11918), .ZN(n1683) );
  INVX0 U11582 ( .INP(n11919), .ZN(n1497) );
  INVX0 U11583 ( .INP(n11920), .ZN(n1335) );
  NOR2X0 U11584 ( .IN1(n11921), .IN2(n11922), .QN(n11920) );
  NOR2X0 U11585 ( .IN1(g1930), .IN2(n10265), .QN(n11922) );
  INVX0 U11586 ( .INP(n11923), .ZN(n1146) );
  NAND2X0 U11587 ( .IN1(n11924), .IN2(n11925), .QN(g30801) );
  INVX0 U11588 ( .INP(n11926), .ZN(n11925) );
  NOR2X0 U11589 ( .IN1(g3109), .IN2(n4334), .QN(n11926) );
  NAND2X0 U11590 ( .IN1(g30072), .IN2(g3109), .QN(n11924) );
  NAND2X0 U11591 ( .IN1(n11927), .IN2(n11928), .QN(g30798) );
  INVX0 U11592 ( .INP(n11929), .ZN(n11928) );
  NOR2X0 U11593 ( .IN1(g8030), .IN2(n4437), .QN(n11929) );
  NAND2X0 U11594 ( .IN1(g30072), .IN2(g8030), .QN(n11927) );
  NAND2X0 U11595 ( .IN1(n11930), .IN2(n11931), .QN(g30796) );
  INVX0 U11596 ( .INP(n11932), .ZN(n11931) );
  NOR2X0 U11597 ( .IN1(g8106), .IN2(n4438), .QN(n11932) );
  NAND2X0 U11598 ( .IN1(g30072), .IN2(g8106), .QN(n11930) );
  NAND2X0 U11599 ( .IN1(n11933), .IN2(n11934), .QN(g30709) );
  NAND2X0 U11600 ( .IN1(n11935), .IN2(g7264), .QN(n11934) );
  INVX0 U11601 ( .INP(n11936), .ZN(n11933) );
  NOR2X0 U11602 ( .IN1(n11937), .IN2(n9535), .QN(n11936) );
  NAND2X0 U11603 ( .IN1(n11938), .IN2(n11939), .QN(g30708) );
  NAND2X0 U11604 ( .IN1(n11940), .IN2(n4618), .QN(n11939) );
  NAND2X0 U11605 ( .IN1(n4511), .IN2(g1698), .QN(n11938) );
  NAND2X0 U11606 ( .IN1(n11941), .IN2(n11942), .QN(g30707) );
  NAND2X0 U11607 ( .IN1(n11935), .IN2(g5555), .QN(n11942) );
  NAND2X0 U11608 ( .IN1(n4516), .IN2(g2390), .QN(n11941) );
  NAND2X0 U11609 ( .IN1(n11943), .IN2(n11944), .QN(g30706) );
  NAND2X0 U11610 ( .IN1(n11940), .IN2(g7014), .QN(n11944) );
  INVX0 U11611 ( .INP(n11945), .ZN(n11943) );
  NOR2X0 U11612 ( .IN1(n11946), .IN2(n9538), .QN(n11945) );
  NAND2X0 U11613 ( .IN1(n11947), .IN2(n11948), .QN(g30705) );
  INVX0 U11614 ( .INP(n11949), .ZN(n11948) );
  NOR2X0 U11615 ( .IN1(g1088), .IN2(n9556), .QN(n11949) );
  NAND2X0 U11616 ( .IN1(n2594), .IN2(g1088), .QN(n11947) );
  NAND2X0 U11617 ( .IN1(n11950), .IN2(n11951), .QN(g30704) );
  NAND2X0 U11618 ( .IN1(n11940), .IN2(g5511), .QN(n11951) );
  NOR2X0 U11619 ( .IN1(n11952), .IN2(n11953), .QN(n11940) );
  NAND2X0 U11620 ( .IN1(n11954), .IN2(n11955), .QN(n11952) );
  NAND2X0 U11621 ( .IN1(n11956), .IN2(n11957), .QN(n11955) );
  INVX0 U11622 ( .INP(n11958), .ZN(n11954) );
  NOR2X0 U11623 ( .IN1(n11956), .IN2(n11957), .QN(n11958) );
  NAND2X0 U11624 ( .IN1(n11959), .IN2(n11960), .QN(n11957) );
  NAND2X0 U11625 ( .IN1(n11961), .IN2(n11962), .QN(n11960) );
  NAND2X0 U11626 ( .IN1(n11963), .IN2(n11964), .QN(n11959) );
  NAND2X0 U11627 ( .IN1(n11965), .IN2(n11966), .QN(n11963) );
  NAND2X0 U11628 ( .IN1(n11967), .IN2(n11956), .QN(n11966) );
  NAND2X0 U11629 ( .IN1(n3070), .IN2(n11968), .QN(n11967) );
  NAND2X0 U11630 ( .IN1(n11969), .IN2(n11970), .QN(n11968) );
  NAND2X0 U11631 ( .IN1(n11971), .IN2(n11972), .QN(n11970) );
  INVX0 U11632 ( .INP(n11973), .ZN(n11972) );
  NOR2X0 U11633 ( .IN1(n11974), .IN2(n11975), .QN(n11971) );
  INVX0 U11634 ( .INP(n11976), .ZN(n11969) );
  NAND2X0 U11635 ( .IN1(n11977), .IN2(n11978), .QN(n11965) );
  NAND2X0 U11636 ( .IN1(n11979), .IN2(n11980), .QN(n11977) );
  NAND2X0 U11637 ( .IN1(n11981), .IN2(n11975), .QN(n11980) );
  NOR2X0 U11638 ( .IN1(n11982), .IN2(n11983), .QN(n11981) );
  NAND2X0 U11639 ( .IN1(n11984), .IN2(n11985), .QN(n11979) );
  NOR2X0 U11640 ( .IN1(n11986), .IN2(n11987), .QN(n11984) );
  NAND2X0 U11641 ( .IN1(n11988), .IN2(n11989), .QN(n11987) );
  NAND2X0 U11642 ( .IN1(n11983), .IN2(n11990), .QN(n11989) );
  NAND2X0 U11643 ( .IN1(n4518), .IN2(g1696), .QN(n11950) );
  NAND2X0 U11644 ( .IN1(n11991), .IN2(n11992), .QN(g30703) );
  NAND2X0 U11645 ( .IN1(n4364), .IN2(g1003), .QN(n11992) );
  NAND2X0 U11646 ( .IN1(n2594), .IN2(g6712), .QN(n11991) );
  NAND2X0 U11647 ( .IN1(n11993), .IN2(n11994), .QN(g30702) );
  NAND2X0 U11648 ( .IN1(n11995), .IN2(n4640), .QN(n11994) );
  NAND2X0 U11649 ( .IN1(n4506), .IN2(g317), .QN(n11993) );
  NAND2X0 U11650 ( .IN1(n11996), .IN2(n11997), .QN(g30701) );
  NAND2X0 U11651 ( .IN1(n4363), .IN2(g1002), .QN(n11997) );
  NAND2X0 U11652 ( .IN1(n2594), .IN2(g5472), .QN(n11996) );
  NAND2X0 U11653 ( .IN1(n11998), .IN2(n11999), .QN(g30700) );
  NAND2X0 U11654 ( .IN1(n11995), .IN2(g6447), .QN(n11999) );
  NAND2X0 U11655 ( .IN1(test_so18), .IN2(n4499), .QN(n11998) );
  NAND2X0 U11656 ( .IN1(n12000), .IN2(n12001), .QN(g30699) );
  NAND2X0 U11657 ( .IN1(n11995), .IN2(g5437), .QN(n12001) );
  NOR2X0 U11658 ( .IN1(n12002), .IN2(n12003), .QN(n11995) );
  NAND2X0 U11659 ( .IN1(n12004), .IN2(n12005), .QN(n12002) );
  NAND2X0 U11660 ( .IN1(n12006), .IN2(n12007), .QN(n12005) );
  INVX0 U11661 ( .INP(n12008), .ZN(n12004) );
  NOR2X0 U11662 ( .IN1(n12006), .IN2(n12007), .QN(n12008) );
  NAND2X0 U11663 ( .IN1(n12009), .IN2(n12010), .QN(n12007) );
  NAND2X0 U11664 ( .IN1(n12011), .IN2(n12012), .QN(n12010) );
  NAND2X0 U11665 ( .IN1(n12013), .IN2(n12014), .QN(n12009) );
  NAND2X0 U11666 ( .IN1(n12015), .IN2(n12016), .QN(n12013) );
  NAND2X0 U11667 ( .IN1(n12017), .IN2(n12006), .QN(n12016) );
  NAND2X0 U11668 ( .IN1(n3130), .IN2(n12018), .QN(n12017) );
  NAND2X0 U11669 ( .IN1(n12019), .IN2(n12020), .QN(n12018) );
  NAND2X0 U11670 ( .IN1(n12021), .IN2(n12022), .QN(n12020) );
  INVX0 U11671 ( .INP(n12023), .ZN(n12022) );
  NOR2X0 U11672 ( .IN1(n12024), .IN2(n12025), .QN(n12021) );
  INVX0 U11673 ( .INP(n12026), .ZN(n12019) );
  NAND2X0 U11674 ( .IN1(n12027), .IN2(n12028), .QN(n12015) );
  NAND2X0 U11675 ( .IN1(n12029), .IN2(n12030), .QN(n12027) );
  NAND2X0 U11676 ( .IN1(n12031), .IN2(n12025), .QN(n12030) );
  NOR2X0 U11677 ( .IN1(n12032), .IN2(n12033), .QN(n12031) );
  NAND2X0 U11678 ( .IN1(n12034), .IN2(n12035), .QN(n12029) );
  NOR2X0 U11679 ( .IN1(n12036), .IN2(n12037), .QN(n12034) );
  NAND2X0 U11680 ( .IN1(n12038), .IN2(n12039), .QN(n12037) );
  NAND2X0 U11681 ( .IN1(n12033), .IN2(n12040), .QN(n12039) );
  INVX0 U11682 ( .INP(n12041), .ZN(n12000) );
  NOR2X0 U11683 ( .IN1(n12042), .IN2(n9564), .QN(n12041) );
  NAND2X0 U11684 ( .IN1(n12043), .IN2(n12044), .QN(g30695) );
  INVX0 U11685 ( .INP(n12045), .ZN(n12044) );
  NOR2X0 U11686 ( .IN1(g2241), .IN2(n9577), .QN(n12045) );
  NAND2X0 U11687 ( .IN1(n12046), .IN2(g2241), .QN(n12043) );
  NAND2X0 U11688 ( .IN1(n12047), .IN2(n12048), .QN(g30694) );
  INVX0 U11689 ( .INP(n12049), .ZN(n12048) );
  NOR2X0 U11690 ( .IN1(g2241), .IN2(n9417), .QN(n12049) );
  NAND2X0 U11691 ( .IN1(n12050), .IN2(g2241), .QN(n12047) );
  NAND2X0 U11692 ( .IN1(n12051), .IN2(n12052), .QN(g30693) );
  NAND2X0 U11693 ( .IN1(g2273), .IN2(n10320), .QN(n12052) );
  NAND2X0 U11694 ( .IN1(test_so73), .IN2(n12046), .QN(n12051) );
  NAND2X0 U11695 ( .IN1(n12053), .IN2(n12054), .QN(g30692) );
  INVX0 U11696 ( .INP(n12055), .ZN(n12054) );
  NOR2X0 U11697 ( .IN1(g1547), .IN2(n9580), .QN(n12055) );
  NAND2X0 U11698 ( .IN1(n12056), .IN2(g1547), .QN(n12053) );
  NAND2X0 U11699 ( .IN1(n12057), .IN2(n12058), .QN(g30691) );
  NAND2X0 U11700 ( .IN1(g2345), .IN2(n10320), .QN(n12058) );
  NAND2X0 U11701 ( .IN1(n12050), .IN2(test_so73), .QN(n12057) );
  NAND2X0 U11702 ( .IN1(n12059), .IN2(n12060), .QN(g30690) );
  INVX0 U11703 ( .INP(n12061), .ZN(n12060) );
  NOR2X0 U11704 ( .IN1(g6837), .IN2(n9480), .QN(n12061) );
  NAND2X0 U11705 ( .IN1(n12046), .IN2(g6837), .QN(n12059) );
  NAND2X0 U11706 ( .IN1(n12062), .IN2(n12063), .QN(n12046) );
  NAND2X0 U11707 ( .IN1(n12064), .IN2(g2175), .QN(n12063) );
  NOR2X0 U11708 ( .IN1(n12065), .IN2(n12066), .QN(n12062) );
  NOR2X0 U11709 ( .IN1(n12067), .IN2(n12068), .QN(n12066) );
  NAND2X0 U11710 ( .IN1(n12069), .IN2(n12070), .QN(n12068) );
  NAND2X0 U11711 ( .IN1(n10962), .IN2(n12071), .QN(n12070) );
  NAND2X0 U11712 ( .IN1(n12072), .IN2(n10961), .QN(n12069) );
  NAND2X0 U11713 ( .IN1(n12073), .IN2(n12074), .QN(g30689) );
  INVX0 U11714 ( .INP(n12075), .ZN(n12074) );
  NOR2X0 U11715 ( .IN1(g1547), .IN2(n9454), .QN(n12075) );
  NAND2X0 U11716 ( .IN1(n12076), .IN2(g1547), .QN(n12073) );
  NAND2X0 U11717 ( .IN1(n12077), .IN2(n12078), .QN(g30688) );
  NAND2X0 U11718 ( .IN1(n4515), .IN2(g1579), .QN(n12078) );
  NAND2X0 U11719 ( .IN1(n12056), .IN2(g6782), .QN(n12077) );
  NAND2X0 U11720 ( .IN1(n12079), .IN2(n12080), .QN(g30687) );
  NAND2X0 U11721 ( .IN1(g888), .IN2(n10321), .QN(n12080) );
  NAND2X0 U11722 ( .IN1(test_so31), .IN2(n12081), .QN(n12079) );
  NAND2X0 U11723 ( .IN1(n12082), .IN2(n12083), .QN(g30686) );
  INVX0 U11724 ( .INP(n12084), .ZN(n12083) );
  NOR2X0 U11725 ( .IN1(g6837), .IN2(n9418), .QN(n12084) );
  NAND2X0 U11726 ( .IN1(n12050), .IN2(g6837), .QN(n12082) );
  INVX0 U11727 ( .INP(n12085), .ZN(n12050) );
  NAND2X0 U11728 ( .IN1(n12086), .IN2(n12087), .QN(n12085) );
  NAND2X0 U11729 ( .IN1(n12064), .IN2(n12088), .QN(n12087) );
  NOR2X0 U11730 ( .IN1(n12089), .IN2(n12090), .QN(n12086) );
  NOR2X0 U11731 ( .IN1(n12067), .IN2(n12091), .QN(n12090) );
  NAND2X0 U11732 ( .IN1(n12092), .IN2(n12093), .QN(n12091) );
  NAND2X0 U11733 ( .IN1(n2669), .IN2(n10986), .QN(n12093) );
  INVX0 U11734 ( .INP(n12094), .ZN(n12092) );
  NOR2X0 U11735 ( .IN1(n10986), .IN2(n2669), .QN(n12094) );
  NAND2X0 U11736 ( .IN1(n12095), .IN2(n12096), .QN(g30684) );
  NAND2X0 U11737 ( .IN1(n4515), .IN2(g1651), .QN(n12096) );
  NAND2X0 U11738 ( .IN1(n12076), .IN2(g6782), .QN(n12095) );
  NAND2X0 U11739 ( .IN1(n12097), .IN2(n12098), .QN(g30683) );
  INVX0 U11740 ( .INP(n12099), .ZN(n12098) );
  NOR2X0 U11741 ( .IN1(g6573), .IN2(n9492), .QN(n12099) );
  NAND2X0 U11742 ( .IN1(n12056), .IN2(g6573), .QN(n12097) );
  NAND2X0 U11743 ( .IN1(n12100), .IN2(n12101), .QN(n12056) );
  NOR2X0 U11744 ( .IN1(n12102), .IN2(n12103), .QN(n12100) );
  NOR2X0 U11745 ( .IN1(n4320), .IN2(n12104), .QN(n12103) );
  NOR2X0 U11746 ( .IN1(n12105), .IN2(n12106), .QN(n12102) );
  NAND2X0 U11747 ( .IN1(n12107), .IN2(n12108), .QN(n12106) );
  NAND2X0 U11748 ( .IN1(n10897), .IN2(n12109), .QN(n12108) );
  NAND2X0 U11749 ( .IN1(n12110), .IN2(n10896), .QN(n12107) );
  NAND2X0 U11750 ( .IN1(n12111), .IN2(n12112), .QN(g30682) );
  NAND2X0 U11751 ( .IN1(g960), .IN2(n10321), .QN(n12112) );
  NAND2X0 U11752 ( .IN1(n12113), .IN2(test_so31), .QN(n12111) );
  NAND2X0 U11753 ( .IN1(n12114), .IN2(n12115), .QN(g30681) );
  INVX0 U11754 ( .INP(n12116), .ZN(n12115) );
  NOR2X0 U11755 ( .IN1(g6518), .IN2(n9506), .QN(n12116) );
  NAND2X0 U11756 ( .IN1(n12081), .IN2(g6518), .QN(n12114) );
  NAND2X0 U11757 ( .IN1(n12117), .IN2(n12118), .QN(g30680) );
  INVX0 U11758 ( .INP(n12119), .ZN(n12118) );
  NOR2X0 U11759 ( .IN1(g165), .IN2(n9586), .QN(n12119) );
  NAND2X0 U11760 ( .IN1(n12120), .IN2(g165), .QN(n12117) );
  NAND2X0 U11761 ( .IN1(n12121), .IN2(n12122), .QN(g30679) );
  INVX0 U11762 ( .INP(n12123), .ZN(n12122) );
  NOR2X0 U11763 ( .IN1(g2241), .IN2(n9460), .QN(n12123) );
  NAND2X0 U11764 ( .IN1(n12124), .IN2(g2241), .QN(n12121) );
  NAND2X0 U11765 ( .IN1(n12125), .IN2(n12126), .QN(g30678) );
  INVX0 U11766 ( .INP(n12127), .ZN(n12126) );
  NOR2X0 U11767 ( .IN1(g6573), .IN2(n9453), .QN(n12127) );
  NAND2X0 U11768 ( .IN1(n12076), .IN2(g6573), .QN(n12125) );
  INVX0 U11769 ( .INP(n12128), .ZN(n12076) );
  NAND2X0 U11770 ( .IN1(n12129), .IN2(n12130), .QN(n12128) );
  NAND2X0 U11771 ( .IN1(n12131), .IN2(n12132), .QN(n12130) );
  NOR2X0 U11772 ( .IN1(n12133), .IN2(n12134), .QN(n12129) );
  NOR2X0 U11773 ( .IN1(n12105), .IN2(n12135), .QN(n12134) );
  NAND2X0 U11774 ( .IN1(n12136), .IN2(n12137), .QN(n12135) );
  NAND2X0 U11775 ( .IN1(n2684), .IN2(n10929), .QN(n12137) );
  INVX0 U11776 ( .INP(n12138), .ZN(n12136) );
  NOR2X0 U11777 ( .IN1(n10929), .IN2(n2684), .QN(n12138) );
  NAND2X0 U11778 ( .IN1(n12139), .IN2(n12140), .QN(g30677) );
  INVX0 U11779 ( .INP(n12141), .ZN(n12140) );
  NOR2X0 U11780 ( .IN1(g6518), .IN2(n9532), .QN(n12141) );
  NAND2X0 U11781 ( .IN1(n12113), .IN2(g6518), .QN(n12139) );
  NAND2X0 U11782 ( .IN1(n12142), .IN2(n12143), .QN(g30676) );
  INVX0 U11783 ( .INP(n12144), .ZN(n12143) );
  NOR2X0 U11784 ( .IN1(g6368), .IN2(n9507), .QN(n12144) );
  NAND2X0 U11785 ( .IN1(n12081), .IN2(g6368), .QN(n12142) );
  NAND2X0 U11786 ( .IN1(n12145), .IN2(n12146), .QN(n12081) );
  NAND2X0 U11787 ( .IN1(n12147), .IN2(g793), .QN(n12146) );
  NOR2X0 U11788 ( .IN1(n12148), .IN2(n12149), .QN(n12145) );
  NOR2X0 U11789 ( .IN1(n12150), .IN2(n12151), .QN(n12149) );
  NAND2X0 U11790 ( .IN1(n12152), .IN2(n12153), .QN(n12151) );
  NAND2X0 U11791 ( .IN1(n10861), .IN2(n12154), .QN(n12153) );
  NAND2X0 U11792 ( .IN1(n12155), .IN2(n10860), .QN(n12152) );
  NAND2X0 U11793 ( .IN1(n12156), .IN2(n12157), .QN(g30675) );
  INVX0 U11794 ( .INP(n12158), .ZN(n12157) );
  NOR2X0 U11795 ( .IN1(g165), .IN2(n9457), .QN(n12158) );
  NAND2X0 U11796 ( .IN1(n12159), .IN2(g165), .QN(n12156) );
  NAND2X0 U11797 ( .IN1(n12160), .IN2(n12161), .QN(g30674) );
  NAND2X0 U11798 ( .IN1(n4512), .IN2(g198), .QN(n12161) );
  NAND2X0 U11799 ( .IN1(n12120), .IN2(g6313), .QN(n12160) );
  NAND2X0 U11800 ( .IN1(n12162), .IN2(n12163), .QN(g30673) );
  NAND2X0 U11801 ( .IN1(g2318), .IN2(n10320), .QN(n12163) );
  NAND2X0 U11802 ( .IN1(n12124), .IN2(test_so73), .QN(n12162) );
  NAND2X0 U11803 ( .IN1(n12164), .IN2(n12165), .QN(g30672) );
  INVX0 U11804 ( .INP(n12166), .ZN(n12165) );
  NOR2X0 U11805 ( .IN1(g2241), .IN2(n9461), .QN(n12166) );
  NAND2X0 U11806 ( .IN1(n12167), .IN2(g2241), .QN(n12164) );
  NAND2X0 U11807 ( .IN1(n12168), .IN2(n12169), .QN(g30671) );
  INVX0 U11808 ( .INP(n12170), .ZN(n12169) );
  NOR2X0 U11809 ( .IN1(g1547), .IN2(n9463), .QN(n12170) );
  NAND2X0 U11810 ( .IN1(n12171), .IN2(g1547), .QN(n12168) );
  NAND2X0 U11811 ( .IN1(n12172), .IN2(n12173), .QN(g30670) );
  INVX0 U11812 ( .INP(n12174), .ZN(n12173) );
  NOR2X0 U11813 ( .IN1(g6368), .IN2(n9496), .QN(n12174) );
  NAND2X0 U11814 ( .IN1(n12113), .IN2(g6368), .QN(n12172) );
  INVX0 U11815 ( .INP(n12175), .ZN(n12113) );
  NAND2X0 U11816 ( .IN1(n12176), .IN2(n12177), .QN(n12175) );
  NAND2X0 U11817 ( .IN1(n12147), .IN2(n12178), .QN(n12177) );
  NOR2X0 U11818 ( .IN1(n12179), .IN2(n12180), .QN(n12176) );
  NOR2X0 U11819 ( .IN1(n12181), .IN2(n12150), .QN(n12180) );
  NOR2X0 U11820 ( .IN1(n12182), .IN2(n12183), .QN(n12181) );
  NOR2X0 U11821 ( .IN1(n10857), .IN2(n12184), .QN(n12183) );
  INVX0 U11822 ( .INP(n12185), .ZN(n12182) );
  NAND2X0 U11823 ( .IN1(n12184), .IN2(n10857), .QN(n12185) );
  NAND2X0 U11824 ( .IN1(n12186), .IN2(n12187), .QN(n12184) );
  NAND2X0 U11825 ( .IN1(n12188), .IN2(n12189), .QN(n12187) );
  NAND2X0 U11826 ( .IN1(n10865), .IN2(n12190), .QN(n12189) );
  NAND2X0 U11827 ( .IN1(n12191), .IN2(n10864), .QN(n12188) );
  NAND2X0 U11828 ( .IN1(n12192), .IN2(n12193), .QN(g30669) );
  NAND2X0 U11829 ( .IN1(n4512), .IN2(g270), .QN(n12193) );
  NAND2X0 U11830 ( .IN1(n12159), .IN2(g6313), .QN(n12192) );
  NAND2X0 U11831 ( .IN1(n12194), .IN2(n12195), .QN(g30668) );
  INVX0 U11832 ( .INP(n12196), .ZN(n12195) );
  NOR2X0 U11833 ( .IN1(g6231), .IN2(n9521), .QN(n12196) );
  NAND2X0 U11834 ( .IN1(n12120), .IN2(g6231), .QN(n12194) );
  NAND2X0 U11835 ( .IN1(n12197), .IN2(n12198), .QN(n12120) );
  NOR2X0 U11836 ( .IN1(n12199), .IN2(n12200), .QN(n12197) );
  NOR2X0 U11837 ( .IN1(n4322), .IN2(n12201), .QN(n12200) );
  NOR2X0 U11838 ( .IN1(n12202), .IN2(n12203), .QN(n12199) );
  NAND2X0 U11839 ( .IN1(n12204), .IN2(n12205), .QN(n12203) );
  NAND2X0 U11840 ( .IN1(n10767), .IN2(n12206), .QN(n12205) );
  NAND2X0 U11841 ( .IN1(n12207), .IN2(n10766), .QN(n12204) );
  NAND2X0 U11842 ( .IN1(n12208), .IN2(n12209), .QN(g30667) );
  INVX0 U11843 ( .INP(n12210), .ZN(n12209) );
  NOR2X0 U11844 ( .IN1(g6837), .IN2(n9478), .QN(n12210) );
  NAND2X0 U11845 ( .IN1(n12124), .IN2(g6837), .QN(n12208) );
  INVX0 U11846 ( .INP(n12211), .ZN(n12124) );
  NAND2X0 U11847 ( .IN1(n12212), .IN2(n12213), .QN(n12211) );
  NAND2X0 U11848 ( .IN1(n12064), .IN2(n4389), .QN(n12213) );
  NOR2X0 U11849 ( .IN1(n12089), .IN2(n12214), .QN(n12212) );
  NOR2X0 U11850 ( .IN1(n12067), .IN2(n12215), .QN(n12214) );
  NAND2X0 U11851 ( .IN1(n12216), .IN2(n12217), .QN(n12215) );
  NAND2X0 U11852 ( .IN1(n12218), .IN2(n10990), .QN(n12217) );
  NAND2X0 U11853 ( .IN1(n12072), .IN2(n12219), .QN(n12218) );
  NAND2X0 U11854 ( .IN1(n12220), .IN2(n12221), .QN(n12219) );
  NAND2X0 U11855 ( .IN1(n10962), .IN2(n11780), .QN(n12221) );
  NAND2X0 U11856 ( .IN1(n4529), .IN2(n10961), .QN(n12220) );
  NAND2X0 U11857 ( .IN1(n12222), .IN2(n10991), .QN(n12216) );
  NOR2X0 U11858 ( .IN1(n12223), .IN2(n12224), .QN(n12222) );
  NOR2X0 U11859 ( .IN1(n10962), .IN2(n4529), .QN(n12223) );
  NAND2X0 U11860 ( .IN1(n12225), .IN2(n12226), .QN(g30666) );
  NAND2X0 U11861 ( .IN1(g2309), .IN2(n10320), .QN(n12226) );
  NAND2X0 U11862 ( .IN1(n12167), .IN2(test_so73), .QN(n12225) );
  NAND2X0 U11863 ( .IN1(n12227), .IN2(n12228), .QN(g30665) );
  INVX0 U11864 ( .INP(n12229), .ZN(n12228) );
  NOR2X0 U11865 ( .IN1(g2241), .IN2(n9425), .QN(n12229) );
  NAND2X0 U11866 ( .IN1(n12230), .IN2(g2241), .QN(n12227) );
  NAND2X0 U11867 ( .IN1(n12231), .IN2(n12232), .QN(g30664) );
  NAND2X0 U11868 ( .IN1(n4515), .IN2(g1624), .QN(n12232) );
  NAND2X0 U11869 ( .IN1(n12171), .IN2(g6782), .QN(n12231) );
  NAND2X0 U11870 ( .IN1(n12233), .IN2(n12234), .QN(g30663) );
  INVX0 U11871 ( .INP(n12235), .ZN(n12234) );
  NOR2X0 U11872 ( .IN1(g1547), .IN2(n9464), .QN(n12235) );
  NAND2X0 U11873 ( .IN1(n12236), .IN2(g1547), .QN(n12233) );
  NAND2X0 U11874 ( .IN1(n12237), .IN2(n12238), .QN(g30662) );
  NAND2X0 U11875 ( .IN1(g933), .IN2(n10321), .QN(n12238) );
  NAND2X0 U11876 ( .IN1(n12239), .IN2(test_so31), .QN(n12237) );
  NAND2X0 U11877 ( .IN1(n12240), .IN2(n12241), .QN(g30661) );
  INVX0 U11878 ( .INP(n12242), .ZN(n12241) );
  NOR2X0 U11879 ( .IN1(g6231), .IN2(n9456), .QN(n12242) );
  NAND2X0 U11880 ( .IN1(n12159), .IN2(g6231), .QN(n12240) );
  INVX0 U11881 ( .INP(n12243), .ZN(n12159) );
  NAND2X0 U11882 ( .IN1(n12244), .IN2(n12245), .QN(n12243) );
  NAND2X0 U11883 ( .IN1(n12246), .IN2(n12247), .QN(n12245) );
  NOR2X0 U11884 ( .IN1(n12248), .IN2(n12249), .QN(n12244) );
  NOR2X0 U11885 ( .IN1(n12202), .IN2(n12250), .QN(n12249) );
  NAND2X0 U11886 ( .IN1(n12251), .IN2(n12252), .QN(n12250) );
  NAND2X0 U11887 ( .IN1(n2717), .IN2(n10792), .QN(n12252) );
  INVX0 U11888 ( .INP(n12253), .ZN(n12251) );
  NOR2X0 U11889 ( .IN1(n10792), .IN2(n2717), .QN(n12253) );
  NAND2X0 U11890 ( .IN1(n12254), .IN2(n12255), .QN(g30660) );
  INVX0 U11891 ( .INP(n12256), .ZN(n12255) );
  NOR2X0 U11892 ( .IN1(g6837), .IN2(n9481), .QN(n12256) );
  NAND2X0 U11893 ( .IN1(n12167), .IN2(g6837), .QN(n12254) );
  INVX0 U11894 ( .INP(n12257), .ZN(n12167) );
  NAND2X0 U11895 ( .IN1(n12258), .IN2(n12259), .QN(n12257) );
  NAND2X0 U11896 ( .IN1(n12064), .IN2(n4373), .QN(n12259) );
  NOR2X0 U11897 ( .IN1(n12089), .IN2(n12260), .QN(n12258) );
  NOR2X0 U11898 ( .IN1(n12261), .IN2(n12067), .QN(n12260) );
  NOR2X0 U11899 ( .IN1(n12262), .IN2(n12263), .QN(n12261) );
  NOR2X0 U11900 ( .IN1(n12264), .IN2(n10978), .QN(n12263) );
  NOR2X0 U11901 ( .IN1(n12265), .IN2(n12266), .QN(n12262) );
  NOR2X0 U11902 ( .IN1(n12267), .IN2(n11780), .QN(n12089) );
  NAND2X0 U11903 ( .IN1(n12268), .IN2(n12269), .QN(g30659) );
  NAND2X0 U11904 ( .IN1(g2300), .IN2(n10320), .QN(n12269) );
  NAND2X0 U11905 ( .IN1(test_so73), .IN2(n12230), .QN(n12268) );
  NAND2X0 U11906 ( .IN1(n12270), .IN2(n12271), .QN(g30658) );
  NAND2X0 U11907 ( .IN1(n12171), .IN2(g6573), .QN(n12271) );
  INVX0 U11908 ( .INP(n12272), .ZN(n12171) );
  NAND2X0 U11909 ( .IN1(n12273), .IN2(n12274), .QN(n12272) );
  NAND2X0 U11910 ( .IN1(n12131), .IN2(n4390), .QN(n12274) );
  NOR2X0 U11911 ( .IN1(n12133), .IN2(n12275), .QN(n12273) );
  NOR2X0 U11912 ( .IN1(n12105), .IN2(n12276), .QN(n12275) );
  NAND2X0 U11913 ( .IN1(n12277), .IN2(n12278), .QN(n12276) );
  NAND2X0 U11914 ( .IN1(n12279), .IN2(n10913), .QN(n12278) );
  NAND2X0 U11915 ( .IN1(n12110), .IN2(n12280), .QN(n12279) );
  NAND2X0 U11916 ( .IN1(n12281), .IN2(n12282), .QN(n12280) );
  NAND2X0 U11917 ( .IN1(n10897), .IN2(n11777), .QN(n12282) );
  NAND2X0 U11918 ( .IN1(n4530), .IN2(n10896), .QN(n12281) );
  NAND2X0 U11919 ( .IN1(n12283), .IN2(n10914), .QN(n12277) );
  NOR2X0 U11920 ( .IN1(n12284), .IN2(n12285), .QN(n12283) );
  NOR2X0 U11921 ( .IN1(n10897), .IN2(n4530), .QN(n12284) );
  NAND2X0 U11922 ( .IN1(test_so55), .IN2(n4317), .QN(n12270) );
  NAND2X0 U11923 ( .IN1(n12286), .IN2(n12287), .QN(g30657) );
  NAND2X0 U11924 ( .IN1(n4515), .IN2(g1615), .QN(n12287) );
  NAND2X0 U11925 ( .IN1(n12236), .IN2(g6782), .QN(n12286) );
  NAND2X0 U11926 ( .IN1(n12288), .IN2(n12289), .QN(g30656) );
  INVX0 U11927 ( .INP(n12290), .ZN(n12289) );
  NOR2X0 U11928 ( .IN1(g1547), .IN2(n9426), .QN(n12290) );
  NAND2X0 U11929 ( .IN1(n12291), .IN2(g1547), .QN(n12288) );
  NAND2X0 U11930 ( .IN1(n12292), .IN2(n12293), .QN(g30655) );
  INVX0 U11931 ( .INP(n12294), .ZN(n12293) );
  NOR2X0 U11932 ( .IN1(g6518), .IN2(n9528), .QN(n12294) );
  NAND2X0 U11933 ( .IN1(n12239), .IN2(g6518), .QN(n12292) );
  NAND2X0 U11934 ( .IN1(n12295), .IN2(n12296), .QN(g30654) );
  NAND2X0 U11935 ( .IN1(test_so34), .IN2(n10321), .QN(n12296) );
  NAND2X0 U11936 ( .IN1(n12297), .IN2(test_so31), .QN(n12295) );
  NAND2X0 U11937 ( .IN1(n12298), .IN2(n12299), .QN(g30653) );
  INVX0 U11938 ( .INP(n12300), .ZN(n12299) );
  NOR2X0 U11939 ( .IN1(g165), .IN2(n9469), .QN(n12300) );
  NAND2X0 U11940 ( .IN1(n12301), .IN2(g165), .QN(n12298) );
  NAND2X0 U11941 ( .IN1(n12302), .IN2(n12303), .QN(g30652) );
  INVX0 U11942 ( .INP(n12304), .ZN(n12303) );
  NOR2X0 U11943 ( .IN1(g6837), .IN2(n9419), .QN(n12304) );
  NAND2X0 U11944 ( .IN1(n12230), .IN2(g6837), .QN(n12302) );
  NAND2X0 U11945 ( .IN1(n12305), .IN2(n12306), .QN(n12230) );
  NAND2X0 U11946 ( .IN1(n12064), .IN2(n12307), .QN(n12306) );
  NOR2X0 U11947 ( .IN1(n12065), .IN2(n12308), .QN(n12305) );
  NOR2X0 U11948 ( .IN1(n12067), .IN2(n12309), .QN(n12308) );
  NAND2X0 U11949 ( .IN1(n12310), .IN2(n12311), .QN(n12309) );
  NAND2X0 U11950 ( .IN1(n10966), .IN2(n2670), .QN(n12311) );
  INVX0 U11951 ( .INP(n12312), .ZN(n12310) );
  NOR2X0 U11952 ( .IN1(n10966), .IN2(n2670), .QN(n12312) );
  NAND2X0 U11953 ( .IN1(n12313), .IN2(n12314), .QN(n2670) );
  NAND2X0 U11954 ( .IN1(n12315), .IN2(n12316), .QN(n12314) );
  NAND2X0 U11955 ( .IN1(n10950), .IN2(n11780), .QN(n12316) );
  NAND2X0 U11956 ( .IN1(n4529), .IN2(n10949), .QN(n12315) );
  NOR2X0 U11957 ( .IN1(n12267), .IN2(n4529), .QN(n12065) );
  INVX0 U11958 ( .INP(n12317), .ZN(n12267) );
  NAND2X0 U11959 ( .IN1(n12318), .IN2(n12319), .QN(g30651) );
  INVX0 U11960 ( .INP(n12320), .ZN(n12319) );
  NOR2X0 U11961 ( .IN1(g6573), .IN2(n9493), .QN(n12320) );
  NAND2X0 U11962 ( .IN1(n12236), .IN2(g6573), .QN(n12318) );
  INVX0 U11963 ( .INP(n12321), .ZN(n12236) );
  NAND2X0 U11964 ( .IN1(n12322), .IN2(n12323), .QN(n12321) );
  NAND2X0 U11965 ( .IN1(n12131), .IN2(n4374), .QN(n12323) );
  NOR2X0 U11966 ( .IN1(n12133), .IN2(n12324), .QN(n12322) );
  NOR2X0 U11967 ( .IN1(n12325), .IN2(n12105), .QN(n12324) );
  NOR2X0 U11968 ( .IN1(n12326), .IN2(n12327), .QN(n12325) );
  NOR2X0 U11969 ( .IN1(n12328), .IN2(n10921), .QN(n12327) );
  NOR2X0 U11970 ( .IN1(n10922), .IN2(n12329), .QN(n12326) );
  INVX0 U11971 ( .INP(n12330), .ZN(n12133) );
  NAND2X0 U11972 ( .IN1(n12331), .IN2(n4530), .QN(n12330) );
  NAND2X0 U11973 ( .IN1(n12332), .IN2(n12333), .QN(g30650) );
  NAND2X0 U11974 ( .IN1(test_so56), .IN2(n4515), .QN(n12333) );
  NAND2X0 U11975 ( .IN1(n12291), .IN2(g6782), .QN(n12332) );
  NAND2X0 U11976 ( .IN1(n12334), .IN2(n12335), .QN(g30649) );
  INVX0 U11977 ( .INP(n12336), .ZN(n12335) );
  NOR2X0 U11978 ( .IN1(g6368), .IN2(n9505), .QN(n12336) );
  NAND2X0 U11979 ( .IN1(n12239), .IN2(g6368), .QN(n12334) );
  INVX0 U11980 ( .INP(n12337), .ZN(n12239) );
  NAND2X0 U11981 ( .IN1(n12338), .IN2(n12339), .QN(n12337) );
  NAND2X0 U11982 ( .IN1(n12147), .IN2(n4391), .QN(n12339) );
  NOR2X0 U11983 ( .IN1(n12179), .IN2(n12340), .QN(n12338) );
  NOR2X0 U11984 ( .IN1(n12341), .IN2(n12150), .QN(n12340) );
  NOR2X0 U11985 ( .IN1(n12342), .IN2(n12343), .QN(n12341) );
  NOR2X0 U11986 ( .IN1(n10840), .IN2(n12344), .QN(n12343) );
  NOR2X0 U11987 ( .IN1(n12345), .IN2(n10839), .QN(n12342) );
  NAND2X0 U11988 ( .IN1(n12346), .IN2(n12347), .QN(g30648) );
  INVX0 U11989 ( .INP(n12348), .ZN(n12347) );
  NOR2X0 U11990 ( .IN1(g6518), .IN2(n9529), .QN(n12348) );
  NAND2X0 U11991 ( .IN1(n12297), .IN2(g6518), .QN(n12346) );
  NAND2X0 U11992 ( .IN1(n12349), .IN2(n12350), .QN(g30647) );
  NAND2X0 U11993 ( .IN1(g915), .IN2(n10321), .QN(n12350) );
  NAND2X0 U11994 ( .IN1(test_so31), .IN2(n12351), .QN(n12349) );
  NAND2X0 U11995 ( .IN1(n12352), .IN2(n12353), .QN(g30646) );
  NAND2X0 U11996 ( .IN1(n4512), .IN2(g243), .QN(n12353) );
  NAND2X0 U11997 ( .IN1(n12301), .IN2(g6313), .QN(n12352) );
  NAND2X0 U11998 ( .IN1(n12354), .IN2(n12355), .QN(g30645) );
  INVX0 U11999 ( .INP(n12356), .ZN(n12355) );
  NOR2X0 U12000 ( .IN1(g165), .IN2(n9470), .QN(n12356) );
  NAND2X0 U12001 ( .IN1(n12357), .IN2(g165), .QN(n12354) );
  NAND2X0 U12002 ( .IN1(n12358), .IN2(n12359), .QN(g30644) );
  INVX0 U12003 ( .INP(n12360), .ZN(n12359) );
  NOR2X0 U12004 ( .IN1(g6573), .IN2(n9420), .QN(n12360) );
  NAND2X0 U12005 ( .IN1(n12291), .IN2(g6573), .QN(n12358) );
  NAND2X0 U12006 ( .IN1(n12361), .IN2(n12101), .QN(n12291) );
  NAND2X0 U12007 ( .IN1(n12331), .IN2(n12362), .QN(n12101) );
  NOR2X0 U12008 ( .IN1(n12363), .IN2(n12364), .QN(n12361) );
  NOR2X0 U12009 ( .IN1(n12365), .IN2(n12104), .QN(n12364) );
  INVX0 U12010 ( .INP(n12131), .ZN(n12104) );
  NOR2X0 U12011 ( .IN1(n12105), .IN2(n12366), .QN(n12363) );
  NAND2X0 U12012 ( .IN1(n12367), .IN2(n12368), .QN(n12366) );
  NAND2X0 U12013 ( .IN1(n10901), .IN2(n2685), .QN(n12368) );
  INVX0 U12014 ( .INP(n12369), .ZN(n12367) );
  NOR2X0 U12015 ( .IN1(n10901), .IN2(n2685), .QN(n12369) );
  NAND2X0 U12016 ( .IN1(n12370), .IN2(n12371), .QN(n2685) );
  NAND2X0 U12017 ( .IN1(n12372), .IN2(n12373), .QN(n12371) );
  NAND2X0 U12018 ( .IN1(n10885), .IN2(n11777), .QN(n12373) );
  NAND2X0 U12019 ( .IN1(n4530), .IN2(n10884), .QN(n12372) );
  NAND2X0 U12020 ( .IN1(n12374), .IN2(n12375), .QN(g30643) );
  INVX0 U12021 ( .INP(n12376), .ZN(n12375) );
  NOR2X0 U12022 ( .IN1(g6368), .IN2(n9508), .QN(n12376) );
  NAND2X0 U12023 ( .IN1(n12297), .IN2(g6368), .QN(n12374) );
  INVX0 U12024 ( .INP(n12377), .ZN(n12297) );
  NAND2X0 U12025 ( .IN1(n12378), .IN2(n12379), .QN(n12377) );
  NAND2X0 U12026 ( .IN1(n12147), .IN2(n4375), .QN(n12379) );
  NOR2X0 U12027 ( .IN1(n12179), .IN2(n12380), .QN(n12378) );
  NOR2X0 U12028 ( .IN1(n12381), .IN2(n12150), .QN(n12380) );
  NOR2X0 U12029 ( .IN1(n12382), .IN2(n12383), .QN(n12381) );
  INVX0 U12030 ( .INP(n12384), .ZN(n12383) );
  NAND2X0 U12031 ( .IN1(n10835), .IN2(n12385), .QN(n12384) );
  NOR2X0 U12032 ( .IN1(n10835), .IN2(n12385), .QN(n12382) );
  NOR2X0 U12033 ( .IN1(n12386), .IN2(n12190), .QN(n12179) );
  NAND2X0 U12034 ( .IN1(n12387), .IN2(n12388), .QN(g30642) );
  INVX0 U12035 ( .INP(n12389), .ZN(n12388) );
  NOR2X0 U12036 ( .IN1(g6518), .IN2(n9533), .QN(n12389) );
  NAND2X0 U12037 ( .IN1(n12351), .IN2(g6518), .QN(n12387) );
  NAND2X0 U12038 ( .IN1(n12390), .IN2(n12391), .QN(g30641) );
  INVX0 U12039 ( .INP(n12392), .ZN(n12391) );
  NOR2X0 U12040 ( .IN1(g6231), .IN2(n9519), .QN(n12392) );
  NAND2X0 U12041 ( .IN1(n12301), .IN2(g6231), .QN(n12390) );
  INVX0 U12042 ( .INP(n12393), .ZN(n12301) );
  NAND2X0 U12043 ( .IN1(n12394), .IN2(n12395), .QN(n12393) );
  NAND2X0 U12044 ( .IN1(n12246), .IN2(n4392), .QN(n12395) );
  NOR2X0 U12045 ( .IN1(n12248), .IN2(n12396), .QN(n12394) );
  NOR2X0 U12046 ( .IN1(n12202), .IN2(n12397), .QN(n12396) );
  NAND2X0 U12047 ( .IN1(n12398), .IN2(n12399), .QN(n12397) );
  NAND2X0 U12048 ( .IN1(n12400), .IN2(n10784), .QN(n12399) );
  NAND2X0 U12049 ( .IN1(n12207), .IN2(n12401), .QN(n12400) );
  NAND2X0 U12050 ( .IN1(n12402), .IN2(n12403), .QN(n12401) );
  NAND2X0 U12051 ( .IN1(n10767), .IN2(n11773), .QN(n12403) );
  NAND2X0 U12052 ( .IN1(n11774), .IN2(n10766), .QN(n12402) );
  NAND2X0 U12053 ( .IN1(n12404), .IN2(n12405), .QN(n12398) );
  NOR2X0 U12054 ( .IN1(n12406), .IN2(n12407), .QN(n12404) );
  NOR2X0 U12055 ( .IN1(n10767), .IN2(n11774), .QN(n12406) );
  NAND2X0 U12056 ( .IN1(n12408), .IN2(n12409), .QN(g30640) );
  NAND2X0 U12057 ( .IN1(n4512), .IN2(g234), .QN(n12409) );
  NAND2X0 U12058 ( .IN1(n12357), .IN2(g6313), .QN(n12408) );
  NAND2X0 U12059 ( .IN1(n12410), .IN2(n12411), .QN(g30639) );
  INVX0 U12060 ( .INP(n12412), .ZN(n12411) );
  NOR2X0 U12061 ( .IN1(g165), .IN2(n9427), .QN(n12412) );
  NAND2X0 U12062 ( .IN1(n12413), .IN2(g165), .QN(n12410) );
  NAND2X0 U12063 ( .IN1(n12414), .IN2(n12415), .QN(g30638) );
  INVX0 U12064 ( .INP(n12416), .ZN(n12415) );
  NOR2X0 U12065 ( .IN1(g6368), .IN2(n9497), .QN(n12416) );
  NAND2X0 U12066 ( .IN1(n12351), .IN2(g6368), .QN(n12414) );
  NAND2X0 U12067 ( .IN1(n12417), .IN2(n12418), .QN(n12351) );
  NAND2X0 U12068 ( .IN1(n12147), .IN2(n12419), .QN(n12418) );
  NOR2X0 U12069 ( .IN1(n12148), .IN2(n12420), .QN(n12417) );
  NOR2X0 U12070 ( .IN1(n12150), .IN2(n12421), .QN(n12420) );
  NAND2X0 U12071 ( .IN1(n12422), .IN2(n12423), .QN(n12421) );
  NAND2X0 U12072 ( .IN1(n10865), .IN2(n12424), .QN(n12423) );
  NAND2X0 U12073 ( .IN1(n12186), .IN2(n10864), .QN(n12422) );
  INVX0 U12074 ( .INP(n12424), .ZN(n12186) );
  NAND2X0 U12075 ( .IN1(n12425), .IN2(n12426), .QN(n12424) );
  NOR2X0 U12076 ( .IN1(n12427), .IN2(n12428), .QN(n12425) );
  NOR2X0 U12077 ( .IN1(n10848), .IN2(n12190), .QN(n12428) );
  NOR2X0 U12078 ( .IN1(n12429), .IN2(n10815), .QN(n12427) );
  INVX0 U12079 ( .INP(n12430), .ZN(n12150) );
  NOR2X0 U12080 ( .IN1(n12386), .IN2(n12191), .QN(n12148) );
  INVX0 U12081 ( .INP(n12431), .ZN(n12386) );
  NAND2X0 U12082 ( .IN1(n12432), .IN2(n12433), .QN(g30637) );
  INVX0 U12083 ( .INP(n12434), .ZN(n12433) );
  NOR2X0 U12084 ( .IN1(g6231), .IN2(n9522), .QN(n12434) );
  NAND2X0 U12085 ( .IN1(n12357), .IN2(g6231), .QN(n12432) );
  INVX0 U12086 ( .INP(n12435), .ZN(n12357) );
  NAND2X0 U12087 ( .IN1(n12436), .IN2(n12437), .QN(n12435) );
  NAND2X0 U12088 ( .IN1(n12246), .IN2(n4376), .QN(n12437) );
  NOR2X0 U12089 ( .IN1(n12248), .IN2(n12438), .QN(n12436) );
  NOR2X0 U12090 ( .IN1(n12439), .IN2(n12202), .QN(n12438) );
  NOR2X0 U12091 ( .IN1(n12440), .IN2(n12441), .QN(n12439) );
  NOR2X0 U12092 ( .IN1(n12442), .IN2(n10754), .QN(n12441) );
  NOR2X0 U12093 ( .IN1(n10755), .IN2(n12443), .QN(n12440) );
  INVX0 U12094 ( .INP(n12444), .ZN(n12248) );
  NAND2X0 U12095 ( .IN1(n12445), .IN2(n11774), .QN(n12444) );
  NAND2X0 U12096 ( .IN1(n12446), .IN2(n12447), .QN(g30636) );
  NAND2X0 U12097 ( .IN1(n4512), .IN2(g225), .QN(n12447) );
  NAND2X0 U12098 ( .IN1(n12413), .IN2(g6313), .QN(n12446) );
  NAND2X0 U12099 ( .IN1(n12448), .IN2(n12449), .QN(g30635) );
  INVX0 U12100 ( .INP(n12450), .ZN(n12449) );
  NOR2X0 U12101 ( .IN1(g6231), .IN2(n9421), .QN(n12450) );
  NAND2X0 U12102 ( .IN1(n12413), .IN2(g6231), .QN(n12448) );
  NAND2X0 U12103 ( .IN1(n12451), .IN2(n12198), .QN(n12413) );
  NAND2X0 U12104 ( .IN1(n12445), .IN2(n11773), .QN(n12198) );
  NOR2X0 U12105 ( .IN1(n12452), .IN2(n12453), .QN(n12451) );
  NOR2X0 U12106 ( .IN1(n12454), .IN2(n12201), .QN(n12453) );
  INVX0 U12107 ( .INP(n12246), .ZN(n12201) );
  NOR2X0 U12108 ( .IN1(n12202), .IN2(n12455), .QN(n12452) );
  NAND2X0 U12109 ( .IN1(n12456), .IN2(n12457), .QN(n12455) );
  NAND2X0 U12110 ( .IN1(n10771), .IN2(n2718), .QN(n12457) );
  INVX0 U12111 ( .INP(n12458), .ZN(n12456) );
  NOR2X0 U12112 ( .IN1(n10771), .IN2(n2718), .QN(n12458) );
  NAND2X0 U12113 ( .IN1(n12459), .IN2(n12460), .QN(n2718) );
  NAND2X0 U12114 ( .IN1(n12461), .IN2(n12462), .QN(n12460) );
  NAND2X0 U12115 ( .IN1(n10759), .IN2(n11773), .QN(n12462) );
  NAND2X0 U12116 ( .IN1(n11774), .IN2(n10758), .QN(n12461) );
  INVX0 U12117 ( .INP(n12463), .ZN(n12202) );
  NAND2X0 U12118 ( .IN1(n12464), .IN2(n12465), .QN(g30566) );
  NAND2X0 U12119 ( .IN1(n11935), .IN2(n4606), .QN(n12465) );
  NOR2X0 U12120 ( .IN1(n12466), .IN2(n12467), .QN(n11935) );
  NAND2X0 U12121 ( .IN1(n12468), .IN2(n12469), .QN(n12466) );
  NAND2X0 U12122 ( .IN1(n12470), .IN2(n12471), .QN(n12469) );
  INVX0 U12123 ( .INP(n12472), .ZN(n12468) );
  NOR2X0 U12124 ( .IN1(n12470), .IN2(n12471), .QN(n12472) );
  NAND2X0 U12125 ( .IN1(n12473), .IN2(n12474), .QN(n12471) );
  NAND2X0 U12126 ( .IN1(n12475), .IN2(n12476), .QN(n12474) );
  NAND2X0 U12127 ( .IN1(n12477), .IN2(n12478), .QN(n12473) );
  NAND2X0 U12128 ( .IN1(n12479), .IN2(n12480), .QN(n12477) );
  NAND2X0 U12129 ( .IN1(n12481), .IN2(n12470), .QN(n12480) );
  NAND2X0 U12130 ( .IN1(n3038), .IN2(n12482), .QN(n12481) );
  INVX0 U12131 ( .INP(n12483), .ZN(n12482) );
  NOR2X0 U12132 ( .IN1(n12484), .IN2(n12485), .QN(n12483) );
  NOR2X0 U12133 ( .IN1(n12486), .IN2(n12487), .QN(n12485) );
  NAND2X0 U12134 ( .IN1(n12488), .IN2(n12489), .QN(n12486) );
  NAND2X0 U12135 ( .IN1(n12490), .IN2(n12491), .QN(n12479) );
  NAND2X0 U12136 ( .IN1(n12492), .IN2(n12493), .QN(n12490) );
  NAND2X0 U12137 ( .IN1(n12494), .IN2(n12487), .QN(n12493) );
  NOR2X0 U12138 ( .IN1(n12495), .IN2(n12496), .QN(n12494) );
  NAND2X0 U12139 ( .IN1(n12497), .IN2(n12498), .QN(n12492) );
  NOR2X0 U12140 ( .IN1(n12499), .IN2(n12500), .QN(n12497) );
  NAND2X0 U12141 ( .IN1(n12501), .IN2(n12488), .QN(n12500) );
  NAND2X0 U12142 ( .IN1(n12502), .IN2(n12496), .QN(n12501) );
  INVX0 U12143 ( .INP(n2792), .ZN(n12496) );
  INVX0 U12144 ( .INP(n12503), .ZN(n12499) );
  NAND2X0 U12145 ( .IN1(n4509), .IN2(g2392), .QN(n12464) );
  NAND2X0 U12146 ( .IN1(n12504), .IN2(n12505), .QN(g30505) );
  NAND2X0 U12147 ( .IN1(n12506), .IN2(g5555), .QN(n12505) );
  NAND2X0 U12148 ( .IN1(n4516), .IN2(g2393), .QN(n12504) );
  NAND2X0 U12149 ( .IN1(n12507), .IN2(n12508), .QN(g30503) );
  NAND2X0 U12150 ( .IN1(n12509), .IN2(g7014), .QN(n12508) );
  INVX0 U12151 ( .INP(n12510), .ZN(n12507) );
  NOR2X0 U12152 ( .IN1(n11946), .IN2(n9537), .QN(n12510) );
  NAND2X0 U12153 ( .IN1(n12511), .IN2(n12512), .QN(g30500) );
  NAND2X0 U12154 ( .IN1(n2798), .IN2(g1088), .QN(n12512) );
  NAND2X0 U12155 ( .IN1(test_so39), .IN2(n4381), .QN(n12511) );
  NAND2X0 U12156 ( .IN1(n12513), .IN2(n12514), .QN(g30487) );
  NAND2X0 U12157 ( .IN1(n12509), .IN2(g5511), .QN(n12514) );
  NAND2X0 U12158 ( .IN1(n4518), .IN2(g1699), .QN(n12513) );
  NAND2X0 U12159 ( .IN1(n12515), .IN2(n12516), .QN(g30485) );
  NAND2X0 U12160 ( .IN1(n4364), .IN2(g1006), .QN(n12516) );
  NAND2X0 U12161 ( .IN1(n2798), .IN2(g6712), .QN(n12515) );
  NAND2X0 U12162 ( .IN1(n12517), .IN2(n12518), .QN(g30482) );
  NAND2X0 U12163 ( .IN1(n12519), .IN2(n4640), .QN(n12518) );
  NAND2X0 U12164 ( .IN1(n4506), .IN2(g320), .QN(n12517) );
  NAND2X0 U12165 ( .IN1(n12520), .IN2(n12521), .QN(g30470) );
  NAND2X0 U12166 ( .IN1(n4363), .IN2(g1005), .QN(n12521) );
  NAND2X0 U12167 ( .IN1(n2798), .IN2(g5472), .QN(n12520) );
  NAND2X0 U12168 ( .IN1(n12522), .IN2(n12523), .QN(g30468) );
  NAND2X0 U12169 ( .IN1(n12519), .IN2(g6447), .QN(n12523) );
  NAND2X0 U12170 ( .IN1(n4499), .IN2(g319), .QN(n12522) );
  NAND2X0 U12171 ( .IN1(n12524), .IN2(n12525), .QN(g30455) );
  NAND2X0 U12172 ( .IN1(n12519), .IN2(g5437), .QN(n12525) );
  NOR2X0 U12173 ( .IN1(n12526), .IN2(n12003), .QN(n12519) );
  NOR2X0 U12174 ( .IN1(n12527), .IN2(n12528), .QN(n12526) );
  INVX0 U12175 ( .INP(n12529), .ZN(n12528) );
  NAND2X0 U12176 ( .IN1(n12530), .IN2(n12035), .QN(n12529) );
  NOR2X0 U12177 ( .IN1(n12530), .IN2(n12035), .QN(n12527) );
  NOR2X0 U12178 ( .IN1(n12531), .IN2(n12532), .QN(n12530) );
  NOR2X0 U12179 ( .IN1(n12025), .IN2(n12533), .QN(n12532) );
  NOR2X0 U12180 ( .IN1(n12534), .IN2(n12011), .QN(n12533) );
  NAND2X0 U12181 ( .IN1(n12535), .IN2(n12536), .QN(n12534) );
  NAND2X0 U12182 ( .IN1(n12028), .IN2(n12537), .QN(n12536) );
  NOR2X0 U12183 ( .IN1(n12538), .IN2(n4388), .QN(n12537) );
  NAND2X0 U12184 ( .IN1(n12006), .IN2(n12036), .QN(n12535) );
  NAND2X0 U12185 ( .IN1(n12539), .IN2(n12540), .QN(n12036) );
  NAND2X0 U12186 ( .IN1(n12024), .IN2(n3130), .QN(n12540) );
  INVX0 U12187 ( .INP(n12032), .ZN(n12539) );
  INVX0 U12188 ( .INP(n12541), .ZN(n12531) );
  NAND2X0 U12189 ( .IN1(n12542), .IN2(n12025), .QN(n12541) );
  NOR2X0 U12190 ( .IN1(n12543), .IN2(n12544), .QN(n12542) );
  NAND2X0 U12191 ( .IN1(n3130), .IN2(n12545), .QN(n12544) );
  NAND2X0 U12192 ( .IN1(n12014), .IN2(n12006), .QN(n12543) );
  INVX0 U12193 ( .INP(n12546), .ZN(n12524) );
  NOR2X0 U12194 ( .IN1(n12042), .IN2(n9562), .QN(n12546) );
  NAND2X0 U12195 ( .IN1(n12547), .IN2(n12548), .QN(g30356) );
  NAND2X0 U12196 ( .IN1(n12506), .IN2(n4606), .QN(n12548) );
  NAND2X0 U12197 ( .IN1(n4509), .IN2(g2395), .QN(n12547) );
  NAND2X0 U12198 ( .IN1(n12549), .IN2(n12550), .QN(g30341) );
  NAND2X0 U12199 ( .IN1(n12506), .IN2(g7264), .QN(n12550) );
  NOR2X0 U12200 ( .IN1(n12551), .IN2(n12467), .QN(n12506) );
  NOR2X0 U12201 ( .IN1(n12552), .IN2(n12553), .QN(n12551) );
  NOR2X0 U12202 ( .IN1(n12554), .IN2(n12487), .QN(n12553) );
  INVX0 U12203 ( .INP(n12555), .ZN(n12552) );
  NAND2X0 U12204 ( .IN1(n12554), .IN2(n12487), .QN(n12555) );
  NAND2X0 U12205 ( .IN1(n12556), .IN2(n12557), .QN(n12554) );
  NAND2X0 U12206 ( .IN1(n12498), .IN2(n12558), .QN(n12557) );
  NAND2X0 U12207 ( .IN1(n12559), .IN2(n12478), .QN(n12558) );
  NOR2X0 U12208 ( .IN1(n12560), .IN2(n12561), .QN(n12559) );
  NOR2X0 U12209 ( .IN1(n12470), .IN2(n12562), .QN(n12561) );
  INVX0 U12210 ( .INP(n12563), .ZN(n12562) );
  NOR2X0 U12211 ( .IN1(n12564), .IN2(n10322), .QN(n12563) );
  NOR2X0 U12212 ( .IN1(n12491), .IN2(n12503), .QN(n12560) );
  NOR2X0 U12213 ( .IN1(n12495), .IN2(n12565), .QN(n12503) );
  NOR2X0 U12214 ( .IN1(n12489), .IN2(n12566), .QN(n12565) );
  NAND2X0 U12215 ( .IN1(n12567), .IN2(n12487), .QN(n12556) );
  NOR2X0 U12216 ( .IN1(n12568), .IN2(n12569), .QN(n12567) );
  NAND2X0 U12217 ( .IN1(n12478), .IN2(n12470), .QN(n12568) );
  INVX0 U12218 ( .INP(n12570), .ZN(n12549) );
  NOR2X0 U12219 ( .IN1(n11937), .IN2(n9534), .QN(n12570) );
  NAND2X0 U12220 ( .IN1(n12571), .IN2(n12572), .QN(g30338) );
  NAND2X0 U12221 ( .IN1(n12509), .IN2(n4618), .QN(n12572) );
  NOR2X0 U12222 ( .IN1(n12573), .IN2(n11953), .QN(n12509) );
  NOR2X0 U12223 ( .IN1(n12574), .IN2(n12575), .QN(n12573) );
  INVX0 U12224 ( .INP(n12576), .ZN(n12575) );
  NAND2X0 U12225 ( .IN1(n12577), .IN2(n11985), .QN(n12576) );
  NOR2X0 U12226 ( .IN1(n12577), .IN2(n11985), .QN(n12574) );
  NOR2X0 U12227 ( .IN1(n12578), .IN2(n12579), .QN(n12577) );
  NOR2X0 U12228 ( .IN1(n11975), .IN2(n12580), .QN(n12579) );
  NOR2X0 U12229 ( .IN1(n12581), .IN2(n11961), .QN(n12580) );
  NAND2X0 U12230 ( .IN1(n12582), .IN2(n12583), .QN(n12581) );
  NAND2X0 U12231 ( .IN1(n11978), .IN2(n12584), .QN(n12583) );
  NOR2X0 U12232 ( .IN1(n12585), .IN2(n4386), .QN(n12584) );
  NAND2X0 U12233 ( .IN1(n11956), .IN2(n11986), .QN(n12582) );
  NAND2X0 U12234 ( .IN1(n12586), .IN2(n12587), .QN(n11986) );
  NAND2X0 U12235 ( .IN1(n11974), .IN2(n3070), .QN(n12587) );
  INVX0 U12236 ( .INP(n11982), .ZN(n12586) );
  INVX0 U12237 ( .INP(n12588), .ZN(n12578) );
  NAND2X0 U12238 ( .IN1(n12589), .IN2(n11975), .QN(n12588) );
  NOR2X0 U12239 ( .IN1(n12590), .IN2(n12591), .QN(n12589) );
  NAND2X0 U12240 ( .IN1(n3070), .IN2(n12592), .QN(n12591) );
  NAND2X0 U12241 ( .IN1(n11964), .IN2(n11956), .QN(n12590) );
  NAND2X0 U12242 ( .IN1(n4511), .IN2(g1701), .QN(n12571) );
  NAND2X0 U12243 ( .IN1(n12593), .IN2(n12594), .QN(g30304) );
  INVX0 U12244 ( .INP(n12595), .ZN(n12594) );
  NOR2X0 U12245 ( .IN1(g2241), .IN2(n9571), .QN(n12595) );
  NAND2X0 U12246 ( .IN1(n12596), .IN2(g2241), .QN(n12593) );
  NAND2X0 U12247 ( .IN1(n12597), .IN2(n12598), .QN(g30303) );
  NAND2X0 U12248 ( .IN1(g2282), .IN2(n10320), .QN(n12598) );
  NAND2X0 U12249 ( .IN1(test_so73), .IN2(n12596), .QN(n12597) );
  NAND2X0 U12250 ( .IN1(n12599), .IN2(n12600), .QN(g30302) );
  INVX0 U12251 ( .INP(n12601), .ZN(n12600) );
  NOR2X0 U12252 ( .IN1(g1547), .IN2(n9572), .QN(n12601) );
  NAND2X0 U12253 ( .IN1(n12602), .IN2(g1547), .QN(n12599) );
  NAND2X0 U12254 ( .IN1(n12603), .IN2(n12604), .QN(g30301) );
  INVX0 U12255 ( .INP(n12605), .ZN(n12604) );
  NOR2X0 U12256 ( .IN1(g6837), .IN2(n9477), .QN(n12605) );
  NAND2X0 U12257 ( .IN1(n12596), .IN2(g6837), .QN(n12603) );
  NAND2X0 U12258 ( .IN1(n12606), .IN2(n12607), .QN(n12596) );
  NAND2X0 U12259 ( .IN1(n12608), .IN2(n12609), .QN(n12607) );
  NOR2X0 U12260 ( .IN1(n12610), .IN2(n12611), .QN(n12608) );
  NOR2X0 U12261 ( .IN1(n10970), .IN2(n12612), .QN(n12611) );
  NOR2X0 U12262 ( .IN1(n12613), .IN2(n10969), .QN(n12610) );
  INVX0 U12263 ( .INP(n12612), .ZN(n12613) );
  NAND2X0 U12264 ( .IN1(n12064), .IN2(g2185), .QN(n12606) );
  NAND2X0 U12265 ( .IN1(n12614), .IN2(n12615), .QN(g30300) );
  INVX0 U12266 ( .INP(n12616), .ZN(n12615) );
  NOR2X0 U12267 ( .IN1(g2241), .IN2(n9578), .QN(n12616) );
  NAND2X0 U12268 ( .IN1(n12617), .IN2(g2241), .QN(n12614) );
  NAND2X0 U12269 ( .IN1(n12618), .IN2(n12619), .QN(g30299) );
  NAND2X0 U12270 ( .IN1(n4515), .IN2(g1588), .QN(n12619) );
  NAND2X0 U12271 ( .IN1(n12602), .IN2(g6782), .QN(n12618) );
  NAND2X0 U12272 ( .IN1(n12620), .IN2(n12621), .QN(g30298) );
  NAND2X0 U12273 ( .IN1(g897), .IN2(n10321), .QN(n12621) );
  NAND2X0 U12274 ( .IN1(test_so31), .IN2(n12622), .QN(n12620) );
  NAND2X0 U12275 ( .IN1(n12623), .IN2(n12624), .QN(g30297) );
  INVX0 U12276 ( .INP(n12625), .ZN(n12624) );
  NOR2X0 U12277 ( .IN1(g2241), .IN2(n9568), .QN(n12625) );
  NAND2X0 U12278 ( .IN1(n12626), .IN2(g2241), .QN(n12623) );
  NAND2X0 U12279 ( .IN1(n12627), .IN2(n12628), .QN(g30296) );
  NAND2X0 U12280 ( .IN1(test_so76), .IN2(n10320), .QN(n12628) );
  NAND2X0 U12281 ( .IN1(test_so73), .IN2(n12617), .QN(n12627) );
  NAND2X0 U12282 ( .IN1(n12629), .IN2(n12630), .QN(g30295) );
  INVX0 U12283 ( .INP(n12631), .ZN(n12630) );
  NOR2X0 U12284 ( .IN1(g6573), .IN2(n9490), .QN(n12631) );
  NAND2X0 U12285 ( .IN1(n12602), .IN2(g6573), .QN(n12629) );
  NAND2X0 U12286 ( .IN1(n12632), .IN2(n12633), .QN(n12602) );
  NAND2X0 U12287 ( .IN1(n12634), .IN2(n12635), .QN(n12633) );
  NOR2X0 U12288 ( .IN1(n12636), .IN2(n12637), .QN(n12634) );
  NOR2X0 U12289 ( .IN1(n10905), .IN2(n12638), .QN(n12637) );
  NOR2X0 U12290 ( .IN1(n12639), .IN2(n10904), .QN(n12636) );
  INVX0 U12291 ( .INP(n12638), .ZN(n12639) );
  NAND2X0 U12292 ( .IN1(n12131), .IN2(g1491), .QN(n12632) );
  NAND2X0 U12293 ( .IN1(n12640), .IN2(n12641), .QN(g30294) );
  INVX0 U12294 ( .INP(n12642), .ZN(n12641) );
  NOR2X0 U12295 ( .IN1(g1547), .IN2(n9581), .QN(n12642) );
  NAND2X0 U12296 ( .IN1(n12643), .IN2(g1547), .QN(n12640) );
  NAND2X0 U12297 ( .IN1(n12644), .IN2(n12645), .QN(g30293) );
  INVX0 U12298 ( .INP(n12646), .ZN(n12645) );
  NOR2X0 U12299 ( .IN1(g6518), .IN2(n9503), .QN(n12646) );
  NAND2X0 U12300 ( .IN1(n12622), .IN2(g6518), .QN(n12644) );
  NAND2X0 U12301 ( .IN1(n12647), .IN2(n12648), .QN(g30292) );
  INVX0 U12302 ( .INP(n12649), .ZN(n12648) );
  NOR2X0 U12303 ( .IN1(g165), .IN2(n9575), .QN(n12649) );
  NAND2X0 U12304 ( .IN1(n12650), .IN2(g165), .QN(n12647) );
  NAND2X0 U12305 ( .IN1(n12651), .IN2(n12652), .QN(g30291) );
  NAND2X0 U12306 ( .IN1(g2336), .IN2(n10320), .QN(n12652) );
  NAND2X0 U12307 ( .IN1(test_so73), .IN2(n12626), .QN(n12651) );
  NAND2X0 U12308 ( .IN1(n12653), .IN2(n12654), .QN(g30290) );
  INVX0 U12309 ( .INP(n12655), .ZN(n12654) );
  NOR2X0 U12310 ( .IN1(g2241), .IN2(n9459), .QN(n12655) );
  NAND2X0 U12311 ( .IN1(n12656), .IN2(g2241), .QN(n12653) );
  NAND2X0 U12312 ( .IN1(n12657), .IN2(n12658), .QN(g30289) );
  INVX0 U12313 ( .INP(n12659), .ZN(n12658) );
  NOR2X0 U12314 ( .IN1(g6837), .IN2(n9482), .QN(n12659) );
  NAND2X0 U12315 ( .IN1(n12617), .IN2(g6837), .QN(n12657) );
  NAND2X0 U12316 ( .IN1(n12660), .IN2(n12661), .QN(n12617) );
  NAND2X0 U12317 ( .IN1(n12609), .IN2(n12662), .QN(n12661) );
  NAND2X0 U12318 ( .IN1(n12663), .IN2(n12664), .QN(n12662) );
  NAND2X0 U12319 ( .IN1(n10954), .IN2(n12665), .QN(n12664) );
  NAND2X0 U12320 ( .IN1(n12666), .IN2(n10953), .QN(n12663) );
  INVX0 U12321 ( .INP(n12665), .ZN(n12666) );
  NAND2X0 U12322 ( .IN1(n12064), .IN2(g2165), .QN(n12660) );
  NAND2X0 U12323 ( .IN1(n12667), .IN2(n12668), .QN(g30288) );
  INVX0 U12324 ( .INP(n12669), .ZN(n12668) );
  NOR2X0 U12325 ( .IN1(g1547), .IN2(n9569), .QN(n12669) );
  NAND2X0 U12326 ( .IN1(n12670), .IN2(g1547), .QN(n12667) );
  NAND2X0 U12327 ( .IN1(n12671), .IN2(n12672), .QN(g30287) );
  NAND2X0 U12328 ( .IN1(n4515), .IN2(g1570), .QN(n12672) );
  NAND2X0 U12329 ( .IN1(n12643), .IN2(g6782), .QN(n12671) );
  NAND2X0 U12330 ( .IN1(n12673), .IN2(n12674), .QN(g30286) );
  INVX0 U12331 ( .INP(n12675), .ZN(n12674) );
  NOR2X0 U12332 ( .IN1(g6368), .IN2(n9504), .QN(n12675) );
  NAND2X0 U12333 ( .IN1(n12622), .IN2(g6368), .QN(n12673) );
  NAND2X0 U12334 ( .IN1(n12676), .IN2(n12677), .QN(n12622) );
  NAND2X0 U12335 ( .IN1(n12678), .IN2(n12430), .QN(n12677) );
  NOR2X0 U12336 ( .IN1(n12679), .IN2(n12680), .QN(n12678) );
  NOR2X0 U12337 ( .IN1(n10824), .IN2(n12681), .QN(n12680) );
  INVX0 U12338 ( .INP(n12682), .ZN(n12679) );
  NAND2X0 U12339 ( .IN1(n12681), .IN2(n10824), .QN(n12682) );
  NAND2X0 U12340 ( .IN1(n12147), .IN2(g801), .QN(n12676) );
  NAND2X0 U12341 ( .IN1(n12683), .IN2(n12684), .QN(g30285) );
  NAND2X0 U12342 ( .IN1(g879), .IN2(n10321), .QN(n12684) );
  NAND2X0 U12343 ( .IN1(test_so31), .IN2(n12685), .QN(n12683) );
  NAND2X0 U12344 ( .IN1(n12686), .IN2(n12687), .QN(g30284) );
  NAND2X0 U12345 ( .IN1(n4512), .IN2(g207), .QN(n12687) );
  NAND2X0 U12346 ( .IN1(n12650), .IN2(g6313), .QN(n12686) );
  NAND2X0 U12347 ( .IN1(n12688), .IN2(n12689), .QN(g30283) );
  INVX0 U12348 ( .INP(n12690), .ZN(n12689) );
  NOR2X0 U12349 ( .IN1(g6837), .IN2(n9472), .QN(n12690) );
  NAND2X0 U12350 ( .IN1(n12626), .IN2(g6837), .QN(n12688) );
  NAND2X0 U12351 ( .IN1(n12691), .IN2(n12692), .QN(n12626) );
  NAND2X0 U12352 ( .IN1(n12064), .IN2(g2200), .QN(n12692) );
  NAND2X0 U12353 ( .IN1(n12693), .IN2(n12694), .QN(n12691) );
  NOR2X0 U12354 ( .IN1(n12695), .IN2(n12696), .QN(n12694) );
  NOR2X0 U12355 ( .IN1(n10950), .IN2(n12697), .QN(n12696) );
  NOR2X0 U12356 ( .IN1(n12313), .IN2(n10949), .QN(n12695) );
  INVX0 U12357 ( .INP(n12697), .ZN(n12313) );
  NAND2X0 U12358 ( .IN1(n12698), .IN2(n12699), .QN(n12697) );
  NAND2X0 U12359 ( .IN1(n12700), .IN2(n12701), .QN(n12699) );
  NAND2X0 U12360 ( .IN1(n10946), .IN2(n11780), .QN(n12701) );
  NAND2X0 U12361 ( .IN1(n4529), .IN2(n10945), .QN(n12700) );
  NAND2X0 U12362 ( .IN1(n12702), .IN2(n12703), .QN(g30282) );
  NAND2X0 U12363 ( .IN1(test_so77), .IN2(n10320), .QN(n12703) );
  NAND2X0 U12364 ( .IN1(test_so73), .IN2(n12656), .QN(n12702) );
  NAND2X0 U12365 ( .IN1(n12704), .IN2(n12705), .QN(g30281) );
  NAND2X0 U12366 ( .IN1(n4515), .IN2(g1642), .QN(n12705) );
  NAND2X0 U12367 ( .IN1(n12670), .IN2(g6782), .QN(n12704) );
  NAND2X0 U12368 ( .IN1(n12706), .IN2(n12707), .QN(g30280) );
  INVX0 U12369 ( .INP(n12708), .ZN(n12707) );
  NOR2X0 U12370 ( .IN1(g1547), .IN2(n9462), .QN(n12708) );
  NAND2X0 U12371 ( .IN1(n12709), .IN2(g1547), .QN(n12706) );
  NAND2X0 U12372 ( .IN1(n12710), .IN2(n12711), .QN(g30279) );
  INVX0 U12373 ( .INP(n12712), .ZN(n12711) );
  NOR2X0 U12374 ( .IN1(g6573), .IN2(n9495), .QN(n12712) );
  NAND2X0 U12375 ( .IN1(n12643), .IN2(g6573), .QN(n12710) );
  NAND2X0 U12376 ( .IN1(n12713), .IN2(n12714), .QN(n12643) );
  NAND2X0 U12377 ( .IN1(n12635), .IN2(n12715), .QN(n12714) );
  NAND2X0 U12378 ( .IN1(n12716), .IN2(n12717), .QN(n12715) );
  NAND2X0 U12379 ( .IN1(n12718), .IN2(n10888), .QN(n12717) );
  NAND2X0 U12380 ( .IN1(n10889), .IN2(n12719), .QN(n12716) );
  NAND2X0 U12381 ( .IN1(n12131), .IN2(g1471), .QN(n12713) );
  NAND2X0 U12382 ( .IN1(n12720), .IN2(n12721), .QN(g30278) );
  NAND2X0 U12383 ( .IN1(g951), .IN2(n10321), .QN(n12721) );
  NAND2X0 U12384 ( .IN1(test_so31), .IN2(n12722), .QN(n12720) );
  NAND2X0 U12385 ( .IN1(n12723), .IN2(n12724), .QN(g30277) );
  INVX0 U12386 ( .INP(n12725), .ZN(n12724) );
  NOR2X0 U12387 ( .IN1(g6518), .IN2(n9509), .QN(n12725) );
  NAND2X0 U12388 ( .IN1(n12685), .IN2(g6518), .QN(n12723) );
  NAND2X0 U12389 ( .IN1(n12726), .IN2(n12727), .QN(g30276) );
  INVX0 U12390 ( .INP(n12728), .ZN(n12727) );
  NOR2X0 U12391 ( .IN1(g6231), .IN2(n9518), .QN(n12728) );
  NAND2X0 U12392 ( .IN1(n12650), .IN2(g6231), .QN(n12726) );
  NAND2X0 U12393 ( .IN1(n12729), .IN2(n12730), .QN(n12650) );
  NAND2X0 U12394 ( .IN1(n12731), .IN2(n12463), .QN(n12730) );
  NOR2X0 U12395 ( .IN1(n12732), .IN2(n12733), .QN(n12731) );
  NOR2X0 U12396 ( .IN1(n10775), .IN2(n12734), .QN(n12733) );
  NOR2X0 U12397 ( .IN1(n12735), .IN2(n10774), .QN(n12732) );
  INVX0 U12398 ( .INP(n12734), .ZN(n12735) );
  NAND2X0 U12399 ( .IN1(n12246), .IN2(g113), .QN(n12729) );
  NAND2X0 U12400 ( .IN1(n12736), .IN2(n12737), .QN(g30275) );
  INVX0 U12401 ( .INP(n12738), .ZN(n12737) );
  NOR2X0 U12402 ( .IN1(g165), .IN2(n9587), .QN(n12738) );
  NAND2X0 U12403 ( .IN1(n12739), .IN2(g165), .QN(n12736) );
  NAND2X0 U12404 ( .IN1(n12740), .IN2(n12741), .QN(g30274) );
  INVX0 U12405 ( .INP(n12742), .ZN(n12741) );
  NOR2X0 U12406 ( .IN1(g6837), .IN2(n9475), .QN(n12742) );
  NAND2X0 U12407 ( .IN1(n12656), .IN2(g6837), .QN(n12740) );
  NAND2X0 U12408 ( .IN1(n12743), .IN2(n12744), .QN(n12656) );
  NAND2X0 U12409 ( .IN1(n12064), .IN2(g2190), .QN(n12744) );
  NAND2X0 U12410 ( .IN1(n12693), .IN2(n12745), .QN(n12743) );
  NOR2X0 U12411 ( .IN1(n12746), .IN2(n12747), .QN(n12745) );
  NOR2X0 U12412 ( .IN1(n10995), .IN2(n12748), .QN(n12747) );
  INVX0 U12413 ( .INP(n12749), .ZN(n12746) );
  NAND2X0 U12414 ( .IN1(n12748), .IN2(n10995), .QN(n12749) );
  NAND2X0 U12415 ( .IN1(n12750), .IN2(n12751), .QN(n12748) );
  NAND2X0 U12416 ( .IN1(n11780), .IN2(n10969), .QN(n12751) );
  NOR2X0 U12417 ( .IN1(n12317), .IN2(n12067), .QN(n12693) );
  INVX0 U12418 ( .INP(n12609), .ZN(n12067) );
  NAND2X0 U12419 ( .IN1(n12752), .IN2(n12753), .QN(g30273) );
  INVX0 U12420 ( .INP(n12754), .ZN(n12753) );
  NOR2X0 U12421 ( .IN1(g6573), .IN2(n9484), .QN(n12754) );
  NAND2X0 U12422 ( .IN1(n12670), .IN2(g6573), .QN(n12752) );
  NAND2X0 U12423 ( .IN1(n12755), .IN2(n12756), .QN(n12670) );
  NAND2X0 U12424 ( .IN1(n12757), .IN2(n12758), .QN(n12756) );
  NOR2X0 U12425 ( .IN1(n12759), .IN2(n12760), .QN(n12758) );
  NOR2X0 U12426 ( .IN1(n10885), .IN2(n12761), .QN(n12760) );
  NOR2X0 U12427 ( .IN1(n12370), .IN2(n10884), .QN(n12759) );
  INVX0 U12428 ( .INP(n12761), .ZN(n12370) );
  NAND2X0 U12429 ( .IN1(n12762), .IN2(n12763), .QN(n12761) );
  NAND2X0 U12430 ( .IN1(n12764), .IN2(n12765), .QN(n12763) );
  NAND2X0 U12431 ( .IN1(n10881), .IN2(n11777), .QN(n12765) );
  NAND2X0 U12432 ( .IN1(n4530), .IN2(n10880), .QN(n12764) );
  NAND2X0 U12433 ( .IN1(n12131), .IN2(g1506), .QN(n12755) );
  NAND2X0 U12434 ( .IN1(n12766), .IN2(n12767), .QN(g30272) );
  NAND2X0 U12435 ( .IN1(n4515), .IN2(g1633), .QN(n12767) );
  NAND2X0 U12436 ( .IN1(n12709), .IN2(g6782), .QN(n12766) );
  NAND2X0 U12437 ( .IN1(n12768), .IN2(n12769), .QN(g30271) );
  INVX0 U12438 ( .INP(n12770), .ZN(n12769) );
  NOR2X0 U12439 ( .IN1(g6518), .IN2(n9498), .QN(n12770) );
  NAND2X0 U12440 ( .IN1(n12722), .IN2(g6518), .QN(n12768) );
  NAND2X0 U12441 ( .IN1(n12771), .IN2(n12772), .QN(g30270) );
  NAND2X0 U12442 ( .IN1(g942), .IN2(n10321), .QN(n12772) );
  NAND2X0 U12443 ( .IN1(test_so31), .IN2(n12773), .QN(n12771) );
  NAND2X0 U12444 ( .IN1(n12774), .IN2(n12775), .QN(g30269) );
  INVX0 U12445 ( .INP(n12776), .ZN(n12775) );
  NOR2X0 U12446 ( .IN1(g6368), .IN2(n9510), .QN(n12776) );
  NAND2X0 U12447 ( .IN1(n12685), .IN2(g6368), .QN(n12774) );
  NAND2X0 U12448 ( .IN1(n12777), .IN2(n12778), .QN(n12685) );
  NAND2X0 U12449 ( .IN1(n12430), .IN2(n12779), .QN(n12778) );
  NAND2X0 U12450 ( .IN1(n12780), .IN2(n12781), .QN(n12779) );
  NAND2X0 U12451 ( .IN1(n10832), .IN2(n12782), .QN(n12781) );
  INVX0 U12452 ( .INP(n12783), .ZN(n12780) );
  NOR2X0 U12453 ( .IN1(n12782), .IN2(n10832), .QN(n12783) );
  NAND2X0 U12454 ( .IN1(n12147), .IN2(g785), .QN(n12777) );
  NAND2X0 U12455 ( .IN1(n12784), .IN2(n12785), .QN(g30268) );
  INVX0 U12456 ( .INP(n12786), .ZN(n12785) );
  NOR2X0 U12457 ( .IN1(g165), .IN2(n9570), .QN(n12786) );
  NAND2X0 U12458 ( .IN1(n12787), .IN2(g165), .QN(n12784) );
  NAND2X0 U12459 ( .IN1(n12788), .IN2(n12789), .QN(g30267) );
  NAND2X0 U12460 ( .IN1(test_so13), .IN2(n4512), .QN(n12789) );
  NAND2X0 U12461 ( .IN1(n12739), .IN2(g6313), .QN(n12788) );
  NAND2X0 U12462 ( .IN1(n12790), .IN2(n12791), .QN(g30266) );
  INVX0 U12463 ( .INP(n12792), .ZN(n12791) );
  NOR2X0 U12464 ( .IN1(g6573), .IN2(n9488), .QN(n12792) );
  NAND2X0 U12465 ( .IN1(n12709), .IN2(g6573), .QN(n12790) );
  NAND2X0 U12466 ( .IN1(n12793), .IN2(n12794), .QN(n12709) );
  NAND2X0 U12467 ( .IN1(n12757), .IN2(n12795), .QN(n12794) );
  NOR2X0 U12468 ( .IN1(n12796), .IN2(n12797), .QN(n12795) );
  NOR2X0 U12469 ( .IN1(n10926), .IN2(n12798), .QN(n12797) );
  INVX0 U12470 ( .INP(n12799), .ZN(n12796) );
  NAND2X0 U12471 ( .IN1(n12798), .IN2(n10926), .QN(n12799) );
  NAND2X0 U12472 ( .IN1(n12800), .IN2(n12801), .QN(n12798) );
  NAND2X0 U12473 ( .IN1(n11777), .IN2(n10904), .QN(n12801) );
  NOR2X0 U12474 ( .IN1(n12331), .IN2(n12105), .QN(n12757) );
  INVX0 U12475 ( .INP(n12635), .ZN(n12105) );
  NAND2X0 U12476 ( .IN1(n12131), .IN2(g1496), .QN(n12793) );
  NAND2X0 U12477 ( .IN1(n12802), .IN2(n12803), .QN(g30265) );
  NAND2X0 U12478 ( .IN1(test_so35), .IN2(n4323), .QN(n12803) );
  NAND2X0 U12479 ( .IN1(n12722), .IN2(g6368), .QN(n12802) );
  NAND2X0 U12480 ( .IN1(n12804), .IN2(n12805), .QN(n12722) );
  NAND2X0 U12481 ( .IN1(n12806), .IN2(n12430), .QN(n12805) );
  NOR2X0 U12482 ( .IN1(n12807), .IN2(n12808), .QN(n12806) );
  NOR2X0 U12483 ( .IN1(n12429), .IN2(n12809), .QN(n12808) );
  INVX0 U12484 ( .INP(n12810), .ZN(n12807) );
  NAND2X0 U12485 ( .IN1(n12809), .IN2(n12429), .QN(n12810) );
  NAND2X0 U12486 ( .IN1(n12426), .IN2(n12811), .QN(n12809) );
  NAND2X0 U12487 ( .IN1(n12191), .IN2(n10816), .QN(n12811) );
  NOR2X0 U12488 ( .IN1(n12812), .IN2(n12813), .QN(n12426) );
  NOR2X0 U12489 ( .IN1(n12191), .IN2(n10816), .QN(n12813) );
  NAND2X0 U12490 ( .IN1(n12147), .IN2(g813), .QN(n12804) );
  NAND2X0 U12491 ( .IN1(n12814), .IN2(n12815), .QN(g30264) );
  INVX0 U12492 ( .INP(n12816), .ZN(n12815) );
  NOR2X0 U12493 ( .IN1(g6518), .IN2(n9501), .QN(n12816) );
  NAND2X0 U12494 ( .IN1(n12773), .IN2(g6518), .QN(n12814) );
  NAND2X0 U12495 ( .IN1(n12817), .IN2(n12818), .QN(g30263) );
  NAND2X0 U12496 ( .IN1(n4512), .IN2(g261), .QN(n12818) );
  NAND2X0 U12497 ( .IN1(n12787), .IN2(g6313), .QN(n12817) );
  NAND2X0 U12498 ( .IN1(n12819), .IN2(n12820), .QN(g30262) );
  NAND2X0 U12499 ( .IN1(n4369), .IN2(test_so14), .QN(n12820) );
  NAND2X0 U12500 ( .IN1(n12821), .IN2(g165), .QN(n12819) );
  NAND2X0 U12501 ( .IN1(n12822), .IN2(n12823), .QN(g30261) );
  INVX0 U12502 ( .INP(n12824), .ZN(n12823) );
  NOR2X0 U12503 ( .IN1(g6231), .IN2(n9523), .QN(n12824) );
  NAND2X0 U12504 ( .IN1(n12739), .IN2(g6231), .QN(n12822) );
  NAND2X0 U12505 ( .IN1(n12825), .IN2(n12826), .QN(n12739) );
  NAND2X0 U12506 ( .IN1(n12463), .IN2(n12827), .QN(n12826) );
  NAND2X0 U12507 ( .IN1(n12828), .IN2(n12829), .QN(n12827) );
  NAND2X0 U12508 ( .IN1(n12830), .IN2(n10796), .QN(n12829) );
  NAND2X0 U12509 ( .IN1(n4513), .IN2(n12831), .QN(n12828) );
  NAND2X0 U12510 ( .IN1(n12246), .IN2(g97), .QN(n12825) );
  NAND2X0 U12511 ( .IN1(n12832), .IN2(n12833), .QN(g30260) );
  INVX0 U12512 ( .INP(n12834), .ZN(n12833) );
  NOR2X0 U12513 ( .IN1(g2241), .IN2(n9576), .QN(n12834) );
  NAND2X0 U12514 ( .IN1(n12835), .IN2(g2241), .QN(n12832) );
  NAND2X0 U12515 ( .IN1(n12836), .IN2(n12837), .QN(g30259) );
  INVX0 U12516 ( .INP(n12838), .ZN(n12837) );
  NOR2X0 U12517 ( .IN1(g6368), .IN2(n9502), .QN(n12838) );
  NAND2X0 U12518 ( .IN1(n12773), .IN2(g6368), .QN(n12836) );
  NAND2X0 U12519 ( .IN1(n12839), .IN2(n12840), .QN(n12773) );
  NAND2X0 U12520 ( .IN1(n12841), .IN2(n12430), .QN(n12840) );
  NOR2X0 U12521 ( .IN1(n12842), .IN2(n12843), .QN(n12841) );
  NOR2X0 U12522 ( .IN1(n10820), .IN2(n12844), .QN(n12843) );
  INVX0 U12523 ( .INP(n12845), .ZN(n12842) );
  NAND2X0 U12524 ( .IN1(n12844), .IN2(n10820), .QN(n12845) );
  NAND2X0 U12525 ( .IN1(n12846), .IN2(n12847), .QN(n12844) );
  NAND2X0 U12526 ( .IN1(n12190), .IN2(n10823), .QN(n12847) );
  NAND2X0 U12527 ( .IN1(n12147), .IN2(g805), .QN(n12839) );
  NAND2X0 U12528 ( .IN1(n12848), .IN2(n12849), .QN(g30258) );
  INVX0 U12529 ( .INP(n12850), .ZN(n12849) );
  NOR2X0 U12530 ( .IN1(g6231), .IN2(n9512), .QN(n12850) );
  NAND2X0 U12531 ( .IN1(n12787), .IN2(g6231), .QN(n12848) );
  NAND2X0 U12532 ( .IN1(n12851), .IN2(n12852), .QN(n12787) );
  NAND2X0 U12533 ( .IN1(n12853), .IN2(n12463), .QN(n12852) );
  NOR2X0 U12534 ( .IN1(n12854), .IN2(n12855), .QN(n12853) );
  NOR2X0 U12535 ( .IN1(n10759), .IN2(n12856), .QN(n12855) );
  NOR2X0 U12536 ( .IN1(n12459), .IN2(n10758), .QN(n12854) );
  INVX0 U12537 ( .INP(n12856), .ZN(n12459) );
  NAND2X0 U12538 ( .IN1(n12857), .IN2(n12858), .QN(n12856) );
  NAND2X0 U12539 ( .IN1(n12859), .IN2(n12860), .QN(n12858) );
  NAND2X0 U12540 ( .IN1(n10751), .IN2(n11773), .QN(n12860) );
  NAND2X0 U12541 ( .IN1(n11774), .IN2(n10750), .QN(n12859) );
  NAND2X0 U12542 ( .IN1(n12246), .IN2(g125), .QN(n12851) );
  NAND2X0 U12543 ( .IN1(n12861), .IN2(n12862), .QN(g30257) );
  NAND2X0 U12544 ( .IN1(n4512), .IN2(g252), .QN(n12862) );
  NAND2X0 U12545 ( .IN1(n12821), .IN2(g6313), .QN(n12861) );
  NAND2X0 U12546 ( .IN1(n12863), .IN2(n12864), .QN(g30256) );
  NAND2X0 U12547 ( .IN1(g2291), .IN2(n10320), .QN(n12864) );
  NAND2X0 U12548 ( .IN1(test_so73), .IN2(n12835), .QN(n12863) );
  NAND2X0 U12549 ( .IN1(n12865), .IN2(n12866), .QN(g30255) );
  INVX0 U12550 ( .INP(n12867), .ZN(n12866) );
  NOR2X0 U12551 ( .IN1(g1547), .IN2(n9579), .QN(n12867) );
  NAND2X0 U12552 ( .IN1(n12868), .IN2(g1547), .QN(n12865) );
  NAND2X0 U12553 ( .IN1(n12869), .IN2(n12870), .QN(g30254) );
  INVX0 U12554 ( .INP(n12871), .ZN(n12870) );
  NOR2X0 U12555 ( .IN1(g6231), .IN2(n9516), .QN(n12871) );
  NAND2X0 U12556 ( .IN1(n12821), .IN2(g6231), .QN(n12869) );
  NAND2X0 U12557 ( .IN1(n12872), .IN2(n12873), .QN(n12821) );
  NAND2X0 U12558 ( .IN1(n12874), .IN2(n12463), .QN(n12873) );
  NOR2X0 U12559 ( .IN1(n12875), .IN2(n12876), .QN(n12874) );
  NOR2X0 U12560 ( .IN1(n10800), .IN2(n12877), .QN(n12876) );
  INVX0 U12561 ( .INP(n12878), .ZN(n12875) );
  NAND2X0 U12562 ( .IN1(n12877), .IN2(n10800), .QN(n12878) );
  NAND2X0 U12563 ( .IN1(n12879), .IN2(n12880), .QN(n12877) );
  NAND2X0 U12564 ( .IN1(n11773), .IN2(n10774), .QN(n12880) );
  NAND2X0 U12565 ( .IN1(n12246), .IN2(g117), .QN(n12872) );
  NAND2X0 U12566 ( .IN1(n12881), .IN2(n12882), .QN(g30253) );
  INVX0 U12567 ( .INP(n12883), .ZN(n12882) );
  NOR2X0 U12568 ( .IN1(g6837), .IN2(n9474), .QN(n12883) );
  NAND2X0 U12569 ( .IN1(n12835), .IN2(g6837), .QN(n12881) );
  NAND2X0 U12570 ( .IN1(n12884), .IN2(n12885), .QN(n12835) );
  NAND2X0 U12571 ( .IN1(n12886), .IN2(n12609), .QN(n12885) );
  NOR2X0 U12572 ( .IN1(n12887), .IN2(n12888), .QN(n12886) );
  NOR2X0 U12573 ( .IN1(n10946), .IN2(n12889), .QN(n12888) );
  NOR2X0 U12574 ( .IN1(n12698), .IN2(n10945), .QN(n12887) );
  INVX0 U12575 ( .INP(n12889), .ZN(n12698) );
  NAND2X0 U12576 ( .IN1(n12890), .IN2(n12750), .QN(n12889) );
  NOR2X0 U12577 ( .IN1(n12612), .IN2(n12891), .QN(n12750) );
  NOR2X0 U12578 ( .IN1(n11780), .IN2(n10969), .QN(n12891) );
  NAND2X0 U12579 ( .IN1(n12892), .IN2(n12893), .QN(n12612) );
  INVX0 U12580 ( .INP(n12224), .ZN(n12893) );
  NAND2X0 U12581 ( .IN1(n12072), .IN2(n12894), .QN(n12224) );
  NAND2X0 U12582 ( .IN1(n4529), .IN2(n10962), .QN(n12894) );
  INVX0 U12583 ( .INP(n12071), .ZN(n12072) );
  NAND2X0 U12584 ( .IN1(n12264), .IN2(n12895), .QN(n12071) );
  NAND2X0 U12585 ( .IN1(n12896), .IN2(n12897), .QN(n12895) );
  NAND2X0 U12586 ( .IN1(n12265), .IN2(n11780), .QN(n12897) );
  NAND2X0 U12587 ( .IN1(n4529), .IN2(n10978), .QN(n12896) );
  INVX0 U12588 ( .INP(n12266), .ZN(n12264) );
  NAND2X0 U12589 ( .IN1(n12898), .IN2(n12665), .QN(n12266) );
  NAND2X0 U12590 ( .IN1(n12899), .IN2(n12900), .QN(n12898) );
  NAND2X0 U12591 ( .IN1(n10954), .IN2(n11780), .QN(n12900) );
  NAND2X0 U12592 ( .IN1(n4529), .IN2(n10953), .QN(n12899) );
  NOR2X0 U12593 ( .IN1(n12901), .IN2(n12902), .QN(n12892) );
  NOR2X0 U12594 ( .IN1(n10991), .IN2(n4529), .QN(n12902) );
  NOR2X0 U12595 ( .IN1(n10962), .IN2(n10990), .QN(n12901) );
  NOR2X0 U12596 ( .IN1(n12903), .IN2(n12904), .QN(n12890) );
  NOR2X0 U12597 ( .IN1(n10995), .IN2(n4529), .QN(n12904) );
  NOR2X0 U12598 ( .IN1(n10970), .IN2(n10994), .QN(n12903) );
  NAND2X0 U12599 ( .IN1(n12064), .IN2(g2195), .QN(n12884) );
  NOR2X0 U12600 ( .IN1(n12609), .IN2(n12317), .QN(n12064) );
  NOR2X0 U12601 ( .IN1(n12905), .IN2(n12906), .QN(n12317) );
  NOR2X0 U12602 ( .IN1(n12905), .IN2(n12907), .QN(n12609) );
  NOR2X0 U12603 ( .IN1(n12906), .IN2(n12908), .QN(n12907) );
  INVX0 U12604 ( .INP(n12909), .ZN(n12908) );
  NAND2X0 U12605 ( .IN1(n4529), .IN2(n12910), .QN(n12909) );
  NAND2X0 U12606 ( .IN1(n12665), .IN2(n12911), .QN(n12906) );
  NAND2X0 U12607 ( .IN1(n12910), .IN2(n10933), .QN(n12911) );
  NAND2X0 U12608 ( .IN1(n12912), .IN2(n12913), .QN(n10933) );
  NOR2X0 U12609 ( .IN1(n10990), .IN2(n12914), .QN(n12913) );
  NAND2X0 U12610 ( .IN1(n10987), .IN2(n12265), .QN(n12914) );
  NOR2X0 U12611 ( .IN1(n12915), .IN2(n12916), .QN(n12912) );
  NAND2X0 U12612 ( .IN1(n10966), .IN2(n10962), .QN(n12916) );
  NAND2X0 U12613 ( .IN1(n12917), .IN2(n12918), .QN(n12910) );
  NOR2X0 U12614 ( .IN1(n12919), .IN2(n12920), .QN(n12918) );
  NAND2X0 U12615 ( .IN1(n10986), .IN2(n10978), .QN(n12920) );
  NAND2X0 U12616 ( .IN1(n10965), .IN2(n10961), .QN(n12919) );
  INVX0 U12617 ( .INP(n12921), .ZN(n12917) );
  NAND2X0 U12618 ( .IN1(n4529), .IN2(n12922), .QN(n12921) );
  NOR2X0 U12619 ( .IN1(n12915), .IN2(n10991), .QN(n12922) );
  NAND2X0 U12620 ( .IN1(n12923), .IN2(n12924), .QN(n12915) );
  NOR2X0 U12621 ( .IN1(n10949), .IN2(n12925), .QN(n12924) );
  NAND2X0 U12622 ( .IN1(n10946), .IN2(n10995), .QN(n12925) );
  NOR2X0 U12623 ( .IN1(n10953), .IN2(n10969), .QN(n12923) );
  NAND2X0 U12624 ( .IN1(n10934), .IN2(n11780), .QN(n12665) );
  INVX0 U12625 ( .INP(n12926), .ZN(n10934) );
  NAND2X0 U12626 ( .IN1(n12927), .IN2(n12928), .QN(n12905) );
  NAND2X0 U12627 ( .IN1(n12495), .IN2(n12478), .QN(n12928) );
  NOR2X0 U12628 ( .IN1(n12467), .IN2(n12929), .QN(n12927) );
  NOR2X0 U12629 ( .IN1(n2792), .IN2(n12930), .QN(n12929) );
  NOR2X0 U12630 ( .IN1(n12931), .IN2(n12932), .QN(n12930) );
  NOR2X0 U12631 ( .IN1(n12564), .IN2(n12933), .QN(n12931) );
  NAND2X0 U12632 ( .IN1(n12491), .IN2(n12478), .QN(n12933) );
  NAND2X0 U12633 ( .IN1(n12934), .IN2(n12935), .QN(n2792) );
  NAND2X0 U12634 ( .IN1(n12936), .IN2(n12937), .QN(n12935) );
  NAND2X0 U12635 ( .IN1(n9588), .IN2(n11937), .QN(n12937) );
  NOR2X0 U12636 ( .IN1(n12938), .IN2(n12939), .QN(n12936) );
  NOR2X0 U12637 ( .IN1(n4516), .IN2(g2397), .QN(n12939) );
  NOR2X0 U12638 ( .IN1(n4509), .IN2(g2396), .QN(n12938) );
  NAND2X0 U12639 ( .IN1(n12940), .IN2(n12941), .QN(g30252) );
  NAND2X0 U12640 ( .IN1(n4515), .IN2(g1597), .QN(n12941) );
  NAND2X0 U12641 ( .IN1(n12868), .IN2(g6782), .QN(n12940) );
  NAND2X0 U12642 ( .IN1(n12942), .IN2(n12943), .QN(g30251) );
  NAND2X0 U12643 ( .IN1(g906), .IN2(n10321), .QN(n12943) );
  NAND2X0 U12644 ( .IN1(test_so31), .IN2(n12944), .QN(n12942) );
  NAND2X0 U12645 ( .IN1(n12945), .IN2(n12946), .QN(g30250) );
  INVX0 U12646 ( .INP(n12947), .ZN(n12946) );
  NOR2X0 U12647 ( .IN1(g6573), .IN2(n9486), .QN(n12947) );
  NAND2X0 U12648 ( .IN1(n12868), .IN2(g6573), .QN(n12945) );
  NAND2X0 U12649 ( .IN1(n12948), .IN2(n12949), .QN(n12868) );
  NAND2X0 U12650 ( .IN1(n12950), .IN2(n12635), .QN(n12949) );
  NOR2X0 U12651 ( .IN1(n12951), .IN2(n12952), .QN(n12950) );
  NOR2X0 U12652 ( .IN1(n10881), .IN2(n12953), .QN(n12952) );
  NOR2X0 U12653 ( .IN1(n12762), .IN2(n10880), .QN(n12951) );
  INVX0 U12654 ( .INP(n12953), .ZN(n12762) );
  NAND2X0 U12655 ( .IN1(n12954), .IN2(n12800), .QN(n12953) );
  NOR2X0 U12656 ( .IN1(n12638), .IN2(n12955), .QN(n12800) );
  NOR2X0 U12657 ( .IN1(n11777), .IN2(n10904), .QN(n12955) );
  NAND2X0 U12658 ( .IN1(n12956), .IN2(n12957), .QN(n12638) );
  INVX0 U12659 ( .INP(n12285), .ZN(n12957) );
  NAND2X0 U12660 ( .IN1(n12110), .IN2(n12958), .QN(n12285) );
  NAND2X0 U12661 ( .IN1(n4530), .IN2(n10897), .QN(n12958) );
  INVX0 U12662 ( .INP(n12109), .ZN(n12110) );
  NAND2X0 U12663 ( .IN1(n12328), .IN2(n12959), .QN(n12109) );
  NAND2X0 U12664 ( .IN1(n12960), .IN2(n12961), .QN(n12959) );
  NAND2X0 U12665 ( .IN1(n10922), .IN2(n11777), .QN(n12961) );
  NAND2X0 U12666 ( .IN1(n4530), .IN2(n10921), .QN(n12960) );
  INVX0 U12667 ( .INP(n12329), .ZN(n12328) );
  NAND2X0 U12668 ( .IN1(n12962), .IN2(n12719), .QN(n12329) );
  NAND2X0 U12669 ( .IN1(n12963), .IN2(n12964), .QN(n12962) );
  NAND2X0 U12670 ( .IN1(n10889), .IN2(n11777), .QN(n12964) );
  NAND2X0 U12671 ( .IN1(n4530), .IN2(n10888), .QN(n12963) );
  NOR2X0 U12672 ( .IN1(n12965), .IN2(n12966), .QN(n12956) );
  NOR2X0 U12673 ( .IN1(n10914), .IN2(n4530), .QN(n12966) );
  NOR2X0 U12674 ( .IN1(n10897), .IN2(n10913), .QN(n12965) );
  NOR2X0 U12675 ( .IN1(n12967), .IN2(n12968), .QN(n12954) );
  NOR2X0 U12676 ( .IN1(n10926), .IN2(n4530), .QN(n12968) );
  NOR2X0 U12677 ( .IN1(n10905), .IN2(n10925), .QN(n12967) );
  NAND2X0 U12678 ( .IN1(n12131), .IN2(g1501), .QN(n12948) );
  NOR2X0 U12679 ( .IN1(n12635), .IN2(n12331), .QN(n12131) );
  NOR2X0 U12680 ( .IN1(n12969), .IN2(n12970), .QN(n12331) );
  NAND2X0 U12681 ( .IN1(n12719), .IN2(n12971), .QN(n12969) );
  NAND2X0 U12682 ( .IN1(n10868), .IN2(n12972), .QN(n12971) );
  NOR2X0 U12683 ( .IN1(n12970), .IN2(n12973), .QN(n12635) );
  NOR2X0 U12684 ( .IN1(n12974), .IN2(n12718), .QN(n12973) );
  INVX0 U12685 ( .INP(n12719), .ZN(n12718) );
  NAND2X0 U12686 ( .IN1(n11777), .IN2(n10869), .QN(n12719) );
  INVX0 U12687 ( .INP(n12975), .ZN(n10869) );
  INVX0 U12688 ( .INP(n12976), .ZN(n12974) );
  NAND2X0 U12689 ( .IN1(n12972), .IN2(n12977), .QN(n12976) );
  NAND2X0 U12690 ( .IN1(n12978), .IN2(n12362), .QN(n12977) );
  INVX0 U12691 ( .INP(n10868), .ZN(n12978) );
  NAND2X0 U12692 ( .IN1(n12979), .IN2(n12980), .QN(n10868) );
  NOR2X0 U12693 ( .IN1(n10929), .IN2(n12981), .QN(n12980) );
  NAND2X0 U12694 ( .IN1(n10922), .IN2(n10914), .QN(n12981) );
  NOR2X0 U12695 ( .IN1(n12982), .IN2(n12983), .QN(n12979) );
  NAND2X0 U12696 ( .IN1(n10901), .IN2(n10897), .QN(n12983) );
  NAND2X0 U12697 ( .IN1(n12984), .IN2(n12985), .QN(n12972) );
  NOR2X0 U12698 ( .IN1(n12986), .IN2(n12987), .QN(n12985) );
  NAND2X0 U12699 ( .IN1(n10929), .IN2(n10921), .QN(n12987) );
  NAND2X0 U12700 ( .IN1(n10900), .IN2(n10896), .QN(n12986) );
  NOR2X0 U12701 ( .IN1(n12362), .IN2(n12988), .QN(n12984) );
  INVX0 U12702 ( .INP(n12989), .ZN(n12988) );
  NOR2X0 U12703 ( .IN1(n12982), .IN2(n10914), .QN(n12989) );
  NAND2X0 U12704 ( .IN1(n12990), .IN2(n12991), .QN(n12982) );
  NOR2X0 U12705 ( .IN1(n10884), .IN2(n12992), .QN(n12991) );
  NAND2X0 U12706 ( .IN1(n10881), .IN2(n10926), .QN(n12992) );
  NOR2X0 U12707 ( .IN1(n10888), .IN2(n10904), .QN(n12990) );
  INVX0 U12708 ( .INP(n4530), .ZN(n12362) );
  NAND2X0 U12709 ( .IN1(n12993), .IN2(n12994), .QN(n12970) );
  NAND2X0 U12710 ( .IN1(n12995), .IN2(n12996), .QN(n12994) );
  NOR2X0 U12711 ( .IN1(n11953), .IN2(n12997), .QN(n12993) );
  NOR2X0 U12712 ( .IN1(n11961), .IN2(n12998), .QN(n12997) );
  NOR2X0 U12713 ( .IN1(n12999), .IN2(n11982), .QN(n12998) );
  NOR2X0 U12714 ( .IN1(n12585), .IN2(n13000), .QN(n12999) );
  NAND2X0 U12715 ( .IN1(n11983), .IN2(n11978), .QN(n13000) );
  NOR2X0 U12716 ( .IN1(n13001), .IN2(n13002), .QN(n11983) );
  INVX0 U12717 ( .INP(n12995), .ZN(n13002) );
  NAND2X0 U12718 ( .IN1(n13003), .IN2(n13004), .QN(n12995) );
  NAND2X0 U12719 ( .IN1(n9589), .IN2(n11946), .QN(n13004) );
  NOR2X0 U12720 ( .IN1(n13005), .IN2(n13006), .QN(n13003) );
  NOR2X0 U12721 ( .IN1(n4518), .IN2(g1703), .QN(n13006) );
  NOR2X0 U12722 ( .IN1(n4511), .IN2(g1702), .QN(n13005) );
  NAND2X0 U12723 ( .IN1(n13007), .IN2(n13008), .QN(g30249) );
  INVX0 U12724 ( .INP(n13009), .ZN(n13008) );
  NOR2X0 U12725 ( .IN1(g6518), .IN2(n9499), .QN(n13009) );
  NAND2X0 U12726 ( .IN1(n12944), .IN2(g6518), .QN(n13007) );
  NAND2X0 U12727 ( .IN1(n13010), .IN2(n13011), .QN(g30248) );
  INVX0 U12728 ( .INP(n13012), .ZN(n13011) );
  NOR2X0 U12729 ( .IN1(g165), .IN2(n9585), .QN(n13012) );
  NAND2X0 U12730 ( .IN1(n13013), .IN2(g165), .QN(n13010) );
  NAND2X0 U12731 ( .IN1(n13014), .IN2(n13015), .QN(g30247) );
  INVX0 U12732 ( .INP(n13016), .ZN(n13015) );
  NOR2X0 U12733 ( .IN1(g6368), .IN2(n9500), .QN(n13016) );
  NAND2X0 U12734 ( .IN1(n12944), .IN2(g6368), .QN(n13014) );
  NAND2X0 U12735 ( .IN1(n13017), .IN2(n13018), .QN(n12944) );
  NAND2X0 U12736 ( .IN1(n13019), .IN2(n12430), .QN(n13018) );
  NOR2X0 U12737 ( .IN1(n13020), .IN2(n13021), .QN(n13019) );
  NOR2X0 U12738 ( .IN1(n10816), .IN2(n12812), .QN(n13021) );
  INVX0 U12739 ( .INP(n13022), .ZN(n13020) );
  NAND2X0 U12740 ( .IN1(n12812), .IN2(n10816), .QN(n13022) );
  NAND2X0 U12741 ( .IN1(n13023), .IN2(n12846), .QN(n12812) );
  NOR2X0 U12742 ( .IN1(n12681), .IN2(n13024), .QN(n12846) );
  NOR2X0 U12743 ( .IN1(n12190), .IN2(n10823), .QN(n13024) );
  NAND2X0 U12744 ( .IN1(n12345), .IN2(n13025), .QN(n12681) );
  NAND2X0 U12745 ( .IN1(n13026), .IN2(n13027), .QN(n13025) );
  NAND2X0 U12746 ( .IN1(n10840), .IN2(n12190), .QN(n13027) );
  NAND2X0 U12747 ( .IN1(n12191), .IN2(n10839), .QN(n13026) );
  INVX0 U12748 ( .INP(n12344), .ZN(n12345) );
  NAND2X0 U12749 ( .IN1(n12155), .IN2(n13028), .QN(n12344) );
  NAND2X0 U12750 ( .IN1(n13029), .IN2(n13030), .QN(n13028) );
  NAND2X0 U12751 ( .IN1(n10861), .IN2(n12190), .QN(n13030) );
  NAND2X0 U12752 ( .IN1(n12191), .IN2(n10860), .QN(n13029) );
  INVX0 U12753 ( .INP(n12154), .ZN(n12155) );
  NAND2X0 U12754 ( .IN1(n12385), .IN2(n13031), .QN(n12154) );
  NAND2X0 U12755 ( .IN1(n13032), .IN2(n13033), .QN(n13031) );
  NAND2X0 U12756 ( .IN1(n10836), .IN2(n12190), .QN(n13033) );
  NAND2X0 U12757 ( .IN1(n12191), .IN2(n10835), .QN(n13032) );
  NAND2X0 U12758 ( .IN1(n13034), .IN2(n13035), .QN(n12385) );
  NAND2X0 U12759 ( .IN1(n12191), .IN2(n10831), .QN(n13035) );
  NAND2X0 U12760 ( .IN1(n13036), .IN2(n10832), .QN(n13034) );
  NOR2X0 U12761 ( .IN1(n13037), .IN2(n13038), .QN(n13023) );
  NOR2X0 U12762 ( .IN1(n10820), .IN2(n12191), .QN(n13038) );
  NOR2X0 U12763 ( .IN1(n10824), .IN2(n10819), .QN(n13037) );
  NAND2X0 U12764 ( .IN1(n12147), .IN2(g809), .QN(n13017) );
  NOR2X0 U12765 ( .IN1(n12430), .IN2(n12431), .QN(n12147) );
  NOR2X0 U12766 ( .IN1(n13039), .IN2(n13040), .QN(n12431) );
  NOR2X0 U12767 ( .IN1(n13039), .IN2(n13041), .QN(n12430) );
  NOR2X0 U12768 ( .IN1(n13040), .IN2(n13042), .QN(n13041) );
  NOR2X0 U12769 ( .IN1(n12190), .IN2(n13043), .QN(n13042) );
  INVX0 U12770 ( .INP(n13044), .ZN(n13043) );
  NAND2X0 U12771 ( .IN1(n12782), .IN2(n13045), .QN(n13040) );
  NAND2X0 U12772 ( .IN1(n13044), .IN2(n10803), .QN(n13045) );
  NAND2X0 U12773 ( .IN1(n13046), .IN2(n13047), .QN(n10803) );
  NOR2X0 U12774 ( .IN1(n10864), .IN2(n13048), .QN(n13047) );
  NAND2X0 U12775 ( .IN1(n10861), .IN2(n10857), .QN(n13048) );
  NOR2X0 U12776 ( .IN1(n13049), .IN2(n13050), .QN(n13046) );
  NAND2X0 U12777 ( .IN1(n10840), .IN2(n10836), .QN(n13050) );
  NAND2X0 U12778 ( .IN1(n13051), .IN2(n13052), .QN(n13044) );
  NOR2X0 U12779 ( .IN1(n13053), .IN2(n13054), .QN(n13052) );
  NAND2X0 U12780 ( .IN1(n10864), .IN2(n10856), .QN(n13054) );
  NAND2X0 U12781 ( .IN1(n10835), .IN2(n10839), .QN(n13053) );
  NOR2X0 U12782 ( .IN1(n12190), .IN2(n13055), .QN(n13051) );
  INVX0 U12783 ( .INP(n13056), .ZN(n13055) );
  NOR2X0 U12784 ( .IN1(n13049), .IN2(n10861), .QN(n13056) );
  NAND2X0 U12785 ( .IN1(n13057), .IN2(n13058), .QN(n13049) );
  NOR2X0 U12786 ( .IN1(n10819), .IN2(n13059), .QN(n13058) );
  NAND2X0 U12787 ( .IN1(n10816), .IN2(n12429), .QN(n13059) );
  NOR2X0 U12788 ( .IN1(n10823), .IN2(n10831), .QN(n13057) );
  NAND2X0 U12789 ( .IN1(n10804), .IN2(n12190), .QN(n12782) );
  NAND2X0 U12790 ( .IN1(n13060), .IN2(n13061), .QN(n13039) );
  NAND2X0 U12791 ( .IN1(n11796), .IN2(n11759), .QN(n13061) );
  NOR2X0 U12792 ( .IN1(n2617), .IN2(n13062), .QN(n13060) );
  NOR2X0 U12793 ( .IN1(n2632), .IN2(n13063), .QN(n13062) );
  NOR2X0 U12794 ( .IN1(n13064), .IN2(n13065), .QN(n13063) );
  NOR2X0 U12795 ( .IN1(n11765), .IN2(n13066), .QN(n13064) );
  NAND2X0 U12796 ( .IN1(n11766), .IN2(n11759), .QN(n13066) );
  NAND2X0 U12797 ( .IN1(n13067), .IN2(n13068), .QN(n2632) );
  NAND2X0 U12798 ( .IN1(n13069), .IN2(n13070), .QN(n13068) );
  NAND2X0 U12799 ( .IN1(n9595), .IN2(g1088), .QN(n13070) );
  NOR2X0 U12800 ( .IN1(n13071), .IN2(n13072), .QN(n13069) );
  NOR2X0 U12801 ( .IN1(n4364), .IN2(g1010), .QN(n13072) );
  NOR2X0 U12802 ( .IN1(n4363), .IN2(g1009), .QN(n13071) );
  NAND2X0 U12803 ( .IN1(n13073), .IN2(n13074), .QN(g30246) );
  NAND2X0 U12804 ( .IN1(n4512), .IN2(g216), .QN(n13074) );
  NAND2X0 U12805 ( .IN1(n13013), .IN2(g6313), .QN(n13073) );
  NAND2X0 U12806 ( .IN1(n13075), .IN2(n13076), .QN(g30245) );
  INVX0 U12807 ( .INP(n13077), .ZN(n13076) );
  NOR2X0 U12808 ( .IN1(g6231), .IN2(n9514), .QN(n13077) );
  NAND2X0 U12809 ( .IN1(n13013), .IN2(g6231), .QN(n13075) );
  NAND2X0 U12810 ( .IN1(n13078), .IN2(n13079), .QN(n13013) );
  NAND2X0 U12811 ( .IN1(n13080), .IN2(n12463), .QN(n13079) );
  NOR2X0 U12812 ( .IN1(n13081), .IN2(n13082), .QN(n13080) );
  NOR2X0 U12813 ( .IN1(n10751), .IN2(n13083), .QN(n13082) );
  NOR2X0 U12814 ( .IN1(n12857), .IN2(n10750), .QN(n13081) );
  INVX0 U12815 ( .INP(n13083), .ZN(n12857) );
  NAND2X0 U12816 ( .IN1(n13084), .IN2(n12879), .QN(n13083) );
  NOR2X0 U12817 ( .IN1(n12734), .IN2(n13085), .QN(n12879) );
  NOR2X0 U12818 ( .IN1(n11773), .IN2(n10774), .QN(n13085) );
  NAND2X0 U12819 ( .IN1(n13086), .IN2(n13087), .QN(n12734) );
  INVX0 U12820 ( .INP(n12407), .ZN(n13087) );
  NAND2X0 U12821 ( .IN1(n12207), .IN2(n13088), .QN(n12407) );
  NAND2X0 U12822 ( .IN1(n11774), .IN2(n10767), .QN(n13088) );
  INVX0 U12823 ( .INP(n12206), .ZN(n12207) );
  NAND2X0 U12824 ( .IN1(n12442), .IN2(n13089), .QN(n12206) );
  NAND2X0 U12825 ( .IN1(n13090), .IN2(n13091), .QN(n13089) );
  NAND2X0 U12826 ( .IN1(n10755), .IN2(n11773), .QN(n13091) );
  NAND2X0 U12827 ( .IN1(n11774), .IN2(n10754), .QN(n13090) );
  INVX0 U12828 ( .INP(n12443), .ZN(n12442) );
  NAND2X0 U12829 ( .IN1(n13092), .IN2(n12831), .QN(n12443) );
  NAND2X0 U12830 ( .IN1(n13093), .IN2(n13094), .QN(n13092) );
  NAND2X0 U12831 ( .IN1(n4513), .IN2(n11773), .QN(n13094) );
  INVX0 U12832 ( .INP(n10796), .ZN(n4513) );
  NAND2X0 U12833 ( .IN1(n11774), .IN2(n10796), .QN(n13093) );
  NAND2X0 U12834 ( .IN1(n13095), .IN2(n13096), .QN(n10796) );
  NAND2X0 U12835 ( .IN1(test_so13), .IN2(g6313), .QN(n13096) );
  NOR2X0 U12836 ( .IN1(n13097), .IN2(n13098), .QN(n13095) );
  NOR2X0 U12837 ( .IN1(n9587), .IN2(n4369), .QN(n13098) );
  NOR2X0 U12838 ( .IN1(n9523), .IN2(n4318), .QN(n13097) );
  NOR2X0 U12839 ( .IN1(n13099), .IN2(n13100), .QN(n13086) );
  NOR2X0 U12840 ( .IN1(n12405), .IN2(n11774), .QN(n13100) );
  NOR2X0 U12841 ( .IN1(n10767), .IN2(n10784), .QN(n13099) );
  NOR2X0 U12842 ( .IN1(n13101), .IN2(n13102), .QN(n13084) );
  NOR2X0 U12843 ( .IN1(n10800), .IN2(n11774), .QN(n13102) );
  NOR2X0 U12844 ( .IN1(n10775), .IN2(n10799), .QN(n13101) );
  NAND2X0 U12845 ( .IN1(n12246), .IN2(g121), .QN(n13078) );
  NOR2X0 U12846 ( .IN1(n12463), .IN2(n12445), .QN(n12246) );
  NOR2X0 U12847 ( .IN1(n13103), .IN2(n13104), .QN(n12445) );
  NAND2X0 U12848 ( .IN1(n12831), .IN2(n13105), .QN(n13103) );
  NAND2X0 U12849 ( .IN1(n10738), .IN2(n13106), .QN(n13105) );
  NOR2X0 U12850 ( .IN1(n13104), .IN2(n13107), .QN(n12463) );
  NOR2X0 U12851 ( .IN1(n13108), .IN2(n12830), .QN(n13107) );
  INVX0 U12852 ( .INP(n12831), .ZN(n12830) );
  NAND2X0 U12853 ( .IN1(n11773), .IN2(n10739), .QN(n12831) );
  INVX0 U12854 ( .INP(n13109), .ZN(n10739) );
  INVX0 U12855 ( .INP(n13110), .ZN(n13108) );
  NAND2X0 U12856 ( .IN1(n13106), .IN2(n13111), .QN(n13110) );
  NAND2X0 U12857 ( .IN1(n13112), .IN2(n11773), .QN(n13111) );
  INVX0 U12858 ( .INP(n10738), .ZN(n13112) );
  NAND2X0 U12859 ( .IN1(n13113), .IN2(n13114), .QN(n10738) );
  NOR2X0 U12860 ( .IN1(n10754), .IN2(n13115), .QN(n13114) );
  NAND2X0 U12861 ( .IN1(n10793), .IN2(n12405), .QN(n13115) );
  NOR2X0 U12862 ( .IN1(n13116), .IN2(n13117), .QN(n13113) );
  NAND2X0 U12863 ( .IN1(n10771), .IN2(n10767), .QN(n13117) );
  NAND2X0 U12864 ( .IN1(n13118), .IN2(n13119), .QN(n13106) );
  NOR2X0 U12865 ( .IN1(n13120), .IN2(n13121), .QN(n13119) );
  NAND2X0 U12866 ( .IN1(n10792), .IN2(n10754), .QN(n13121) );
  NAND2X0 U12867 ( .IN1(n10770), .IN2(n10766), .QN(n13120) );
  NOR2X0 U12868 ( .IN1(n11773), .IN2(n13122), .QN(n13118) );
  INVX0 U12869 ( .INP(n13123), .ZN(n13122) );
  NOR2X0 U12870 ( .IN1(n13116), .IN2(n12405), .QN(n13123) );
  NAND2X0 U12871 ( .IN1(n13124), .IN2(n13125), .QN(n13116) );
  NOR2X0 U12872 ( .IN1(n10758), .IN2(n13126), .QN(n13125) );
  NAND2X0 U12873 ( .IN1(n10751), .IN2(n10800), .QN(n13126) );
  NOR2X0 U12874 ( .IN1(n10774), .IN2(n13127), .QN(n13124) );
  NAND2X0 U12875 ( .IN1(n13128), .IN2(n13129), .QN(n13104) );
  NAND2X0 U12876 ( .IN1(n13130), .IN2(n13131), .QN(n13129) );
  NOR2X0 U12877 ( .IN1(n12003), .IN2(n13132), .QN(n13128) );
  NOR2X0 U12878 ( .IN1(n12011), .IN2(n13133), .QN(n13132) );
  NOR2X0 U12879 ( .IN1(n13134), .IN2(n12032), .QN(n13133) );
  NOR2X0 U12880 ( .IN1(n12538), .IN2(n13135), .QN(n13134) );
  NAND2X0 U12881 ( .IN1(n12033), .IN2(n12028), .QN(n13135) );
  NOR2X0 U12882 ( .IN1(n13136), .IN2(n13137), .QN(n12033) );
  INVX0 U12883 ( .INP(n13130), .ZN(n13137) );
  NAND2X0 U12884 ( .IN1(n13138), .IN2(n13139), .QN(n13130) );
  NAND2X0 U12885 ( .IN1(n9599), .IN2(n12042), .QN(n13139) );
  NOR2X0 U12886 ( .IN1(n13140), .IN2(n13141), .QN(n13138) );
  NOR2X0 U12887 ( .IN1(n4506), .IN2(g321), .QN(n13141) );
  NOR2X0 U12888 ( .IN1(n4499), .IN2(g323), .QN(n13140) );
  NAND2X0 U12889 ( .IN1(n13142), .IN2(n13143), .QN(g30072) );
  NAND2X0 U12890 ( .IN1(g2574), .IN2(n7930), .QN(n13143) );
  NAND2X0 U12891 ( .IN1(n4543), .IN2(n13144), .QN(n13142) );
  NAND2X0 U12892 ( .IN1(n13145), .IN2(n13146), .QN(n13144) );
  NAND2X0 U12893 ( .IN1(n618), .IN2(n13147), .QN(n13146) );
  NAND2X0 U12894 ( .IN1(n13148), .IN2(n7929), .QN(n13145) );
  NAND2X0 U12895 ( .IN1(n13149), .IN2(n13150), .QN(g30061) );
  NAND2X0 U12896 ( .IN1(g2580), .IN2(n7926), .QN(n13150) );
  NAND2X0 U12897 ( .IN1(n9796), .IN2(n13151), .QN(n13149) );
  NAND2X0 U12898 ( .IN1(n13152), .IN2(n13153), .QN(n13151) );
  NAND2X0 U12899 ( .IN1(n4370), .IN2(g16437), .QN(n13153) );
  NAND2X0 U12900 ( .IN1(n626), .IN2(g7390), .QN(n13152) );
  INVX0 U12901 ( .INP(n13154), .ZN(n626) );
  NAND2X0 U12902 ( .IN1(n13155), .IN2(n13156), .QN(n13154) );
  NAND2X0 U12903 ( .IN1(g1886), .IN2(DFF_1133_n1), .QN(n13156) );
  NAND2X0 U12904 ( .IN1(n4493), .IN2(n13157), .QN(n13155) );
  NAND2X0 U12905 ( .IN1(n13158), .IN2(n13159), .QN(n13157) );
  NAND2X0 U12906 ( .IN1(n4315), .IN2(DFF_1142_n1), .QN(n13159) );
  NAND2X0 U12907 ( .IN1(n10723), .IN2(g7194), .QN(n13158) );
  NAND2X0 U12908 ( .IN1(n13160), .IN2(n13161), .QN(n10723) );
  NAND2X0 U12909 ( .IN1(g1192), .IN2(DFF_783_n1), .QN(n13161) );
  NAND2X0 U12910 ( .IN1(n4454), .IN2(n13162), .QN(n13160) );
  NAND2X0 U12911 ( .IN1(n13163), .IN2(n13164), .QN(n13162) );
  NAND2X0 U12912 ( .IN1(n4316), .IN2(DFF_792_n1), .QN(n13164) );
  NAND2X0 U12913 ( .IN1(n10722), .IN2(g6944), .QN(n13163) );
  NAND2X0 U12914 ( .IN1(n13165), .IN2(n13166), .QN(n10722) );
  NAND2X0 U12915 ( .IN1(n9713), .IN2(g506), .QN(n13166) );
  NAND2X0 U12916 ( .IN1(n13167), .IN2(n4570), .QN(n13165) );
  NOR2X0 U12917 ( .IN1(g16297), .IN2(g6642), .QN(n13167) );
  NAND2X0 U12918 ( .IN1(n13168), .IN2(n13169), .QN(g30055) );
  NAND2X0 U12919 ( .IN1(n4487), .IN2(DFF_1378_n1), .QN(n13169) );
  NAND2X0 U12920 ( .IN1(n13170), .IN2(g2374), .QN(n13168) );
  NAND2X0 U12921 ( .IN1(n13171), .IN2(n13172), .QN(n13170) );
  NAND2X0 U12922 ( .IN1(n530), .IN2(g7264), .QN(n13172) );
  INVX0 U12923 ( .INP(n13173), .ZN(n530) );
  NAND2X0 U12924 ( .IN1(n13174), .IN2(n13175), .QN(n13173) );
  NAND2X0 U12925 ( .IN1(n4488), .IN2(n7978), .QN(n13175) );
  NAND2X0 U12926 ( .IN1(n13176), .IN2(g1680), .QN(n13174) );
  NOR2X0 U12927 ( .IN1(n13177), .IN2(n13178), .QN(n13176) );
  NOR2X0 U12928 ( .IN1(n10027), .IN2(n11946), .QN(n13178) );
  NOR2X0 U12929 ( .IN1(n10726), .IN2(n13179), .QN(n13177) );
  NAND2X0 U12930 ( .IN1(n13180), .IN2(n13181), .QN(n10726) );
  NAND2X0 U12931 ( .IN1(n4432), .IN2(n8017), .QN(n13181) );
  NAND2X0 U12932 ( .IN1(n13182), .IN2(g986), .QN(n13180) );
  NAND2X0 U12933 ( .IN1(n13183), .IN2(n13184), .QN(n13182) );
  NAND2X0 U12934 ( .IN1(n4364), .IN2(n10028), .QN(n13184) );
  INVX0 U12935 ( .INP(n13185), .ZN(n13183) );
  NOR2X0 U12936 ( .IN1(g21346), .IN2(n4364), .QN(n13185) );
  NAND2X0 U12937 ( .IN1(n4524), .IN2(g2380), .QN(n13171) );
  NAND2X0 U12938 ( .IN1(n13186), .IN2(n13187), .QN(g29941) );
  NAND2X0 U12939 ( .IN1(n4494), .IN2(g3105), .QN(n13187) );
  NAND2X0 U12940 ( .IN1(n618), .IN2(g3109), .QN(n13186) );
  NAND2X0 U12941 ( .IN1(n13188), .IN2(n13189), .QN(g29939) );
  INVX0 U12942 ( .INP(n13190), .ZN(n13189) );
  NOR2X0 U12943 ( .IN1(g8030), .IN2(n4452), .QN(n13190) );
  NAND2X0 U12944 ( .IN1(n618), .IN2(g8030), .QN(n13188) );
  NAND2X0 U12945 ( .IN1(n13191), .IN2(n13192), .QN(g29936) );
  INVX0 U12946 ( .INP(n13193), .ZN(n13192) );
  NOR2X0 U12947 ( .IN1(g8106), .IN2(n4447), .QN(n13193) );
  NAND2X0 U12948 ( .IN1(n618), .IN2(g8106), .QN(n13191) );
  INVX0 U12949 ( .INP(n13194), .ZN(n618) );
  NAND2X0 U12950 ( .IN1(n13195), .IN2(n13196), .QN(n13194) );
  NAND2X0 U12951 ( .IN1(g1880), .IN2(DFF_1099_n1), .QN(n13196) );
  NAND2X0 U12952 ( .IN1(n13197), .IN2(n4545), .QN(n13195) );
  NOR2X0 U12953 ( .IN1(n13198), .IN2(n13199), .QN(n13197) );
  NOR2X0 U12954 ( .IN1(g7052), .IN2(DFF_1100_n1), .QN(n13199) );
  NOR2X0 U12955 ( .IN1(n4296), .IN2(n13200), .QN(n13198) );
  NAND2X0 U12956 ( .IN1(n13201), .IN2(n13202), .QN(g29623) );
  NAND2X0 U12957 ( .IN1(n13203), .IN2(n4606), .QN(n13202) );
  NAND2X0 U12958 ( .IN1(n4509), .IN2(g2389), .QN(n13201) );
  NAND2X0 U12959 ( .IN1(n13204), .IN2(n13205), .QN(g29621) );
  NAND2X0 U12960 ( .IN1(n13203), .IN2(g7264), .QN(n13205) );
  INVX0 U12961 ( .INP(n13206), .ZN(n13204) );
  NOR2X0 U12962 ( .IN1(n11937), .IN2(n9536), .QN(n13206) );
  NAND2X0 U12963 ( .IN1(n13207), .IN2(n13208), .QN(g29620) );
  NAND2X0 U12964 ( .IN1(n13209), .IN2(n4618), .QN(n13208) );
  NAND2X0 U12965 ( .IN1(n4511), .IN2(g1695), .QN(n13207) );
  NAND2X0 U12966 ( .IN1(n13210), .IN2(n13211), .QN(g29618) );
  NAND2X0 U12967 ( .IN1(n13203), .IN2(g5555), .QN(n13211) );
  NOR2X0 U12968 ( .IN1(n13212), .IN2(n12467), .QN(n13203) );
  INVX0 U12969 ( .INP(n13213), .ZN(n12467) );
  NAND2X0 U12970 ( .IN1(n12934), .IN2(n13214), .QN(n13213) );
  NOR2X0 U12971 ( .IN1(n4529), .IN2(n13215), .QN(n13212) );
  NOR2X0 U12972 ( .IN1(n13216), .IN2(n12932), .QN(n13215) );
  NAND2X0 U12973 ( .IN1(n12564), .IN2(n12478), .QN(n13216) );
  INVX0 U12974 ( .INP(n11780), .ZN(n4529) );
  NAND2X0 U12975 ( .IN1(n13217), .IN2(n12498), .QN(n11780) );
  NOR2X0 U12976 ( .IN1(n12491), .IN2(n12478), .QN(n13217) );
  NAND2X0 U12977 ( .IN1(n4516), .IN2(g2387), .QN(n13210) );
  NAND2X0 U12978 ( .IN1(n13218), .IN2(n13219), .QN(g29617) );
  NAND2X0 U12979 ( .IN1(n13209), .IN2(g7014), .QN(n13219) );
  INVX0 U12980 ( .INP(n13220), .ZN(n13218) );
  NOR2X0 U12981 ( .IN1(n11946), .IN2(n9539), .QN(n13220) );
  NAND2X0 U12982 ( .IN1(n13221), .IN2(n13222), .QN(g29616) );
  INVX0 U12983 ( .INP(n13223), .ZN(n13222) );
  NOR2X0 U12984 ( .IN1(g1088), .IN2(n9558), .QN(n13223) );
  NAND2X0 U12985 ( .IN1(n13224), .IN2(g1088), .QN(n13221) );
  NAND2X0 U12986 ( .IN1(n13225), .IN2(n13226), .QN(g29613) );
  NAND2X0 U12987 ( .IN1(n13209), .IN2(g5511), .QN(n13226) );
  NOR2X0 U12988 ( .IN1(n13227), .IN2(n11953), .QN(n13209) );
  INVX0 U12989 ( .INP(n13228), .ZN(n11953) );
  NAND2X0 U12990 ( .IN1(n13229), .IN2(n13230), .QN(n13228) );
  NOR2X0 U12991 ( .IN1(n4530), .IN2(n13231), .QN(n13227) );
  INVX0 U12992 ( .INP(n13232), .ZN(n13231) );
  NAND2X0 U12993 ( .IN1(n13233), .IN2(n12585), .QN(n13232) );
  NOR2X0 U12994 ( .IN1(n11961), .IN2(n13234), .QN(n13233) );
  INVX0 U12995 ( .INP(n11777), .ZN(n4530) );
  NAND2X0 U12996 ( .IN1(n13235), .IN2(n11985), .QN(n11777) );
  NOR2X0 U12997 ( .IN1(n11978), .IN2(n11964), .QN(n13235) );
  NAND2X0 U12998 ( .IN1(n4518), .IN2(g1693), .QN(n13225) );
  NAND2X0 U12999 ( .IN1(n13236), .IN2(n13237), .QN(g29612) );
  NAND2X0 U13000 ( .IN1(n4364), .IN2(g1000), .QN(n13237) );
  NAND2X0 U13001 ( .IN1(n13224), .IN2(g6712), .QN(n13236) );
  NAND2X0 U13002 ( .IN1(n13238), .IN2(n13239), .QN(g29611) );
  NAND2X0 U13003 ( .IN1(n13240), .IN2(n4640), .QN(n13239) );
  NAND2X0 U13004 ( .IN1(n4506), .IN2(g314), .QN(n13238) );
  NAND2X0 U13005 ( .IN1(n13241), .IN2(n13242), .QN(g29609) );
  NAND2X0 U13006 ( .IN1(n4363), .IN2(g999), .QN(n13242) );
  NAND2X0 U13007 ( .IN1(n13224), .IN2(g5472), .QN(n13241) );
  NOR2X0 U13008 ( .IN1(n13243), .IN2(n2617), .QN(n13224) );
  INVX0 U13009 ( .INP(n13244), .ZN(n2617) );
  NAND2X0 U13010 ( .IN1(n13067), .IN2(n13245), .QN(n13244) );
  NOR2X0 U13011 ( .IN1(n12191), .IN2(n13246), .QN(n13243) );
  NOR2X0 U13012 ( .IN1(n13247), .IN2(n13065), .QN(n13246) );
  NAND2X0 U13013 ( .IN1(n11765), .IN2(n11759), .QN(n13247) );
  INVX0 U13014 ( .INP(n12190), .ZN(n12191) );
  NAND2X0 U13015 ( .IN1(n13248), .IN2(n11756), .QN(n12190) );
  NOR2X0 U13016 ( .IN1(n11766), .IN2(n11759), .QN(n13248) );
  NAND2X0 U13017 ( .IN1(n13249), .IN2(n13250), .QN(g29608) );
  NAND2X0 U13018 ( .IN1(n13240), .IN2(g6447), .QN(n13250) );
  NAND2X0 U13019 ( .IN1(n4499), .IN2(g313), .QN(n13249) );
  NAND2X0 U13020 ( .IN1(n13251), .IN2(n13252), .QN(g29606) );
  NAND2X0 U13021 ( .IN1(n13240), .IN2(g5437), .QN(n13252) );
  NOR2X0 U13022 ( .IN1(n13253), .IN2(n12003), .QN(n13240) );
  INVX0 U13023 ( .INP(n13254), .ZN(n12003) );
  NAND2X0 U13024 ( .IN1(n13255), .IN2(n13256), .QN(n13254) );
  NOR2X0 U13025 ( .IN1(n11774), .IN2(n13257), .QN(n13253) );
  INVX0 U13026 ( .INP(n13258), .ZN(n13257) );
  NAND2X0 U13027 ( .IN1(n13259), .IN2(n12538), .QN(n13258) );
  NOR2X0 U13028 ( .IN1(n12011), .IN2(n13260), .QN(n13259) );
  INVX0 U13029 ( .INP(n11773), .ZN(n11774) );
  NAND2X0 U13030 ( .IN1(n13261), .IN2(n12035), .QN(n11773) );
  NOR2X0 U13031 ( .IN1(n12028), .IN2(n12014), .QN(n13261) );
  INVX0 U13032 ( .INP(n13262), .ZN(n13251) );
  NOR2X0 U13033 ( .IN1(n12042), .IN2(n9567), .QN(n13262) );
  NOR2X0 U13034 ( .IN1(n13263), .IN2(n13264), .QN(g29582) );
  NOR2X0 U13035 ( .IN1(n13265), .IN2(n13266), .QN(n13264) );
  INVX0 U13036 ( .INP(n13267), .ZN(n13266) );
  NAND2X0 U13037 ( .IN1(g2120), .IN2(n2981), .QN(n13267) );
  NOR2X0 U13038 ( .IN1(n2981), .IN2(g2120), .QN(n13265) );
  NOR2X0 U13039 ( .IN1(n13268), .IN2(n13269), .QN(g29581) );
  NOR2X0 U13040 ( .IN1(n13270), .IN2(n13271), .QN(n13269) );
  INVX0 U13041 ( .INP(n13272), .ZN(n13271) );
  NAND2X0 U13042 ( .IN1(g1426), .IN2(n2984), .QN(n13272) );
  NOR2X0 U13043 ( .IN1(n2984), .IN2(g1426), .QN(n13270) );
  NOR2X0 U13044 ( .IN1(n13273), .IN2(n13274), .QN(g29580) );
  NOR2X0 U13045 ( .IN1(n13275), .IN2(n13276), .QN(n13274) );
  INVX0 U13046 ( .INP(n13277), .ZN(n13276) );
  NAND2X0 U13047 ( .IN1(g740), .IN2(n2987), .QN(n13277) );
  NOR2X0 U13048 ( .IN1(n2987), .IN2(g740), .QN(n13275) );
  NOR2X0 U13049 ( .IN1(n13278), .IN2(n13279), .QN(g29579) );
  NOR2X0 U13050 ( .IN1(n13280), .IN2(n13281), .QN(n13279) );
  INVX0 U13051 ( .INP(n13282), .ZN(n13281) );
  NAND2X0 U13052 ( .IN1(g52), .IN2(n2990), .QN(n13282) );
  NOR2X0 U13053 ( .IN1(n2990), .IN2(g52), .QN(n13280) );
  NAND2X0 U13054 ( .IN1(n13283), .IN2(n13284), .QN(g29357) );
  NAND2X0 U13055 ( .IN1(n13285), .IN2(g2124), .QN(n13284) );
  INVX0 U13056 ( .INP(n13286), .ZN(n13285) );
  NAND2X0 U13057 ( .IN1(n13287), .IN2(n9600), .QN(n13283) );
  NOR2X0 U13058 ( .IN1(n13263), .IN2(n2982), .QN(n13287) );
  NAND2X0 U13059 ( .IN1(n13288), .IN2(n13289), .QN(g29355) );
  NAND2X0 U13060 ( .IN1(n13290), .IN2(g1430), .QN(n13289) );
  INVX0 U13061 ( .INP(n13291), .ZN(n13290) );
  NAND2X0 U13062 ( .IN1(n13292), .IN2(n9601), .QN(n13288) );
  NOR2X0 U13063 ( .IN1(n13268), .IN2(n2985), .QN(n13292) );
  NAND2X0 U13064 ( .IN1(n13293), .IN2(n13294), .QN(g29354) );
  NAND2X0 U13065 ( .IN1(n13295), .IN2(g744), .QN(n13294) );
  INVX0 U13066 ( .INP(n13296), .ZN(n13295) );
  NAND2X0 U13067 ( .IN1(n13297), .IN2(n9602), .QN(n13293) );
  NOR2X0 U13068 ( .IN1(n13273), .IN2(n2988), .QN(n13297) );
  NAND2X0 U13069 ( .IN1(n13298), .IN2(n13299), .QN(g29353) );
  NAND2X0 U13070 ( .IN1(n13300), .IN2(g56), .QN(n13299) );
  INVX0 U13071 ( .INP(n13301), .ZN(n13300) );
  NAND2X0 U13072 ( .IN1(n13302), .IN2(n9603), .QN(n13298) );
  NOR2X0 U13073 ( .IN1(n13278), .IN2(n2991), .QN(n13302) );
  NAND2X0 U13074 ( .IN1(n13303), .IN2(n13304), .QN(g29226) );
  NAND2X0 U13075 ( .IN1(n13305), .IN2(n4606), .QN(n13304) );
  INVX0 U13076 ( .INP(n13306), .ZN(n13303) );
  NOR2X0 U13077 ( .IN1(n13307), .IN2(n9756), .QN(n13306) );
  NAND2X0 U13078 ( .IN1(n13308), .IN2(n13309), .QN(g29221) );
  NAND2X0 U13079 ( .IN1(n13305), .IN2(g7264), .QN(n13309) );
  INVX0 U13080 ( .INP(n13310), .ZN(n13308) );
  NOR2X0 U13081 ( .IN1(n11937), .IN2(n9743), .QN(n13310) );
  NAND2X0 U13082 ( .IN1(n13311), .IN2(n13312), .QN(g29218) );
  NAND2X0 U13083 ( .IN1(n13313), .IN2(n4618), .QN(n13312) );
  INVX0 U13084 ( .INP(n13314), .ZN(n13311) );
  NOR2X0 U13085 ( .IN1(n13315), .IN2(n9762), .QN(n13314) );
  NAND2X0 U13086 ( .IN1(n13316), .IN2(n13317), .QN(g29213) );
  NAND2X0 U13087 ( .IN1(n13305), .IN2(g5555), .QN(n13317) );
  NOR2X0 U13088 ( .IN1(n13318), .IN2(n13319), .QN(n13305) );
  INVX0 U13089 ( .INP(n13320), .ZN(n13319) );
  NAND2X0 U13090 ( .IN1(n13321), .IN2(n13322), .QN(n13320) );
  NOR2X0 U13091 ( .IN1(n13321), .IN2(n13322), .QN(n13318) );
  NAND2X0 U13092 ( .IN1(n13323), .IN2(n13324), .QN(n13321) );
  NOR2X0 U13093 ( .IN1(n13325), .IN2(n13326), .QN(n13324) );
  NOR2X0 U13094 ( .IN1(n4285), .IN2(n13327), .QN(n13326) );
  NOR2X0 U13095 ( .IN1(n13322), .IN2(n11748), .QN(n13325) );
  NOR2X0 U13096 ( .IN1(n13328), .IN2(n10322), .QN(n13323) );
  INVX0 U13097 ( .INP(n13329), .ZN(n13328) );
  NAND2X0 U13098 ( .IN1(n11746), .IN2(n13330), .QN(n13329) );
  NAND2X0 U13099 ( .IN1(n11747), .IN2(n13331), .QN(n13330) );
  NAND2X0 U13100 ( .IN1(n12495), .IN2(n13322), .QN(n11746) );
  NAND2X0 U13101 ( .IN1(n4516), .IN2(g2492), .QN(n13316) );
  NAND2X0 U13102 ( .IN1(n13332), .IN2(n13333), .QN(g29212) );
  NAND2X0 U13103 ( .IN1(n13313), .IN2(g7014), .QN(n13333) );
  INVX0 U13104 ( .INP(n13334), .ZN(n13332) );
  NOR2X0 U13105 ( .IN1(n11946), .IN2(n9747), .QN(n13334) );
  NAND2X0 U13106 ( .IN1(n13335), .IN2(n13336), .QN(g29209) );
  NAND2X0 U13107 ( .IN1(n4381), .IN2(g1110), .QN(n13336) );
  NAND2X0 U13108 ( .IN1(n13337), .IN2(g1088), .QN(n13335) );
  NAND2X0 U13109 ( .IN1(n13338), .IN2(n13339), .QN(g29205) );
  NAND2X0 U13110 ( .IN1(n13313), .IN2(g5511), .QN(n13339) );
  NOR2X0 U13111 ( .IN1(n13340), .IN2(n13341), .QN(n13313) );
  INVX0 U13112 ( .INP(n13342), .ZN(n13341) );
  NAND2X0 U13113 ( .IN1(n13343), .IN2(n13344), .QN(n13342) );
  NOR2X0 U13114 ( .IN1(n13343), .IN2(n13344), .QN(n13340) );
  NAND2X0 U13115 ( .IN1(n13345), .IN2(n13346), .QN(n13343) );
  NOR2X0 U13116 ( .IN1(n13347), .IN2(n13348), .QN(n13346) );
  NOR2X0 U13117 ( .IN1(n4284), .IN2(n13349), .QN(n13348) );
  NOR2X0 U13118 ( .IN1(n13344), .IN2(n11743), .QN(n13347) );
  NOR2X0 U13119 ( .IN1(n4386), .IN2(n13350), .QN(n13345) );
  INVX0 U13120 ( .INP(n13351), .ZN(n13350) );
  NAND2X0 U13121 ( .IN1(n11741), .IN2(n13352), .QN(n13351) );
  NAND2X0 U13122 ( .IN1(n11742), .IN2(n13353), .QN(n13352) );
  NAND2X0 U13123 ( .IN1(n11982), .IN2(n13344), .QN(n11741) );
  NAND2X0 U13124 ( .IN1(n4518), .IN2(g1798), .QN(n13338) );
  NAND2X0 U13125 ( .IN1(n13354), .IN2(n13355), .QN(g29204) );
  INVX0 U13126 ( .INP(n13356), .ZN(n13355) );
  NOR2X0 U13127 ( .IN1(g6712), .IN2(n9750), .QN(n13356) );
  NAND2X0 U13128 ( .IN1(n13337), .IN2(g6712), .QN(n13354) );
  NAND2X0 U13129 ( .IN1(n13357), .IN2(n13358), .QN(g29201) );
  NAND2X0 U13130 ( .IN1(n13359), .IN2(n4640), .QN(n13358) );
  INVX0 U13131 ( .INP(n13360), .ZN(n13357) );
  NOR2X0 U13132 ( .IN1(n13361), .IN2(n9780), .QN(n13360) );
  NAND2X0 U13133 ( .IN1(n13362), .IN2(n13363), .QN(g29198) );
  INVX0 U13134 ( .INP(n13364), .ZN(n13363) );
  NOR2X0 U13135 ( .IN1(g5472), .IN2(n9771), .QN(n13364) );
  NAND2X0 U13136 ( .IN1(n13337), .IN2(g5472), .QN(n13362) );
  NOR2X0 U13137 ( .IN1(n13365), .IN2(n13366), .QN(n13337) );
  INVX0 U13138 ( .INP(n13367), .ZN(n13366) );
  NAND2X0 U13139 ( .IN1(n13368), .IN2(n13369), .QN(n13367) );
  NOR2X0 U13140 ( .IN1(n13368), .IN2(n13369), .QN(n13365) );
  NAND2X0 U13141 ( .IN1(n13370), .IN2(n13371), .QN(n13368) );
  NOR2X0 U13142 ( .IN1(n13372), .IN2(n13373), .QN(n13371) );
  NOR2X0 U13143 ( .IN1(n4283), .IN2(n13374), .QN(n13373) );
  NOR2X0 U13144 ( .IN1(n13369), .IN2(n11738), .QN(n13372) );
  NOR2X0 U13145 ( .IN1(n4387), .IN2(n13375), .QN(n13370) );
  INVX0 U13146 ( .INP(n13376), .ZN(n13375) );
  NAND2X0 U13147 ( .IN1(n11736), .IN2(n13377), .QN(n13376) );
  NAND2X0 U13148 ( .IN1(n11737), .IN2(n13378), .QN(n13377) );
  NAND2X0 U13149 ( .IN1(n11796), .IN2(n13369), .QN(n11736) );
  NAND2X0 U13150 ( .IN1(n13379), .IN2(n13380), .QN(g29197) );
  NAND2X0 U13151 ( .IN1(n13359), .IN2(g6447), .QN(n13380) );
  INVX0 U13152 ( .INP(n13381), .ZN(n13379) );
  NOR2X0 U13153 ( .IN1(n13382), .IN2(n9781), .QN(n13381) );
  NAND2X0 U13154 ( .IN1(n13383), .IN2(n13384), .QN(g29194) );
  NAND2X0 U13155 ( .IN1(n13359), .IN2(g5437), .QN(n13384) );
  NOR2X0 U13156 ( .IN1(n13385), .IN2(n13386), .QN(n13359) );
  INVX0 U13157 ( .INP(n13387), .ZN(n13386) );
  NAND2X0 U13158 ( .IN1(n13388), .IN2(n13389), .QN(n13387) );
  NOR2X0 U13159 ( .IN1(n13388), .IN2(n13389), .QN(n13385) );
  NAND2X0 U13160 ( .IN1(n13390), .IN2(n13391), .QN(n13388) );
  NOR2X0 U13161 ( .IN1(n13392), .IN2(n13393), .QN(n13391) );
  NOR2X0 U13162 ( .IN1(n4282), .IN2(n13394), .QN(n13393) );
  NOR2X0 U13163 ( .IN1(n13389), .IN2(n11733), .QN(n13392) );
  NOR2X0 U13164 ( .IN1(n4388), .IN2(n13395), .QN(n13390) );
  NOR2X0 U13165 ( .IN1(n13396), .IN2(n13397), .QN(n13395) );
  NOR2X0 U13166 ( .IN1(n13398), .IN2(n13399), .QN(n13397) );
  INVX0 U13167 ( .INP(n11731), .ZN(n13396) );
  NAND2X0 U13168 ( .IN1(n12032), .IN2(n13389), .QN(n11731) );
  NAND2X0 U13169 ( .IN1(n4520), .IN2(g417), .QN(n13383) );
  NAND2X0 U13170 ( .IN1(n13400), .IN2(n13401), .QN(g29187) );
  NAND2X0 U13171 ( .IN1(n13402), .IN2(g2396), .QN(n13401) );
  NAND2X0 U13172 ( .IN1(n13403), .IN2(n13307), .QN(n13402) );
  NAND2X0 U13173 ( .IN1(n13404), .IN2(n13307), .QN(n13400) );
  NAND2X0 U13174 ( .IN1(n13405), .IN2(n13406), .QN(g29185) );
  NAND2X0 U13175 ( .IN1(n13407), .IN2(g2398), .QN(n13406) );
  NAND2X0 U13176 ( .IN1(n13403), .IN2(n11937), .QN(n13407) );
  NAND2X0 U13177 ( .IN1(n13404), .IN2(n11937), .QN(n13405) );
  NAND2X0 U13178 ( .IN1(n13408), .IN2(n13409), .QN(g29184) );
  NAND2X0 U13179 ( .IN1(n13410), .IN2(g1702), .QN(n13409) );
  NAND2X0 U13180 ( .IN1(n13411), .IN2(n13315), .QN(n13410) );
  NAND2X0 U13181 ( .IN1(n13412), .IN2(n13315), .QN(n13408) );
  NAND2X0 U13182 ( .IN1(n13413), .IN2(n13414), .QN(g29182) );
  NAND2X0 U13183 ( .IN1(n13415), .IN2(g2397), .QN(n13414) );
  NAND2X0 U13184 ( .IN1(n13403), .IN2(n13416), .QN(n13415) );
  NAND2X0 U13185 ( .IN1(n13404), .IN2(n13416), .QN(n13413) );
  NOR2X0 U13186 ( .IN1(n13417), .IN2(n13403), .QN(n13404) );
  NOR2X0 U13187 ( .IN1(n13417), .IN2(n13418), .QN(n13403) );
  INVX0 U13188 ( .INP(n13419), .ZN(n13418) );
  NAND2X0 U13189 ( .IN1(n3036), .IN2(n13420), .QN(n13419) );
  NAND2X0 U13190 ( .IN1(n13421), .IN2(n13422), .QN(n13420) );
  NOR2X0 U13191 ( .IN1(n12475), .IN2(n12487), .QN(n13422) );
  NOR2X0 U13192 ( .IN1(n13423), .IN2(n12564), .QN(n13421) );
  NAND2X0 U13193 ( .IN1(n12502), .IN2(n12488), .QN(n12564) );
  NAND2X0 U13194 ( .IN1(n3038), .IN2(n13424), .QN(n12488) );
  NAND2X0 U13195 ( .IN1(n13425), .IN2(n13426), .QN(n13424) );
  NAND2X0 U13196 ( .IN1(n13427), .IN2(n13428), .QN(n13426) );
  NOR2X0 U13197 ( .IN1(n13429), .IN2(n13430), .QN(n13427) );
  NOR2X0 U13198 ( .IN1(n13431), .IN2(n13432), .QN(n13430) );
  NOR2X0 U13199 ( .IN1(n13433), .IN2(n13434), .QN(n13429) );
  NOR2X0 U13200 ( .IN1(n13435), .IN2(n13436), .QN(n13425) );
  NOR2X0 U13201 ( .IN1(n13437), .IN2(n13438), .QN(n13436) );
  NAND2X0 U13202 ( .IN1(n13439), .IN2(n13440), .QN(n13438) );
  NAND2X0 U13203 ( .IN1(n13441), .IN2(n13442), .QN(n13440) );
  NAND2X0 U13204 ( .IN1(n13443), .IN2(n13444), .QN(n13439) );
  NOR2X0 U13205 ( .IN1(n13443), .IN2(n13445), .QN(n13435) );
  NAND2X0 U13206 ( .IN1(n13446), .IN2(n13447), .QN(n13445) );
  NAND2X0 U13207 ( .IN1(n13442), .IN2(n13437), .QN(n13447) );
  INVX0 U13208 ( .INP(n13431), .ZN(n13437) );
  INVX0 U13209 ( .INP(n13433), .ZN(n13442) );
  NAND2X0 U13210 ( .IN1(n13441), .IN2(n13444), .QN(n13446) );
  NAND2X0 U13211 ( .IN1(n3038), .IN2(n12484), .QN(n12502) );
  NAND2X0 U13212 ( .IN1(n13448), .IN2(n13449), .QN(n12484) );
  NAND2X0 U13213 ( .IN1(n13450), .IN2(n13451), .QN(n13449) );
  NOR2X0 U13214 ( .IN1(n13452), .IN2(n13453), .QN(n13450) );
  NOR2X0 U13215 ( .IN1(n13454), .IN2(n13455), .QN(n13453) );
  NOR2X0 U13216 ( .IN1(n13456), .IN2(n13457), .QN(n13452) );
  NOR2X0 U13217 ( .IN1(n13458), .IN2(n13459), .QN(n13448) );
  NOR2X0 U13218 ( .IN1(n13460), .IN2(n13461), .QN(n13459) );
  NAND2X0 U13219 ( .IN1(n13462), .IN2(n13463), .QN(n13461) );
  NAND2X0 U13220 ( .IN1(n13464), .IN2(n13465), .QN(n13463) );
  NAND2X0 U13221 ( .IN1(n13466), .IN2(n13467), .QN(n13462) );
  NOR2X0 U13222 ( .IN1(n13464), .IN2(n13468), .QN(n13458) );
  NAND2X0 U13223 ( .IN1(n13469), .IN2(n13470), .QN(n13468) );
  NAND2X0 U13224 ( .IN1(n13466), .IN2(n13460), .QN(n13470) );
  NAND2X0 U13225 ( .IN1(n13467), .IN2(n13465), .QN(n13469) );
  INVX0 U13226 ( .INP(n13456), .ZN(n13465) );
  INVX0 U13227 ( .INP(n13451), .ZN(n13467) );
  NAND2X0 U13228 ( .IN1(n12932), .IN2(n12934), .QN(n3036) );
  INVX0 U13229 ( .INP(n13423), .ZN(n12934) );
  NOR2X0 U13230 ( .IN1(n13471), .IN2(n13472), .QN(n13417) );
  NOR2X0 U13231 ( .IN1(n12569), .IN2(n12932), .QN(n13472) );
  NAND2X0 U13232 ( .IN1(n12489), .IN2(n3038), .QN(n12569) );
  NAND2X0 U13233 ( .IN1(n13473), .IN2(n13474), .QN(n12489) );
  NOR2X0 U13234 ( .IN1(n13475), .IN2(n13476), .QN(n13474) );
  NAND2X0 U13235 ( .IN1(n13443), .IN2(n13441), .QN(n13476) );
  INVX0 U13236 ( .INP(n13428), .ZN(n13441) );
  NAND2X0 U13237 ( .IN1(n13477), .IN2(n13478), .QN(n13428) );
  NAND2X0 U13238 ( .IN1(n4555), .IN2(n10994), .QN(n13478) );
  NAND2X0 U13239 ( .IN1(n10995), .IN2(g2190), .QN(n13477) );
  INVX0 U13240 ( .INP(n10994), .ZN(n10995) );
  NAND2X0 U13241 ( .IN1(n13479), .IN2(n13480), .QN(n10994) );
  NAND2X0 U13242 ( .IN1(test_so77), .IN2(test_so73), .QN(n13480) );
  NOR2X0 U13243 ( .IN1(n13481), .IN2(n13482), .QN(n13479) );
  NOR2X0 U13244 ( .IN1(n9459), .IN2(n4367), .QN(n13482) );
  NOR2X0 U13245 ( .IN1(n9475), .IN2(n4324), .QN(n13481) );
  INVX0 U13246 ( .INP(n13434), .ZN(n13443) );
  NAND2X0 U13247 ( .IN1(n13483), .IN2(n13484), .QN(n13434) );
  NAND2X0 U13248 ( .IN1(n10987), .IN2(n13485), .QN(n13484) );
  INVX0 U13249 ( .INP(n10986), .ZN(n10987) );
  NAND2X0 U13250 ( .IN1(n12088), .IN2(n10986), .QN(n13483) );
  NAND2X0 U13251 ( .IN1(n13486), .IN2(n13487), .QN(n10986) );
  NAND2X0 U13252 ( .IN1(test_so73), .IN2(g2345), .QN(n13487) );
  NOR2X0 U13253 ( .IN1(n13488), .IN2(n13489), .QN(n13486) );
  NOR2X0 U13254 ( .IN1(n9417), .IN2(n4367), .QN(n13489) );
  NOR2X0 U13255 ( .IN1(n9418), .IN2(n4324), .QN(n13488) );
  NAND2X0 U13256 ( .IN1(n13490), .IN2(n13444), .QN(n13475) );
  INVX0 U13257 ( .INP(n13432), .ZN(n13444) );
  NAND2X0 U13258 ( .IN1(n13491), .IN2(n13492), .QN(n13432) );
  NAND2X0 U13259 ( .IN1(n4287), .IN2(n10949), .QN(n13492) );
  NAND2X0 U13260 ( .IN1(n10950), .IN2(g2200), .QN(n13491) );
  INVX0 U13261 ( .INP(n10949), .ZN(n10950) );
  NAND2X0 U13262 ( .IN1(n13493), .IN2(n13494), .QN(n10949) );
  NAND2X0 U13263 ( .IN1(test_so73), .IN2(g2336), .QN(n13494) );
  NOR2X0 U13264 ( .IN1(n13495), .IN2(n13496), .QN(n13493) );
  NOR2X0 U13265 ( .IN1(n9568), .IN2(n4367), .QN(n13496) );
  NOR2X0 U13266 ( .IN1(n9472), .IN2(n4324), .QN(n13495) );
  NOR2X0 U13267 ( .IN1(n13431), .IN2(n13433), .QN(n13490) );
  NAND2X0 U13268 ( .IN1(n13497), .IN2(n13498), .QN(n13433) );
  NAND2X0 U13269 ( .IN1(n4389), .IN2(n10990), .QN(n13498) );
  NAND2X0 U13270 ( .IN1(n10991), .IN2(g2180), .QN(n13497) );
  INVX0 U13271 ( .INP(n10990), .ZN(n10991) );
  NAND2X0 U13272 ( .IN1(n13499), .IN2(n13500), .QN(n10990) );
  NAND2X0 U13273 ( .IN1(test_so73), .IN2(g2318), .QN(n13500) );
  NOR2X0 U13274 ( .IN1(n13501), .IN2(n13502), .QN(n13499) );
  NOR2X0 U13275 ( .IN1(n9460), .IN2(n4367), .QN(n13502) );
  NOR2X0 U13276 ( .IN1(n9478), .IN2(n4324), .QN(n13501) );
  NAND2X0 U13277 ( .IN1(n13503), .IN2(n13504), .QN(n13431) );
  NAND2X0 U13278 ( .IN1(n4373), .IN2(n10978), .QN(n13504) );
  NAND2X0 U13279 ( .IN1(n12265), .IN2(g2170), .QN(n13503) );
  INVX0 U13280 ( .INP(n10978), .ZN(n12265) );
  NAND2X0 U13281 ( .IN1(n13505), .IN2(n13506), .QN(n10978) );
  NAND2X0 U13282 ( .IN1(test_so73), .IN2(g2309), .QN(n13506) );
  NOR2X0 U13283 ( .IN1(n13507), .IN2(n13508), .QN(n13505) );
  NOR2X0 U13284 ( .IN1(n9461), .IN2(n4367), .QN(n13508) );
  NOR2X0 U13285 ( .IN1(n9481), .IN2(n4324), .QN(n13507) );
  NOR2X0 U13286 ( .IN1(n13509), .IN2(n13510), .QN(n13473) );
  NAND2X0 U13287 ( .IN1(n13464), .IN2(n13466), .QN(n13510) );
  INVX0 U13288 ( .INP(n13454), .ZN(n13466) );
  NAND2X0 U13289 ( .IN1(n13511), .IN2(n13512), .QN(n13454) );
  NAND2X0 U13290 ( .IN1(n4319), .IN2(n10961), .QN(n13512) );
  NAND2X0 U13291 ( .IN1(n10962), .IN2(g2175), .QN(n13511) );
  INVX0 U13292 ( .INP(n10961), .ZN(n10962) );
  NAND2X0 U13293 ( .IN1(n13513), .IN2(n13514), .QN(n10961) );
  NAND2X0 U13294 ( .IN1(test_so73), .IN2(g2273), .QN(n13514) );
  NOR2X0 U13295 ( .IN1(n13515), .IN2(n13516), .QN(n13513) );
  NOR2X0 U13296 ( .IN1(n9577), .IN2(n4367), .QN(n13516) );
  NOR2X0 U13297 ( .IN1(n9480), .IN2(n4324), .QN(n13515) );
  INVX0 U13298 ( .INP(n13455), .ZN(n13464) );
  NAND2X0 U13299 ( .IN1(n13517), .IN2(n13518), .QN(n13455) );
  NAND2X0 U13300 ( .IN1(n10966), .IN2(n12307), .QN(n13518) );
  INVX0 U13301 ( .INP(n10965), .ZN(n10966) );
  NAND2X0 U13302 ( .IN1(n13519), .IN2(n10965), .QN(n13517) );
  NAND2X0 U13303 ( .IN1(n13520), .IN2(n13521), .QN(n10965) );
  NAND2X0 U13304 ( .IN1(test_so73), .IN2(g2300), .QN(n13521) );
  NOR2X0 U13305 ( .IN1(n13522), .IN2(n13523), .QN(n13520) );
  NOR2X0 U13306 ( .IN1(n9425), .IN2(n4367), .QN(n13523) );
  NOR2X0 U13307 ( .IN1(n9419), .IN2(n4324), .QN(n13522) );
  NAND2X0 U13308 ( .IN1(n13524), .IN2(n13460), .QN(n13509) );
  INVX0 U13309 ( .INP(n13457), .ZN(n13460) );
  NAND2X0 U13310 ( .IN1(n13525), .IN2(n13526), .QN(n13457) );
  NAND2X0 U13311 ( .IN1(n4377), .IN2(n10953), .QN(n13526) );
  NAND2X0 U13312 ( .IN1(n10954), .IN2(g2165), .QN(n13525) );
  INVX0 U13313 ( .INP(n10953), .ZN(n10954) );
  NAND2X0 U13314 ( .IN1(n13527), .IN2(n13528), .QN(n10953) );
  NAND2X0 U13315 ( .IN1(test_so76), .IN2(test_so73), .QN(n13528) );
  NOR2X0 U13316 ( .IN1(n13529), .IN2(n13530), .QN(n13527) );
  NOR2X0 U13317 ( .IN1(n9578), .IN2(n4367), .QN(n13530) );
  NOR2X0 U13318 ( .IN1(n9482), .IN2(n4324), .QN(n13529) );
  NOR2X0 U13319 ( .IN1(n13456), .IN2(n13451), .QN(n13524) );
  NAND2X0 U13320 ( .IN1(n13531), .IN2(n13532), .QN(n13451) );
  NAND2X0 U13321 ( .IN1(n4325), .IN2(n10969), .QN(n13532) );
  NAND2X0 U13322 ( .IN1(n10970), .IN2(g2185), .QN(n13531) );
  INVX0 U13323 ( .INP(n10969), .ZN(n10970) );
  NAND2X0 U13324 ( .IN1(n13533), .IN2(n13534), .QN(n10969) );
  NAND2X0 U13325 ( .IN1(test_so73), .IN2(g2282), .QN(n13534) );
  NOR2X0 U13326 ( .IN1(n13535), .IN2(n13536), .QN(n13533) );
  NOR2X0 U13327 ( .IN1(n9571), .IN2(n4367), .QN(n13536) );
  NOR2X0 U13328 ( .IN1(n9477), .IN2(n4324), .QN(n13535) );
  NAND2X0 U13329 ( .IN1(n13537), .IN2(n13538), .QN(n13456) );
  NAND2X0 U13330 ( .IN1(n4563), .IN2(n10945), .QN(n13538) );
  NAND2X0 U13331 ( .IN1(n10946), .IN2(g2195), .QN(n13537) );
  INVX0 U13332 ( .INP(n10945), .ZN(n10946) );
  NAND2X0 U13333 ( .IN1(n13539), .IN2(n13540), .QN(n10945) );
  NAND2X0 U13334 ( .IN1(test_so73), .IN2(g2291), .QN(n13540) );
  NOR2X0 U13335 ( .IN1(n13541), .IN2(n13542), .QN(n13539) );
  NOR2X0 U13336 ( .IN1(n9576), .IN2(n4367), .QN(n13542) );
  NOR2X0 U13337 ( .IN1(n9474), .IN2(n4324), .QN(n13541) );
  INVX0 U13338 ( .INP(n13543), .ZN(n13471) );
  NAND2X0 U13339 ( .IN1(n12932), .IN2(test_so79), .QN(n13543) );
  NAND2X0 U13340 ( .IN1(n13544), .IN2(n13545), .QN(g29181) );
  NAND2X0 U13341 ( .IN1(n13546), .IN2(g1704), .QN(n13545) );
  NAND2X0 U13342 ( .IN1(n13411), .IN2(n11946), .QN(n13546) );
  NAND2X0 U13343 ( .IN1(n13412), .IN2(n11946), .QN(n13544) );
  NAND2X0 U13344 ( .IN1(n13547), .IN2(n13548), .QN(g29179) );
  NAND2X0 U13345 ( .IN1(n13549), .IN2(g1008), .QN(n13548) );
  NAND2X0 U13346 ( .IN1(n13550), .IN2(g1088), .QN(n13549) );
  NAND2X0 U13347 ( .IN1(n13551), .IN2(g1088), .QN(n13547) );
  NAND2X0 U13348 ( .IN1(n13552), .IN2(n13553), .QN(g29178) );
  NAND2X0 U13349 ( .IN1(n13554), .IN2(g1703), .QN(n13553) );
  NAND2X0 U13350 ( .IN1(n13411), .IN2(n13555), .QN(n13554) );
  NAND2X0 U13351 ( .IN1(n13412), .IN2(n13555), .QN(n13552) );
  NOR2X0 U13352 ( .IN1(n13556), .IN2(n13411), .QN(n13412) );
  INVX0 U13353 ( .INP(n13557), .ZN(n13411) );
  NAND2X0 U13354 ( .IN1(n13558), .IN2(n13559), .QN(n13557) );
  NAND2X0 U13355 ( .IN1(n3068), .IN2(n13560), .QN(n13559) );
  NAND2X0 U13356 ( .IN1(n13561), .IN2(n13562), .QN(n13560) );
  NOR2X0 U13357 ( .IN1(n11961), .IN2(n11975), .QN(n13562) );
  NOR2X0 U13358 ( .IN1(n13001), .IN2(n12585), .QN(n13561) );
  NAND2X0 U13359 ( .IN1(n11990), .IN2(n11988), .QN(n12585) );
  NAND2X0 U13360 ( .IN1(n3070), .IN2(n11973), .QN(n11988) );
  NAND2X0 U13361 ( .IN1(n13563), .IN2(n13564), .QN(n11973) );
  NAND2X0 U13362 ( .IN1(n13565), .IN2(n13566), .QN(n13564) );
  NOR2X0 U13363 ( .IN1(n13567), .IN2(n13568), .QN(n13565) );
  NOR2X0 U13364 ( .IN1(n13569), .IN2(n13570), .QN(n13567) );
  NOR2X0 U13365 ( .IN1(n13571), .IN2(n13572), .QN(n13563) );
  NOR2X0 U13366 ( .IN1(n13573), .IN2(n13574), .QN(n13572) );
  NAND2X0 U13367 ( .IN1(n13575), .IN2(n13576), .QN(n13574) );
  NAND2X0 U13368 ( .IN1(n13577), .IN2(n13578), .QN(n13576) );
  NAND2X0 U13369 ( .IN1(n13579), .IN2(n13580), .QN(n13575) );
  NOR2X0 U13370 ( .IN1(n13579), .IN2(n13581), .QN(n13571) );
  NAND2X0 U13371 ( .IN1(n13582), .IN2(n13583), .QN(n13581) );
  NAND2X0 U13372 ( .IN1(n13578), .IN2(n13573), .QN(n13583) );
  INVX0 U13373 ( .INP(n13584), .ZN(n13573) );
  NAND2X0 U13374 ( .IN1(n13577), .IN2(n13580), .QN(n13582) );
  INVX0 U13375 ( .INP(n13585), .ZN(n13580) );
  NAND2X0 U13376 ( .IN1(n3070), .IN2(n11976), .QN(n11990) );
  NAND2X0 U13377 ( .IN1(n13586), .IN2(n13587), .QN(n11976) );
  NAND2X0 U13378 ( .IN1(n13588), .IN2(n13589), .QN(n13587) );
  NOR2X0 U13379 ( .IN1(n13590), .IN2(n13591), .QN(n13588) );
  NOR2X0 U13380 ( .IN1(n13592), .IN2(n13593), .QN(n13591) );
  NOR2X0 U13381 ( .IN1(n13594), .IN2(n13595), .QN(n13590) );
  NOR2X0 U13382 ( .IN1(n13596), .IN2(n13597), .QN(n13586) );
  NOR2X0 U13383 ( .IN1(n13598), .IN2(n13599), .QN(n13597) );
  NAND2X0 U13384 ( .IN1(n13600), .IN2(n13601), .QN(n13599) );
  NAND2X0 U13385 ( .IN1(n13602), .IN2(n13603), .QN(n13601) );
  NAND2X0 U13386 ( .IN1(n13604), .IN2(n13605), .QN(n13600) );
  NOR2X0 U13387 ( .IN1(n13602), .IN2(n13606), .QN(n13596) );
  NAND2X0 U13388 ( .IN1(n13607), .IN2(n13608), .QN(n13606) );
  NAND2X0 U13389 ( .IN1(n13604), .IN2(n13598), .QN(n13608) );
  NAND2X0 U13390 ( .IN1(n13605), .IN2(n13603), .QN(n13607) );
  INVX0 U13391 ( .INP(n13594), .ZN(n13603) );
  INVX0 U13392 ( .INP(n13589), .ZN(n13605) );
  INVX0 U13393 ( .INP(n12996), .ZN(n3068) );
  NOR2X0 U13394 ( .IN1(n13609), .IN2(n13001), .QN(n12996) );
  INVX0 U13395 ( .INP(n13558), .ZN(n13556) );
  NAND2X0 U13396 ( .IN1(n13610), .IN2(n13611), .QN(n13558) );
  NAND2X0 U13397 ( .IN1(n13234), .IN2(g1690), .QN(n13611) );
  NAND2X0 U13398 ( .IN1(n13612), .IN2(n13609), .QN(n13610) );
  NOR2X0 U13399 ( .IN1(n11974), .IN2(n13613), .QN(n13612) );
  INVX0 U13400 ( .INP(n12592), .ZN(n11974) );
  NAND2X0 U13401 ( .IN1(n13614), .IN2(n13615), .QN(n12592) );
  NOR2X0 U13402 ( .IN1(n13616), .IN2(n13617), .QN(n13615) );
  NAND2X0 U13403 ( .IN1(n13579), .IN2(n13577), .QN(n13617) );
  INVX0 U13404 ( .INP(n13566), .ZN(n13577) );
  NAND2X0 U13405 ( .IN1(n13618), .IN2(n13619), .QN(n13566) );
  NAND2X0 U13406 ( .IN1(n4557), .IN2(n10925), .QN(n13619) );
  NAND2X0 U13407 ( .IN1(n10926), .IN2(g1496), .QN(n13618) );
  INVX0 U13408 ( .INP(n10925), .ZN(n10926) );
  NAND2X0 U13409 ( .IN1(n13620), .IN2(n13621), .QN(n10925) );
  NAND2X0 U13410 ( .IN1(g6782), .IN2(g1633), .QN(n13621) );
  NOR2X0 U13411 ( .IN1(n13622), .IN2(n13623), .QN(n13620) );
  NOR2X0 U13412 ( .IN1(n9462), .IN2(n4368), .QN(n13623) );
  NOR2X0 U13413 ( .IN1(n9488), .IN2(n4317), .QN(n13622) );
  INVX0 U13414 ( .INP(n13570), .ZN(n13579) );
  NAND2X0 U13415 ( .IN1(n13624), .IN2(n13625), .QN(n13570) );
  NAND2X0 U13416 ( .IN1(n10930), .IN2(n13626), .QN(n13625) );
  INVX0 U13417 ( .INP(n10929), .ZN(n10930) );
  NAND2X0 U13418 ( .IN1(n12132), .IN2(n10929), .QN(n13624) );
  NAND2X0 U13419 ( .IN1(n13627), .IN2(n13628), .QN(n10929) );
  NAND2X0 U13420 ( .IN1(g6782), .IN2(g1651), .QN(n13628) );
  NOR2X0 U13421 ( .IN1(n13629), .IN2(n13630), .QN(n13627) );
  NOR2X0 U13422 ( .IN1(n9454), .IN2(n4368), .QN(n13630) );
  NOR2X0 U13423 ( .IN1(n9453), .IN2(n4317), .QN(n13629) );
  NAND2X0 U13424 ( .IN1(n13568), .IN2(n13578), .QN(n13616) );
  INVX0 U13425 ( .INP(n13569), .ZN(n13578) );
  NAND2X0 U13426 ( .IN1(n13631), .IN2(n13632), .QN(n13569) );
  NAND2X0 U13427 ( .IN1(n4390), .IN2(n10913), .QN(n13632) );
  NAND2X0 U13428 ( .IN1(n10914), .IN2(g1486), .QN(n13631) );
  INVX0 U13429 ( .INP(n10913), .ZN(n10914) );
  NAND2X0 U13430 ( .IN1(n13633), .IN2(n13634), .QN(n10913) );
  NAND2X0 U13431 ( .IN1(g6782), .IN2(g1624), .QN(n13634) );
  NOR2X0 U13432 ( .IN1(n13635), .IN2(n13636), .QN(n13633) );
  NOR2X0 U13433 ( .IN1(n9463), .IN2(n4368), .QN(n13636) );
  INVX0 U13434 ( .INP(n13637), .ZN(n13635) );
  NAND2X0 U13435 ( .IN1(g6573), .IN2(test_so55), .QN(n13637) );
  NOR2X0 U13436 ( .IN1(n13585), .IN2(n13584), .QN(n13568) );
  NAND2X0 U13437 ( .IN1(n13638), .IN2(n13639), .QN(n13584) );
  NAND2X0 U13438 ( .IN1(n4374), .IN2(n10921), .QN(n13639) );
  NAND2X0 U13439 ( .IN1(n10922), .IN2(g1476), .QN(n13638) );
  INVX0 U13440 ( .INP(n10921), .ZN(n10922) );
  NAND2X0 U13441 ( .IN1(n13640), .IN2(n13641), .QN(n10921) );
  NAND2X0 U13442 ( .IN1(g6782), .IN2(g1615), .QN(n13641) );
  NOR2X0 U13443 ( .IN1(n13642), .IN2(n13643), .QN(n13640) );
  NOR2X0 U13444 ( .IN1(n9464), .IN2(n4368), .QN(n13643) );
  NOR2X0 U13445 ( .IN1(n9493), .IN2(n4317), .QN(n13642) );
  NAND2X0 U13446 ( .IN1(n13644), .IN2(n13645), .QN(n13585) );
  NAND2X0 U13447 ( .IN1(n4288), .IN2(n10884), .QN(n13645) );
  NAND2X0 U13448 ( .IN1(n10885), .IN2(g1506), .QN(n13644) );
  INVX0 U13449 ( .INP(n10884), .ZN(n10885) );
  NAND2X0 U13450 ( .IN1(n13646), .IN2(n13647), .QN(n10884) );
  NAND2X0 U13451 ( .IN1(g6782), .IN2(g1642), .QN(n13647) );
  NOR2X0 U13452 ( .IN1(n13648), .IN2(n13649), .QN(n13646) );
  NOR2X0 U13453 ( .IN1(n9569), .IN2(n4368), .QN(n13649) );
  NOR2X0 U13454 ( .IN1(n9484), .IN2(n4317), .QN(n13648) );
  NOR2X0 U13455 ( .IN1(n13650), .IN2(n13651), .QN(n13614) );
  NAND2X0 U13456 ( .IN1(n13602), .IN2(n13604), .QN(n13651) );
  INVX0 U13457 ( .INP(n13592), .ZN(n13604) );
  NAND2X0 U13458 ( .IN1(n13652), .IN2(n13653), .QN(n13592) );
  NAND2X0 U13459 ( .IN1(n4320), .IN2(n10896), .QN(n13653) );
  NAND2X0 U13460 ( .IN1(n10897), .IN2(g1481), .QN(n13652) );
  INVX0 U13461 ( .INP(n10896), .ZN(n10897) );
  NAND2X0 U13462 ( .IN1(n13654), .IN2(n13655), .QN(n10896) );
  NAND2X0 U13463 ( .IN1(g6782), .IN2(g1579), .QN(n13655) );
  NOR2X0 U13464 ( .IN1(n13656), .IN2(n13657), .QN(n13654) );
  NOR2X0 U13465 ( .IN1(n9580), .IN2(n4368), .QN(n13657) );
  NOR2X0 U13466 ( .IN1(n9492), .IN2(n4317), .QN(n13656) );
  INVX0 U13467 ( .INP(n13593), .ZN(n13602) );
  NAND2X0 U13468 ( .IN1(n13658), .IN2(n13659), .QN(n13593) );
  NAND2X0 U13469 ( .IN1(n10901), .IN2(n13660), .QN(n13659) );
  INVX0 U13470 ( .INP(n10900), .ZN(n10901) );
  NAND2X0 U13471 ( .IN1(n12365), .IN2(n10900), .QN(n13658) );
  NAND2X0 U13472 ( .IN1(n13661), .IN2(n13662), .QN(n10900) );
  NAND2X0 U13473 ( .IN1(test_so56), .IN2(g6782), .QN(n13662) );
  NOR2X0 U13474 ( .IN1(n13663), .IN2(n13664), .QN(n13661) );
  NOR2X0 U13475 ( .IN1(n9426), .IN2(n4368), .QN(n13664) );
  NOR2X0 U13476 ( .IN1(n9420), .IN2(n4317), .QN(n13663) );
  NAND2X0 U13477 ( .IN1(n13665), .IN2(n13598), .QN(n13650) );
  INVX0 U13478 ( .INP(n13595), .ZN(n13598) );
  NAND2X0 U13479 ( .IN1(n13666), .IN2(n13667), .QN(n13595) );
  NAND2X0 U13480 ( .IN1(n4378), .IN2(n10888), .QN(n13667) );
  NAND2X0 U13481 ( .IN1(n10889), .IN2(g1471), .QN(n13666) );
  INVX0 U13482 ( .INP(n10888), .ZN(n10889) );
  NAND2X0 U13483 ( .IN1(n13668), .IN2(n13669), .QN(n10888) );
  NAND2X0 U13484 ( .IN1(g6782), .IN2(g1570), .QN(n13669) );
  NOR2X0 U13485 ( .IN1(n13670), .IN2(n13671), .QN(n13668) );
  NOR2X0 U13486 ( .IN1(n9581), .IN2(n4368), .QN(n13671) );
  NOR2X0 U13487 ( .IN1(n9495), .IN2(n4317), .QN(n13670) );
  NOR2X0 U13488 ( .IN1(n13594), .IN2(n13589), .QN(n13665) );
  NAND2X0 U13489 ( .IN1(n13672), .IN2(n13673), .QN(n13589) );
  NAND2X0 U13490 ( .IN1(n4326), .IN2(n10904), .QN(n13673) );
  NAND2X0 U13491 ( .IN1(n10905), .IN2(g1491), .QN(n13672) );
  INVX0 U13492 ( .INP(n10904), .ZN(n10905) );
  NAND2X0 U13493 ( .IN1(n13674), .IN2(n13675), .QN(n10904) );
  NAND2X0 U13494 ( .IN1(g6782), .IN2(g1588), .QN(n13675) );
  NOR2X0 U13495 ( .IN1(n13676), .IN2(n13677), .QN(n13674) );
  NOR2X0 U13496 ( .IN1(n9572), .IN2(n4368), .QN(n13677) );
  NOR2X0 U13497 ( .IN1(n9490), .IN2(n4317), .QN(n13676) );
  NAND2X0 U13498 ( .IN1(n13678), .IN2(n13679), .QN(n13594) );
  NAND2X0 U13499 ( .IN1(n4565), .IN2(n10880), .QN(n13679) );
  NAND2X0 U13500 ( .IN1(n10881), .IN2(g1501), .QN(n13678) );
  INVX0 U13501 ( .INP(n10880), .ZN(n10881) );
  NAND2X0 U13502 ( .IN1(n13680), .IN2(n13681), .QN(n10880) );
  NAND2X0 U13503 ( .IN1(g6782), .IN2(g1597), .QN(n13681) );
  NOR2X0 U13504 ( .IN1(n13682), .IN2(n13683), .QN(n13680) );
  NOR2X0 U13505 ( .IN1(n9579), .IN2(n4368), .QN(n13683) );
  NOR2X0 U13506 ( .IN1(n9486), .IN2(n4317), .QN(n13682) );
  NAND2X0 U13507 ( .IN1(n13684), .IN2(n13685), .QN(g29173) );
  NAND2X0 U13508 ( .IN1(n13686), .IN2(g1010), .QN(n13685) );
  NAND2X0 U13509 ( .IN1(n13550), .IN2(g6712), .QN(n13686) );
  NAND2X0 U13510 ( .IN1(n13551), .IN2(g6712), .QN(n13684) );
  NAND2X0 U13511 ( .IN1(n13687), .IN2(n13688), .QN(g29172) );
  NAND2X0 U13512 ( .IN1(n13689), .IN2(g321), .QN(n13688) );
  NAND2X0 U13513 ( .IN1(n13690), .IN2(n13361), .QN(n13689) );
  NAND2X0 U13514 ( .IN1(n13691), .IN2(n13361), .QN(n13687) );
  NAND2X0 U13515 ( .IN1(n13692), .IN2(n13693), .QN(g29170) );
  NAND2X0 U13516 ( .IN1(n13694), .IN2(g1009), .QN(n13693) );
  NAND2X0 U13517 ( .IN1(n13550), .IN2(g5472), .QN(n13694) );
  NAND2X0 U13518 ( .IN1(n13551), .IN2(g5472), .QN(n13692) );
  NOR2X0 U13519 ( .IN1(n13695), .IN2(n13550), .QN(n13551) );
  INVX0 U13520 ( .INP(n145), .ZN(n13550) );
  NAND2X0 U13521 ( .IN1(n13696), .IN2(n13067), .QN(n145) );
  NOR2X0 U13522 ( .IN1(n13697), .IN2(n13695), .QN(n13696) );
  NOR2X0 U13523 ( .IN1(n13698), .IN2(n13065), .QN(n13697) );
  NOR2X0 U13524 ( .IN1(n11765), .IN2(n13699), .QN(n13698) );
  NAND2X0 U13525 ( .IN1(n11756), .IN2(n11759), .QN(n13699) );
  NAND2X0 U13526 ( .IN1(n11801), .IN2(n11811), .QN(n11765) );
  NAND2X0 U13527 ( .IN1(n3102), .IN2(n13700), .QN(n11811) );
  NAND2X0 U13528 ( .IN1(n13701), .IN2(n13702), .QN(n13700) );
  NAND2X0 U13529 ( .IN1(n13703), .IN2(n13704), .QN(n13702) );
  NOR2X0 U13530 ( .IN1(n13705), .IN2(n13706), .QN(n13703) );
  NOR2X0 U13531 ( .IN1(n13707), .IN2(n13708), .QN(n13706) );
  NOR2X0 U13532 ( .IN1(n13709), .IN2(n13710), .QN(n13705) );
  NOR2X0 U13533 ( .IN1(n13711), .IN2(n13712), .QN(n13701) );
  NOR2X0 U13534 ( .IN1(n13713), .IN2(n13714), .QN(n13712) );
  NAND2X0 U13535 ( .IN1(n13715), .IN2(n13716), .QN(n13714) );
  NAND2X0 U13536 ( .IN1(n13717), .IN2(n13718), .QN(n13716) );
  NAND2X0 U13537 ( .IN1(n13719), .IN2(n13720), .QN(n13715) );
  NOR2X0 U13538 ( .IN1(n13717), .IN2(n13721), .QN(n13711) );
  NAND2X0 U13539 ( .IN1(n13722), .IN2(n13723), .QN(n13721) );
  NAND2X0 U13540 ( .IN1(n13719), .IN2(n13718), .QN(n13723) );
  INVX0 U13541 ( .INP(n13704), .ZN(n13719) );
  NAND2X0 U13542 ( .IN1(n13713), .IN2(n13720), .QN(n13722) );
  INVX0 U13543 ( .INP(n13709), .ZN(n13720) );
  NAND2X0 U13544 ( .IN1(n3102), .IN2(n11812), .QN(n11801) );
  NAND2X0 U13545 ( .IN1(n13724), .IN2(n13725), .QN(n11812) );
  NAND2X0 U13546 ( .IN1(n13726), .IN2(n13727), .QN(n13725) );
  NOR2X0 U13547 ( .IN1(n13728), .IN2(n13729), .QN(n13726) );
  NOR2X0 U13548 ( .IN1(n13730), .IN2(n13731), .QN(n13729) );
  NOR2X0 U13549 ( .IN1(n13732), .IN2(n13733), .QN(n13728) );
  NOR2X0 U13550 ( .IN1(n13734), .IN2(n13735), .QN(n13724) );
  NOR2X0 U13551 ( .IN1(n13736), .IN2(n13737), .QN(n13735) );
  NAND2X0 U13552 ( .IN1(n13738), .IN2(n13739), .QN(n13737) );
  NAND2X0 U13553 ( .IN1(n13740), .IN2(n13741), .QN(n13739) );
  NAND2X0 U13554 ( .IN1(n13742), .IN2(n13743), .QN(n13738) );
  NOR2X0 U13555 ( .IN1(n13742), .IN2(n13744), .QN(n13734) );
  NAND2X0 U13556 ( .IN1(n13745), .IN2(n13746), .QN(n13744) );
  NAND2X0 U13557 ( .IN1(n13740), .IN2(n13736), .QN(n13746) );
  INVX0 U13558 ( .INP(n13730), .ZN(n13736) );
  NAND2X0 U13559 ( .IN1(n13741), .IN2(n13743), .QN(n13745) );
  INVX0 U13560 ( .INP(n13727), .ZN(n13741) );
  NOR2X0 U13561 ( .IN1(n13747), .IN2(n13748), .QN(n13695) );
  NOR2X0 U13562 ( .IN1(n13749), .IN2(n4387), .QN(n13748) );
  NOR2X0 U13563 ( .IN1(n11770), .IN2(n13065), .QN(n13747) );
  NAND2X0 U13564 ( .IN1(n11798), .IN2(n3102), .QN(n11770) );
  NAND2X0 U13565 ( .IN1(n13750), .IN2(n13751), .QN(n11798) );
  NOR2X0 U13566 ( .IN1(n13752), .IN2(n13753), .QN(n13751) );
  NAND2X0 U13567 ( .IN1(n13713), .IN2(n13743), .QN(n13753) );
  INVX0 U13568 ( .INP(n13731), .ZN(n13743) );
  NAND2X0 U13569 ( .IN1(n13754), .IN2(n13755), .QN(n13731) );
  NAND2X0 U13570 ( .IN1(n4567), .IN2(n10815), .QN(n13755) );
  NAND2X0 U13571 ( .IN1(n10816), .IN2(g809), .QN(n13754) );
  INVX0 U13572 ( .INP(n10815), .ZN(n10816) );
  NAND2X0 U13573 ( .IN1(n13756), .IN2(n13757), .QN(n10815) );
  NAND2X0 U13574 ( .IN1(test_so31), .IN2(g906), .QN(n13757) );
  NOR2X0 U13575 ( .IN1(n13758), .IN2(n13759), .QN(n13756) );
  NOR2X0 U13576 ( .IN1(n9500), .IN2(n4323), .QN(n13759) );
  NOR2X0 U13577 ( .IN1(n9499), .IN2(n4312), .QN(n13758) );
  INVX0 U13578 ( .INP(n13708), .ZN(n13713) );
  NAND2X0 U13579 ( .IN1(n13760), .IN2(n13761), .QN(n13708) );
  NAND2X0 U13580 ( .IN1(n4375), .IN2(n10835), .QN(n13761) );
  NAND2X0 U13581 ( .IN1(n10836), .IN2(g789), .QN(n13760) );
  INVX0 U13582 ( .INP(n10835), .ZN(n10836) );
  NAND2X0 U13583 ( .IN1(n13762), .IN2(n13763), .QN(n10835) );
  NAND2X0 U13584 ( .IN1(test_so34), .IN2(test_so31), .QN(n13763) );
  NOR2X0 U13585 ( .IN1(n13764), .IN2(n13765), .QN(n13762) );
  NOR2X0 U13586 ( .IN1(n9508), .IN2(n4323), .QN(n13765) );
  NOR2X0 U13587 ( .IN1(n9529), .IN2(n4312), .QN(n13764) );
  NAND2X0 U13588 ( .IN1(n13766), .IN2(n13718), .QN(n13752) );
  INVX0 U13589 ( .INP(n13707), .ZN(n13718) );
  NAND2X0 U13590 ( .IN1(n13767), .IN2(n13768), .QN(n13707) );
  NAND2X0 U13591 ( .IN1(n4289), .IN2(n10848), .QN(n13768) );
  NAND2X0 U13592 ( .IN1(n12429), .IN2(g813), .QN(n13767) );
  INVX0 U13593 ( .INP(n10848), .ZN(n12429) );
  NAND2X0 U13594 ( .IN1(n13769), .IN2(n13770), .QN(n10848) );
  NAND2X0 U13595 ( .IN1(test_so31), .IN2(g951), .QN(n13770) );
  NOR2X0 U13596 ( .IN1(n13771), .IN2(n13772), .QN(n13769) );
  INVX0 U13597 ( .INP(n13773), .ZN(n13772) );
  NAND2X0 U13598 ( .IN1(g6368), .IN2(test_so35), .QN(n13773) );
  NOR2X0 U13599 ( .IN1(n9498), .IN2(n4312), .QN(n13771) );
  NOR2X0 U13600 ( .IN1(n13730), .IN2(n13709), .QN(n13766) );
  NAND2X0 U13601 ( .IN1(n13774), .IN2(n13775), .QN(n13709) );
  NAND2X0 U13602 ( .IN1(n4391), .IN2(n10839), .QN(n13775) );
  NAND2X0 U13603 ( .IN1(n10840), .IN2(g797), .QN(n13774) );
  INVX0 U13604 ( .INP(n10839), .ZN(n10840) );
  NAND2X0 U13605 ( .IN1(n13776), .IN2(n13777), .QN(n10839) );
  NAND2X0 U13606 ( .IN1(test_so31), .IN2(g933), .QN(n13777) );
  NOR2X0 U13607 ( .IN1(n13778), .IN2(n13779), .QN(n13776) );
  NOR2X0 U13608 ( .IN1(n9505), .IN2(n4323), .QN(n13779) );
  NOR2X0 U13609 ( .IN1(n9528), .IN2(n4312), .QN(n13778) );
  NAND2X0 U13610 ( .IN1(n13780), .IN2(n13781), .QN(n13730) );
  NAND2X0 U13611 ( .IN1(n4379), .IN2(n10831), .QN(n13781) );
  NAND2X0 U13612 ( .IN1(n10832), .IN2(g785), .QN(n13780) );
  INVX0 U13613 ( .INP(n10831), .ZN(n10832) );
  NAND2X0 U13614 ( .IN1(n13782), .IN2(n13783), .QN(n10831) );
  NAND2X0 U13615 ( .IN1(test_so31), .IN2(g879), .QN(n13783) );
  NOR2X0 U13616 ( .IN1(n13784), .IN2(n13785), .QN(n13782) );
  NOR2X0 U13617 ( .IN1(n9510), .IN2(n4323), .QN(n13785) );
  NOR2X0 U13618 ( .IN1(n9509), .IN2(n4312), .QN(n13784) );
  NOR2X0 U13619 ( .IN1(n13786), .IN2(n13787), .QN(n13750) );
  NAND2X0 U13620 ( .IN1(n13717), .IN2(n13740), .QN(n13787) );
  INVX0 U13621 ( .INP(n13733), .ZN(n13740) );
  NAND2X0 U13622 ( .IN1(n13788), .IN2(n13789), .QN(n13733) );
  NAND2X0 U13623 ( .IN1(n4321), .IN2(n10860), .QN(n13789) );
  NAND2X0 U13624 ( .IN1(n10861), .IN2(g793), .QN(n13788) );
  INVX0 U13625 ( .INP(n10860), .ZN(n10861) );
  NAND2X0 U13626 ( .IN1(n13790), .IN2(n13791), .QN(n10860) );
  NAND2X0 U13627 ( .IN1(test_so31), .IN2(g888), .QN(n13791) );
  NOR2X0 U13628 ( .IN1(n13792), .IN2(n13793), .QN(n13790) );
  NOR2X0 U13629 ( .IN1(n9507), .IN2(n4323), .QN(n13793) );
  NOR2X0 U13630 ( .IN1(n9506), .IN2(n4312), .QN(n13792) );
  INVX0 U13631 ( .INP(n13710), .ZN(n13717) );
  NAND2X0 U13632 ( .IN1(n13794), .IN2(n13795), .QN(n13710) );
  NAND2X0 U13633 ( .IN1(n10857), .IN2(n13796), .QN(n13795) );
  INVX0 U13634 ( .INP(n10856), .ZN(n10857) );
  NAND2X0 U13635 ( .IN1(n12178), .IN2(n10856), .QN(n13794) );
  NAND2X0 U13636 ( .IN1(n13797), .IN2(n13798), .QN(n10856) );
  NAND2X0 U13637 ( .IN1(test_so31), .IN2(g960), .QN(n13798) );
  NOR2X0 U13638 ( .IN1(n13799), .IN2(n13800), .QN(n13797) );
  NOR2X0 U13639 ( .IN1(n9496), .IN2(n4323), .QN(n13800) );
  NOR2X0 U13640 ( .IN1(n9532), .IN2(n4312), .QN(n13799) );
  NAND2X0 U13641 ( .IN1(n13801), .IN2(n13742), .QN(n13786) );
  INVX0 U13642 ( .INP(n13732), .ZN(n13742) );
  NAND2X0 U13643 ( .IN1(n13802), .IN2(n13803), .QN(n13732) );
  NAND2X0 U13644 ( .IN1(n10865), .IN2(n12419), .QN(n13803) );
  INVX0 U13645 ( .INP(n10864), .ZN(n10865) );
  NAND2X0 U13646 ( .IN1(n13804), .IN2(n10864), .QN(n13802) );
  NAND2X0 U13647 ( .IN1(n13805), .IN2(n13806), .QN(n10864) );
  NAND2X0 U13648 ( .IN1(test_so31), .IN2(g915), .QN(n13806) );
  NOR2X0 U13649 ( .IN1(n13807), .IN2(n13808), .QN(n13805) );
  NOR2X0 U13650 ( .IN1(n9497), .IN2(n4323), .QN(n13808) );
  NOR2X0 U13651 ( .IN1(n9533), .IN2(n4312), .QN(n13807) );
  NOR2X0 U13652 ( .IN1(n13727), .IN2(n13704), .QN(n13801) );
  NAND2X0 U13653 ( .IN1(n13809), .IN2(n13810), .QN(n13704) );
  NAND2X0 U13654 ( .IN1(n4559), .IN2(n10819), .QN(n13810) );
  NAND2X0 U13655 ( .IN1(n10820), .IN2(g805), .QN(n13809) );
  INVX0 U13656 ( .INP(n10819), .ZN(n10820) );
  NAND2X0 U13657 ( .IN1(n13811), .IN2(n13812), .QN(n10819) );
  NAND2X0 U13658 ( .IN1(test_so31), .IN2(g942), .QN(n13812) );
  NOR2X0 U13659 ( .IN1(n13813), .IN2(n13814), .QN(n13811) );
  NOR2X0 U13660 ( .IN1(n9502), .IN2(n4323), .QN(n13814) );
  NOR2X0 U13661 ( .IN1(n9501), .IN2(n4312), .QN(n13813) );
  NAND2X0 U13662 ( .IN1(n13815), .IN2(n13816), .QN(n13727) );
  NAND2X0 U13663 ( .IN1(n4327), .IN2(n10823), .QN(n13816) );
  NAND2X0 U13664 ( .IN1(n10824), .IN2(g801), .QN(n13815) );
  INVX0 U13665 ( .INP(n10823), .ZN(n10824) );
  NAND2X0 U13666 ( .IN1(n13817), .IN2(n13818), .QN(n10823) );
  NAND2X0 U13667 ( .IN1(test_so31), .IN2(g897), .QN(n13818) );
  NOR2X0 U13668 ( .IN1(n13819), .IN2(n13820), .QN(n13817) );
  NOR2X0 U13669 ( .IN1(n9504), .IN2(n4323), .QN(n13820) );
  NOR2X0 U13670 ( .IN1(n9503), .IN2(n4312), .QN(n13819) );
  NAND2X0 U13671 ( .IN1(n13821), .IN2(n13822), .QN(g29169) );
  NAND2X0 U13672 ( .IN1(n13823), .IN2(g323), .QN(n13822) );
  NAND2X0 U13673 ( .IN1(n13690), .IN2(n13382), .QN(n13823) );
  NAND2X0 U13674 ( .IN1(n13691), .IN2(n13382), .QN(n13821) );
  NAND2X0 U13675 ( .IN1(n13824), .IN2(n13825), .QN(g29167) );
  NAND2X0 U13676 ( .IN1(n13826), .IN2(g322), .QN(n13825) );
  NAND2X0 U13677 ( .IN1(n13690), .IN2(n12042), .QN(n13826) );
  NAND2X0 U13678 ( .IN1(n13691), .IN2(n12042), .QN(n13824) );
  NOR2X0 U13679 ( .IN1(n13827), .IN2(n13690), .QN(n13691) );
  INVX0 U13680 ( .INP(n13828), .ZN(n13690) );
  NAND2X0 U13681 ( .IN1(n13829), .IN2(n13830), .QN(n13828) );
  NAND2X0 U13682 ( .IN1(n3128), .IN2(n13831), .QN(n13830) );
  NAND2X0 U13683 ( .IN1(n13832), .IN2(n13833), .QN(n13831) );
  NOR2X0 U13684 ( .IN1(n12011), .IN2(n12025), .QN(n13833) );
  NOR2X0 U13685 ( .IN1(n13136), .IN2(n12538), .QN(n13832) );
  NAND2X0 U13686 ( .IN1(n12040), .IN2(n12038), .QN(n12538) );
  NAND2X0 U13687 ( .IN1(n3130), .IN2(n12023), .QN(n12038) );
  NAND2X0 U13688 ( .IN1(n13834), .IN2(n13835), .QN(n12023) );
  NAND2X0 U13689 ( .IN1(n13836), .IN2(n13837), .QN(n13835) );
  NOR2X0 U13690 ( .IN1(n13838), .IN2(n13839), .QN(n13836) );
  NOR2X0 U13691 ( .IN1(n13840), .IN2(n13841), .QN(n13838) );
  NOR2X0 U13692 ( .IN1(n13842), .IN2(n13843), .QN(n13834) );
  NOR2X0 U13693 ( .IN1(n13844), .IN2(n13845), .QN(n13843) );
  NAND2X0 U13694 ( .IN1(n13846), .IN2(n13847), .QN(n13845) );
  NAND2X0 U13695 ( .IN1(n13848), .IN2(n13849), .QN(n13847) );
  NAND2X0 U13696 ( .IN1(n13850), .IN2(n13851), .QN(n13846) );
  NOR2X0 U13697 ( .IN1(n13850), .IN2(n13852), .QN(n13842) );
  NAND2X0 U13698 ( .IN1(n13853), .IN2(n13854), .QN(n13852) );
  NAND2X0 U13699 ( .IN1(n13849), .IN2(n13844), .QN(n13854) );
  INVX0 U13700 ( .INP(n13855), .ZN(n13844) );
  NAND2X0 U13701 ( .IN1(n13848), .IN2(n13851), .QN(n13853) );
  INVX0 U13702 ( .INP(n13856), .ZN(n13851) );
  NAND2X0 U13703 ( .IN1(n3130), .IN2(n12026), .QN(n12040) );
  NAND2X0 U13704 ( .IN1(n13857), .IN2(n13858), .QN(n12026) );
  NAND2X0 U13705 ( .IN1(n13859), .IN2(n13860), .QN(n13858) );
  NOR2X0 U13706 ( .IN1(n13861), .IN2(n13862), .QN(n13859) );
  NOR2X0 U13707 ( .IN1(n13863), .IN2(n13864), .QN(n13862) );
  NOR2X0 U13708 ( .IN1(n13865), .IN2(n13866), .QN(n13861) );
  NOR2X0 U13709 ( .IN1(n13867), .IN2(n13868), .QN(n13857) );
  NOR2X0 U13710 ( .IN1(n13869), .IN2(n13870), .QN(n13868) );
  NAND2X0 U13711 ( .IN1(n13871), .IN2(n13872), .QN(n13870) );
  NAND2X0 U13712 ( .IN1(n13873), .IN2(n13874), .QN(n13872) );
  NAND2X0 U13713 ( .IN1(n13875), .IN2(n13876), .QN(n13871) );
  NOR2X0 U13714 ( .IN1(n13873), .IN2(n13877), .QN(n13867) );
  NAND2X0 U13715 ( .IN1(n13878), .IN2(n13879), .QN(n13877) );
  NAND2X0 U13716 ( .IN1(n13875), .IN2(n13869), .QN(n13879) );
  NAND2X0 U13717 ( .IN1(n13876), .IN2(n13874), .QN(n13878) );
  INVX0 U13718 ( .INP(n13865), .ZN(n13874) );
  INVX0 U13719 ( .INP(n13860), .ZN(n13876) );
  INVX0 U13720 ( .INP(n13131), .ZN(n3128) );
  NOR2X0 U13721 ( .IN1(n13880), .IN2(n13136), .QN(n13131) );
  INVX0 U13722 ( .INP(n13829), .ZN(n13827) );
  NAND2X0 U13723 ( .IN1(n13881), .IN2(n13882), .QN(n13829) );
  NAND2X0 U13724 ( .IN1(n13260), .IN2(g309), .QN(n13882) );
  NAND2X0 U13725 ( .IN1(n13883), .IN2(n13880), .QN(n13881) );
  NOR2X0 U13726 ( .IN1(n12024), .IN2(n13884), .QN(n13883) );
  INVX0 U13727 ( .INP(n12545), .ZN(n12024) );
  NAND2X0 U13728 ( .IN1(n13885), .IN2(n13886), .QN(n12545) );
  NOR2X0 U13729 ( .IN1(n13887), .IN2(n13888), .QN(n13886) );
  NAND2X0 U13730 ( .IN1(n13850), .IN2(n13848), .QN(n13888) );
  INVX0 U13731 ( .INP(n13837), .ZN(n13848) );
  NAND2X0 U13732 ( .IN1(n13889), .IN2(n13890), .QN(n13837) );
  NAND2X0 U13733 ( .IN1(n4561), .IN2(n10799), .QN(n13890) );
  NAND2X0 U13734 ( .IN1(n10800), .IN2(g117), .QN(n13889) );
  INVX0 U13735 ( .INP(n10799), .ZN(n10800) );
  NAND2X0 U13736 ( .IN1(n13891), .IN2(n13892), .QN(n10799) );
  NAND2X0 U13737 ( .IN1(g6313), .IN2(g252), .QN(n13892) );
  NOR2X0 U13738 ( .IN1(n13893), .IN2(n13894), .QN(n13891) );
  INVX0 U13739 ( .INP(n13895), .ZN(n13894) );
  NAND2X0 U13740 ( .IN1(g165), .IN2(test_so14), .QN(n13895) );
  NOR2X0 U13741 ( .IN1(n9516), .IN2(n4318), .QN(n13893) );
  INVX0 U13742 ( .INP(n13841), .ZN(n13850) );
  NAND2X0 U13743 ( .IN1(n13896), .IN2(n13897), .QN(n13841) );
  NAND2X0 U13744 ( .IN1(n10793), .IN2(n13898), .QN(n13897) );
  INVX0 U13745 ( .INP(n10792), .ZN(n10793) );
  NAND2X0 U13746 ( .IN1(n12247), .IN2(n10792), .QN(n13896) );
  NAND2X0 U13747 ( .IN1(n13899), .IN2(n13900), .QN(n10792) );
  NAND2X0 U13748 ( .IN1(g6313), .IN2(g270), .QN(n13900) );
  NOR2X0 U13749 ( .IN1(n13901), .IN2(n13902), .QN(n13899) );
  NOR2X0 U13750 ( .IN1(n9457), .IN2(n4369), .QN(n13902) );
  NOR2X0 U13751 ( .IN1(n9456), .IN2(n4318), .QN(n13901) );
  NAND2X0 U13752 ( .IN1(n13839), .IN2(n13849), .QN(n13887) );
  INVX0 U13753 ( .INP(n13840), .ZN(n13849) );
  NAND2X0 U13754 ( .IN1(n13903), .IN2(n13904), .QN(n13840) );
  NAND2X0 U13755 ( .IN1(n4392), .IN2(n10784), .QN(n13904) );
  NAND2X0 U13756 ( .IN1(n12405), .IN2(g109), .QN(n13903) );
  INVX0 U13757 ( .INP(n10784), .ZN(n12405) );
  NAND2X0 U13758 ( .IN1(n13905), .IN2(n13906), .QN(n10784) );
  NAND2X0 U13759 ( .IN1(g6313), .IN2(g243), .QN(n13906) );
  NOR2X0 U13760 ( .IN1(n13907), .IN2(n13908), .QN(n13905) );
  NOR2X0 U13761 ( .IN1(n9469), .IN2(n4369), .QN(n13908) );
  NOR2X0 U13762 ( .IN1(n9519), .IN2(n4318), .QN(n13907) );
  NOR2X0 U13763 ( .IN1(n13856), .IN2(n13855), .QN(n13839) );
  NAND2X0 U13764 ( .IN1(n13909), .IN2(n13910), .QN(n13855) );
  NAND2X0 U13765 ( .IN1(n4376), .IN2(n10754), .QN(n13910) );
  NAND2X0 U13766 ( .IN1(n10755), .IN2(g101), .QN(n13909) );
  INVX0 U13767 ( .INP(n10754), .ZN(n10755) );
  NAND2X0 U13768 ( .IN1(n13911), .IN2(n13912), .QN(n10754) );
  NAND2X0 U13769 ( .IN1(g6313), .IN2(g234), .QN(n13912) );
  NOR2X0 U13770 ( .IN1(n13913), .IN2(n13914), .QN(n13911) );
  NOR2X0 U13771 ( .IN1(n9470), .IN2(n4369), .QN(n13914) );
  NOR2X0 U13772 ( .IN1(n9522), .IN2(n4318), .QN(n13913) );
  NAND2X0 U13773 ( .IN1(n13915), .IN2(n13916), .QN(n13856) );
  NAND2X0 U13774 ( .IN1(n4290), .IN2(n10758), .QN(n13916) );
  NAND2X0 U13775 ( .IN1(n10759), .IN2(g125), .QN(n13915) );
  INVX0 U13776 ( .INP(n10758), .ZN(n10759) );
  NAND2X0 U13777 ( .IN1(n13917), .IN2(n13918), .QN(n10758) );
  NAND2X0 U13778 ( .IN1(g6313), .IN2(g261), .QN(n13918) );
  NOR2X0 U13779 ( .IN1(n13919), .IN2(n13920), .QN(n13917) );
  NOR2X0 U13780 ( .IN1(n9570), .IN2(n4369), .QN(n13920) );
  NOR2X0 U13781 ( .IN1(n9512), .IN2(n4318), .QN(n13919) );
  NOR2X0 U13782 ( .IN1(n13921), .IN2(n13922), .QN(n13885) );
  NAND2X0 U13783 ( .IN1(n13873), .IN2(n13875), .QN(n13922) );
  INVX0 U13784 ( .INP(n13863), .ZN(n13875) );
  NAND2X0 U13785 ( .IN1(n13923), .IN2(n13924), .QN(n13863) );
  NAND2X0 U13786 ( .IN1(n4322), .IN2(n10766), .QN(n13924) );
  NAND2X0 U13787 ( .IN1(n10767), .IN2(g105), .QN(n13923) );
  INVX0 U13788 ( .INP(n10766), .ZN(n10767) );
  NAND2X0 U13789 ( .IN1(n13925), .IN2(n13926), .QN(n10766) );
  NAND2X0 U13790 ( .IN1(g6313), .IN2(g198), .QN(n13926) );
  NOR2X0 U13791 ( .IN1(n13927), .IN2(n13928), .QN(n13925) );
  NOR2X0 U13792 ( .IN1(n9586), .IN2(n4369), .QN(n13928) );
  NOR2X0 U13793 ( .IN1(n9521), .IN2(n4318), .QN(n13927) );
  INVX0 U13794 ( .INP(n13864), .ZN(n13873) );
  NAND2X0 U13795 ( .IN1(n13929), .IN2(n13930), .QN(n13864) );
  NAND2X0 U13796 ( .IN1(n10771), .IN2(n13931), .QN(n13930) );
  INVX0 U13797 ( .INP(n10770), .ZN(n10771) );
  NAND2X0 U13798 ( .IN1(n12454), .IN2(n10770), .QN(n13929) );
  NAND2X0 U13799 ( .IN1(n13932), .IN2(n13933), .QN(n10770) );
  NAND2X0 U13800 ( .IN1(g6313), .IN2(g225), .QN(n13933) );
  NOR2X0 U13801 ( .IN1(n13934), .IN2(n13935), .QN(n13932) );
  NOR2X0 U13802 ( .IN1(n9427), .IN2(n4369), .QN(n13935) );
  NOR2X0 U13803 ( .IN1(n9421), .IN2(n4318), .QN(n13934) );
  NAND2X0 U13804 ( .IN1(n13936), .IN2(n13869), .QN(n13921) );
  INVX0 U13805 ( .INP(n13866), .ZN(n13869) );
  NAND2X0 U13806 ( .IN1(n13937), .IN2(n13938), .QN(n13866) );
  NAND2X0 U13807 ( .IN1(n4513), .IN2(g97), .QN(n13938) );
  NAND2X0 U13808 ( .IN1(n4380), .IN2(n13127), .QN(n13937) );
  INVX0 U13809 ( .INP(n4513), .ZN(n13127) );
  NOR2X0 U13810 ( .IN1(n13865), .IN2(n13860), .QN(n13936) );
  NAND2X0 U13811 ( .IN1(n13939), .IN2(n13940), .QN(n13860) );
  NAND2X0 U13812 ( .IN1(n4328), .IN2(n10774), .QN(n13940) );
  NAND2X0 U13813 ( .IN1(n10775), .IN2(g113), .QN(n13939) );
  INVX0 U13814 ( .INP(n10774), .ZN(n10775) );
  NAND2X0 U13815 ( .IN1(n13941), .IN2(n13942), .QN(n10774) );
  NAND2X0 U13816 ( .IN1(g6313), .IN2(g207), .QN(n13942) );
  NOR2X0 U13817 ( .IN1(n13943), .IN2(n13944), .QN(n13941) );
  NOR2X0 U13818 ( .IN1(n9575), .IN2(n4369), .QN(n13944) );
  NOR2X0 U13819 ( .IN1(n9518), .IN2(n4318), .QN(n13943) );
  NAND2X0 U13820 ( .IN1(n13945), .IN2(n13946), .QN(n13865) );
  NAND2X0 U13821 ( .IN1(n4569), .IN2(n10750), .QN(n13946) );
  NAND2X0 U13822 ( .IN1(n10751), .IN2(g121), .QN(n13945) );
  INVX0 U13823 ( .INP(n10750), .ZN(n10751) );
  NAND2X0 U13824 ( .IN1(n13947), .IN2(n13948), .QN(n10750) );
  NAND2X0 U13825 ( .IN1(g6313), .IN2(g216), .QN(n13948) );
  NOR2X0 U13826 ( .IN1(n13949), .IN2(n13950), .QN(n13947) );
  NOR2X0 U13827 ( .IN1(n9585), .IN2(n4369), .QN(n13950) );
  NOR2X0 U13828 ( .IN1(n9514), .IN2(n4318), .QN(n13949) );
  NOR2X0 U13829 ( .IN1(n13951), .IN2(n13286), .QN(g29112) );
  NAND2X0 U13830 ( .IN1(n2982), .IN2(n13952), .QN(n13286) );
  NAND2X0 U13831 ( .IN1(n3159), .IN2(g2129), .QN(n2982) );
  NOR2X0 U13832 ( .IN1(n3159), .IN2(g2129), .QN(n13951) );
  NOR2X0 U13833 ( .IN1(n13953), .IN2(n13291), .QN(g29111) );
  NAND2X0 U13834 ( .IN1(n2985), .IN2(n13954), .QN(n13291) );
  NAND2X0 U13835 ( .IN1(n3163), .IN2(g1435), .QN(n2985) );
  NOR2X0 U13836 ( .IN1(n3163), .IN2(g1435), .QN(n13953) );
  NOR2X0 U13837 ( .IN1(n13955), .IN2(n13296), .QN(g29110) );
  NAND2X0 U13838 ( .IN1(n2988), .IN2(n13956), .QN(n13296) );
  NAND2X0 U13839 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NOR2X0 U13840 ( .IN1(n3167), .IN2(test_so36), .QN(n13955) );
  NOR2X0 U13841 ( .IN1(n13957), .IN2(n13301), .QN(g29109) );
  NAND2X0 U13842 ( .IN1(n2991), .IN2(n13958), .QN(n13301) );
  NAND2X0 U13843 ( .IN1(n3171), .IN2(g61), .QN(n2991) );
  NOR2X0 U13844 ( .IN1(n3171), .IN2(g61), .QN(n13957) );
  NAND2X0 U13845 ( .IN1(n13959), .IN2(n13960), .QN(g28788) );
  NAND2X0 U13846 ( .IN1(n13961), .IN2(g2501), .QN(n13960) );
  NAND2X0 U13847 ( .IN1(n13962), .IN2(n13307), .QN(n13961) );
  NAND2X0 U13848 ( .IN1(n13963), .IN2(n13307), .QN(n13959) );
  NAND2X0 U13849 ( .IN1(n13964), .IN2(n13965), .QN(g28783) );
  NAND2X0 U13850 ( .IN1(n13966), .IN2(g2503), .QN(n13965) );
  NAND2X0 U13851 ( .IN1(n13962), .IN2(n11937), .QN(n13966) );
  NAND2X0 U13852 ( .IN1(n13963), .IN2(n11937), .QN(n13964) );
  NAND2X0 U13853 ( .IN1(n13967), .IN2(n13968), .QN(g28782) );
  NAND2X0 U13854 ( .IN1(n4606), .IN2(n13969), .QN(n13968) );
  NAND2X0 U13855 ( .IN1(n4509), .IN2(test_so80), .QN(n13967) );
  NAND2X0 U13856 ( .IN1(n13970), .IN2(n13971), .QN(g28778) );
  NAND2X0 U13857 ( .IN1(n13972), .IN2(g1807), .QN(n13971) );
  NAND2X0 U13858 ( .IN1(n13973), .IN2(n13315), .QN(n13972) );
  NAND2X0 U13859 ( .IN1(n13974), .IN2(n13315), .QN(n13970) );
  NAND2X0 U13860 ( .IN1(n13975), .IN2(n13976), .QN(g28774) );
  NAND2X0 U13861 ( .IN1(n13977), .IN2(g2502), .QN(n13976) );
  NAND2X0 U13862 ( .IN1(n13962), .IN2(n13416), .QN(n13977) );
  NOR2X0 U13863 ( .IN1(n13978), .IN2(n13331), .QN(n13962) );
  NAND2X0 U13864 ( .IN1(n13963), .IN2(n13416), .QN(n13975) );
  NAND2X0 U13865 ( .IN1(n13979), .IN2(n13980), .QN(g28773) );
  NAND2X0 U13866 ( .IN1(g7264), .IN2(n13969), .QN(n13980) );
  INVX0 U13867 ( .INP(n13981), .ZN(n13979) );
  NOR2X0 U13868 ( .IN1(n11937), .IN2(n9744), .QN(n13981) );
  NAND2X0 U13869 ( .IN1(n13982), .IN2(n13983), .QN(g28772) );
  NAND2X0 U13870 ( .IN1(n13984), .IN2(g1809), .QN(n13983) );
  NAND2X0 U13871 ( .IN1(n13973), .IN2(n11946), .QN(n13984) );
  NAND2X0 U13872 ( .IN1(n13974), .IN2(n11946), .QN(n13982) );
  NAND2X0 U13873 ( .IN1(n13985), .IN2(n13986), .QN(g28771) );
  NAND2X0 U13874 ( .IN1(n4618), .IN2(n13987), .QN(n13986) );
  INVX0 U13875 ( .INP(n13988), .ZN(n13985) );
  NOR2X0 U13876 ( .IN1(n13315), .IN2(n9764), .QN(n13988) );
  NAND2X0 U13877 ( .IN1(n13989), .IN2(n13990), .QN(g28767) );
  NAND2X0 U13878 ( .IN1(n13991), .IN2(g1113), .QN(n13990) );
  NAND2X0 U13879 ( .IN1(n13992), .IN2(g1088), .QN(n13991) );
  NAND2X0 U13880 ( .IN1(n13993), .IN2(g1088), .QN(n13989) );
  NAND2X0 U13881 ( .IN1(n13994), .IN2(n13995), .QN(g28763) );
  NAND2X0 U13882 ( .IN1(g5555), .IN2(n13969), .QN(n13995) );
  NAND2X0 U13883 ( .IN1(n13996), .IN2(n13997), .QN(n13969) );
  NAND2X0 U13884 ( .IN1(n13998), .IN2(n11747), .QN(n13997) );
  NAND2X0 U13885 ( .IN1(test_so79), .IN2(n13999), .QN(n13998) );
  NAND2X0 U13886 ( .IN1(n14000), .IN2(n14001), .QN(n13999) );
  INVX0 U13887 ( .INP(n13331), .ZN(n14000) );
  NAND2X0 U13888 ( .IN1(n14002), .IN2(n14003), .QN(n13331) );
  NAND2X0 U13889 ( .IN1(n9979), .IN2(n11937), .QN(n14003) );
  NOR2X0 U13890 ( .IN1(n14004), .IN2(n14005), .QN(n14002) );
  NOR2X0 U13891 ( .IN1(n4516), .IN2(g2502), .QN(n14005) );
  NOR2X0 U13892 ( .IN1(n4509), .IN2(g2501), .QN(n14004) );
  INVX0 U13893 ( .INP(n13963), .ZN(n13996) );
  NOR2X0 U13894 ( .IN1(n13978), .IN2(n11747), .QN(n13963) );
  NAND2X0 U13895 ( .IN1(n14006), .IN2(n14007), .QN(n11747) );
  NAND2X0 U13896 ( .IN1(g5555), .IN2(g2483), .QN(n14007) );
  NOR2X0 U13897 ( .IN1(n14008), .IN2(n14009), .QN(n14006) );
  NOR2X0 U13898 ( .IN1(n9744), .IN2(n14010), .QN(n14009) );
  INVX0 U13899 ( .INP(n14011), .ZN(n14008) );
  NAND2X0 U13900 ( .IN1(n4606), .IN2(test_so80), .QN(n14011) );
  NAND2X0 U13901 ( .IN1(n14001), .IN2(test_so79), .QN(n13978) );
  NAND2X0 U13902 ( .IN1(n14012), .IN2(n14013), .QN(n14001) );
  NAND2X0 U13903 ( .IN1(n4285), .IN2(n11748), .QN(n14013) );
  NAND2X0 U13904 ( .IN1(n14014), .IN2(n13327), .QN(n14012) );
  INVX0 U13905 ( .INP(n11748), .ZN(n13327) );
  NAND2X0 U13906 ( .IN1(n14015), .IN2(n14016), .QN(n11748) );
  NOR2X0 U13907 ( .IN1(n13519), .IN2(n12088), .QN(n14015) );
  NOR2X0 U13908 ( .IN1(n12495), .IN2(n4285), .QN(n14014) );
  NOR2X0 U13909 ( .IN1(n11919), .IN2(n10029), .QN(n12495) );
  NAND2X0 U13910 ( .IN1(n14017), .IN2(n14018), .QN(n11919) );
  NAND2X0 U13911 ( .IN1(n9900), .IN2(test_so73), .QN(n14018) );
  NOR2X0 U13912 ( .IN1(n14019), .IN2(n14020), .QN(n14017) );
  NOR2X0 U13913 ( .IN1(n4367), .IN2(g2244), .QN(n14020) );
  NOR2X0 U13914 ( .IN1(n4324), .IN2(g2245), .QN(n14019) );
  NAND2X0 U13915 ( .IN1(n4516), .IN2(g2483), .QN(n13994) );
  NAND2X0 U13916 ( .IN1(n14021), .IN2(n14022), .QN(g28761) );
  NAND2X0 U13917 ( .IN1(n14023), .IN2(g1808), .QN(n14022) );
  NAND2X0 U13918 ( .IN1(n13973), .IN2(n13555), .QN(n14023) );
  NOR2X0 U13919 ( .IN1(n14024), .IN2(n13353), .QN(n13973) );
  NAND2X0 U13920 ( .IN1(n13974), .IN2(n13555), .QN(n14021) );
  NAND2X0 U13921 ( .IN1(n14025), .IN2(n14026), .QN(g28760) );
  NAND2X0 U13922 ( .IN1(g7014), .IN2(n13987), .QN(n14026) );
  INVX0 U13923 ( .INP(n14027), .ZN(n14025) );
  NOR2X0 U13924 ( .IN1(n11946), .IN2(n9748), .QN(n14027) );
  NAND2X0 U13925 ( .IN1(n14028), .IN2(n14029), .QN(g28759) );
  NAND2X0 U13926 ( .IN1(n14030), .IN2(g1115), .QN(n14029) );
  NAND2X0 U13927 ( .IN1(n13992), .IN2(g6712), .QN(n14030) );
  NAND2X0 U13928 ( .IN1(n13993), .IN2(g6712), .QN(n14028) );
  NAND2X0 U13929 ( .IN1(n14031), .IN2(n14032), .QN(g28758) );
  NAND2X0 U13930 ( .IN1(n4381), .IN2(g1101), .QN(n14032) );
  NAND2X0 U13931 ( .IN1(n14033), .IN2(g1088), .QN(n14031) );
  NAND2X0 U13932 ( .IN1(n14034), .IN2(n14035), .QN(g28754) );
  NAND2X0 U13933 ( .IN1(n14036), .IN2(g426), .QN(n14035) );
  NAND2X0 U13934 ( .IN1(n14037), .IN2(n13361), .QN(n14036) );
  NAND2X0 U13935 ( .IN1(n14038), .IN2(n13361), .QN(n14034) );
  NAND2X0 U13936 ( .IN1(n14039), .IN2(n14040), .QN(g28749) );
  NAND2X0 U13937 ( .IN1(g5511), .IN2(n13987), .QN(n14040) );
  NAND2X0 U13938 ( .IN1(n14041), .IN2(n14042), .QN(n13987) );
  NAND2X0 U13939 ( .IN1(n14043), .IN2(n11742), .QN(n14042) );
  NAND2X0 U13940 ( .IN1(g1690), .IN2(n14044), .QN(n14043) );
  NAND2X0 U13941 ( .IN1(n14045), .IN2(n14046), .QN(n14044) );
  INVX0 U13942 ( .INP(n13353), .ZN(n14045) );
  NAND2X0 U13943 ( .IN1(n14047), .IN2(n14048), .QN(n13353) );
  NAND2X0 U13944 ( .IN1(n9982), .IN2(n11946), .QN(n14048) );
  NOR2X0 U13945 ( .IN1(n14049), .IN2(n14050), .QN(n14047) );
  NOR2X0 U13946 ( .IN1(n4518), .IN2(g1808), .QN(n14050) );
  NOR2X0 U13947 ( .IN1(n4511), .IN2(g1807), .QN(n14049) );
  INVX0 U13948 ( .INP(n13974), .ZN(n14041) );
  NOR2X0 U13949 ( .IN1(n14024), .IN2(n11742), .QN(n13974) );
  NAND2X0 U13950 ( .IN1(n14051), .IN2(n14052), .QN(n11742) );
  NAND2X0 U13951 ( .IN1(g5511), .IN2(g1789), .QN(n14052) );
  NOR2X0 U13952 ( .IN1(n14053), .IN2(n14054), .QN(n14051) );
  NOR2X0 U13953 ( .IN1(n9748), .IN2(n13179), .QN(n14054) );
  NOR2X0 U13954 ( .IN1(n9764), .IN2(n14055), .QN(n14053) );
  NAND2X0 U13955 ( .IN1(g1690), .IN2(n14046), .QN(n14024) );
  NAND2X0 U13956 ( .IN1(n14056), .IN2(n14057), .QN(n14046) );
  NAND2X0 U13957 ( .IN1(n4284), .IN2(n11743), .QN(n14057) );
  NAND2X0 U13958 ( .IN1(n14058), .IN2(n13349), .QN(n14056) );
  INVX0 U13959 ( .INP(n11743), .ZN(n13349) );
  NAND2X0 U13960 ( .IN1(n14059), .IN2(n14060), .QN(n11743) );
  NOR2X0 U13961 ( .IN1(n12365), .IN2(n12132), .QN(n14059) );
  NOR2X0 U13962 ( .IN1(n11982), .IN2(n4284), .QN(n14058) );
  NOR2X0 U13963 ( .IN1(n11923), .IN2(n10030), .QN(n11982) );
  NAND2X0 U13964 ( .IN1(n14061), .IN2(n14062), .QN(n11923) );
  NAND2X0 U13965 ( .IN1(n9911), .IN2(g6782), .QN(n14062) );
  NOR2X0 U13966 ( .IN1(n14063), .IN2(n14064), .QN(n14061) );
  NOR2X0 U13967 ( .IN1(n4368), .IN2(g1550), .QN(n14064) );
  NOR2X0 U13968 ( .IN1(n4317), .IN2(g1551), .QN(n14063) );
  NAND2X0 U13969 ( .IN1(n4518), .IN2(g1789), .QN(n14039) );
  NAND2X0 U13970 ( .IN1(n14065), .IN2(n14066), .QN(g28747) );
  NAND2X0 U13971 ( .IN1(n14067), .IN2(g1114), .QN(n14066) );
  NAND2X0 U13972 ( .IN1(n13992), .IN2(g5472), .QN(n14067) );
  NOR2X0 U13973 ( .IN1(n14068), .IN2(n13378), .QN(n13992) );
  NAND2X0 U13974 ( .IN1(n13993), .IN2(g5472), .QN(n14065) );
  NAND2X0 U13975 ( .IN1(n14069), .IN2(n14070), .QN(g28746) );
  INVX0 U13976 ( .INP(n14071), .ZN(n14070) );
  NOR2X0 U13977 ( .IN1(g6712), .IN2(n9751), .QN(n14071) );
  NAND2X0 U13978 ( .IN1(n14033), .IN2(g6712), .QN(n14069) );
  NAND2X0 U13979 ( .IN1(n14072), .IN2(n14073), .QN(g28745) );
  NAND2X0 U13980 ( .IN1(n14074), .IN2(g428), .QN(n14073) );
  NAND2X0 U13981 ( .IN1(n14037), .IN2(n13382), .QN(n14074) );
  NAND2X0 U13982 ( .IN1(n14038), .IN2(n13382), .QN(n14072) );
  NAND2X0 U13983 ( .IN1(n14075), .IN2(n14076), .QN(g28744) );
  NAND2X0 U13984 ( .IN1(n4640), .IN2(n14077), .QN(n14076) );
  INVX0 U13985 ( .INP(n14078), .ZN(n14075) );
  NOR2X0 U13986 ( .IN1(n13361), .IN2(n9783), .QN(n14078) );
  NAND2X0 U13987 ( .IN1(n14079), .IN2(n14080), .QN(g28738) );
  INVX0 U13988 ( .INP(n14081), .ZN(n14080) );
  NOR2X0 U13989 ( .IN1(g5472), .IN2(n9773), .QN(n14081) );
  NAND2X0 U13990 ( .IN1(n14033), .IN2(g5472), .QN(n14079) );
  NAND2X0 U13991 ( .IN1(n14082), .IN2(n14083), .QN(n14033) );
  NAND2X0 U13992 ( .IN1(n14084), .IN2(n11737), .QN(n14083) );
  NAND2X0 U13993 ( .IN1(g996), .IN2(n14085), .QN(n14084) );
  NAND2X0 U13994 ( .IN1(n14086), .IN2(n14087), .QN(n14085) );
  INVX0 U13995 ( .INP(n13378), .ZN(n14086) );
  NAND2X0 U13996 ( .IN1(n14088), .IN2(n14089), .QN(n13378) );
  NAND2X0 U13997 ( .IN1(n9999), .IN2(g1088), .QN(n14089) );
  NOR2X0 U13998 ( .IN1(n14090), .IN2(n14091), .QN(n14088) );
  NOR2X0 U13999 ( .IN1(n4364), .IN2(g1115), .QN(n14091) );
  NOR2X0 U14000 ( .IN1(n4363), .IN2(g1114), .QN(n14090) );
  INVX0 U14001 ( .INP(n13993), .ZN(n14082) );
  NOR2X0 U14002 ( .IN1(n14068), .IN2(n11737), .QN(n13993) );
  NAND2X0 U14003 ( .IN1(n14092), .IN2(n14093), .QN(n11737) );
  NAND2X0 U14004 ( .IN1(g1088), .IN2(g1101), .QN(n14093) );
  NOR2X0 U14005 ( .IN1(n14094), .IN2(n14095), .QN(n14092) );
  NOR2X0 U14006 ( .IN1(n9751), .IN2(n4364), .QN(n14095) );
  NOR2X0 U14007 ( .IN1(n9773), .IN2(n4363), .QN(n14094) );
  NAND2X0 U14008 ( .IN1(g996), .IN2(n14087), .QN(n14068) );
  NAND2X0 U14009 ( .IN1(n14096), .IN2(n14097), .QN(n14087) );
  NAND2X0 U14010 ( .IN1(n4283), .IN2(n11738), .QN(n14097) );
  NAND2X0 U14011 ( .IN1(n14098), .IN2(n13374), .QN(n14096) );
  INVX0 U14012 ( .INP(n11738), .ZN(n13374) );
  NAND2X0 U14013 ( .IN1(n14099), .IN2(n14100), .QN(n11738) );
  NOR2X0 U14014 ( .IN1(n13804), .IN2(n12178), .QN(n14099) );
  NOR2X0 U14015 ( .IN1(n11796), .IN2(n4283), .QN(n14098) );
  NOR2X0 U14016 ( .IN1(n10718), .IN2(n10031), .QN(n11796) );
  NAND2X0 U14017 ( .IN1(n14101), .IN2(n14102), .QN(n10718) );
  NAND2X0 U14018 ( .IN1(test_so31), .IN2(n9922), .QN(n14102) );
  NOR2X0 U14019 ( .IN1(n14103), .IN2(n14104), .QN(n14101) );
  NOR2X0 U14020 ( .IN1(n4323), .IN2(g857), .QN(n14104) );
  NOR2X0 U14021 ( .IN1(test_so33), .IN2(n4312), .QN(n14103) );
  NAND2X0 U14022 ( .IN1(n14105), .IN2(n14106), .QN(g28736) );
  NAND2X0 U14023 ( .IN1(test_so17), .IN2(n14107), .QN(n14106) );
  NAND2X0 U14024 ( .IN1(n14037), .IN2(n12042), .QN(n14107) );
  INVX0 U14025 ( .INP(n14108), .ZN(n14037) );
  NAND2X0 U14026 ( .IN1(n14109), .IN2(n13399), .QN(n14108) );
  NAND2X0 U14027 ( .IN1(n14038), .IN2(n12042), .QN(n14105) );
  INVX0 U14028 ( .INP(n14110), .ZN(n14038) );
  NAND2X0 U14029 ( .IN1(n14111), .IN2(n14112), .QN(g28735) );
  NAND2X0 U14030 ( .IN1(g6447), .IN2(n14077), .QN(n14112) );
  INVX0 U14031 ( .INP(n14113), .ZN(n14111) );
  NOR2X0 U14032 ( .IN1(n13382), .IN2(n9784), .QN(n14113) );
  NAND2X0 U14033 ( .IN1(n14114), .IN2(n14115), .QN(g28732) );
  NAND2X0 U14034 ( .IN1(g5437), .IN2(n14077), .QN(n14115) );
  NAND2X0 U14035 ( .IN1(n14110), .IN2(n14116), .QN(n14077) );
  NAND2X0 U14036 ( .IN1(n14117), .IN2(n11732), .QN(n14116) );
  NAND2X0 U14037 ( .IN1(g309), .IN2(n14118), .QN(n14117) );
  NAND2X0 U14038 ( .IN1(n13399), .IN2(n14119), .QN(n14118) );
  NOR2X0 U14039 ( .IN1(n14120), .IN2(n14121), .QN(n13399) );
  NOR2X0 U14040 ( .IN1(n4520), .IN2(test_so17), .QN(n14121) );
  INVX0 U14041 ( .INP(n14122), .ZN(n14120) );
  NOR2X0 U14042 ( .IN1(n14123), .IN2(n14124), .QN(n14122) );
  NOR2X0 U14043 ( .IN1(n4499), .IN2(g428), .QN(n14124) );
  NOR2X0 U14044 ( .IN1(n4506), .IN2(g426), .QN(n14123) );
  NAND2X0 U14045 ( .IN1(n14109), .IN2(n13398), .QN(n14110) );
  INVX0 U14046 ( .INP(n11732), .ZN(n13398) );
  NAND2X0 U14047 ( .IN1(n14125), .IN2(n14126), .QN(n11732) );
  NAND2X0 U14048 ( .IN1(g5437), .IN2(g408), .QN(n14126) );
  NOR2X0 U14049 ( .IN1(n14127), .IN2(n14128), .QN(n14125) );
  NOR2X0 U14050 ( .IN1(n9784), .IN2(n14129), .QN(n14128) );
  NOR2X0 U14051 ( .IN1(n9783), .IN2(n14130), .QN(n14127) );
  NOR2X0 U14052 ( .IN1(n4388), .IN2(n14131), .QN(n14109) );
  INVX0 U14053 ( .INP(n14119), .ZN(n14131) );
  NAND2X0 U14054 ( .IN1(n14132), .IN2(n14133), .QN(n14119) );
  NAND2X0 U14055 ( .IN1(n4282), .IN2(n11733), .QN(n14133) );
  NAND2X0 U14056 ( .IN1(n14134), .IN2(n13394), .QN(n14132) );
  INVX0 U14057 ( .INP(n11733), .ZN(n13394) );
  NAND2X0 U14058 ( .IN1(n14135), .IN2(n14136), .QN(n11733) );
  NOR2X0 U14059 ( .IN1(n12454), .IN2(n12247), .QN(n14135) );
  NOR2X0 U14060 ( .IN1(n12032), .IN2(n4282), .QN(n14134) );
  NOR2X0 U14061 ( .IN1(n11721), .IN2(n10032), .QN(n12032) );
  NAND2X0 U14062 ( .IN1(n14137), .IN2(n14138), .QN(n11721) );
  NAND2X0 U14063 ( .IN1(n9934), .IN2(g6313), .QN(n14138) );
  NOR2X0 U14064 ( .IN1(n14139), .IN2(n14140), .QN(n14137) );
  NOR2X0 U14065 ( .IN1(n4369), .IN2(g168), .QN(n14140) );
  NOR2X0 U14066 ( .IN1(n4318), .IN2(g169), .QN(n14139) );
  NAND2X0 U14067 ( .IN1(n4520), .IN2(g408), .QN(n14114) );
  NOR2X0 U14068 ( .IN1(n14141), .IN2(n14142), .QN(g28668) );
  NAND2X0 U14069 ( .IN1(n14143), .IN2(n14144), .QN(n14142) );
  NAND2X0 U14070 ( .IN1(n4418), .IN2(n14145), .QN(n14144) );
  NAND2X0 U14071 ( .IN1(n14146), .IN2(g692), .QN(n14143) );
  NAND2X0 U14072 ( .IN1(n14147), .IN2(n14148), .QN(g28637) );
  NAND2X0 U14073 ( .IN1(n14149), .IN2(g2133), .QN(n14148) );
  INVX0 U14074 ( .INP(n14150), .ZN(n14149) );
  NAND2X0 U14075 ( .IN1(n14151), .IN2(n10010), .QN(n14147) );
  NOR2X0 U14076 ( .IN1(n13263), .IN2(n3160), .QN(n14151) );
  NAND2X0 U14077 ( .IN1(n14152), .IN2(n14153), .QN(g28636) );
  NAND2X0 U14078 ( .IN1(n14154), .IN2(g1439), .QN(n14153) );
  INVX0 U14079 ( .INP(n14155), .ZN(n14154) );
  NAND2X0 U14080 ( .IN1(n14156), .IN2(n10014), .QN(n14152) );
  NOR2X0 U14081 ( .IN1(n13268), .IN2(n3164), .QN(n14156) );
  NAND2X0 U14082 ( .IN1(n14157), .IN2(n14158), .QN(g28635) );
  NAND2X0 U14083 ( .IN1(n14159), .IN2(g753), .QN(n14158) );
  INVX0 U14084 ( .INP(n14160), .ZN(n14159) );
  NAND2X0 U14085 ( .IN1(n14161), .IN2(n10018), .QN(n14157) );
  NOR2X0 U14086 ( .IN1(n13273), .IN2(n3168), .QN(n14161) );
  NAND2X0 U14087 ( .IN1(n14162), .IN2(n14163), .QN(g28634) );
  NAND2X0 U14088 ( .IN1(n14164), .IN2(g65), .QN(n14163) );
  INVX0 U14089 ( .INP(n14165), .ZN(n14164) );
  NAND2X0 U14090 ( .IN1(n14166), .IN2(n10022), .QN(n14162) );
  NOR2X0 U14091 ( .IN1(n13278), .IN2(n3172), .QN(n14166) );
  NAND2X0 U14092 ( .IN1(n14167), .IN2(n14168), .QN(g28425) );
  INVX0 U14093 ( .INP(n14169), .ZN(n14168) );
  NOR2X0 U14094 ( .IN1(g3109), .IN2(n4343), .QN(n14169) );
  NAND2X0 U14095 ( .IN1(n588), .IN2(g3109), .QN(n14167) );
  NAND2X0 U14096 ( .IN1(n14170), .IN2(n14171), .QN(g28421) );
  NAND2X0 U14097 ( .IN1(n4383), .IN2(test_so7), .QN(n14171) );
  NAND2X0 U14098 ( .IN1(n588), .IN2(g8030), .QN(n14170) );
  NAND2X0 U14099 ( .IN1(n14172), .IN2(n14173), .QN(g28420) );
  INVX0 U14100 ( .INP(n14174), .ZN(n14173) );
  NOR2X0 U14101 ( .IN1(g8106), .IN2(n4342), .QN(n14174) );
  NAND2X0 U14102 ( .IN1(n588), .IN2(g8106), .QN(n14172) );
  INVX0 U14103 ( .INP(n13200), .ZN(n588) );
  NAND2X0 U14104 ( .IN1(n14175), .IN2(n14176), .QN(n13200) );
  NAND2X0 U14105 ( .IN1(n9414), .IN2(g1186), .QN(n14176) );
  NAND2X0 U14106 ( .IN1(n14177), .IN2(n4548), .QN(n14175) );
  NOR2X0 U14107 ( .IN1(n14178), .IN2(n14179), .QN(n14177) );
  NOR2X0 U14108 ( .IN1(n9415), .IN2(n14180), .QN(n14179) );
  INVX0 U14109 ( .INP(n14181), .ZN(n14178) );
  NAND2X0 U14110 ( .IN1(g21851), .IN2(g6750), .QN(n14181) );
  NAND2X0 U14111 ( .IN1(n14182), .IN2(n14183), .QN(g28371) );
  INVX0 U14112 ( .INP(n14184), .ZN(n14183) );
  NOR2X0 U14113 ( .IN1(g2624), .IN2(n9720), .QN(n14184) );
  NAND2X0 U14114 ( .IN1(n14185), .IN2(g2624), .QN(n14182) );
  NAND2X0 U14115 ( .IN1(n14186), .IN2(n14187), .QN(g28368) );
  NAND2X0 U14116 ( .IN1(n4370), .IN2(g2691), .QN(n14187) );
  NAND2X0 U14117 ( .IN1(n14185), .IN2(g7390), .QN(n14186) );
  NAND2X0 U14118 ( .IN1(n14188), .IN2(n14189), .QN(g28367) );
  INVX0 U14119 ( .INP(n14190), .ZN(n14189) );
  NOR2X0 U14120 ( .IN1(g2624), .IN2(n9729), .QN(n14190) );
  NAND2X0 U14121 ( .IN1(n14191), .IN2(g2624), .QN(n14188) );
  NAND2X0 U14122 ( .IN1(n14192), .IN2(n14193), .QN(g28366) );
  NAND2X0 U14123 ( .IN1(n4366), .IN2(g2000), .QN(n14193) );
  NAND2X0 U14124 ( .IN1(n14194), .IN2(g1930), .QN(n14192) );
  NAND2X0 U14125 ( .IN1(n14195), .IN2(n14196), .QN(g28364) );
  INVX0 U14126 ( .INP(n14197), .ZN(n14196) );
  NOR2X0 U14127 ( .IN1(n13147), .IN2(n9719), .QN(n14197) );
  NAND2X0 U14128 ( .IN1(n14185), .IN2(n13147), .QN(n14195) );
  NAND2X0 U14129 ( .IN1(n14198), .IN2(n14199), .QN(n14185) );
  NAND2X0 U14130 ( .IN1(n3252), .IN2(n14200), .QN(n14199) );
  NAND2X0 U14131 ( .IN1(n11354), .IN2(n14201), .QN(n14198) );
  NAND2X0 U14132 ( .IN1(n14202), .IN2(n14203), .QN(g28363) );
  NAND2X0 U14133 ( .IN1(n14191), .IN2(g7390), .QN(n14203) );
  NAND2X0 U14134 ( .IN1(n4370), .IN2(test_so90), .QN(n14202) );
  NAND2X0 U14135 ( .IN1(n14204), .IN2(n14205), .QN(g28362) );
  INVX0 U14136 ( .INP(n14206), .ZN(n14205) );
  NOR2X0 U14137 ( .IN1(g7194), .IN2(n9724), .QN(n14206) );
  NAND2X0 U14138 ( .IN1(n14194), .IN2(g7194), .QN(n14204) );
  NAND2X0 U14139 ( .IN1(n14207), .IN2(n14208), .QN(g28361) );
  NAND2X0 U14140 ( .IN1(n4366), .IN2(g1991), .QN(n14208) );
  NAND2X0 U14141 ( .IN1(n14209), .IN2(g1930), .QN(n14207) );
  NAND2X0 U14142 ( .IN1(n14210), .IN2(n14211), .QN(g28360) );
  INVX0 U14143 ( .INP(n14212), .ZN(n14211) );
  NOR2X0 U14144 ( .IN1(g1236), .IN2(n9726), .QN(n14212) );
  NAND2X0 U14145 ( .IN1(n14213), .IN2(g1236), .QN(n14210) );
  NAND2X0 U14146 ( .IN1(n14214), .IN2(n14215), .QN(g28358) );
  NAND2X0 U14147 ( .IN1(g7302), .IN2(n14191), .QN(n14215) );
  NAND2X0 U14148 ( .IN1(n14216), .IN2(n14217), .QN(n14191) );
  NAND2X0 U14149 ( .IN1(n11846), .IN2(n14201), .QN(n14217) );
  NAND2X0 U14150 ( .IN1(n14218), .IN2(n14200), .QN(n14216) );
  NOR2X0 U14151 ( .IN1(n14219), .IN2(n11727), .QN(n14218) );
  NAND2X0 U14152 ( .IN1(n14220), .IN2(n14221), .QN(n11727) );
  NOR2X0 U14153 ( .IN1(n14222), .IN2(n14223), .QN(n14221) );
  NOR2X0 U14154 ( .IN1(n14224), .IN2(n14225), .QN(n14223) );
  NAND2X0 U14155 ( .IN1(n14226), .IN2(n14227), .QN(n14225) );
  NAND2X0 U14156 ( .IN1(n14228), .IN2(n14229), .QN(n14227) );
  NAND2X0 U14157 ( .IN1(n14230), .IN2(n14231), .QN(n14229) );
  NOR2X0 U14158 ( .IN1(n14232), .IN2(n14233), .QN(n14222) );
  NOR2X0 U14159 ( .IN1(n14234), .IN2(n14235), .QN(n14232) );
  INVX0 U14160 ( .INP(n14236), .ZN(n14235) );
  NAND2X0 U14161 ( .IN1(n14230), .IN2(n14237), .QN(n14236) );
  NAND2X0 U14162 ( .IN1(n14238), .IN2(n14239), .QN(n14230) );
  NAND2X0 U14163 ( .IN1(n14240), .IN2(n14241), .QN(n14239) );
  NOR2X0 U14164 ( .IN1(n14228), .IN2(n14242), .QN(n14234) );
  INVX0 U14165 ( .INP(n14243), .ZN(n14228) );
  NAND2X0 U14166 ( .IN1(n14244), .IN2(n14245), .QN(n14243) );
  NAND2X0 U14167 ( .IN1(n14246), .IN2(n14247), .QN(n14245) );
  NAND2X0 U14168 ( .IN1(n14248), .IN2(n14241), .QN(n14244) );
  NOR2X0 U14169 ( .IN1(n14249), .IN2(n14250), .QN(n14220) );
  NOR2X0 U14170 ( .IN1(n14247), .IN2(n14251), .QN(n14250) );
  NAND2X0 U14171 ( .IN1(n14252), .IN2(n14253), .QN(n14251) );
  NAND2X0 U14172 ( .IN1(n14254), .IN2(n14255), .QN(n14252) );
  NAND2X0 U14173 ( .IN1(n14256), .IN2(n14257), .QN(n14255) );
  NAND2X0 U14174 ( .IN1(n14226), .IN2(n14248), .QN(n14257) );
  NOR2X0 U14175 ( .IN1(n14258), .IN2(n14241), .QN(n14249) );
  NOR2X0 U14176 ( .IN1(n14259), .IN2(n14260), .QN(n14258) );
  NOR2X0 U14177 ( .IN1(n14240), .IN2(n14261), .QN(n14260) );
  NOR2X0 U14178 ( .IN1(n14262), .IN2(n14256), .QN(n14261) );
  NOR2X0 U14179 ( .IN1(n14224), .IN2(n14237), .QN(n14262) );
  NOR2X0 U14180 ( .IN1(n14263), .IN2(n14264), .QN(n14259) );
  NAND2X0 U14181 ( .IN1(n14256), .IN2(n14246), .QN(n14264) );
  INVX0 U14182 ( .INP(n14253), .ZN(n14246) );
  NAND2X0 U14183 ( .IN1(n14238), .IN2(n14265), .QN(n14263) );
  NAND2X0 U14184 ( .IN1(n14266), .IN2(n11724), .QN(n14219) );
  NAND2X0 U14185 ( .IN1(n11726), .IN2(n14267), .QN(n11724) );
  NAND2X0 U14186 ( .IN1(n1658), .IN2(n14268), .QN(n14266) );
  INVX0 U14187 ( .INP(n14269), .ZN(n1658) );
  NAND2X0 U14188 ( .IN1(n14270), .IN2(n14271), .QN(n14269) );
  NAND2X0 U14189 ( .IN1(n14272), .IN2(n14233), .QN(n14271) );
  NAND2X0 U14190 ( .IN1(n14273), .IN2(n14274), .QN(n14272) );
  NAND2X0 U14191 ( .IN1(n14275), .IN2(n14237), .QN(n14274) );
  NAND2X0 U14192 ( .IN1(n14247), .IN2(n14276), .QN(n14273) );
  NAND2X0 U14193 ( .IN1(n14277), .IN2(n14278), .QN(n14276) );
  NAND2X0 U14194 ( .IN1(n14256), .IN2(n14253), .QN(n14278) );
  NOR2X0 U14195 ( .IN1(n14279), .IN2(n14280), .QN(n14277) );
  NOR2X0 U14196 ( .IN1(n14242), .IN2(n14281), .QN(n14280) );
  INVX0 U14197 ( .INP(n14282), .ZN(n14281) );
  NOR2X0 U14198 ( .IN1(n14237), .IN2(n14283), .QN(n14279) );
  NAND2X0 U14199 ( .IN1(n14248), .IN2(n14265), .QN(n14283) );
  NOR2X0 U14200 ( .IN1(n14284), .IN2(n14285), .QN(n14270) );
  NOR2X0 U14201 ( .IN1(n14247), .IN2(n14286), .QN(n14285) );
  NOR2X0 U14202 ( .IN1(n14287), .IN2(n14288), .QN(n14286) );
  NOR2X0 U14203 ( .IN1(n14289), .IN2(n14233), .QN(n14288) );
  NOR2X0 U14204 ( .IN1(n14290), .IN2(n14291), .QN(n14289) );
  NAND2X0 U14205 ( .IN1(n14292), .IN2(n14293), .QN(n14291) );
  NAND2X0 U14206 ( .IN1(n14282), .IN2(n14256), .QN(n14293) );
  INVX0 U14207 ( .INP(n14231), .ZN(n14256) );
  INVX0 U14208 ( .INP(n14294), .ZN(n14292) );
  NOR2X0 U14209 ( .IN1(n14254), .IN2(n14253), .QN(n14294) );
  NAND2X0 U14210 ( .IN1(n14295), .IN2(n14238), .QN(n14254) );
  NOR2X0 U14211 ( .IN1(n14226), .IN2(n14237), .QN(n14295) );
  INVX0 U14212 ( .INP(n14296), .ZN(n14237) );
  NAND2X0 U14213 ( .IN1(n14297), .IN2(n14298), .QN(n14296) );
  NAND2X0 U14214 ( .IN1(test_so85), .IN2(g2412), .QN(n14298) );
  NOR2X0 U14215 ( .IN1(n14299), .IN2(n14300), .QN(n14297) );
  NOR2X0 U14216 ( .IN1(n18860), .IN2(n9651), .QN(n14300) );
  NOR2X0 U14217 ( .IN1(n9654), .IN2(n9452), .QN(n14299) );
  INVX0 U14218 ( .INP(n14265), .ZN(n14226) );
  NOR2X0 U14219 ( .IN1(n14238), .IN2(n14265), .QN(n14290) );
  NOR2X0 U14220 ( .IN1(n14240), .IN2(n14242), .QN(n14287) );
  NAND2X0 U14221 ( .IN1(n14231), .IN2(n14265), .QN(n14242) );
  NOR2X0 U14222 ( .IN1(n14265), .IN2(n14301), .QN(n14284) );
  NAND2X0 U14223 ( .IN1(n14302), .IN2(n14253), .QN(n14301) );
  NAND2X0 U14224 ( .IN1(n14303), .IN2(n14304), .QN(n14302) );
  NAND2X0 U14225 ( .IN1(n14247), .IN2(n14238), .QN(n14304) );
  INVX0 U14226 ( .INP(n14241), .ZN(n14247) );
  NAND2X0 U14227 ( .IN1(n14305), .IN2(n14306), .QN(n14241) );
  NAND2X0 U14228 ( .IN1(g5796), .IN2(g2426), .QN(n14306) );
  NOR2X0 U14229 ( .IN1(n14307), .IN2(n14308), .QN(n14305) );
  NOR2X0 U14230 ( .IN1(n9653), .IN2(n9652), .QN(n14308) );
  NOR2X0 U14231 ( .IN1(n18859), .IN2(n9651), .QN(n14307) );
  NAND2X0 U14232 ( .IN1(n14224), .IN2(n14231), .QN(n14303) );
  NAND2X0 U14233 ( .IN1(n14309), .IN2(n14310), .QN(n14231) );
  NAND2X0 U14234 ( .IN1(g5747), .IN2(g2454), .QN(n14310) );
  NOR2X0 U14235 ( .IN1(n14311), .IN2(n14312), .QN(n14309) );
  NOR2X0 U14236 ( .IN1(n9654), .IN2(n9618), .QN(n14312) );
  NOR2X0 U14237 ( .IN1(n9652), .IN2(n9617), .QN(n14311) );
  NAND2X0 U14238 ( .IN1(n14313), .IN2(n14314), .QN(n14265) );
  NAND2X0 U14239 ( .IN1(g5747), .IN2(g2439), .QN(n14314) );
  NOR2X0 U14240 ( .IN1(n14315), .IN2(n14316), .QN(n14313) );
  NOR2X0 U14241 ( .IN1(n9654), .IN2(n9444), .QN(n14316) );
  NOR2X0 U14242 ( .IN1(n9652), .IN2(n9443), .QN(n14315) );
  INVX0 U14243 ( .INP(n14317), .ZN(n14214) );
  NOR2X0 U14244 ( .IN1(n13147), .IN2(n9728), .QN(n14317) );
  NAND2X0 U14245 ( .IN1(n14318), .IN2(n14319), .QN(g28357) );
  INVX0 U14246 ( .INP(n14320), .ZN(n14319) );
  NOR2X0 U14247 ( .IN1(n14321), .IN2(n9722), .QN(n14320) );
  NAND2X0 U14248 ( .IN1(n14194), .IN2(n14321), .QN(n14318) );
  NAND2X0 U14249 ( .IN1(n14322), .IN2(n14323), .QN(n14194) );
  NAND2X0 U14250 ( .IN1(n11527), .IN2(n14201), .QN(n14323) );
  NAND2X0 U14251 ( .IN1(n14324), .IN2(n14200), .QN(n14322) );
  NOR2X0 U14252 ( .IN1(n14325), .IN2(n14326), .QN(n14324) );
  NAND2X0 U14253 ( .IN1(n14327), .IN2(n14328), .QN(n14325) );
  INVX0 U14254 ( .INP(n14329), .ZN(n14327) );
  NOR2X0 U14255 ( .IN1(n14330), .IN2(n14331), .QN(n14329) );
  NAND2X0 U14256 ( .IN1(n14332), .IN2(n14333), .QN(g28356) );
  INVX0 U14257 ( .INP(n14334), .ZN(n14333) );
  NOR2X0 U14258 ( .IN1(g7194), .IN2(n9732), .QN(n14334) );
  NAND2X0 U14259 ( .IN1(n14209), .IN2(g7194), .QN(n14332) );
  NAND2X0 U14260 ( .IN1(n14335), .IN2(n14336), .QN(g28355) );
  INVX0 U14261 ( .INP(n14337), .ZN(n14336) );
  NOR2X0 U14262 ( .IN1(g6944), .IN2(n9727), .QN(n14337) );
  NAND2X0 U14263 ( .IN1(n14213), .IN2(g6944), .QN(n14335) );
  NAND2X0 U14264 ( .IN1(n14338), .IN2(n14339), .QN(g28354) );
  INVX0 U14265 ( .INP(n14340), .ZN(n14339) );
  NOR2X0 U14266 ( .IN1(g1236), .IN2(n9734), .QN(n14340) );
  NAND2X0 U14267 ( .IN1(n14341), .IN2(g1236), .QN(n14338) );
  NAND2X0 U14268 ( .IN1(n14342), .IN2(n14343), .QN(g28353) );
  NAND2X0 U14269 ( .IN1(n14344), .IN2(g550), .QN(n14343) );
  NAND2X0 U14270 ( .IN1(test_so26), .IN2(n4313), .QN(n14342) );
  NAND2X0 U14271 ( .IN1(n14345), .IN2(n14346), .QN(g28352) );
  NAND2X0 U14272 ( .IN1(g7052), .IN2(n14209), .QN(n14346) );
  NAND2X0 U14273 ( .IN1(n14347), .IN2(n14348), .QN(n14209) );
  NAND2X0 U14274 ( .IN1(n11508), .IN2(n14201), .QN(n14348) );
  NAND2X0 U14275 ( .IN1(n14349), .IN2(n14200), .QN(n14347) );
  NOR2X0 U14276 ( .IN1(n14350), .IN2(n14331), .QN(n14349) );
  NAND2X0 U14277 ( .IN1(n14351), .IN2(n14352), .QN(n14331) );
  NOR2X0 U14278 ( .IN1(n14353), .IN2(n14354), .QN(n14352) );
  NOR2X0 U14279 ( .IN1(n14355), .IN2(n14356), .QN(n14354) );
  NAND2X0 U14280 ( .IN1(n14357), .IN2(n14358), .QN(n14356) );
  NAND2X0 U14281 ( .IN1(n14359), .IN2(n14360), .QN(n14358) );
  NAND2X0 U14282 ( .IN1(n14361), .IN2(n14362), .QN(n14360) );
  NOR2X0 U14283 ( .IN1(n14363), .IN2(n14364), .QN(n14353) );
  NOR2X0 U14284 ( .IN1(n14365), .IN2(n14366), .QN(n14363) );
  INVX0 U14285 ( .INP(n14367), .ZN(n14366) );
  NAND2X0 U14286 ( .IN1(n14361), .IN2(n14368), .QN(n14367) );
  NAND2X0 U14287 ( .IN1(n14369), .IN2(n14370), .QN(n14361) );
  NAND2X0 U14288 ( .IN1(n14371), .IN2(n14372), .QN(n14370) );
  NOR2X0 U14289 ( .IN1(n14359), .IN2(n14373), .QN(n14365) );
  INVX0 U14290 ( .INP(n14374), .ZN(n14359) );
  NAND2X0 U14291 ( .IN1(n14375), .IN2(n14376), .QN(n14374) );
  NAND2X0 U14292 ( .IN1(n14377), .IN2(n14378), .QN(n14376) );
  NAND2X0 U14293 ( .IN1(n14379), .IN2(n14372), .QN(n14375) );
  NOR2X0 U14294 ( .IN1(n14380), .IN2(n14381), .QN(n14351) );
  NOR2X0 U14295 ( .IN1(n14378), .IN2(n14382), .QN(n14381) );
  NAND2X0 U14296 ( .IN1(n14383), .IN2(n14384), .QN(n14382) );
  NAND2X0 U14297 ( .IN1(n14385), .IN2(n14386), .QN(n14383) );
  NAND2X0 U14298 ( .IN1(n14387), .IN2(n14388), .QN(n14386) );
  NAND2X0 U14299 ( .IN1(n14357), .IN2(n14379), .QN(n14388) );
  NOR2X0 U14300 ( .IN1(n14389), .IN2(n14372), .QN(n14380) );
  NOR2X0 U14301 ( .IN1(n14390), .IN2(n14391), .QN(n14389) );
  NOR2X0 U14302 ( .IN1(n14371), .IN2(n14392), .QN(n14391) );
  NOR2X0 U14303 ( .IN1(n14393), .IN2(n14387), .QN(n14392) );
  NOR2X0 U14304 ( .IN1(n14355), .IN2(n14368), .QN(n14393) );
  NOR2X0 U14305 ( .IN1(n14394), .IN2(n14395), .QN(n14390) );
  NAND2X0 U14306 ( .IN1(n14387), .IN2(n14377), .QN(n14395) );
  INVX0 U14307 ( .INP(n14384), .ZN(n14377) );
  NAND2X0 U14308 ( .IN1(n14369), .IN2(n14396), .QN(n14394) );
  NAND2X0 U14309 ( .IN1(n14328), .IN2(n14397), .QN(n14350) );
  INVX0 U14310 ( .INP(n14398), .ZN(n14397) );
  NOR2X0 U14311 ( .IN1(n14399), .IN2(n14326), .QN(n14398) );
  NAND2X0 U14312 ( .IN1(n14400), .IN2(n14401), .QN(n14326) );
  NAND2X0 U14313 ( .IN1(n14402), .IN2(n14364), .QN(n14401) );
  NAND2X0 U14314 ( .IN1(n14403), .IN2(n14404), .QN(n14402) );
  NAND2X0 U14315 ( .IN1(n14405), .IN2(n14368), .QN(n14404) );
  NAND2X0 U14316 ( .IN1(n14378), .IN2(n14406), .QN(n14403) );
  NAND2X0 U14317 ( .IN1(n14407), .IN2(n14408), .QN(n14406) );
  NAND2X0 U14318 ( .IN1(n14387), .IN2(n14384), .QN(n14408) );
  NOR2X0 U14319 ( .IN1(n14409), .IN2(n14410), .QN(n14407) );
  NOR2X0 U14320 ( .IN1(n14373), .IN2(n14411), .QN(n14410) );
  INVX0 U14321 ( .INP(n14412), .ZN(n14411) );
  NOR2X0 U14322 ( .IN1(n14368), .IN2(n14413), .QN(n14409) );
  NAND2X0 U14323 ( .IN1(n14379), .IN2(n14396), .QN(n14413) );
  NOR2X0 U14324 ( .IN1(n14414), .IN2(n14415), .QN(n14400) );
  NOR2X0 U14325 ( .IN1(n14378), .IN2(n14416), .QN(n14415) );
  NOR2X0 U14326 ( .IN1(n14417), .IN2(n14418), .QN(n14416) );
  NOR2X0 U14327 ( .IN1(n14419), .IN2(n14364), .QN(n14418) );
  NOR2X0 U14328 ( .IN1(n14420), .IN2(n14421), .QN(n14419) );
  NAND2X0 U14329 ( .IN1(n14422), .IN2(n14423), .QN(n14421) );
  NAND2X0 U14330 ( .IN1(n14412), .IN2(n14387), .QN(n14423) );
  INVX0 U14331 ( .INP(n14362), .ZN(n14387) );
  INVX0 U14332 ( .INP(n14424), .ZN(n14422) );
  NOR2X0 U14333 ( .IN1(n14385), .IN2(n14384), .QN(n14424) );
  NAND2X0 U14334 ( .IN1(n14425), .IN2(n14369), .QN(n14385) );
  NOR2X0 U14335 ( .IN1(n14357), .IN2(n14368), .QN(n14425) );
  INVX0 U14336 ( .INP(n14426), .ZN(n14368) );
  NAND2X0 U14337 ( .IN1(n14427), .IN2(n14428), .QN(n14426) );
  NAND2X0 U14338 ( .IN1(test_so63), .IN2(g1775), .QN(n14428) );
  NOR2X0 U14339 ( .IN1(n14429), .IN2(n14430), .QN(n14427) );
  NOR2X0 U14340 ( .IN1(n9665), .IN2(n9664), .QN(n14430) );
  NOR2X0 U14341 ( .IN1(n9663), .IN2(n9662), .QN(n14429) );
  INVX0 U14342 ( .INP(n14396), .ZN(n14357) );
  NOR2X0 U14343 ( .IN1(n14369), .IN2(n14396), .QN(n14420) );
  NOR2X0 U14344 ( .IN1(n14371), .IN2(n14373), .QN(n14417) );
  NAND2X0 U14345 ( .IN1(n14362), .IN2(n14396), .QN(n14373) );
  NOR2X0 U14346 ( .IN1(n14396), .IN2(n14431), .QN(n14414) );
  NAND2X0 U14347 ( .IN1(n14432), .IN2(n14384), .QN(n14431) );
  NAND2X0 U14348 ( .IN1(n14433), .IN2(n14434), .QN(n14432) );
  NAND2X0 U14349 ( .IN1(n14378), .IN2(n14369), .QN(n14434) );
  INVX0 U14350 ( .INP(n14372), .ZN(n14378) );
  NAND2X0 U14351 ( .IN1(n14435), .IN2(n14436), .QN(n14372) );
  NAND2X0 U14352 ( .IN1(test_so63), .IN2(g1730), .QN(n14436) );
  NOR2X0 U14353 ( .IN1(n14437), .IN2(n14438), .QN(n14435) );
  NOR2X0 U14354 ( .IN1(n9664), .IN2(n9657), .QN(n14438) );
  NOR2X0 U14355 ( .IN1(n9662), .IN2(n9656), .QN(n14437) );
  NAND2X0 U14356 ( .IN1(n14355), .IN2(n14362), .QN(n14433) );
  NAND2X0 U14357 ( .IN1(n14439), .IN2(n14440), .QN(n14362) );
  NAND2X0 U14358 ( .IN1(test_so63), .IN2(g1760), .QN(n14440) );
  NOR2X0 U14359 ( .IN1(n14441), .IN2(n14442), .QN(n14439) );
  NOR2X0 U14360 ( .IN1(n9664), .IN2(n9620), .QN(n14442) );
  NOR2X0 U14361 ( .IN1(n9662), .IN2(n9619), .QN(n14441) );
  NAND2X0 U14362 ( .IN1(n14443), .IN2(n14444), .QN(n14396) );
  NAND2X0 U14363 ( .IN1(test_so63), .IN2(g1745), .QN(n14444) );
  NOR2X0 U14364 ( .IN1(n14445), .IN2(n14446), .QN(n14443) );
  NOR2X0 U14365 ( .IN1(n9664), .IN2(n9446), .QN(n14446) );
  NOR2X0 U14366 ( .IN1(n9662), .IN2(n9445), .QN(n14445) );
  NAND2X0 U14367 ( .IN1(n14330), .IN2(n14399), .QN(n14328) );
  INVX0 U14368 ( .INP(n14447), .ZN(n14345) );
  NOR2X0 U14369 ( .IN1(n14321), .IN2(n9730), .QN(n14447) );
  NAND2X0 U14370 ( .IN1(n14448), .IN2(n14449), .QN(g28351) );
  NAND2X0 U14371 ( .IN1(n4371), .IN2(g1300), .QN(n14449) );
  NAND2X0 U14372 ( .IN1(n14213), .IN2(n14180), .QN(n14448) );
  NAND2X0 U14373 ( .IN1(n14450), .IN2(n14451), .QN(n14213) );
  NAND2X0 U14374 ( .IN1(n11703), .IN2(n14201), .QN(n14451) );
  NAND2X0 U14375 ( .IN1(n14452), .IN2(n14200), .QN(n14450) );
  NOR2X0 U14376 ( .IN1(n14453), .IN2(n14454), .QN(n14452) );
  NAND2X0 U14377 ( .IN1(n14455), .IN2(n14456), .QN(n14453) );
  INVX0 U14378 ( .INP(n14457), .ZN(n14455) );
  NOR2X0 U14379 ( .IN1(n14458), .IN2(n14459), .QN(n14457) );
  NAND2X0 U14380 ( .IN1(n14460), .IN2(n14461), .QN(g28350) );
  NAND2X0 U14381 ( .IN1(n4316), .IN2(g1294), .QN(n14461) );
  NAND2X0 U14382 ( .IN1(n14341), .IN2(g6944), .QN(n14460) );
  NAND2X0 U14383 ( .IN1(n14462), .IN2(n14463), .QN(g28349) );
  NAND2X0 U14384 ( .IN1(n4372), .IN2(g617), .QN(n14463) );
  NAND2X0 U14385 ( .IN1(n14344), .IN2(g6642), .QN(n14462) );
  NAND2X0 U14386 ( .IN1(n14464), .IN2(n14465), .QN(g28348) );
  INVX0 U14387 ( .INP(n14466), .ZN(n14465) );
  NOR2X0 U14388 ( .IN1(g550), .IN2(n9717), .QN(n14466) );
  NAND2X0 U14389 ( .IN1(n14467), .IN2(g550), .QN(n14464) );
  NAND2X0 U14390 ( .IN1(n14468), .IN2(n14469), .QN(g28346) );
  NAND2X0 U14391 ( .IN1(g6750), .IN2(n14341), .QN(n14469) );
  NAND2X0 U14392 ( .IN1(n14470), .IN2(n14471), .QN(n14341) );
  NAND2X0 U14393 ( .IN1(n11684), .IN2(n14201), .QN(n14471) );
  NAND2X0 U14394 ( .IN1(n14472), .IN2(n14200), .QN(n14470) );
  NOR2X0 U14395 ( .IN1(n14473), .IN2(n14459), .QN(n14472) );
  NAND2X0 U14396 ( .IN1(n14474), .IN2(n14475), .QN(n14459) );
  NOR2X0 U14397 ( .IN1(n14476), .IN2(n14477), .QN(n14475) );
  NOR2X0 U14398 ( .IN1(n14478), .IN2(n14479), .QN(n14477) );
  NAND2X0 U14399 ( .IN1(n14480), .IN2(n14481), .QN(n14479) );
  NAND2X0 U14400 ( .IN1(n14482), .IN2(n14483), .QN(n14481) );
  NAND2X0 U14401 ( .IN1(n14484), .IN2(n14485), .QN(n14483) );
  NOR2X0 U14402 ( .IN1(n14486), .IN2(n14487), .QN(n14476) );
  NOR2X0 U14403 ( .IN1(n14488), .IN2(n14489), .QN(n14486) );
  INVX0 U14404 ( .INP(n14490), .ZN(n14489) );
  NAND2X0 U14405 ( .IN1(n14484), .IN2(n14491), .QN(n14490) );
  NAND2X0 U14406 ( .IN1(n14492), .IN2(n14493), .QN(n14484) );
  NAND2X0 U14407 ( .IN1(n14494), .IN2(n14495), .QN(n14493) );
  NOR2X0 U14408 ( .IN1(n14482), .IN2(n14496), .QN(n14488) );
  INVX0 U14409 ( .INP(n14497), .ZN(n14482) );
  NAND2X0 U14410 ( .IN1(n14498), .IN2(n14499), .QN(n14497) );
  NAND2X0 U14411 ( .IN1(n14500), .IN2(n14501), .QN(n14499) );
  NAND2X0 U14412 ( .IN1(n14502), .IN2(n14495), .QN(n14498) );
  NOR2X0 U14413 ( .IN1(n14503), .IN2(n14504), .QN(n14474) );
  NOR2X0 U14414 ( .IN1(n14501), .IN2(n14505), .QN(n14504) );
  NAND2X0 U14415 ( .IN1(n14506), .IN2(n14507), .QN(n14505) );
  NAND2X0 U14416 ( .IN1(n14508), .IN2(n14509), .QN(n14506) );
  NAND2X0 U14417 ( .IN1(n14510), .IN2(n14511), .QN(n14509) );
  NAND2X0 U14418 ( .IN1(n14480), .IN2(n14502), .QN(n14511) );
  NOR2X0 U14419 ( .IN1(n14512), .IN2(n14495), .QN(n14503) );
  NOR2X0 U14420 ( .IN1(n14513), .IN2(n14514), .QN(n14512) );
  NOR2X0 U14421 ( .IN1(n14494), .IN2(n14515), .QN(n14514) );
  NOR2X0 U14422 ( .IN1(n14516), .IN2(n14510), .QN(n14515) );
  NOR2X0 U14423 ( .IN1(n14478), .IN2(n14491), .QN(n14516) );
  NOR2X0 U14424 ( .IN1(n14517), .IN2(n14518), .QN(n14513) );
  NAND2X0 U14425 ( .IN1(n14510), .IN2(n14500), .QN(n14518) );
  INVX0 U14426 ( .INP(n14507), .ZN(n14500) );
  NAND2X0 U14427 ( .IN1(n14492), .IN2(n14519), .QN(n14517) );
  NAND2X0 U14428 ( .IN1(n14456), .IN2(n14520), .QN(n14473) );
  INVX0 U14429 ( .INP(n14521), .ZN(n14520) );
  NOR2X0 U14430 ( .IN1(n14522), .IN2(n14454), .QN(n14521) );
  NAND2X0 U14431 ( .IN1(n14523), .IN2(n14524), .QN(n14454) );
  NAND2X0 U14432 ( .IN1(n14525), .IN2(n14487), .QN(n14524) );
  NAND2X0 U14433 ( .IN1(n14526), .IN2(n14527), .QN(n14525) );
  NAND2X0 U14434 ( .IN1(n14528), .IN2(n14491), .QN(n14527) );
  NAND2X0 U14435 ( .IN1(n14501), .IN2(n14529), .QN(n14526) );
  NAND2X0 U14436 ( .IN1(n14530), .IN2(n14531), .QN(n14529) );
  NAND2X0 U14437 ( .IN1(n14510), .IN2(n14507), .QN(n14531) );
  NOR2X0 U14438 ( .IN1(n14532), .IN2(n14533), .QN(n14530) );
  NOR2X0 U14439 ( .IN1(n14496), .IN2(n14534), .QN(n14533) );
  INVX0 U14440 ( .INP(n14535), .ZN(n14534) );
  NOR2X0 U14441 ( .IN1(n14491), .IN2(n14536), .QN(n14532) );
  NAND2X0 U14442 ( .IN1(n14502), .IN2(n14519), .QN(n14536) );
  NOR2X0 U14443 ( .IN1(n14537), .IN2(n14538), .QN(n14523) );
  NOR2X0 U14444 ( .IN1(n14501), .IN2(n14539), .QN(n14538) );
  NOR2X0 U14445 ( .IN1(n14540), .IN2(n14541), .QN(n14539) );
  NOR2X0 U14446 ( .IN1(n14542), .IN2(n14487), .QN(n14541) );
  NOR2X0 U14447 ( .IN1(n14543), .IN2(n14544), .QN(n14542) );
  NAND2X0 U14448 ( .IN1(n14545), .IN2(n14546), .QN(n14544) );
  NAND2X0 U14449 ( .IN1(n14535), .IN2(n14510), .QN(n14546) );
  INVX0 U14450 ( .INP(n14485), .ZN(n14510) );
  INVX0 U14451 ( .INP(n14547), .ZN(n14545) );
  NOR2X0 U14452 ( .IN1(n14508), .IN2(n14507), .QN(n14547) );
  NAND2X0 U14453 ( .IN1(n14548), .IN2(n14492), .QN(n14508) );
  NOR2X0 U14454 ( .IN1(n14480), .IN2(n14491), .QN(n14548) );
  INVX0 U14455 ( .INP(n14549), .ZN(n14491) );
  NAND2X0 U14456 ( .IN1(n14550), .IN2(n14551), .QN(n14549) );
  NAND2X0 U14457 ( .IN1(g5686), .IN2(g1083), .QN(n14551) );
  NOR2X0 U14458 ( .IN1(n14552), .IN2(n14553), .QN(n14550) );
  NOR2X0 U14459 ( .IN1(n9668), .IN2(n9667), .QN(n14553) );
  NOR2X0 U14460 ( .IN1(n18861), .IN2(n9666), .QN(n14552) );
  INVX0 U14461 ( .INP(n14519), .ZN(n14480) );
  NOR2X0 U14462 ( .IN1(n14492), .IN2(n14519), .QN(n14543) );
  NOR2X0 U14463 ( .IN1(n14494), .IN2(n14496), .QN(n14540) );
  NAND2X0 U14464 ( .IN1(n14485), .IN2(n14519), .QN(n14496) );
  NOR2X0 U14465 ( .IN1(n14519), .IN2(n14554), .QN(n14537) );
  NAND2X0 U14466 ( .IN1(n14555), .IN2(n14507), .QN(n14554) );
  NAND2X0 U14467 ( .IN1(n14556), .IN2(n14557), .QN(n14555) );
  NAND2X0 U14468 ( .IN1(n14501), .IN2(n14492), .QN(n14557) );
  INVX0 U14469 ( .INP(n14495), .ZN(n14501) );
  NAND2X0 U14470 ( .IN1(n14558), .IN2(n14559), .QN(n14495) );
  NAND2X0 U14471 ( .IN1(g5657), .IN2(g1036), .QN(n14559) );
  NOR2X0 U14472 ( .IN1(n14560), .IN2(n14561), .QN(n14558) );
  NOR2X0 U14473 ( .IN1(n9669), .IN2(n9659), .QN(n14561) );
  NOR2X0 U14474 ( .IN1(n9667), .IN2(n9658), .QN(n14560) );
  NAND2X0 U14475 ( .IN1(n14478), .IN2(n14485), .QN(n14556) );
  NAND2X0 U14476 ( .IN1(n14562), .IN2(n14563), .QN(n14485) );
  NAND2X0 U14477 ( .IN1(g5657), .IN2(g1066), .QN(n14563) );
  NOR2X0 U14478 ( .IN1(n14564), .IN2(n14565), .QN(n14562) );
  NOR2X0 U14479 ( .IN1(n9669), .IN2(n9622), .QN(n14565) );
  NOR2X0 U14480 ( .IN1(n9667), .IN2(n9621), .QN(n14564) );
  NAND2X0 U14481 ( .IN1(n14566), .IN2(n14567), .QN(n14519) );
  NAND2X0 U14482 ( .IN1(g5657), .IN2(g1051), .QN(n14567) );
  NOR2X0 U14483 ( .IN1(n14568), .IN2(n14569), .QN(n14566) );
  NOR2X0 U14484 ( .IN1(n9669), .IN2(n9448), .QN(n14569) );
  NOR2X0 U14485 ( .IN1(n9667), .IN2(n9447), .QN(n14568) );
  NAND2X0 U14486 ( .IN1(n14458), .IN2(n14522), .QN(n14456) );
  INVX0 U14487 ( .INP(n14570), .ZN(n14468) );
  NOR2X0 U14488 ( .IN1(n14180), .IN2(n9733), .QN(n14570) );
  NAND2X0 U14489 ( .IN1(n14571), .IN2(n14572), .QN(g28345) );
  INVX0 U14490 ( .INP(n14573), .ZN(n14572) );
  NOR2X0 U14491 ( .IN1(n14574), .IN2(n9714), .QN(n14573) );
  NAND2X0 U14492 ( .IN1(n14344), .IN2(n14574), .QN(n14571) );
  NAND2X0 U14493 ( .IN1(n14575), .IN2(n14576), .QN(n14344) );
  NAND2X0 U14494 ( .IN1(n11183), .IN2(n14201), .QN(n14576) );
  NAND2X0 U14495 ( .IN1(n14577), .IN2(n14200), .QN(n14575) );
  NOR2X0 U14496 ( .IN1(n14578), .IN2(n14579), .QN(n14577) );
  NAND2X0 U14497 ( .IN1(n14580), .IN2(n14581), .QN(n14578) );
  INVX0 U14498 ( .INP(n14582), .ZN(n14580) );
  NOR2X0 U14499 ( .IN1(n14583), .IN2(n14584), .QN(n14582) );
  NAND2X0 U14500 ( .IN1(n14585), .IN2(n14586), .QN(g28344) );
  NAND2X0 U14501 ( .IN1(n4372), .IN2(g608), .QN(n14586) );
  NAND2X0 U14502 ( .IN1(n14467), .IN2(g6642), .QN(n14585) );
  NAND2X0 U14503 ( .IN1(n14587), .IN2(n14588), .QN(g28342) );
  NAND2X0 U14504 ( .IN1(g6485), .IN2(n14467), .QN(n14588) );
  NAND2X0 U14505 ( .IN1(n14589), .IN2(n14590), .QN(n14467) );
  NAND2X0 U14506 ( .IN1(n11174), .IN2(n14201), .QN(n14590) );
  NAND2X0 U14507 ( .IN1(n14591), .IN2(n14200), .QN(n14589) );
  NOR2X0 U14508 ( .IN1(n14592), .IN2(n14584), .QN(n14591) );
  NAND2X0 U14509 ( .IN1(n14593), .IN2(n14594), .QN(n14584) );
  NOR2X0 U14510 ( .IN1(n14595), .IN2(n14596), .QN(n14594) );
  NOR2X0 U14511 ( .IN1(n14597), .IN2(n14598), .QN(n14596) );
  NAND2X0 U14512 ( .IN1(n14599), .IN2(n14600), .QN(n14598) );
  NAND2X0 U14513 ( .IN1(n14601), .IN2(n14602), .QN(n14600) );
  NAND2X0 U14514 ( .IN1(n14603), .IN2(n14604), .QN(n14602) );
  NOR2X0 U14515 ( .IN1(n14605), .IN2(n14606), .QN(n14595) );
  NOR2X0 U14516 ( .IN1(n14607), .IN2(n14608), .QN(n14605) );
  INVX0 U14517 ( .INP(n14609), .ZN(n14608) );
  NAND2X0 U14518 ( .IN1(n14603), .IN2(n14610), .QN(n14609) );
  NAND2X0 U14519 ( .IN1(n14611), .IN2(n14612), .QN(n14603) );
  NAND2X0 U14520 ( .IN1(n14613), .IN2(n14614), .QN(n14612) );
  NOR2X0 U14521 ( .IN1(n14601), .IN2(n14615), .QN(n14607) );
  INVX0 U14522 ( .INP(n14616), .ZN(n14601) );
  NAND2X0 U14523 ( .IN1(n14617), .IN2(n14618), .QN(n14616) );
  NAND2X0 U14524 ( .IN1(n14619), .IN2(n14620), .QN(n14618) );
  NAND2X0 U14525 ( .IN1(n14621), .IN2(n14614), .QN(n14617) );
  NOR2X0 U14526 ( .IN1(n14622), .IN2(n14623), .QN(n14593) );
  NOR2X0 U14527 ( .IN1(n14620), .IN2(n14624), .QN(n14623) );
  NAND2X0 U14528 ( .IN1(n14625), .IN2(n14626), .QN(n14624) );
  NAND2X0 U14529 ( .IN1(n14627), .IN2(n14628), .QN(n14625) );
  NAND2X0 U14530 ( .IN1(n14629), .IN2(n14630), .QN(n14628) );
  NAND2X0 U14531 ( .IN1(n14599), .IN2(n14621), .QN(n14630) );
  NOR2X0 U14532 ( .IN1(n14631), .IN2(n14614), .QN(n14622) );
  NOR2X0 U14533 ( .IN1(n14632), .IN2(n14633), .QN(n14631) );
  NOR2X0 U14534 ( .IN1(n14613), .IN2(n14634), .QN(n14633) );
  NOR2X0 U14535 ( .IN1(n14635), .IN2(n14629), .QN(n14634) );
  NOR2X0 U14536 ( .IN1(n14597), .IN2(n14610), .QN(n14635) );
  NOR2X0 U14537 ( .IN1(n14636), .IN2(n14637), .QN(n14632) );
  NAND2X0 U14538 ( .IN1(n14629), .IN2(n14619), .QN(n14637) );
  INVX0 U14539 ( .INP(n14626), .ZN(n14619) );
  NAND2X0 U14540 ( .IN1(n14611), .IN2(n14638), .QN(n14636) );
  NAND2X0 U14541 ( .IN1(n14581), .IN2(n14639), .QN(n14592) );
  INVX0 U14542 ( .INP(n14640), .ZN(n14639) );
  NOR2X0 U14543 ( .IN1(n14641), .IN2(n14579), .QN(n14640) );
  NAND2X0 U14544 ( .IN1(n14642), .IN2(n14643), .QN(n14579) );
  NAND2X0 U14545 ( .IN1(n14644), .IN2(n14606), .QN(n14643) );
  NAND2X0 U14546 ( .IN1(n14645), .IN2(n14646), .QN(n14644) );
  NAND2X0 U14547 ( .IN1(n14647), .IN2(n14610), .QN(n14646) );
  NAND2X0 U14548 ( .IN1(n14620), .IN2(n14648), .QN(n14645) );
  NAND2X0 U14549 ( .IN1(n14649), .IN2(n14650), .QN(n14648) );
  NAND2X0 U14550 ( .IN1(n14629), .IN2(n14626), .QN(n14650) );
  NOR2X0 U14551 ( .IN1(n14651), .IN2(n14652), .QN(n14649) );
  NOR2X0 U14552 ( .IN1(n14615), .IN2(n14653), .QN(n14652) );
  INVX0 U14553 ( .INP(n14654), .ZN(n14653) );
  NOR2X0 U14554 ( .IN1(n14610), .IN2(n14655), .QN(n14651) );
  NAND2X0 U14555 ( .IN1(n14621), .IN2(n14638), .QN(n14655) );
  NOR2X0 U14556 ( .IN1(n14656), .IN2(n14657), .QN(n14642) );
  NOR2X0 U14557 ( .IN1(n14620), .IN2(n14658), .QN(n14657) );
  NOR2X0 U14558 ( .IN1(n14659), .IN2(n14660), .QN(n14658) );
  NOR2X0 U14559 ( .IN1(n14661), .IN2(n14606), .QN(n14660) );
  NOR2X0 U14560 ( .IN1(n14662), .IN2(n14663), .QN(n14661) );
  NAND2X0 U14561 ( .IN1(n14664), .IN2(n14665), .QN(n14663) );
  NAND2X0 U14562 ( .IN1(n14654), .IN2(n14629), .QN(n14665) );
  INVX0 U14563 ( .INP(n14604), .ZN(n14629) );
  INVX0 U14564 ( .INP(n14666), .ZN(n14664) );
  NOR2X0 U14565 ( .IN1(n14627), .IN2(n14626), .QN(n14666) );
  NAND2X0 U14566 ( .IN1(n14667), .IN2(n14611), .QN(n14627) );
  NOR2X0 U14567 ( .IN1(n14599), .IN2(n14610), .QN(n14667) );
  INVX0 U14568 ( .INP(n14668), .ZN(n14610) );
  NAND2X0 U14569 ( .IN1(n14669), .IN2(n14670), .QN(n14668) );
  NAND2X0 U14570 ( .IN1(g5648), .IN2(g396), .QN(n14670) );
  NOR2X0 U14571 ( .IN1(n14671), .IN2(n14672), .QN(n14669) );
  NOR2X0 U14572 ( .IN1(n9673), .IN2(n9672), .QN(n14672) );
  NOR2X0 U14573 ( .IN1(n18862), .IN2(n9671), .QN(n14671) );
  INVX0 U14574 ( .INP(n14638), .ZN(n14599) );
  NOR2X0 U14575 ( .IN1(n14611), .IN2(n14638), .QN(n14662) );
  NOR2X0 U14576 ( .IN1(n14613), .IN2(n14615), .QN(n14659) );
  NAND2X0 U14577 ( .IN1(n14604), .IN2(n14638), .QN(n14615) );
  NOR2X0 U14578 ( .IN1(n14638), .IN2(n14673), .QN(n14656) );
  NAND2X0 U14579 ( .IN1(n14674), .IN2(n14626), .QN(n14673) );
  NAND2X0 U14580 ( .IN1(n14675), .IN2(n14676), .QN(n14674) );
  NAND2X0 U14581 ( .IN1(n14620), .IN2(n14611), .QN(n14676) );
  INVX0 U14582 ( .INP(n14614), .ZN(n14620) );
  NAND2X0 U14583 ( .IN1(n14677), .IN2(n14678), .QN(n14614) );
  NAND2X0 U14584 ( .IN1(g5629), .IN2(g349), .QN(n14678) );
  NOR2X0 U14585 ( .IN1(n14679), .IN2(n14680), .QN(n14677) );
  NOR2X0 U14586 ( .IN1(n9674), .IN2(n9661), .QN(n14680) );
  NOR2X0 U14587 ( .IN1(n9672), .IN2(n9660), .QN(n14679) );
  NAND2X0 U14588 ( .IN1(n14597), .IN2(n14604), .QN(n14675) );
  NAND2X0 U14589 ( .IN1(n14681), .IN2(n14682), .QN(n14604) );
  NAND2X0 U14590 ( .IN1(g5629), .IN2(g379), .QN(n14682) );
  NOR2X0 U14591 ( .IN1(n14683), .IN2(n14684), .QN(n14681) );
  NOR2X0 U14592 ( .IN1(n9674), .IN2(n9624), .QN(n14684) );
  NOR2X0 U14593 ( .IN1(n9672), .IN2(n9623), .QN(n14683) );
  NAND2X0 U14594 ( .IN1(n14685), .IN2(n14686), .QN(n14638) );
  NAND2X0 U14595 ( .IN1(g5629), .IN2(g364), .QN(n14686) );
  NOR2X0 U14596 ( .IN1(n14687), .IN2(n14688), .QN(n14685) );
  NOR2X0 U14597 ( .IN1(n9674), .IN2(n9450), .QN(n14688) );
  NOR2X0 U14598 ( .IN1(n9672), .IN2(n9449), .QN(n14687) );
  NAND2X0 U14599 ( .IN1(n14583), .IN2(n14641), .QN(n14581) );
  INVX0 U14600 ( .INP(n14689), .ZN(n14587) );
  NOR2X0 U14601 ( .IN1(n14574), .IN2(n9716), .QN(n14689) );
  NOR2X0 U14602 ( .IN1(n14690), .IN2(n14691), .QN(g28328) );
  NAND2X0 U14603 ( .IN1(n14692), .IN2(n14693), .QN(n14691) );
  NAND2X0 U14604 ( .IN1(n4415), .IN2(n14694), .QN(n14693) );
  NAND2X0 U14605 ( .IN1(n14695), .IN2(g2766), .QN(n14692) );
  NAND2X0 U14606 ( .IN1(n14696), .IN2(n14697), .QN(g28325) );
  NAND2X0 U14607 ( .IN1(n14698), .IN2(g2072), .QN(n14697) );
  INVX0 U14608 ( .INP(n14699), .ZN(n14698) );
  NAND2X0 U14609 ( .IN1(n14700), .IN2(n4416), .QN(n14696) );
  NOR2X0 U14610 ( .IN1(n10323), .IN2(n14701), .QN(n14700) );
  NAND2X0 U14611 ( .IN1(n14702), .IN2(n14703), .QN(n14701) );
  NOR2X0 U14612 ( .IN1(n14704), .IN2(n14705), .QN(g28321) );
  NAND2X0 U14613 ( .IN1(n14706), .IN2(n14707), .QN(n14705) );
  NAND2X0 U14614 ( .IN1(n4417), .IN2(n14708), .QN(n14707) );
  NAND2X0 U14615 ( .IN1(n14709), .IN2(g1378), .QN(n14706) );
  NOR2X0 U14616 ( .IN1(n14710), .IN2(n14711), .QN(g28199) );
  NAND2X0 U14617 ( .IN1(n14145), .IN2(n14712), .QN(n14711) );
  INVX0 U14618 ( .INP(n14146), .ZN(n14145) );
  NOR2X0 U14619 ( .IN1(n14713), .IN2(n4396), .QN(n14146) );
  NOR2X0 U14620 ( .IN1(n14714), .IN2(g686), .QN(n14710) );
  INVX0 U14621 ( .INP(n14713), .ZN(n14714) );
  NOR2X0 U14622 ( .IN1(n14715), .IN2(n14150), .QN(g28148) );
  NAND2X0 U14623 ( .IN1(n3160), .IN2(n13952), .QN(n14150) );
  NAND2X0 U14624 ( .IN1(n3424), .IN2(g2138), .QN(n3160) );
  NOR2X0 U14625 ( .IN1(n3424), .IN2(g2138), .QN(n14715) );
  NOR2X0 U14626 ( .IN1(n14716), .IN2(n14155), .QN(g28147) );
  NAND2X0 U14627 ( .IN1(n3164), .IN2(n13954), .QN(n14155) );
  NAND2X0 U14628 ( .IN1(n3427), .IN2(g1444), .QN(n3164) );
  NOR2X0 U14629 ( .IN1(n3427), .IN2(g1444), .QN(n14716) );
  NOR2X0 U14630 ( .IN1(n14717), .IN2(n14160), .QN(g28146) );
  NAND2X0 U14631 ( .IN1(n3168), .IN2(n13956), .QN(n14160) );
  NAND2X0 U14632 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NOR2X0 U14633 ( .IN1(n3430), .IN2(g758), .QN(n14717) );
  NOR2X0 U14634 ( .IN1(n14718), .IN2(n14165), .QN(g28145) );
  NAND2X0 U14635 ( .IN1(n3172), .IN2(n13958), .QN(n14165) );
  NAND2X0 U14636 ( .IN1(n3433), .IN2(g70), .QN(n3172) );
  NOR2X0 U14637 ( .IN1(n3433), .IN2(g70), .QN(n14718) );
  NAND2X0 U14638 ( .IN1(n14719), .IN2(n14720), .QN(g27771) );
  NAND2X0 U14639 ( .IN1(test_so81), .IN2(n14721), .QN(n14720) );
  NAND2X0 U14640 ( .IN1(n14722), .IN2(n13307), .QN(n14721) );
  NAND2X0 U14641 ( .IN1(n14723), .IN2(n13307), .QN(n14719) );
  NAND2X0 U14642 ( .IN1(n14724), .IN2(n14725), .QN(g27769) );
  NAND2X0 U14643 ( .IN1(n14726), .IN2(g2524), .QN(n14725) );
  NAND2X0 U14644 ( .IN1(n14722), .IN2(n11937), .QN(n14726) );
  NAND2X0 U14645 ( .IN1(n14723), .IN2(n11937), .QN(n14724) );
  NAND2X0 U14646 ( .IN1(n14727), .IN2(n14728), .QN(g27768) );
  NAND2X0 U14647 ( .IN1(n14729), .IN2(g1828), .QN(n14728) );
  NAND2X0 U14648 ( .IN1(n14730), .IN2(n13315), .QN(n14729) );
  NAND2X0 U14649 ( .IN1(n14731), .IN2(n13315), .QN(n14727) );
  NAND2X0 U14650 ( .IN1(n14732), .IN2(n14733), .QN(g27767) );
  NAND2X0 U14651 ( .IN1(n14734), .IN2(g2523), .QN(n14733) );
  NAND2X0 U14652 ( .IN1(n14722), .IN2(n13416), .QN(n14734) );
  INVX0 U14653 ( .INP(n14735), .ZN(n14722) );
  NAND2X0 U14654 ( .IN1(n14736), .IN2(n14737), .QN(n14735) );
  NOR2X0 U14655 ( .IN1(n14738), .IN2(n14739), .QN(n14737) );
  NOR2X0 U14656 ( .IN1(n10322), .IN2(n14740), .QN(n14736) );
  NAND2X0 U14657 ( .IN1(n14723), .IN2(n13416), .QN(n14732) );
  INVX0 U14658 ( .INP(n14741), .ZN(n14723) );
  NAND2X0 U14659 ( .IN1(n14742), .IN2(n14743), .QN(n14741) );
  NOR2X0 U14660 ( .IN1(n14744), .IN2(n14745), .QN(n14743) );
  NOR2X0 U14661 ( .IN1(n14746), .IN2(n14747), .QN(n14745) );
  NOR2X0 U14662 ( .IN1(n14748), .IN2(n14749), .QN(n14744) );
  NOR2X0 U14663 ( .IN1(n14750), .IN2(n10322), .QN(n14742) );
  NAND2X0 U14664 ( .IN1(n14751), .IN2(n14752), .QN(g27766) );
  NAND2X0 U14665 ( .IN1(n14753), .IN2(g1830), .QN(n14752) );
  NAND2X0 U14666 ( .IN1(n14730), .IN2(n11946), .QN(n14753) );
  NAND2X0 U14667 ( .IN1(n14731), .IN2(n11946), .QN(n14751) );
  NAND2X0 U14668 ( .IN1(n14754), .IN2(n14755), .QN(g27765) );
  NAND2X0 U14669 ( .IN1(n14756), .IN2(g1134), .QN(n14755) );
  NAND2X0 U14670 ( .IN1(n14757), .IN2(g1088), .QN(n14756) );
  NAND2X0 U14671 ( .IN1(n14758), .IN2(g1088), .QN(n14754) );
  NAND2X0 U14672 ( .IN1(n14759), .IN2(n14760), .QN(g27764) );
  NAND2X0 U14673 ( .IN1(n14761), .IN2(g1829), .QN(n14760) );
  NAND2X0 U14674 ( .IN1(n14730), .IN2(n13555), .QN(n14761) );
  NOR2X0 U14675 ( .IN1(n14762), .IN2(n14763), .QN(n14730) );
  NAND2X0 U14676 ( .IN1(n14764), .IN2(n14765), .QN(n14762) );
  INVX0 U14677 ( .INP(n14766), .ZN(n14765) );
  NAND2X0 U14678 ( .IN1(n11946), .IN2(n9981), .QN(n14764) );
  NAND2X0 U14679 ( .IN1(n14731), .IN2(n13555), .QN(n14759) );
  INVX0 U14680 ( .INP(n14767), .ZN(n14731) );
  NAND2X0 U14681 ( .IN1(n14768), .IN2(n14769), .QN(n14767) );
  NOR2X0 U14682 ( .IN1(n14770), .IN2(n14771), .QN(n14769) );
  NOR2X0 U14683 ( .IN1(n14772), .IN2(n14773), .QN(n14771) );
  NOR2X0 U14684 ( .IN1(n4386), .IN2(n14774), .QN(n14768) );
  NOR2X0 U14685 ( .IN1(n14775), .IN2(n14776), .QN(n14774) );
  NAND2X0 U14686 ( .IN1(n14777), .IN2(n14778), .QN(g27763) );
  NAND2X0 U14687 ( .IN1(n14779), .IN2(g1136), .QN(n14778) );
  NAND2X0 U14688 ( .IN1(n14757), .IN2(g6712), .QN(n14779) );
  NAND2X0 U14689 ( .IN1(n14758), .IN2(g6712), .QN(n14777) );
  NAND2X0 U14690 ( .IN1(n14780), .IN2(n14781), .QN(g27762) );
  NAND2X0 U14691 ( .IN1(n14782), .IN2(g447), .QN(n14781) );
  NAND2X0 U14692 ( .IN1(n14783), .IN2(n13361), .QN(n14782) );
  NAND2X0 U14693 ( .IN1(n14784), .IN2(n13361), .QN(n14780) );
  NAND2X0 U14694 ( .IN1(n14785), .IN2(n14786), .QN(g27761) );
  NAND2X0 U14695 ( .IN1(n14787), .IN2(g1135), .QN(n14786) );
  NAND2X0 U14696 ( .IN1(n14757), .IN2(g5472), .QN(n14787) );
  NOR2X0 U14697 ( .IN1(n14788), .IN2(n14789), .QN(n14757) );
  NAND2X0 U14698 ( .IN1(n14790), .IN2(n14791), .QN(n14788) );
  INVX0 U14699 ( .INP(n14792), .ZN(n14791) );
  NAND2X0 U14700 ( .IN1(g6712), .IN2(n9984), .QN(n14790) );
  NAND2X0 U14701 ( .IN1(n14758), .IN2(g5472), .QN(n14785) );
  INVX0 U14702 ( .INP(n14793), .ZN(n14758) );
  NAND2X0 U14703 ( .IN1(n14794), .IN2(n14795), .QN(n14793) );
  NOR2X0 U14704 ( .IN1(n14796), .IN2(n14797), .QN(n14795) );
  NOR2X0 U14705 ( .IN1(n14798), .IN2(n14799), .QN(n14797) );
  NOR2X0 U14706 ( .IN1(n4387), .IN2(n14800), .QN(n14794) );
  NOR2X0 U14707 ( .IN1(n14801), .IN2(n14802), .QN(n14800) );
  NAND2X0 U14708 ( .IN1(n14803), .IN2(n14804), .QN(g27760) );
  NAND2X0 U14709 ( .IN1(n14805), .IN2(g449), .QN(n14804) );
  NAND2X0 U14710 ( .IN1(n14783), .IN2(n13382), .QN(n14805) );
  NAND2X0 U14711 ( .IN1(n14784), .IN2(n13382), .QN(n14803) );
  NAND2X0 U14712 ( .IN1(n14806), .IN2(n14807), .QN(g27759) );
  NAND2X0 U14713 ( .IN1(n14808), .IN2(g448), .QN(n14807) );
  NAND2X0 U14714 ( .IN1(n14783), .IN2(n12042), .QN(n14808) );
  NOR2X0 U14715 ( .IN1(n14809), .IN2(n14810), .QN(n14783) );
  NAND2X0 U14716 ( .IN1(n14811), .IN2(n14812), .QN(n14809) );
  INVX0 U14717 ( .INP(n14813), .ZN(n14812) );
  NAND2X0 U14718 ( .IN1(n13361), .IN2(n10004), .QN(n14811) );
  NAND2X0 U14719 ( .IN1(n14784), .IN2(n12042), .QN(n14806) );
  INVX0 U14720 ( .INP(n14814), .ZN(n14784) );
  NAND2X0 U14721 ( .IN1(n14815), .IN2(n14816), .QN(n14814) );
  NOR2X0 U14722 ( .IN1(n14817), .IN2(n14818), .QN(n14816) );
  NOR2X0 U14723 ( .IN1(n14819), .IN2(n14820), .QN(n14818) );
  NOR2X0 U14724 ( .IN1(n4388), .IN2(n14821), .QN(n14815) );
  NOR2X0 U14725 ( .IN1(n14822), .IN2(n14823), .QN(n14821) );
  NOR2X0 U14726 ( .IN1(n14824), .IN2(n14825), .QN(g27724) );
  NAND2X0 U14727 ( .IN1(n14694), .IN2(n14826), .QN(n14825) );
  INVX0 U14728 ( .INP(n14695), .ZN(n14694) );
  NOR2X0 U14729 ( .IN1(n14827), .IN2(n4393), .QN(n14695) );
  NOR2X0 U14730 ( .IN1(n14828), .IN2(g2760), .QN(n14824) );
  INVX0 U14731 ( .INP(n14827), .ZN(n14828) );
  NOR2X0 U14732 ( .IN1(n14829), .IN2(n14699), .QN(g27722) );
  NAND2X0 U14733 ( .IN1(n14703), .IN2(n14830), .QN(n14699) );
  NAND2X0 U14734 ( .IN1(test_so70), .IN2(n14702), .QN(n14830) );
  NOR2X0 U14735 ( .IN1(n14702), .IN2(test_so70), .QN(n14829) );
  INVX0 U14736 ( .INP(n14831), .ZN(n14702) );
  NOR2X0 U14737 ( .IN1(n14832), .IN2(n14833), .QN(g27718) );
  NAND2X0 U14738 ( .IN1(n14708), .IN2(n14834), .QN(n14833) );
  INVX0 U14739 ( .INP(n14709), .ZN(n14708) );
  NOR2X0 U14740 ( .IN1(n14835), .IN2(n4395), .QN(n14709) );
  NOR2X0 U14741 ( .IN1(n14836), .IN2(g1372), .QN(n14832) );
  INVX0 U14742 ( .INP(n14835), .ZN(n14836) );
  NOR2X0 U14743 ( .IN1(n14837), .IN2(n14838), .QN(g27682) );
  NAND2X0 U14744 ( .IN1(n14831), .IN2(n14703), .QN(n14838) );
  NAND2X0 U14745 ( .IN1(n14839), .IN2(n14840), .QN(n14831) );
  NOR2X0 U14746 ( .IN1(n4473), .IN2(n4468), .QN(n14839) );
  NOR2X0 U14747 ( .IN1(n14841), .IN2(g2059), .QN(n14837) );
  NOR2X0 U14748 ( .IN1(n4468), .IN2(n14842), .QN(n14841) );
  NOR2X0 U14749 ( .IN1(n14843), .IN2(n14844), .QN(g27678) );
  NAND2X0 U14750 ( .IN1(n14835), .IN2(n14834), .QN(n14844) );
  NAND2X0 U14751 ( .IN1(n14845), .IN2(n14846), .QN(n14835) );
  NOR2X0 U14752 ( .IN1(n4475), .IN2(n4469), .QN(n14845) );
  NOR2X0 U14753 ( .IN1(n14847), .IN2(g1365), .QN(n14843) );
  NOR2X0 U14754 ( .IN1(n4469), .IN2(n14848), .QN(n14847) );
  NOR2X0 U14755 ( .IN1(n14849), .IN2(n14850), .QN(g27672) );
  NAND2X0 U14756 ( .IN1(n14713), .IN2(n14712), .QN(n14850) );
  NAND2X0 U14757 ( .IN1(n14851), .IN2(test_so28), .QN(n14713) );
  NOR2X0 U14758 ( .IN1(n4477), .IN2(n14852), .QN(n14851) );
  NOR2X0 U14759 ( .IN1(n14853), .IN2(g679), .QN(n14849) );
  NOR2X0 U14760 ( .IN1(n14852), .IN2(n10325), .QN(n14853) );
  NOR2X0 U14761 ( .IN1(n13263), .IN2(n14854), .QN(g27621) );
  NOR2X0 U14762 ( .IN1(n14855), .IN2(n14856), .QN(n14854) );
  NOR2X0 U14763 ( .IN1(n4522), .IN2(g2142), .QN(n14856) );
  NOR2X0 U14764 ( .IN1(n10011), .IN2(n14857), .QN(n14855) );
  NOR2X0 U14765 ( .IN1(n13268), .IN2(n14858), .QN(g27612) );
  NOR2X0 U14766 ( .IN1(n14859), .IN2(n14860), .QN(n14858) );
  NOR2X0 U14767 ( .IN1(n4523), .IN2(g1448), .QN(n14860) );
  NOR2X0 U14768 ( .IN1(n10015), .IN2(n14861), .QN(n14859) );
  NAND2X0 U14769 ( .IN1(n14862), .IN2(n14863), .QN(g27603) );
  NAND2X0 U14770 ( .IN1(n14864), .IN2(g762), .QN(n14863) );
  INVX0 U14771 ( .INP(n14865), .ZN(n14864) );
  NAND2X0 U14772 ( .IN1(n14866), .IN2(n10019), .QN(n14862) );
  NOR2X0 U14773 ( .IN1(n13273), .IN2(n3431), .QN(n14866) );
  NOR2X0 U14774 ( .IN1(n13278), .IN2(n14867), .QN(g27594) );
  NOR2X0 U14775 ( .IN1(n14868), .IN2(n14869), .QN(n14867) );
  NOR2X0 U14776 ( .IN1(n4521), .IN2(g74), .QN(n14869) );
  NOR2X0 U14777 ( .IN1(n10023), .IN2(n14870), .QN(n14868) );
  NAND2X0 U14778 ( .IN1(n14871), .IN2(n14872), .QN(g27380) );
  NOR2X0 U14779 ( .IN1(n14873), .IN2(n14874), .QN(n14872) );
  NAND2X0 U14780 ( .IN1(n14875), .IN2(n14876), .QN(n14874) );
  NAND2X0 U14781 ( .IN1(n14877), .IN2(n14878), .QN(n14876) );
  NAND2X0 U14782 ( .IN1(n14879), .IN2(n14880), .QN(n14878) );
  NAND2X0 U14783 ( .IN1(n14881), .IN2(n4384), .QN(n14880) );
  NOR2X0 U14784 ( .IN1(n4405), .IN2(n14882), .QN(n14881) );
  INVX0 U14785 ( .INP(n14883), .ZN(n14875) );
  NOR2X0 U14786 ( .IN1(n14884), .IN2(n4424), .QN(n14883) );
  NAND2X0 U14787 ( .IN1(n14885), .IN2(n14886), .QN(n14873) );
  NAND2X0 U14788 ( .IN1(n14887), .IN2(n14888), .QN(n14885) );
  NOR2X0 U14789 ( .IN1(n14889), .IN2(n14890), .QN(n14888) );
  NOR2X0 U14790 ( .IN1(n18868), .IN2(n14891), .QN(n14890) );
  NOR2X0 U14791 ( .IN1(n18869), .IN2(n14892), .QN(n14889) );
  NOR2X0 U14792 ( .IN1(n14893), .IN2(n14882), .QN(n14887) );
  NOR2X0 U14793 ( .IN1(n14894), .IN2(n14895), .QN(n14871) );
  NAND2X0 U14794 ( .IN1(n14896), .IN2(n14897), .QN(n14895) );
  INVX0 U14795 ( .INP(n14898), .ZN(n14897) );
  NOR2X0 U14796 ( .IN1(n14899), .IN2(n18870), .QN(n14898) );
  NAND2X0 U14797 ( .IN1(n9737), .IN2(n14900), .QN(n14896) );
  INVX0 U14798 ( .INP(n3700), .ZN(n14894) );
  NAND2X0 U14799 ( .IN1(n14901), .IN2(n14902), .QN(g27354) );
  NAND2X0 U14800 ( .IN1(n14903), .IN2(g2658), .QN(n14902) );
  NAND2X0 U14801 ( .IN1(n14904), .IN2(n14905), .QN(n14901) );
  NAND2X0 U14802 ( .IN1(n14906), .IN2(n14907), .QN(g27348) );
  NAND2X0 U14803 ( .IN1(n14908), .IN2(n14905), .QN(n14907) );
  INVX0 U14804 ( .INP(n14909), .ZN(n14906) );
  NOR2X0 U14805 ( .IN1(n14908), .IN2(n9642), .QN(n14909) );
  NAND2X0 U14806 ( .IN1(n14910), .IN2(n14911), .QN(g27347) );
  NAND2X0 U14807 ( .IN1(n14903), .IN2(g2655), .QN(n14911) );
  NAND2X0 U14808 ( .IN1(n14904), .IN2(n14912), .QN(n14910) );
  NAND2X0 U14809 ( .IN1(n14913), .IN2(n14914), .QN(g27346) );
  INVX0 U14810 ( .INP(n14915), .ZN(n14914) );
  NOR2X0 U14811 ( .IN1(n14916), .IN2(n9643), .QN(n14915) );
  NAND2X0 U14812 ( .IN1(n14916), .IN2(n14917), .QN(n14913) );
  NAND2X0 U14813 ( .IN1(n14918), .IN2(n14919), .QN(g27345) );
  NAND2X0 U14814 ( .IN1(n14920), .IN2(n14905), .QN(n14919) );
  NAND2X0 U14815 ( .IN1(n14275), .IN2(n14921), .QN(n14905) );
  NOR2X0 U14816 ( .IN1(n14248), .IN2(n14253), .QN(n14275) );
  NAND2X0 U14817 ( .IN1(n14922), .IN2(g2659), .QN(n14918) );
  NAND2X0 U14818 ( .IN1(n14923), .IN2(n14924), .QN(g27344) );
  NAND2X0 U14819 ( .IN1(test_so89), .IN2(n14925), .QN(n14924) );
  NAND2X0 U14820 ( .IN1(n14908), .IN2(n14912), .QN(n14923) );
  NAND2X0 U14821 ( .IN1(n14926), .IN2(n14927), .QN(g27343) );
  NAND2X0 U14822 ( .IN1(n14903), .IN2(g2652), .QN(n14927) );
  NAND2X0 U14823 ( .IN1(n14928), .IN2(n14904), .QN(n14926) );
  NAND2X0 U14824 ( .IN1(n14929), .IN2(n14930), .QN(g27342) );
  NAND2X0 U14825 ( .IN1(n14931), .IN2(g2466), .QN(n14930) );
  NAND2X0 U14826 ( .IN1(n14932), .IN2(n14933), .QN(n14929) );
  NAND2X0 U14827 ( .IN1(n14934), .IN2(n14935), .QN(g27341) );
  NAND2X0 U14828 ( .IN1(n14936), .IN2(n14917), .QN(n14935) );
  NAND2X0 U14829 ( .IN1(n14937), .IN2(g1966), .QN(n14934) );
  NAND2X0 U14830 ( .IN1(n14938), .IN2(n14939), .QN(g27340) );
  INVX0 U14831 ( .INP(n14940), .ZN(n14939) );
  NOR2X0 U14832 ( .IN1(n14916), .IN2(n9436), .QN(n14940) );
  NAND2X0 U14833 ( .IN1(n14916), .IN2(n14941), .QN(n14938) );
  NAND2X0 U14834 ( .IN1(n14942), .IN2(n14943), .QN(g27339) );
  NAND2X0 U14835 ( .IN1(n14944), .IN2(g1270), .QN(n14943) );
  NAND2X0 U14836 ( .IN1(n14945), .IN2(n14946), .QN(n14942) );
  NAND2X0 U14837 ( .IN1(n14947), .IN2(n14948), .QN(g27338) );
  NAND2X0 U14838 ( .IN1(n14922), .IN2(g2656), .QN(n14948) );
  NAND2X0 U14839 ( .IN1(n14920), .IN2(n14912), .QN(n14947) );
  INVX0 U14840 ( .INP(n14949), .ZN(n14912) );
  NAND2X0 U14841 ( .IN1(n14950), .IN2(n14951), .QN(n14949) );
  NAND2X0 U14842 ( .IN1(n14952), .IN2(n14282), .QN(n14951) );
  NOR2X0 U14843 ( .IN1(n14253), .IN2(n14953), .QN(n14282) );
  NAND2X0 U14844 ( .IN1(n14921), .IN2(n14253), .QN(n14950) );
  NAND2X0 U14845 ( .IN1(n14954), .IN2(n14955), .QN(g27337) );
  INVX0 U14846 ( .INP(n14956), .ZN(n14955) );
  NOR2X0 U14847 ( .IN1(n14908), .IN2(n9627), .QN(n14956) );
  NAND2X0 U14848 ( .IN1(n14928), .IN2(n14908), .QN(n14954) );
  NAND2X0 U14849 ( .IN1(n14957), .IN2(n14958), .QN(g27336) );
  NAND2X0 U14850 ( .IN1(n14903), .IN2(g2649), .QN(n14958) );
  NAND2X0 U14851 ( .IN1(n14959), .IN2(n14904), .QN(n14957) );
  INVX0 U14852 ( .INP(n14903), .ZN(n14904) );
  NAND2X0 U14853 ( .IN1(g2624), .IN2(g22687), .QN(n14903) );
  NAND2X0 U14854 ( .IN1(n14960), .IN2(n14961), .QN(g27335) );
  NAND2X0 U14855 ( .IN1(n14962), .IN2(n14933), .QN(n14961) );
  INVX0 U14856 ( .INP(n14963), .ZN(n14960) );
  NOR2X0 U14857 ( .IN1(n14962), .IN2(n9956), .QN(n14963) );
  NAND2X0 U14858 ( .IN1(n14964), .IN2(n14965), .QN(g27334) );
  NAND2X0 U14859 ( .IN1(n14931), .IN2(g2451), .QN(n14965) );
  NAND2X0 U14860 ( .IN1(n14932), .IN2(n14966), .QN(n14964) );
  NAND2X0 U14861 ( .IN1(n14967), .IN2(n14968), .QN(g27333) );
  NAND2X0 U14862 ( .IN1(n14969), .IN2(n14917), .QN(n14968) );
  NAND2X0 U14863 ( .IN1(n14405), .IN2(n14970), .QN(n14917) );
  NOR2X0 U14864 ( .IN1(n14379), .IN2(n14384), .QN(n14405) );
  NAND2X0 U14865 ( .IN1(test_so67), .IN2(n14971), .QN(n14967) );
  NAND2X0 U14866 ( .IN1(n14972), .IN2(n14973), .QN(g27332) );
  NAND2X0 U14867 ( .IN1(n14937), .IN2(g1963), .QN(n14973) );
  NAND2X0 U14868 ( .IN1(n14936), .IN2(n14941), .QN(n14972) );
  NAND2X0 U14869 ( .IN1(n14974), .IN2(n14975), .QN(g27331) );
  INVX0 U14870 ( .INP(n14976), .ZN(n14975) );
  NOR2X0 U14871 ( .IN1(n14916), .IN2(n9629), .QN(n14976) );
  NAND2X0 U14872 ( .IN1(n14977), .IN2(n14916), .QN(n14974) );
  NAND2X0 U14873 ( .IN1(n14978), .IN2(n14979), .QN(g27330) );
  NAND2X0 U14874 ( .IN1(n14980), .IN2(g1772), .QN(n14979) );
  NAND2X0 U14875 ( .IN1(n14981), .IN2(n14982), .QN(n14978) );
  NAND2X0 U14876 ( .IN1(n14983), .IN2(n14984), .QN(g27329) );
  NAND2X0 U14877 ( .IN1(n14985), .IN2(n14946), .QN(n14984) );
  NAND2X0 U14878 ( .IN1(n14986), .IN2(g1272), .QN(n14983) );
  NAND2X0 U14879 ( .IN1(n14987), .IN2(n14988), .QN(g27328) );
  NAND2X0 U14880 ( .IN1(test_so46), .IN2(n14944), .QN(n14988) );
  NAND2X0 U14881 ( .IN1(n14945), .IN2(n14989), .QN(n14987) );
  NAND2X0 U14882 ( .IN1(n14990), .IN2(n14991), .QN(g27327) );
  NAND2X0 U14883 ( .IN1(n14992), .IN2(g584), .QN(n14991) );
  NAND2X0 U14884 ( .IN1(n14993), .IN2(n14994), .QN(n14990) );
  NAND2X0 U14885 ( .IN1(n14995), .IN2(n14996), .QN(g27326) );
  NAND2X0 U14886 ( .IN1(n14922), .IN2(g2653), .QN(n14996) );
  NAND2X0 U14887 ( .IN1(n14928), .IN2(n14920), .QN(n14995) );
  NOR2X0 U14888 ( .IN1(n14997), .IN2(n14998), .QN(n14928) );
  NOR2X0 U14889 ( .IN1(n14921), .IN2(n14238), .QN(n14998) );
  INVX0 U14890 ( .INP(n14952), .ZN(n14921) );
  NAND2X0 U14891 ( .IN1(n14999), .IN2(n15000), .QN(n14952) );
  NAND2X0 U14892 ( .IN1(g3229), .IN2(n14233), .QN(n15000) );
  NAND2X0 U14893 ( .IN1(n14224), .IN2(n11195), .QN(n14999) );
  INVX0 U14894 ( .INP(n14233), .ZN(n14224) );
  NAND2X0 U14895 ( .IN1(n15001), .IN2(n15002), .QN(g27325) );
  INVX0 U14896 ( .INP(n15003), .ZN(n15002) );
  NOR2X0 U14897 ( .IN1(n14908), .IN2(n9607), .QN(n15003) );
  NAND2X0 U14898 ( .IN1(n14959), .IN2(n14908), .QN(n15001) );
  INVX0 U14899 ( .INP(n14925), .ZN(n14908) );
  NAND2X0 U14900 ( .IN1(g7390), .IN2(g22687), .QN(n14925) );
  NAND2X0 U14901 ( .IN1(n15004), .IN2(n15005), .QN(g27324) );
  NAND2X0 U14902 ( .IN1(n15006), .IN2(n14933), .QN(n15005) );
  NAND2X0 U14903 ( .IN1(n15007), .IN2(n15008), .QN(n14933) );
  NOR2X0 U14904 ( .IN1(n15009), .IN2(n15010), .QN(n15007) );
  NAND2X0 U14905 ( .IN1(n15011), .IN2(g2473), .QN(n15004) );
  NAND2X0 U14906 ( .IN1(n15012), .IN2(n15013), .QN(g27323) );
  INVX0 U14907 ( .INP(n15014), .ZN(n15013) );
  NOR2X0 U14908 ( .IN1(n14962), .IN2(n9678), .QN(n15014) );
  NAND2X0 U14909 ( .IN1(n14962), .IN2(n14966), .QN(n15012) );
  NAND2X0 U14910 ( .IN1(n15015), .IN2(n15016), .QN(g27322) );
  NAND2X0 U14911 ( .IN1(n15017), .IN2(n14932), .QN(n15016) );
  NAND2X0 U14912 ( .IN1(n14931), .IN2(g2436), .QN(n15015) );
  NAND2X0 U14913 ( .IN1(n15018), .IN2(n15019), .QN(g27321) );
  NAND2X0 U14914 ( .IN1(n14971), .IN2(g1962), .QN(n15019) );
  NAND2X0 U14915 ( .IN1(n14969), .IN2(n14941), .QN(n15018) );
  INVX0 U14916 ( .INP(n15020), .ZN(n14941) );
  NAND2X0 U14917 ( .IN1(n15021), .IN2(n15022), .QN(n15020) );
  NAND2X0 U14918 ( .IN1(n15023), .IN2(n14412), .QN(n15022) );
  NOR2X0 U14919 ( .IN1(n14384), .IN2(n15024), .QN(n14412) );
  NAND2X0 U14920 ( .IN1(n14970), .IN2(n14384), .QN(n15021) );
  NAND2X0 U14921 ( .IN1(n15025), .IN2(n15026), .QN(g27320) );
  NAND2X0 U14922 ( .IN1(n14937), .IN2(g1960), .QN(n15026) );
  NAND2X0 U14923 ( .IN1(n14977), .IN2(n14936), .QN(n15025) );
  NAND2X0 U14924 ( .IN1(n15027), .IN2(n15028), .QN(g27319) );
  INVX0 U14925 ( .INP(n15029), .ZN(n15028) );
  NOR2X0 U14926 ( .IN1(n14916), .IN2(n9609), .QN(n15029) );
  NAND2X0 U14927 ( .IN1(n15030), .IN2(n14916), .QN(n15027) );
  INVX0 U14928 ( .INP(n15031), .ZN(n14916) );
  NAND2X0 U14929 ( .IN1(g1930), .IN2(g22651), .QN(n15031) );
  NAND2X0 U14930 ( .IN1(n15032), .IN2(n15033), .QN(g27318) );
  NAND2X0 U14931 ( .IN1(n15034), .IN2(n14982), .QN(n15033) );
  NAND2X0 U14932 ( .IN1(test_so58), .IN2(n15035), .QN(n15032) );
  NAND2X0 U14933 ( .IN1(n15036), .IN2(n15037), .QN(g27317) );
  NAND2X0 U14934 ( .IN1(n14980), .IN2(g1757), .QN(n15037) );
  NAND2X0 U14935 ( .IN1(n14981), .IN2(n15038), .QN(n15036) );
  NAND2X0 U14936 ( .IN1(n15039), .IN2(n15040), .QN(g27316) );
  NAND2X0 U14937 ( .IN1(n15041), .IN2(n14946), .QN(n15040) );
  NAND2X0 U14938 ( .IN1(n14528), .IN2(n15042), .QN(n14946) );
  NOR2X0 U14939 ( .IN1(n14502), .IN2(n14507), .QN(n14528) );
  INVX0 U14940 ( .INP(n15043), .ZN(n15039) );
  NOR2X0 U14941 ( .IN1(n15041), .IN2(n9645), .QN(n15043) );
  NAND2X0 U14942 ( .IN1(n15044), .IN2(n15045), .QN(g27315) );
  NAND2X0 U14943 ( .IN1(n14986), .IN2(g1269), .QN(n15045) );
  NAND2X0 U14944 ( .IN1(n14985), .IN2(n14989), .QN(n15044) );
  NAND2X0 U14945 ( .IN1(n15046), .IN2(n15047), .QN(g27314) );
  NAND2X0 U14946 ( .IN1(n14944), .IN2(g1264), .QN(n15047) );
  NAND2X0 U14947 ( .IN1(n15048), .IN2(n14945), .QN(n15046) );
  NAND2X0 U14948 ( .IN1(n15049), .IN2(n15050), .QN(g27313) );
  INVX0 U14949 ( .INP(n15051), .ZN(n15050) );
  NOR2X0 U14950 ( .IN1(n15052), .IN2(n9960), .QN(n15051) );
  NAND2X0 U14951 ( .IN1(n15052), .IN2(n15053), .QN(n15049) );
  NAND2X0 U14952 ( .IN1(n15054), .IN2(n15055), .QN(g27312) );
  NAND2X0 U14953 ( .IN1(n15056), .IN2(n14994), .QN(n15055) );
  INVX0 U14954 ( .INP(n15057), .ZN(n15054) );
  NOR2X0 U14955 ( .IN1(n15056), .IN2(n9650), .QN(n15057) );
  NAND2X0 U14956 ( .IN1(n15058), .IN2(n15059), .QN(g27311) );
  NAND2X0 U14957 ( .IN1(n14992), .IN2(g581), .QN(n15059) );
  NAND2X0 U14958 ( .IN1(n14993), .IN2(n15060), .QN(n15058) );
  NAND2X0 U14959 ( .IN1(n15061), .IN2(n15062), .QN(g27310) );
  NAND2X0 U14960 ( .IN1(n14922), .IN2(g2650), .QN(n15062) );
  NAND2X0 U14961 ( .IN1(n14959), .IN2(n14920), .QN(n15061) );
  INVX0 U14962 ( .INP(n14922), .ZN(n14920) );
  NAND2X0 U14963 ( .IN1(g7302), .IN2(g22687), .QN(n14922) );
  INVX0 U14964 ( .INP(n15063), .ZN(n14959) );
  NAND2X0 U14965 ( .IN1(n15064), .IN2(n15065), .QN(n15063) );
  NAND2X0 U14966 ( .IN1(g3229), .IN2(n14953), .QN(n15065) );
  NOR2X0 U14967 ( .IN1(n15066), .IN2(n15067), .QN(n15064) );
  NOR2X0 U14968 ( .IN1(n14997), .IN2(n15068), .QN(n15067) );
  NAND2X0 U14969 ( .IN1(n14240), .IN2(n14233), .QN(n15068) );
  NAND2X0 U14970 ( .IN1(n15069), .IN2(n15070), .QN(n14233) );
  NAND2X0 U14971 ( .IN1(n9607), .IN2(g7390), .QN(n15070) );
  NOR2X0 U14972 ( .IN1(n15071), .IN2(n15072), .QN(n15069) );
  NOR2X0 U14973 ( .IN1(n4314), .IN2(g2650), .QN(n15072) );
  NOR2X0 U14974 ( .IN1(n4299), .IN2(g2649), .QN(n15071) );
  INVX0 U14975 ( .INP(n14953), .ZN(n14240) );
  NAND2X0 U14976 ( .IN1(n15073), .IN2(n15074), .QN(n14953) );
  NAND2X0 U14977 ( .IN1(n9642), .IN2(g7390), .QN(n15074) );
  NOR2X0 U14978 ( .IN1(n15075), .IN2(n15076), .QN(n15073) );
  NOR2X0 U14979 ( .IN1(n4314), .IN2(g2659), .QN(n15076) );
  NOR2X0 U14980 ( .IN1(n4299), .IN2(g2658), .QN(n15075) );
  INVX0 U14981 ( .INP(n15077), .ZN(n14997) );
  NOR2X0 U14982 ( .IN1(g3229), .IN2(n15077), .QN(n15066) );
  NAND2X0 U14983 ( .IN1(n14238), .IN2(n14253), .QN(n15077) );
  NAND2X0 U14984 ( .IN1(n15078), .IN2(n15079), .QN(n14253) );
  NAND2X0 U14985 ( .IN1(n9627), .IN2(g7390), .QN(n15079) );
  NOR2X0 U14986 ( .IN1(n15080), .IN2(n15081), .QN(n15078) );
  NOR2X0 U14987 ( .IN1(n4314), .IN2(g2653), .QN(n15081) );
  NOR2X0 U14988 ( .IN1(n4299), .IN2(g2652), .QN(n15080) );
  INVX0 U14989 ( .INP(n14248), .ZN(n14238) );
  NAND2X0 U14990 ( .IN1(n15082), .IN2(n15083), .QN(n14248) );
  NAND2X0 U14991 ( .IN1(g7390), .IN2(n10332), .QN(n15083) );
  NOR2X0 U14992 ( .IN1(n15084), .IN2(n15085), .QN(n15082) );
  NOR2X0 U14993 ( .IN1(n4314), .IN2(g2656), .QN(n15085) );
  NOR2X0 U14994 ( .IN1(n4299), .IN2(g2655), .QN(n15084) );
  NAND2X0 U14995 ( .IN1(n15086), .IN2(n15087), .QN(g27309) );
  NAND2X0 U14996 ( .IN1(n15011), .IN2(g2459), .QN(n15087) );
  NAND2X0 U14997 ( .IN1(n15006), .IN2(n14966), .QN(n15086) );
  INVX0 U14998 ( .INP(n15088), .ZN(n14966) );
  NAND2X0 U14999 ( .IN1(n15089), .IN2(n15090), .QN(n15088) );
  NAND2X0 U15000 ( .IN1(n15091), .IN2(n15009), .QN(n15090) );
  NAND2X0 U15001 ( .IN1(n15092), .IN2(n15093), .QN(n15089) );
  NOR2X0 U15002 ( .IN1(n15091), .IN2(n15094), .QN(n15092) );
  INVX0 U15003 ( .INP(n15010), .ZN(n15091) );
  NAND2X0 U15004 ( .IN1(n15095), .IN2(n15096), .QN(n15010) );
  NAND2X0 U15005 ( .IN1(g3229), .IN2(n15097), .QN(n15096) );
  NAND2X0 U15006 ( .IN1(n15098), .IN2(n11195), .QN(n15095) );
  NAND2X0 U15007 ( .IN1(n15099), .IN2(n15100), .QN(g27308) );
  NAND2X0 U15008 ( .IN1(n15017), .IN2(n14962), .QN(n15100) );
  INVX0 U15009 ( .INP(n15101), .ZN(n15099) );
  NOR2X0 U15010 ( .IN1(n14962), .IN2(n9944), .QN(n15101) );
  NAND2X0 U15011 ( .IN1(n15102), .IN2(n15103), .QN(g27307) );
  NAND2X0 U15012 ( .IN1(n14931), .IN2(g2421), .QN(n15103) );
  NAND2X0 U15013 ( .IN1(n15104), .IN2(n14932), .QN(n15102) );
  INVX0 U15014 ( .INP(n14931), .ZN(n14932) );
  NAND2X0 U15015 ( .IN1(n15105), .IN2(n13307), .QN(n14931) );
  NAND2X0 U15016 ( .IN1(n15106), .IN2(n15107), .QN(g27306) );
  NAND2X0 U15017 ( .IN1(n14971), .IN2(g1959), .QN(n15107) );
  NAND2X0 U15018 ( .IN1(n14977), .IN2(n14969), .QN(n15106) );
  NOR2X0 U15019 ( .IN1(n15108), .IN2(n15109), .QN(n14977) );
  NOR2X0 U15020 ( .IN1(n14970), .IN2(n14369), .QN(n15109) );
  INVX0 U15021 ( .INP(n15023), .ZN(n14970) );
  NAND2X0 U15022 ( .IN1(n15110), .IN2(n15111), .QN(n15023) );
  NAND2X0 U15023 ( .IN1(g3229), .IN2(n14364), .QN(n15111) );
  NAND2X0 U15024 ( .IN1(n14355), .IN2(n11195), .QN(n15110) );
  INVX0 U15025 ( .INP(n14364), .ZN(n14355) );
  NAND2X0 U15026 ( .IN1(n15112), .IN2(n15113), .QN(g27305) );
  NAND2X0 U15027 ( .IN1(n14937), .IN2(g1957), .QN(n15113) );
  NAND2X0 U15028 ( .IN1(n15030), .IN2(n14936), .QN(n15112) );
  INVX0 U15029 ( .INP(n14937), .ZN(n14936) );
  NAND2X0 U15030 ( .IN1(g7194), .IN2(g22651), .QN(n14937) );
  NAND2X0 U15031 ( .IN1(n15114), .IN2(n15115), .QN(g27304) );
  NAND2X0 U15032 ( .IN1(n15116), .IN2(n14982), .QN(n15115) );
  NAND2X0 U15033 ( .IN1(n15117), .IN2(n15118), .QN(n14982) );
  NOR2X0 U15034 ( .IN1(n15119), .IN2(n15120), .QN(n15117) );
  NAND2X0 U15035 ( .IN1(n15121), .IN2(g1779), .QN(n15114) );
  NAND2X0 U15036 ( .IN1(n15122), .IN2(n15123), .QN(g27303) );
  INVX0 U15037 ( .INP(n15124), .ZN(n15123) );
  NOR2X0 U15038 ( .IN1(n15034), .IN2(n9681), .QN(n15124) );
  NAND2X0 U15039 ( .IN1(n15034), .IN2(n15038), .QN(n15122) );
  NAND2X0 U15040 ( .IN1(n15125), .IN2(n15126), .QN(g27302) );
  NAND2X0 U15041 ( .IN1(n15127), .IN2(n14981), .QN(n15126) );
  NAND2X0 U15042 ( .IN1(n14980), .IN2(g1742), .QN(n15125) );
  NAND2X0 U15043 ( .IN1(n15128), .IN2(n15129), .QN(g27301) );
  INVX0 U15044 ( .INP(n15130), .ZN(n15129) );
  NOR2X0 U15045 ( .IN1(n15041), .IN2(n9438), .QN(n15130) );
  NAND2X0 U15046 ( .IN1(n15041), .IN2(n14989), .QN(n15128) );
  INVX0 U15047 ( .INP(n15131), .ZN(n14989) );
  NAND2X0 U15048 ( .IN1(n15132), .IN2(n15133), .QN(n15131) );
  NAND2X0 U15049 ( .IN1(n15134), .IN2(n14535), .QN(n15133) );
  NOR2X0 U15050 ( .IN1(n14507), .IN2(n15135), .QN(n14535) );
  NAND2X0 U15051 ( .IN1(n15042), .IN2(n14507), .QN(n15132) );
  NAND2X0 U15052 ( .IN1(n15136), .IN2(n15137), .QN(g27300) );
  NAND2X0 U15053 ( .IN1(n14986), .IN2(g1266), .QN(n15137) );
  NAND2X0 U15054 ( .IN1(n15048), .IN2(n14985), .QN(n15136) );
  NAND2X0 U15055 ( .IN1(n15138), .IN2(n15139), .QN(g27299) );
  NAND2X0 U15056 ( .IN1(n14944), .IN2(g1261), .QN(n15139) );
  NAND2X0 U15057 ( .IN1(n15140), .IN2(n14945), .QN(n15138) );
  INVX0 U15058 ( .INP(n14944), .ZN(n14945) );
  NAND2X0 U15059 ( .IN1(g1236), .IN2(g22615), .QN(n14944) );
  NAND2X0 U15060 ( .IN1(n15141), .IN2(n15142), .QN(g27298) );
  NAND2X0 U15061 ( .IN1(n15143), .IN2(n15053), .QN(n15142) );
  NAND2X0 U15062 ( .IN1(n15144), .IN2(g1075), .QN(n15141) );
  NAND2X0 U15063 ( .IN1(n15145), .IN2(n15146), .QN(g27297) );
  INVX0 U15064 ( .INP(n15147), .ZN(n15146) );
  NOR2X0 U15065 ( .IN1(n15052), .IN2(n9683), .QN(n15147) );
  NAND2X0 U15066 ( .IN1(n15052), .IN2(n15148), .QN(n15145) );
  NAND2X0 U15067 ( .IN1(n15149), .IN2(n15150), .QN(g27296) );
  NAND2X0 U15068 ( .IN1(n15151), .IN2(n14994), .QN(n15150) );
  NAND2X0 U15069 ( .IN1(n14647), .IN2(n15152), .QN(n14994) );
  NOR2X0 U15070 ( .IN1(n14621), .IN2(n14626), .QN(n14647) );
  NAND2X0 U15071 ( .IN1(n15153), .IN2(g585), .QN(n15149) );
  NAND2X0 U15072 ( .IN1(n15154), .IN2(n15155), .QN(g27295) );
  INVX0 U15073 ( .INP(n15156), .ZN(n15155) );
  NOR2X0 U15074 ( .IN1(n15056), .IN2(n9442), .QN(n15156) );
  NAND2X0 U15075 ( .IN1(n15056), .IN2(n15060), .QN(n15154) );
  NAND2X0 U15076 ( .IN1(n15157), .IN2(n15158), .QN(g27294) );
  NAND2X0 U15077 ( .IN1(n14992), .IN2(g578), .QN(n15158) );
  NAND2X0 U15078 ( .IN1(n15159), .IN2(n14993), .QN(n15157) );
  NAND2X0 U15079 ( .IN1(n15160), .IN2(n15161), .QN(g27293) );
  NAND2X0 U15080 ( .IN1(n15162), .IN2(g391), .QN(n15161) );
  NAND2X0 U15081 ( .IN1(n15163), .IN2(n15164), .QN(n15160) );
  NAND2X0 U15082 ( .IN1(n15165), .IN2(n15166), .QN(g27292) );
  NAND2X0 U15083 ( .IN1(n15017), .IN2(n15006), .QN(n15166) );
  INVX0 U15084 ( .INP(n15167), .ZN(n15017) );
  NAND2X0 U15085 ( .IN1(n15168), .IN2(n15169), .QN(n15167) );
  NAND2X0 U15086 ( .IN1(n15170), .IN2(n15098), .QN(n15169) );
  INVX0 U15087 ( .INP(n15097), .ZN(n15098) );
  NOR2X0 U15088 ( .IN1(g3229), .IN2(n15008), .QN(n15170) );
  INVX0 U15089 ( .INP(n15171), .ZN(n15008) );
  NOR2X0 U15090 ( .IN1(n15172), .IN2(n15173), .QN(n15168) );
  NAND2X0 U15091 ( .IN1(n15011), .IN2(g2444), .QN(n15165) );
  NAND2X0 U15092 ( .IN1(n15174), .IN2(n15175), .QN(g27291) );
  INVX0 U15093 ( .INP(n15176), .ZN(n15175) );
  NOR2X0 U15094 ( .IN1(n14962), .IN2(n9967), .QN(n15176) );
  NAND2X0 U15095 ( .IN1(n15104), .IN2(n14962), .QN(n15174) );
  INVX0 U15096 ( .INP(n15177), .ZN(n14962) );
  NAND2X0 U15097 ( .IN1(n15105), .IN2(g7264), .QN(n15177) );
  NAND2X0 U15098 ( .IN1(n15178), .IN2(n15179), .QN(g27290) );
  NAND2X0 U15099 ( .IN1(n14971), .IN2(g1956), .QN(n15179) );
  NAND2X0 U15100 ( .IN1(n15030), .IN2(n14969), .QN(n15178) );
  INVX0 U15101 ( .INP(n14971), .ZN(n14969) );
  NAND2X0 U15102 ( .IN1(g7052), .IN2(g22651), .QN(n14971) );
  INVX0 U15103 ( .INP(n15180), .ZN(n15030) );
  NAND2X0 U15104 ( .IN1(n15181), .IN2(n15182), .QN(n15180) );
  NAND2X0 U15105 ( .IN1(g3229), .IN2(n15024), .QN(n15182) );
  NOR2X0 U15106 ( .IN1(n15183), .IN2(n15184), .QN(n15181) );
  NOR2X0 U15107 ( .IN1(n15108), .IN2(n15185), .QN(n15184) );
  NAND2X0 U15108 ( .IN1(n14371), .IN2(n14364), .QN(n15185) );
  NAND2X0 U15109 ( .IN1(n15186), .IN2(n15187), .QN(n14364) );
  NAND2X0 U15110 ( .IN1(n9609), .IN2(g1930), .QN(n15187) );
  NOR2X0 U15111 ( .IN1(n15188), .IN2(n15189), .QN(n15186) );
  NOR2X0 U15112 ( .IN1(n4315), .IN2(g1957), .QN(n15189) );
  NOR2X0 U15113 ( .IN1(n4296), .IN2(g1956), .QN(n15188) );
  INVX0 U15114 ( .INP(n15024), .ZN(n14371) );
  NAND2X0 U15115 ( .IN1(n15190), .IN2(n15191), .QN(n15024) );
  NAND2X0 U15116 ( .IN1(n9643), .IN2(g1930), .QN(n15191) );
  NOR2X0 U15117 ( .IN1(n15192), .IN2(n15193), .QN(n15190) );
  NOR2X0 U15118 ( .IN1(n4315), .IN2(g1966), .QN(n15193) );
  NOR2X0 U15119 ( .IN1(test_so67), .IN2(n4296), .QN(n15192) );
  INVX0 U15120 ( .INP(n15194), .ZN(n15108) );
  NOR2X0 U15121 ( .IN1(g3229), .IN2(n15194), .QN(n15183) );
  NAND2X0 U15122 ( .IN1(n14369), .IN2(n14384), .QN(n15194) );
  NAND2X0 U15123 ( .IN1(n15195), .IN2(n15196), .QN(n14384) );
  NAND2X0 U15124 ( .IN1(n9629), .IN2(g1930), .QN(n15196) );
  NOR2X0 U15125 ( .IN1(n15197), .IN2(n15198), .QN(n15195) );
  NOR2X0 U15126 ( .IN1(n4315), .IN2(g1960), .QN(n15198) );
  NOR2X0 U15127 ( .IN1(n4296), .IN2(g1959), .QN(n15197) );
  INVX0 U15128 ( .INP(n14379), .ZN(n14369) );
  NAND2X0 U15129 ( .IN1(n15199), .IN2(n15200), .QN(n14379) );
  NAND2X0 U15130 ( .IN1(n9436), .IN2(g1930), .QN(n15200) );
  NOR2X0 U15131 ( .IN1(n15201), .IN2(n15202), .QN(n15199) );
  NOR2X0 U15132 ( .IN1(n4315), .IN2(g1963), .QN(n15202) );
  NOR2X0 U15133 ( .IN1(n4296), .IN2(g1962), .QN(n15201) );
  NAND2X0 U15134 ( .IN1(n15203), .IN2(n15204), .QN(g27289) );
  NAND2X0 U15135 ( .IN1(n15121), .IN2(g1765), .QN(n15204) );
  NAND2X0 U15136 ( .IN1(n15116), .IN2(n15038), .QN(n15203) );
  INVX0 U15137 ( .INP(n15205), .ZN(n15038) );
  NAND2X0 U15138 ( .IN1(n15206), .IN2(n15207), .QN(n15205) );
  NAND2X0 U15139 ( .IN1(n15208), .IN2(n15119), .QN(n15207) );
  NAND2X0 U15140 ( .IN1(n15209), .IN2(n15210), .QN(n15206) );
  INVX0 U15141 ( .INP(n15119), .ZN(n15210) );
  NOR2X0 U15142 ( .IN1(n15208), .IN2(n15211), .QN(n15209) );
  INVX0 U15143 ( .INP(n15120), .ZN(n15208) );
  NAND2X0 U15144 ( .IN1(n15212), .IN2(n15213), .QN(n15120) );
  NAND2X0 U15145 ( .IN1(g3229), .IN2(n15214), .QN(n15213) );
  NAND2X0 U15146 ( .IN1(n15215), .IN2(n11195), .QN(n15212) );
  NAND2X0 U15147 ( .IN1(n15216), .IN2(n15217), .QN(g27288) );
  NAND2X0 U15148 ( .IN1(n15127), .IN2(n15034), .QN(n15217) );
  INVX0 U15149 ( .INP(n15218), .ZN(n15216) );
  NOR2X0 U15150 ( .IN1(n15034), .IN2(n9947), .QN(n15218) );
  NAND2X0 U15151 ( .IN1(n15219), .IN2(n15220), .QN(g27287) );
  NAND2X0 U15152 ( .IN1(n14980), .IN2(g1727), .QN(n15220) );
  NAND2X0 U15153 ( .IN1(n15221), .IN2(n14981), .QN(n15219) );
  INVX0 U15154 ( .INP(n14980), .ZN(n14981) );
  NAND2X0 U15155 ( .IN1(n15222), .IN2(n13315), .QN(n14980) );
  NAND2X0 U15156 ( .IN1(n15223), .IN2(n15224), .QN(g27286) );
  INVX0 U15157 ( .INP(n15225), .ZN(n15224) );
  NOR2X0 U15158 ( .IN1(n15041), .IN2(n9631), .QN(n15225) );
  NAND2X0 U15159 ( .IN1(n15048), .IN2(n15041), .QN(n15223) );
  NOR2X0 U15160 ( .IN1(n15226), .IN2(n15227), .QN(n15048) );
  NOR2X0 U15161 ( .IN1(n15042), .IN2(n14492), .QN(n15227) );
  INVX0 U15162 ( .INP(n15134), .ZN(n15042) );
  NAND2X0 U15163 ( .IN1(n15228), .IN2(n15229), .QN(n15134) );
  NAND2X0 U15164 ( .IN1(g3229), .IN2(n14487), .QN(n15229) );
  NAND2X0 U15165 ( .IN1(n14478), .IN2(n11195), .QN(n15228) );
  INVX0 U15166 ( .INP(n14487), .ZN(n14478) );
  NAND2X0 U15167 ( .IN1(n15230), .IN2(n15231), .QN(g27285) );
  NAND2X0 U15168 ( .IN1(n14986), .IN2(g1263), .QN(n15231) );
  NAND2X0 U15169 ( .IN1(n15140), .IN2(n14985), .QN(n15230) );
  INVX0 U15170 ( .INP(n14986), .ZN(n14985) );
  NAND2X0 U15171 ( .IN1(g6944), .IN2(g22615), .QN(n14986) );
  NAND2X0 U15172 ( .IN1(n15232), .IN2(n15233), .QN(g27284) );
  NAND2X0 U15173 ( .IN1(n15234), .IN2(n15053), .QN(n15233) );
  NAND2X0 U15174 ( .IN1(n15235), .IN2(n15236), .QN(n15053) );
  NOR2X0 U15175 ( .IN1(n15237), .IN2(n15238), .QN(n15235) );
  NAND2X0 U15176 ( .IN1(n15239), .IN2(g1085), .QN(n15232) );
  NAND2X0 U15177 ( .IN1(n15240), .IN2(n15241), .QN(g27283) );
  NAND2X0 U15178 ( .IN1(n15144), .IN2(g1060), .QN(n15241) );
  NAND2X0 U15179 ( .IN1(n15143), .IN2(n15148), .QN(n15240) );
  NAND2X0 U15180 ( .IN1(n15242), .IN2(n15243), .QN(g27282) );
  NAND2X0 U15181 ( .IN1(n15244), .IN2(n15052), .QN(n15243) );
  INVX0 U15182 ( .INP(n15245), .ZN(n15242) );
  NOR2X0 U15183 ( .IN1(n15052), .IN2(n9949), .QN(n15245) );
  NAND2X0 U15184 ( .IN1(n15246), .IN2(n15247), .QN(g27281) );
  NAND2X0 U15185 ( .IN1(n15153), .IN2(g582), .QN(n15247) );
  NAND2X0 U15186 ( .IN1(n15151), .IN2(n15060), .QN(n15246) );
  INVX0 U15187 ( .INP(n15248), .ZN(n15060) );
  NAND2X0 U15188 ( .IN1(n15249), .IN2(n15250), .QN(n15248) );
  NAND2X0 U15189 ( .IN1(n15251), .IN2(n14654), .QN(n15250) );
  NOR2X0 U15190 ( .IN1(n14626), .IN2(n15252), .QN(n14654) );
  NAND2X0 U15191 ( .IN1(n15152), .IN2(n14626), .QN(n15249) );
  NAND2X0 U15192 ( .IN1(n15253), .IN2(n15254), .QN(g27280) );
  NAND2X0 U15193 ( .IN1(test_so25), .IN2(n15255), .QN(n15254) );
  NAND2X0 U15194 ( .IN1(n15159), .IN2(n15056), .QN(n15253) );
  NAND2X0 U15195 ( .IN1(n15256), .IN2(n15257), .QN(g27279) );
  NAND2X0 U15196 ( .IN1(n14992), .IN2(g575), .QN(n15257) );
  NAND2X0 U15197 ( .IN1(n15258), .IN2(n14993), .QN(n15256) );
  INVX0 U15198 ( .INP(n14992), .ZN(n14993) );
  NAND2X0 U15199 ( .IN1(g550), .IN2(g22578), .QN(n14992) );
  NAND2X0 U15200 ( .IN1(n15259), .IN2(n15260), .QN(g27278) );
  NAND2X0 U15201 ( .IN1(n15261), .IN2(n15164), .QN(n15260) );
  NAND2X0 U15202 ( .IN1(n15262), .IN2(g388), .QN(n15259) );
  NAND2X0 U15203 ( .IN1(n15263), .IN2(n15264), .QN(g27277) );
  NAND2X0 U15204 ( .IN1(n15162), .IN2(g376), .QN(n15264) );
  NAND2X0 U15205 ( .IN1(n15163), .IN2(n15265), .QN(n15263) );
  NAND2X0 U15206 ( .IN1(n15266), .IN2(n15267), .QN(g27276) );
  NAND2X0 U15207 ( .IN1(n15011), .IN2(g2429), .QN(n15267) );
  NAND2X0 U15208 ( .IN1(n15104), .IN2(n15006), .QN(n15266) );
  INVX0 U15209 ( .INP(n15011), .ZN(n15006) );
  NAND2X0 U15210 ( .IN1(n15105), .IN2(g5555), .QN(n15011) );
  NOR2X0 U15211 ( .IN1(n15268), .IN2(n15269), .QN(n15105) );
  NOR2X0 U15212 ( .IN1(n10780), .IN2(n12926), .QN(n15269) );
  NOR2X0 U15213 ( .IN1(n15270), .IN2(n15271), .QN(n15104) );
  NAND2X0 U15214 ( .IN1(n15272), .IN2(n15273), .QN(n15271) );
  NAND2X0 U15215 ( .IN1(n11195), .IN2(n15172), .QN(n15273) );
  NOR2X0 U15216 ( .IN1(n15171), .IN2(n15093), .QN(n15172) );
  INVX0 U15217 ( .INP(n15009), .ZN(n15093) );
  NAND2X0 U15218 ( .IN1(n15094), .IN2(g3229), .QN(n15272) );
  INVX0 U15219 ( .INP(n15274), .ZN(n15270) );
  NOR2X0 U15220 ( .IN1(n15173), .IN2(n15275), .QN(n15274) );
  NOR2X0 U15221 ( .IN1(n15094), .IN2(n15276), .QN(n15275) );
  NAND2X0 U15222 ( .IN1(n15277), .IN2(n15097), .QN(n15276) );
  NAND2X0 U15223 ( .IN1(g3229), .IN2(n15009), .QN(n15277) );
  NAND2X0 U15224 ( .IN1(n15278), .IN2(n15279), .QN(n15009) );
  NAND2X0 U15225 ( .IN1(n9944), .IN2(n11937), .QN(n15279) );
  NOR2X0 U15226 ( .IN1(n15280), .IN2(n15281), .QN(n15278) );
  NOR2X0 U15227 ( .IN1(n4516), .IN2(g2444), .QN(n15281) );
  NOR2X0 U15228 ( .IN1(n4509), .IN2(g2436), .QN(n15280) );
  NAND2X0 U15229 ( .IN1(n15282), .IN2(n15283), .QN(n15094) );
  NAND2X0 U15230 ( .IN1(n9956), .IN2(n11937), .QN(n15283) );
  NOR2X0 U15231 ( .IN1(n15284), .IN2(n15285), .QN(n15282) );
  NOR2X0 U15232 ( .IN1(n4516), .IN2(g2473), .QN(n15285) );
  NOR2X0 U15233 ( .IN1(n4509), .IN2(g2466), .QN(n15284) );
  NOR2X0 U15234 ( .IN1(n15286), .IN2(n11195), .QN(n15173) );
  NAND2X0 U15235 ( .IN1(n15171), .IN2(n15097), .QN(n15286) );
  NAND2X0 U15236 ( .IN1(n15287), .IN2(n15288), .QN(n15097) );
  NAND2X0 U15237 ( .IN1(n9967), .IN2(n11937), .QN(n15288) );
  NOR2X0 U15238 ( .IN1(n15289), .IN2(n15290), .QN(n15287) );
  NOR2X0 U15239 ( .IN1(n4516), .IN2(g2429), .QN(n15290) );
  NOR2X0 U15240 ( .IN1(n4509), .IN2(g2421), .QN(n15289) );
  NAND2X0 U15241 ( .IN1(n15291), .IN2(n15292), .QN(n15171) );
  NAND2X0 U15242 ( .IN1(n9678), .IN2(n11937), .QN(n15292) );
  NOR2X0 U15243 ( .IN1(n15293), .IN2(n15294), .QN(n15291) );
  NOR2X0 U15244 ( .IN1(n4516), .IN2(g2459), .QN(n15294) );
  NOR2X0 U15245 ( .IN1(n4509), .IN2(g2451), .QN(n15293) );
  NAND2X0 U15246 ( .IN1(n15295), .IN2(n15296), .QN(g27275) );
  NAND2X0 U15247 ( .IN1(n15127), .IN2(n15116), .QN(n15296) );
  INVX0 U15248 ( .INP(n15297), .ZN(n15127) );
  NAND2X0 U15249 ( .IN1(n15298), .IN2(n15299), .QN(n15297) );
  NAND2X0 U15250 ( .IN1(n15300), .IN2(n15215), .QN(n15299) );
  INVX0 U15251 ( .INP(n15214), .ZN(n15215) );
  NOR2X0 U15252 ( .IN1(g3229), .IN2(n15118), .QN(n15300) );
  NOR2X0 U15253 ( .IN1(n15301), .IN2(n15302), .QN(n15298) );
  INVX0 U15254 ( .INP(n15303), .ZN(n15301) );
  NAND2X0 U15255 ( .IN1(n15121), .IN2(g1750), .QN(n15295) );
  NAND2X0 U15256 ( .IN1(n15304), .IN2(n15305), .QN(g27274) );
  INVX0 U15257 ( .INP(n15306), .ZN(n15305) );
  NOR2X0 U15258 ( .IN1(n15034), .IN2(n9970), .QN(n15306) );
  NAND2X0 U15259 ( .IN1(n15221), .IN2(n15034), .QN(n15304) );
  INVX0 U15260 ( .INP(n15035), .ZN(n15034) );
  NAND2X0 U15261 ( .IN1(n15222), .IN2(g7014), .QN(n15035) );
  NAND2X0 U15262 ( .IN1(n15307), .IN2(n15308), .QN(g27273) );
  INVX0 U15263 ( .INP(n15309), .ZN(n15308) );
  NOR2X0 U15264 ( .IN1(n15041), .IN2(n9611), .QN(n15309) );
  NAND2X0 U15265 ( .IN1(n15140), .IN2(n15041), .QN(n15307) );
  INVX0 U15266 ( .INP(n15310), .ZN(n15041) );
  NAND2X0 U15267 ( .IN1(g6750), .IN2(g22615), .QN(n15310) );
  INVX0 U15268 ( .INP(n15311), .ZN(n15140) );
  NAND2X0 U15269 ( .IN1(n15312), .IN2(n15313), .QN(n15311) );
  NAND2X0 U15270 ( .IN1(g3229), .IN2(n15135), .QN(n15313) );
  NOR2X0 U15271 ( .IN1(n15314), .IN2(n15315), .QN(n15312) );
  NOR2X0 U15272 ( .IN1(n15226), .IN2(n15316), .QN(n15315) );
  NAND2X0 U15273 ( .IN1(n14494), .IN2(n14487), .QN(n15316) );
  NAND2X0 U15274 ( .IN1(n15317), .IN2(n15318), .QN(n14487) );
  NAND2X0 U15275 ( .IN1(n9611), .IN2(n14180), .QN(n15318) );
  NOR2X0 U15276 ( .IN1(n15319), .IN2(n15320), .QN(n15317) );
  NOR2X0 U15277 ( .IN1(n4316), .IN2(g1263), .QN(n15320) );
  NOR2X0 U15278 ( .IN1(n4300), .IN2(g1261), .QN(n15319) );
  INVX0 U15279 ( .INP(n15135), .ZN(n14494) );
  NAND2X0 U15280 ( .IN1(n15321), .IN2(n15322), .QN(n15135) );
  NAND2X0 U15281 ( .IN1(n9645), .IN2(n14180), .QN(n15322) );
  NOR2X0 U15282 ( .IN1(n15323), .IN2(n15324), .QN(n15321) );
  NOR2X0 U15283 ( .IN1(n4316), .IN2(g1272), .QN(n15324) );
  NOR2X0 U15284 ( .IN1(n4300), .IN2(g1270), .QN(n15323) );
  INVX0 U15285 ( .INP(n15325), .ZN(n15226) );
  NOR2X0 U15286 ( .IN1(g3229), .IN2(n15325), .QN(n15314) );
  NAND2X0 U15287 ( .IN1(n14492), .IN2(n14507), .QN(n15325) );
  NAND2X0 U15288 ( .IN1(n15326), .IN2(n15327), .QN(n14507) );
  NAND2X0 U15289 ( .IN1(n9631), .IN2(n14180), .QN(n15327) );
  NOR2X0 U15290 ( .IN1(n15328), .IN2(n15329), .QN(n15326) );
  NOR2X0 U15291 ( .IN1(n4316), .IN2(g1266), .QN(n15329) );
  NOR2X0 U15292 ( .IN1(n4300), .IN2(g1264), .QN(n15328) );
  INVX0 U15293 ( .INP(n14502), .ZN(n14492) );
  NAND2X0 U15294 ( .IN1(n15330), .IN2(n15331), .QN(n14502) );
  NAND2X0 U15295 ( .IN1(n9438), .IN2(n14180), .QN(n15331) );
  NOR2X0 U15296 ( .IN1(n15332), .IN2(n15333), .QN(n15330) );
  NOR2X0 U15297 ( .IN1(n4316), .IN2(g1269), .QN(n15333) );
  NOR2X0 U15298 ( .IN1(test_so46), .IN2(n4300), .QN(n15332) );
  NAND2X0 U15299 ( .IN1(n15334), .IN2(n15335), .QN(g27272) );
  NAND2X0 U15300 ( .IN1(test_so37), .IN2(n15239), .QN(n15335) );
  NAND2X0 U15301 ( .IN1(n15234), .IN2(n15148), .QN(n15334) );
  INVX0 U15302 ( .INP(n15336), .ZN(n15148) );
  NAND2X0 U15303 ( .IN1(n15337), .IN2(n15338), .QN(n15336) );
  NAND2X0 U15304 ( .IN1(n15339), .IN2(n15237), .QN(n15338) );
  NAND2X0 U15305 ( .IN1(n15340), .IN2(n15341), .QN(n15337) );
  NOR2X0 U15306 ( .IN1(n15339), .IN2(n15342), .QN(n15340) );
  INVX0 U15307 ( .INP(n15238), .ZN(n15339) );
  NAND2X0 U15308 ( .IN1(n15343), .IN2(n15344), .QN(n15238) );
  NAND2X0 U15309 ( .IN1(g3229), .IN2(n15345), .QN(n15344) );
  NAND2X0 U15310 ( .IN1(n15346), .IN2(n11195), .QN(n15343) );
  NAND2X0 U15311 ( .IN1(n15347), .IN2(n15348), .QN(g27271) );
  NAND2X0 U15312 ( .IN1(n15244), .IN2(n15143), .QN(n15348) );
  NAND2X0 U15313 ( .IN1(n15144), .IN2(g1045), .QN(n15347) );
  NAND2X0 U15314 ( .IN1(n15349), .IN2(n15350), .QN(g27270) );
  INVX0 U15315 ( .INP(n15351), .ZN(n15350) );
  NOR2X0 U15316 ( .IN1(n15052), .IN2(n9972), .QN(n15351) );
  NAND2X0 U15317 ( .IN1(n15352), .IN2(n15052), .QN(n15349) );
  NOR2X0 U15318 ( .IN1(n15353), .IN2(n4381), .QN(n15052) );
  NAND2X0 U15319 ( .IN1(n15354), .IN2(n15355), .QN(g27269) );
  NAND2X0 U15320 ( .IN1(n15153), .IN2(g579), .QN(n15355) );
  NAND2X0 U15321 ( .IN1(n15159), .IN2(n15151), .QN(n15354) );
  NOR2X0 U15322 ( .IN1(n15356), .IN2(n15357), .QN(n15159) );
  NOR2X0 U15323 ( .IN1(n15152), .IN2(n14611), .QN(n15357) );
  INVX0 U15324 ( .INP(n15251), .ZN(n15152) );
  NAND2X0 U15325 ( .IN1(n15358), .IN2(n15359), .QN(n15251) );
  NAND2X0 U15326 ( .IN1(g3229), .IN2(n14606), .QN(n15359) );
  NAND2X0 U15327 ( .IN1(n14597), .IN2(n11195), .QN(n15358) );
  INVX0 U15328 ( .INP(n14606), .ZN(n14597) );
  NAND2X0 U15329 ( .IN1(n15360), .IN2(n15361), .QN(g27268) );
  INVX0 U15330 ( .INP(n15362), .ZN(n15361) );
  NOR2X0 U15331 ( .IN1(n15056), .IN2(n9616), .QN(n15362) );
  NAND2X0 U15332 ( .IN1(n15258), .IN2(n15056), .QN(n15360) );
  INVX0 U15333 ( .INP(n15255), .ZN(n15056) );
  NAND2X0 U15334 ( .IN1(g6642), .IN2(g22578), .QN(n15255) );
  NAND2X0 U15335 ( .IN1(n15363), .IN2(n15364), .QN(g27267) );
  NAND2X0 U15336 ( .IN1(n15365), .IN2(n15164), .QN(n15364) );
  NAND2X0 U15337 ( .IN1(n15366), .IN2(n15367), .QN(n15164) );
  NOR2X0 U15338 ( .IN1(n15368), .IN2(n15369), .QN(n15366) );
  INVX0 U15339 ( .INP(n15370), .ZN(n15363) );
  NOR2X0 U15340 ( .IN1(n15365), .IN2(n9965), .QN(n15370) );
  NAND2X0 U15341 ( .IN1(n15371), .IN2(n15372), .QN(g27266) );
  NAND2X0 U15342 ( .IN1(n15262), .IN2(g373), .QN(n15372) );
  NAND2X0 U15343 ( .IN1(n15261), .IN2(n15265), .QN(n15371) );
  NAND2X0 U15344 ( .IN1(n15373), .IN2(n15374), .QN(g27265) );
  NAND2X0 U15345 ( .IN1(n15375), .IN2(n15163), .QN(n15374) );
  NAND2X0 U15346 ( .IN1(n15162), .IN2(g361), .QN(n15373) );
  NAND2X0 U15347 ( .IN1(n15376), .IN2(n15377), .QN(g27264) );
  NAND2X0 U15348 ( .IN1(n15121), .IN2(g1735), .QN(n15377) );
  NAND2X0 U15349 ( .IN1(n15221), .IN2(n15116), .QN(n15376) );
  INVX0 U15350 ( .INP(n15121), .ZN(n15116) );
  NAND2X0 U15351 ( .IN1(n15222), .IN2(g5511), .QN(n15121) );
  NOR2X0 U15352 ( .IN1(n15378), .IN2(n15379), .QN(n15222) );
  NOR2X0 U15353 ( .IN1(n10780), .IN2(n12975), .QN(n15379) );
  INVX0 U15354 ( .INP(n15380), .ZN(n15221) );
  NAND2X0 U15355 ( .IN1(n15381), .IN2(n15382), .QN(n15380) );
  NOR2X0 U15356 ( .IN1(n15383), .IN2(n15384), .QN(n15382) );
  NOR2X0 U15357 ( .IN1(g3229), .IN2(n15303), .QN(n15384) );
  NAND2X0 U15358 ( .IN1(n15118), .IN2(n15119), .QN(n15303) );
  INVX0 U15359 ( .INP(n15385), .ZN(n15118) );
  NOR2X0 U15360 ( .IN1(n15386), .IN2(n11195), .QN(n15383) );
  INVX0 U15361 ( .INP(n15211), .ZN(n15386) );
  NOR2X0 U15362 ( .IN1(n15302), .IN2(n15387), .QN(n15381) );
  NOR2X0 U15363 ( .IN1(n15211), .IN2(n15388), .QN(n15387) );
  NAND2X0 U15364 ( .IN1(n15389), .IN2(n15214), .QN(n15388) );
  NAND2X0 U15365 ( .IN1(g3229), .IN2(n15119), .QN(n15389) );
  NAND2X0 U15366 ( .IN1(n15390), .IN2(n15391), .QN(n15119) );
  NAND2X0 U15367 ( .IN1(n9947), .IN2(n11946), .QN(n15391) );
  NOR2X0 U15368 ( .IN1(n15392), .IN2(n15393), .QN(n15390) );
  NOR2X0 U15369 ( .IN1(n4518), .IN2(g1750), .QN(n15393) );
  NOR2X0 U15370 ( .IN1(n4511), .IN2(g1742), .QN(n15392) );
  NAND2X0 U15371 ( .IN1(n15394), .IN2(n15395), .QN(n15211) );
  NAND2X0 U15372 ( .IN1(n11946), .IN2(n10331), .QN(n15395) );
  NOR2X0 U15373 ( .IN1(n15396), .IN2(n15397), .QN(n15394) );
  NOR2X0 U15374 ( .IN1(n4518), .IN2(g1779), .QN(n15397) );
  NOR2X0 U15375 ( .IN1(n4511), .IN2(g1772), .QN(n15396) );
  NOR2X0 U15376 ( .IN1(n15398), .IN2(n11195), .QN(n15302) );
  NAND2X0 U15377 ( .IN1(n15385), .IN2(n15214), .QN(n15398) );
  NAND2X0 U15378 ( .IN1(n15399), .IN2(n15400), .QN(n15214) );
  NAND2X0 U15379 ( .IN1(n9970), .IN2(n11946), .QN(n15400) );
  NOR2X0 U15380 ( .IN1(n15401), .IN2(n15402), .QN(n15399) );
  NOR2X0 U15381 ( .IN1(n4518), .IN2(g1735), .QN(n15402) );
  NOR2X0 U15382 ( .IN1(n4511), .IN2(g1727), .QN(n15401) );
  NAND2X0 U15383 ( .IN1(n15403), .IN2(n15404), .QN(n15385) );
  NAND2X0 U15384 ( .IN1(n9681), .IN2(n11946), .QN(n15404) );
  NOR2X0 U15385 ( .IN1(n15405), .IN2(n15406), .QN(n15403) );
  NOR2X0 U15386 ( .IN1(n4518), .IN2(g1765), .QN(n15406) );
  NOR2X0 U15387 ( .IN1(n4511), .IN2(g1757), .QN(n15405) );
  NAND2X0 U15388 ( .IN1(n15407), .IN2(n15408), .QN(g27263) );
  NAND2X0 U15389 ( .IN1(n15244), .IN2(n15234), .QN(n15408) );
  INVX0 U15390 ( .INP(n15409), .ZN(n15244) );
  NAND2X0 U15391 ( .IN1(n15410), .IN2(n15411), .QN(n15409) );
  NAND2X0 U15392 ( .IN1(n15412), .IN2(n15346), .QN(n15411) );
  INVX0 U15393 ( .INP(n15345), .ZN(n15346) );
  NOR2X0 U15394 ( .IN1(g3229), .IN2(n15236), .QN(n15412) );
  INVX0 U15395 ( .INP(n15413), .ZN(n15236) );
  NOR2X0 U15396 ( .IN1(n15414), .IN2(n15415), .QN(n15410) );
  NAND2X0 U15397 ( .IN1(n15239), .IN2(g1056), .QN(n15407) );
  NAND2X0 U15398 ( .IN1(n15416), .IN2(n15417), .QN(g27262) );
  NAND2X0 U15399 ( .IN1(n15144), .IN2(g1030), .QN(n15417) );
  INVX0 U15400 ( .INP(n15143), .ZN(n15144) );
  NAND2X0 U15401 ( .IN1(n15352), .IN2(n15143), .QN(n15416) );
  NOR2X0 U15402 ( .IN1(n15353), .IN2(n4364), .QN(n15143) );
  NAND2X0 U15403 ( .IN1(n15418), .IN2(n15419), .QN(g27261) );
  NAND2X0 U15404 ( .IN1(n15153), .IN2(g576), .QN(n15419) );
  NAND2X0 U15405 ( .IN1(n15258), .IN2(n15151), .QN(n15418) );
  INVX0 U15406 ( .INP(n15153), .ZN(n15151) );
  NAND2X0 U15407 ( .IN1(g6485), .IN2(g22578), .QN(n15153) );
  INVX0 U15408 ( .INP(n15420), .ZN(n15258) );
  NAND2X0 U15409 ( .IN1(n15421), .IN2(n15422), .QN(n15420) );
  NAND2X0 U15410 ( .IN1(g3229), .IN2(n15252), .QN(n15422) );
  NOR2X0 U15411 ( .IN1(n15423), .IN2(n15424), .QN(n15421) );
  NOR2X0 U15412 ( .IN1(n15356), .IN2(n15425), .QN(n15424) );
  NAND2X0 U15413 ( .IN1(n14613), .IN2(n14606), .QN(n15425) );
  NAND2X0 U15414 ( .IN1(n15426), .IN2(n15427), .QN(n14606) );
  NAND2X0 U15415 ( .IN1(n9616), .IN2(g6642), .QN(n15427) );
  NOR2X0 U15416 ( .IN1(n15428), .IN2(n15429), .QN(n15426) );
  NOR2X0 U15417 ( .IN1(n4313), .IN2(g575), .QN(n15429) );
  NOR2X0 U15418 ( .IN1(n4298), .IN2(g576), .QN(n15428) );
  INVX0 U15419 ( .INP(n15252), .ZN(n14613) );
  NAND2X0 U15420 ( .IN1(n15430), .IN2(n15431), .QN(n15252) );
  NAND2X0 U15421 ( .IN1(n9650), .IN2(g6642), .QN(n15431) );
  NOR2X0 U15422 ( .IN1(n15432), .IN2(n15433), .QN(n15430) );
  NOR2X0 U15423 ( .IN1(n4313), .IN2(g584), .QN(n15433) );
  NOR2X0 U15424 ( .IN1(n4298), .IN2(g585), .QN(n15432) );
  INVX0 U15425 ( .INP(n15434), .ZN(n15356) );
  NOR2X0 U15426 ( .IN1(g3229), .IN2(n15434), .QN(n15423) );
  NAND2X0 U15427 ( .IN1(n14611), .IN2(n14626), .QN(n15434) );
  NAND2X0 U15428 ( .IN1(n15435), .IN2(n15436), .QN(n14626) );
  NAND2X0 U15429 ( .IN1(g6642), .IN2(n10333), .QN(n15436) );
  NOR2X0 U15430 ( .IN1(n15437), .IN2(n15438), .QN(n15435) );
  NOR2X0 U15431 ( .IN1(n4313), .IN2(g578), .QN(n15438) );
  NOR2X0 U15432 ( .IN1(n4298), .IN2(g579), .QN(n15437) );
  INVX0 U15433 ( .INP(n14621), .ZN(n14611) );
  NAND2X0 U15434 ( .IN1(n15439), .IN2(n15440), .QN(n14621) );
  NAND2X0 U15435 ( .IN1(n9442), .IN2(g6642), .QN(n15440) );
  NOR2X0 U15436 ( .IN1(n15441), .IN2(n15442), .QN(n15439) );
  NOR2X0 U15437 ( .IN1(n4313), .IN2(g581), .QN(n15442) );
  NOR2X0 U15438 ( .IN1(n4298), .IN2(g582), .QN(n15441) );
  NAND2X0 U15439 ( .IN1(n15443), .IN2(n15444), .QN(g27260) );
  INVX0 U15440 ( .INP(n15445), .ZN(n15444) );
  NOR2X0 U15441 ( .IN1(n15365), .IN2(n9684), .QN(n15445) );
  NAND2X0 U15442 ( .IN1(n15365), .IN2(n15265), .QN(n15443) );
  INVX0 U15443 ( .INP(n15446), .ZN(n15265) );
  NAND2X0 U15444 ( .IN1(n15447), .IN2(n15448), .QN(n15446) );
  NAND2X0 U15445 ( .IN1(n15449), .IN2(n15368), .QN(n15448) );
  NAND2X0 U15446 ( .IN1(n15450), .IN2(n15451), .QN(n15447) );
  NOR2X0 U15447 ( .IN1(n15449), .IN2(n15452), .QN(n15450) );
  INVX0 U15448 ( .INP(n15369), .ZN(n15449) );
  NAND2X0 U15449 ( .IN1(n15453), .IN2(n15454), .QN(n15369) );
  NAND2X0 U15450 ( .IN1(g3229), .IN2(n15455), .QN(n15454) );
  NAND2X0 U15451 ( .IN1(n15456), .IN2(n11195), .QN(n15453) );
  NAND2X0 U15452 ( .IN1(n15457), .IN2(n15458), .QN(g27259) );
  NAND2X0 U15453 ( .IN1(n15375), .IN2(n15261), .QN(n15458) );
  NAND2X0 U15454 ( .IN1(n15262), .IN2(g358), .QN(n15457) );
  NAND2X0 U15455 ( .IN1(n15459), .IN2(n15460), .QN(g27258) );
  NAND2X0 U15456 ( .IN1(test_so16), .IN2(n15162), .QN(n15460) );
  NAND2X0 U15457 ( .IN1(n15461), .IN2(n15163), .QN(n15459) );
  INVX0 U15458 ( .INP(n15162), .ZN(n15163) );
  NAND2X0 U15459 ( .IN1(n15462), .IN2(n13361), .QN(n15162) );
  NAND2X0 U15460 ( .IN1(n15463), .IN2(n15464), .QN(g27257) );
  NAND2X0 U15461 ( .IN1(n15239), .IN2(g1041), .QN(n15464) );
  INVX0 U15462 ( .INP(n15234), .ZN(n15239) );
  NAND2X0 U15463 ( .IN1(n15352), .IN2(n15234), .QN(n15463) );
  NOR2X0 U15464 ( .IN1(n15353), .IN2(n4363), .QN(n15234) );
  NAND2X0 U15465 ( .IN1(n10845), .IN2(n15465), .QN(n15353) );
  NAND2X0 U15466 ( .IN1(n15466), .IN2(n10804), .QN(n15465) );
  NOR2X0 U15467 ( .IN1(n15467), .IN2(n15468), .QN(n15352) );
  NAND2X0 U15468 ( .IN1(n15469), .IN2(n15470), .QN(n15468) );
  NAND2X0 U15469 ( .IN1(n11195), .IN2(n15414), .QN(n15470) );
  NOR2X0 U15470 ( .IN1(n15413), .IN2(n15341), .QN(n15414) );
  INVX0 U15471 ( .INP(n15237), .ZN(n15341) );
  NAND2X0 U15472 ( .IN1(n15342), .IN2(g3229), .QN(n15469) );
  INVX0 U15473 ( .INP(n15471), .ZN(n15467) );
  NOR2X0 U15474 ( .IN1(n15415), .IN2(n15472), .QN(n15471) );
  NOR2X0 U15475 ( .IN1(n15342), .IN2(n15473), .QN(n15472) );
  NAND2X0 U15476 ( .IN1(n15474), .IN2(n15345), .QN(n15473) );
  NAND2X0 U15477 ( .IN1(g3229), .IN2(n15237), .QN(n15474) );
  NAND2X0 U15478 ( .IN1(n15475), .IN2(n15476), .QN(n15237) );
  NAND2X0 U15479 ( .IN1(n9949), .IN2(g1088), .QN(n15476) );
  NOR2X0 U15480 ( .IN1(n15477), .IN2(n15478), .QN(n15475) );
  NOR2X0 U15481 ( .IN1(n4364), .IN2(g1045), .QN(n15478) );
  NOR2X0 U15482 ( .IN1(n4363), .IN2(g1056), .QN(n15477) );
  NAND2X0 U15483 ( .IN1(n15479), .IN2(n15480), .QN(n15342) );
  NAND2X0 U15484 ( .IN1(n9960), .IN2(g1088), .QN(n15480) );
  NOR2X0 U15485 ( .IN1(n15481), .IN2(n15482), .QN(n15479) );
  NOR2X0 U15486 ( .IN1(n4364), .IN2(g1075), .QN(n15482) );
  NOR2X0 U15487 ( .IN1(n4363), .IN2(g1085), .QN(n15481) );
  NOR2X0 U15488 ( .IN1(n15483), .IN2(n11195), .QN(n15415) );
  NAND2X0 U15489 ( .IN1(n15413), .IN2(n15345), .QN(n15483) );
  NAND2X0 U15490 ( .IN1(n15484), .IN2(n15485), .QN(n15345) );
  NAND2X0 U15491 ( .IN1(n9972), .IN2(g1088), .QN(n15485) );
  NOR2X0 U15492 ( .IN1(n15486), .IN2(n15487), .QN(n15484) );
  NOR2X0 U15493 ( .IN1(n4364), .IN2(g1030), .QN(n15487) );
  NOR2X0 U15494 ( .IN1(n4363), .IN2(g1041), .QN(n15486) );
  NAND2X0 U15495 ( .IN1(n15488), .IN2(n15489), .QN(n15413) );
  NAND2X0 U15496 ( .IN1(n9683), .IN2(g1088), .QN(n15489) );
  NOR2X0 U15497 ( .IN1(n15490), .IN2(n15491), .QN(n15488) );
  NOR2X0 U15498 ( .IN1(n4364), .IN2(g1060), .QN(n15491) );
  NOR2X0 U15499 ( .IN1(test_so37), .IN2(n4363), .QN(n15490) );
  NAND2X0 U15500 ( .IN1(n15492), .IN2(n15493), .QN(g27256) );
  NAND2X0 U15501 ( .IN1(n15375), .IN2(n15365), .QN(n15493) );
  INVX0 U15502 ( .INP(n15494), .ZN(n15375) );
  NAND2X0 U15503 ( .IN1(n15495), .IN2(n15496), .QN(n15494) );
  NAND2X0 U15504 ( .IN1(n15497), .IN2(n15456), .QN(n15496) );
  INVX0 U15505 ( .INP(n15455), .ZN(n15456) );
  NOR2X0 U15506 ( .IN1(g3229), .IN2(n15367), .QN(n15497) );
  INVX0 U15507 ( .INP(n15498), .ZN(n15367) );
  NOR2X0 U15508 ( .IN1(n15499), .IN2(n15500), .QN(n15495) );
  INVX0 U15509 ( .INP(n15501), .ZN(n15492) );
  NOR2X0 U15510 ( .IN1(n15365), .IN2(n9954), .QN(n15501) );
  NAND2X0 U15511 ( .IN1(n15502), .IN2(n15503), .QN(g27255) );
  NAND2X0 U15512 ( .IN1(n15262), .IN2(g343), .QN(n15503) );
  NAND2X0 U15513 ( .IN1(n15461), .IN2(n15261), .QN(n15502) );
  INVX0 U15514 ( .INP(n15262), .ZN(n15261) );
  NAND2X0 U15515 ( .IN1(n15462), .IN2(g6447), .QN(n15262) );
  NAND2X0 U15516 ( .IN1(n15504), .IN2(n15505), .QN(g27253) );
  INVX0 U15517 ( .INP(n15506), .ZN(n15505) );
  NOR2X0 U15518 ( .IN1(n15365), .IN2(n9976), .QN(n15506) );
  NAND2X0 U15519 ( .IN1(n15461), .IN2(n15365), .QN(n15504) );
  INVX0 U15520 ( .INP(n15507), .ZN(n15365) );
  NAND2X0 U15521 ( .IN1(n15462), .IN2(g5437), .QN(n15507) );
  NOR2X0 U15522 ( .IN1(n15508), .IN2(n15509), .QN(n15462) );
  NOR2X0 U15523 ( .IN1(n10780), .IN2(n13109), .QN(n15509) );
  NOR2X0 U15524 ( .IN1(n15510), .IN2(n15511), .QN(n15461) );
  NAND2X0 U15525 ( .IN1(n15512), .IN2(n15513), .QN(n15511) );
  NAND2X0 U15526 ( .IN1(n11195), .IN2(n15499), .QN(n15513) );
  NOR2X0 U15527 ( .IN1(n15498), .IN2(n15451), .QN(n15499) );
  INVX0 U15528 ( .INP(n15368), .ZN(n15451) );
  NAND2X0 U15529 ( .IN1(n15452), .IN2(g3229), .QN(n15512) );
  INVX0 U15530 ( .INP(n15514), .ZN(n15510) );
  NOR2X0 U15531 ( .IN1(n15500), .IN2(n15515), .QN(n15514) );
  NOR2X0 U15532 ( .IN1(n15452), .IN2(n15516), .QN(n15515) );
  NAND2X0 U15533 ( .IN1(n15517), .IN2(n15455), .QN(n15516) );
  NAND2X0 U15534 ( .IN1(g3229), .IN2(n15368), .QN(n15517) );
  NAND2X0 U15535 ( .IN1(n15518), .IN2(n15519), .QN(n15368) );
  NAND2X0 U15536 ( .IN1(n9954), .IN2(n12042), .QN(n15519) );
  NOR2X0 U15537 ( .IN1(n15520), .IN2(n15521), .QN(n15518) );
  NOR2X0 U15538 ( .IN1(n4506), .IN2(g361), .QN(n15521) );
  NOR2X0 U15539 ( .IN1(n4499), .IN2(g358), .QN(n15520) );
  NAND2X0 U15540 ( .IN1(n15522), .IN2(n15523), .QN(n15452) );
  NAND2X0 U15541 ( .IN1(n9965), .IN2(n12042), .QN(n15523) );
  NOR2X0 U15542 ( .IN1(n15524), .IN2(n15525), .QN(n15522) );
  NOR2X0 U15543 ( .IN1(n4506), .IN2(g391), .QN(n15525) );
  NOR2X0 U15544 ( .IN1(n4499), .IN2(g388), .QN(n15524) );
  NOR2X0 U15545 ( .IN1(n15526), .IN2(n11195), .QN(n15500) );
  NAND2X0 U15546 ( .IN1(n15498), .IN2(n15455), .QN(n15526) );
  NAND2X0 U15547 ( .IN1(n15527), .IN2(n15528), .QN(n15455) );
  NAND2X0 U15548 ( .IN1(n9976), .IN2(n12042), .QN(n15528) );
  NOR2X0 U15549 ( .IN1(n15529), .IN2(n15530), .QN(n15527) );
  NOR2X0 U15550 ( .IN1(test_so16), .IN2(n4506), .QN(n15530) );
  NOR2X0 U15551 ( .IN1(n4499), .IN2(g343), .QN(n15529) );
  NAND2X0 U15552 ( .IN1(n15531), .IN2(n15532), .QN(n15498) );
  NAND2X0 U15553 ( .IN1(n9684), .IN2(n12042), .QN(n15532) );
  NOR2X0 U15554 ( .IN1(n15533), .IN2(n15534), .QN(n15531) );
  NOR2X0 U15555 ( .IN1(n4506), .IN2(g376), .QN(n15534) );
  NOR2X0 U15556 ( .IN1(n4499), .IN2(g373), .QN(n15533) );
  NOR2X0 U15557 ( .IN1(n15535), .IN2(n15536), .QN(g27243) );
  NAND2X0 U15558 ( .IN1(n14827), .IN2(n14826), .QN(n15536) );
  NAND2X0 U15559 ( .IN1(n15537), .IN2(test_so92), .QN(n14827) );
  NOR2X0 U15560 ( .IN1(n4471), .IN2(n15538), .QN(n15537) );
  NOR2X0 U15561 ( .IN1(n15539), .IN2(g2753), .QN(n15535) );
  NOR2X0 U15562 ( .IN1(n15538), .IN2(n10324), .QN(n15539) );
  NOR2X0 U15563 ( .IN1(n14857), .IN2(n15540), .QN(g27131) );
  NAND2X0 U15564 ( .IN1(n15541), .IN2(n13952), .QN(n15540) );
  INVX0 U15565 ( .INP(n15542), .ZN(n15541) );
  NOR2X0 U15566 ( .IN1(g2147), .IN2(n3683), .QN(n15542) );
  INVX0 U15567 ( .INP(n4522), .ZN(n14857) );
  NOR2X0 U15568 ( .IN1(n14861), .IN2(n15543), .QN(g27129) );
  NAND2X0 U15569 ( .IN1(n15544), .IN2(n13954), .QN(n15543) );
  INVX0 U15570 ( .INP(n15545), .ZN(n15544) );
  NOR2X0 U15571 ( .IN1(g1453), .IN2(n3686), .QN(n15545) );
  INVX0 U15572 ( .INP(n4523), .ZN(n14861) );
  NOR2X0 U15573 ( .IN1(n15546), .IN2(n14865), .QN(g27123) );
  NAND2X0 U15574 ( .IN1(n3431), .IN2(n13956), .QN(n14865) );
  NAND2X0 U15575 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NOR2X0 U15576 ( .IN1(n3689), .IN2(g767), .QN(n15546) );
  NOR2X0 U15577 ( .IN1(n14870), .IN2(n15547), .QN(g27120) );
  NAND2X0 U15578 ( .IN1(n15548), .IN2(n13958), .QN(n15547) );
  INVX0 U15579 ( .INP(n15549), .ZN(n15548) );
  NOR2X0 U15580 ( .IN1(test_so15), .IN2(n3692), .QN(n15549) );
  INVX0 U15581 ( .INP(n4521), .ZN(n14870) );
  NAND2X0 U15582 ( .IN1(n15550), .IN2(n15551), .QN(g26827) );
  NAND2X0 U15583 ( .IN1(n15552), .IN2(n4606), .QN(n15551) );
  INVX0 U15584 ( .INP(n15553), .ZN(n15550) );
  NOR2X0 U15585 ( .IN1(n13307), .IN2(n9752), .QN(n15553) );
  NAND2X0 U15586 ( .IN1(n15554), .IN2(n15555), .QN(g26826) );
  NAND2X0 U15587 ( .IN1(n15552), .IN2(g7264), .QN(n15555) );
  INVX0 U15588 ( .INP(n15556), .ZN(n15554) );
  NOR2X0 U15589 ( .IN1(n11937), .IN2(n9741), .QN(n15556) );
  NAND2X0 U15590 ( .IN1(n15557), .IN2(n15558), .QN(g26825) );
  NAND2X0 U15591 ( .IN1(n4606), .IN2(n15559), .QN(n15558) );
  INVX0 U15592 ( .INP(n15560), .ZN(n15557) );
  NOR2X0 U15593 ( .IN1(n13307), .IN2(n9754), .QN(n15560) );
  NAND2X0 U15594 ( .IN1(n15561), .IN2(n15562), .QN(g26824) );
  NAND2X0 U15595 ( .IN1(n15563), .IN2(n4618), .QN(n15562) );
  NAND2X0 U15596 ( .IN1(test_so59), .IN2(n4511), .QN(n15561) );
  NAND2X0 U15597 ( .IN1(n15564), .IN2(n15565), .QN(g26823) );
  NAND2X0 U15598 ( .IN1(n15552), .IN2(g5555), .QN(n15565) );
  NOR2X0 U15599 ( .IN1(n15566), .IN2(n15567), .QN(n15552) );
  INVX0 U15600 ( .INP(n15568), .ZN(n15567) );
  NAND2X0 U15601 ( .IN1(n15569), .IN2(n15570), .QN(n15568) );
  NOR2X0 U15602 ( .IN1(n15570), .IN2(n15569), .QN(n15566) );
  NAND2X0 U15603 ( .IN1(n15571), .IN2(test_so79), .QN(n15570) );
  NOR2X0 U15604 ( .IN1(n15572), .IN2(n14739), .QN(n15571) );
  INVX0 U15605 ( .INP(n15573), .ZN(n14739) );
  NAND2X0 U15606 ( .IN1(n15574), .IN2(n15575), .QN(n15573) );
  NAND2X0 U15607 ( .IN1(n14750), .IN2(n14749), .QN(n15575) );
  NOR2X0 U15608 ( .IN1(n15569), .IN2(n15576), .QN(n14750) );
  INVX0 U15609 ( .INP(n14747), .ZN(n15569) );
  NAND2X0 U15610 ( .IN1(n15577), .IN2(n14746), .QN(n15574) );
  NOR2X0 U15611 ( .IN1(n14748), .IN2(n14747), .QN(n15577) );
  INVX0 U15612 ( .INP(n15576), .ZN(n14748) );
  NOR2X0 U15613 ( .IN1(n14738), .IN2(n14740), .QN(n15572) );
  NAND2X0 U15614 ( .IN1(n15578), .IN2(n15579), .QN(n14740) );
  NAND2X0 U15615 ( .IN1(n9987), .IN2(n13416), .QN(n15579) );
  NAND2X0 U15616 ( .IN1(n9978), .IN2(n11937), .QN(n15578) );
  NOR2X0 U15617 ( .IN1(n4509), .IN2(test_so81), .QN(n14738) );
  NAND2X0 U15618 ( .IN1(n4516), .IN2(g2513), .QN(n15564) );
  NAND2X0 U15619 ( .IN1(n15580), .IN2(n15581), .QN(g26822) );
  NAND2X0 U15620 ( .IN1(g7264), .IN2(n15559), .QN(n15581) );
  INVX0 U15621 ( .INP(n15582), .ZN(n15580) );
  NOR2X0 U15622 ( .IN1(n11937), .IN2(n9742), .QN(n15582) );
  NAND2X0 U15623 ( .IN1(n15583), .IN2(n15584), .QN(g26821) );
  NAND2X0 U15624 ( .IN1(n15563), .IN2(g7014), .QN(n15584) );
  INVX0 U15625 ( .INP(n15585), .ZN(n15583) );
  NOR2X0 U15626 ( .IN1(n11946), .IN2(n9745), .QN(n15585) );
  NAND2X0 U15627 ( .IN1(n15586), .IN2(n15587), .QN(g26820) );
  NAND2X0 U15628 ( .IN1(n4618), .IN2(n15588), .QN(n15587) );
  INVX0 U15629 ( .INP(n15589), .ZN(n15586) );
  NOR2X0 U15630 ( .IN1(n13315), .IN2(n9760), .QN(n15589) );
  NAND2X0 U15631 ( .IN1(n15590), .IN2(n15591), .QN(g26818) );
  NAND2X0 U15632 ( .IN1(n4381), .IN2(g1131), .QN(n15591) );
  NAND2X0 U15633 ( .IN1(n15592), .IN2(g1088), .QN(n15590) );
  NAND2X0 U15634 ( .IN1(n15593), .IN2(n15594), .QN(g26817) );
  NAND2X0 U15635 ( .IN1(g5555), .IN2(n15559), .QN(n15594) );
  NAND2X0 U15636 ( .IN1(n15595), .IN2(n15596), .QN(n15559) );
  NAND2X0 U15637 ( .IN1(n14746), .IN2(test_so79), .QN(n15596) );
  INVX0 U15638 ( .INP(n14749), .ZN(n14746) );
  NAND2X0 U15639 ( .IN1(n14016), .IN2(n15597), .QN(n14749) );
  NAND2X0 U15640 ( .IN1(n15598), .IN2(n15599), .QN(n15597) );
  NAND2X0 U15641 ( .IN1(n9891), .IN2(test_so73), .QN(n15599) );
  NOR2X0 U15642 ( .IN1(n15600), .IN2(n15601), .QN(n15598) );
  NOR2X0 U15643 ( .IN1(n4367), .IN2(g2253), .QN(n15601) );
  NOR2X0 U15644 ( .IN1(n4324), .IN2(g2254), .QN(n15600) );
  INVX0 U15645 ( .INP(n15602), .ZN(n14016) );
  NAND2X0 U15646 ( .IN1(n15576), .IN2(n10322), .QN(n15595) );
  NAND2X0 U15647 ( .IN1(n15603), .IN2(n15604), .QN(n15576) );
  NAND2X0 U15648 ( .IN1(g5555), .IN2(g2504), .QN(n15604) );
  NOR2X0 U15649 ( .IN1(n15605), .IN2(n15606), .QN(n15603) );
  NOR2X0 U15650 ( .IN1(n9742), .IN2(n14010), .QN(n15606) );
  NOR2X0 U15651 ( .IN1(n9754), .IN2(n15607), .QN(n15605) );
  NAND2X0 U15652 ( .IN1(n4516), .IN2(g2504), .QN(n15593) );
  NAND2X0 U15653 ( .IN1(n15608), .IN2(n15609), .QN(g26816) );
  NAND2X0 U15654 ( .IN1(n15563), .IN2(g5511), .QN(n15609) );
  NOR2X0 U15655 ( .IN1(n15610), .IN2(n15611), .QN(n15563) );
  NOR2X0 U15656 ( .IN1(n14773), .IN2(n15612), .QN(n15611) );
  INVX0 U15657 ( .INP(n15613), .ZN(n15610) );
  NAND2X0 U15658 ( .IN1(n15612), .IN2(n14773), .QN(n15613) );
  NOR2X0 U15659 ( .IN1(n14763), .IN2(n15614), .QN(n15612) );
  NOR2X0 U15660 ( .IN1(n14766), .IN2(n15615), .QN(n15614) );
  NOR2X0 U15661 ( .IN1(g1830), .IN2(n4525), .QN(n15615) );
  NAND2X0 U15662 ( .IN1(n15616), .IN2(n15617), .QN(n14766) );
  NAND2X0 U15663 ( .IN1(n9991), .IN2(n13315), .QN(n15617) );
  NAND2X0 U15664 ( .IN1(n9992), .IN2(n13555), .QN(n15616) );
  NAND2X0 U15665 ( .IN1(n15618), .IN2(g1690), .QN(n14763) );
  NOR2X0 U15666 ( .IN1(n15619), .IN2(n15620), .QN(n15618) );
  NOR2X0 U15667 ( .IN1(n14770), .IN2(n14773), .QN(n15620) );
  NOR2X0 U15668 ( .IN1(n15621), .IN2(n15622), .QN(n14770) );
  INVX0 U15669 ( .INP(n14776), .ZN(n15621) );
  NOR2X0 U15670 ( .IN1(n14775), .IN2(n15623), .QN(n15619) );
  NOR2X0 U15671 ( .IN1(n14772), .IN2(n14776), .QN(n15623) );
  INVX0 U15672 ( .INP(n14773), .ZN(n14775) );
  NAND2X0 U15673 ( .IN1(n4518), .IN2(g1819), .QN(n15608) );
  NAND2X0 U15674 ( .IN1(n15624), .IN2(n15625), .QN(g26815) );
  NAND2X0 U15675 ( .IN1(g7014), .IN2(n15588), .QN(n15625) );
  INVX0 U15676 ( .INP(n15626), .ZN(n15624) );
  NOR2X0 U15677 ( .IN1(n11946), .IN2(n9746), .QN(n15626) );
  NAND2X0 U15678 ( .IN1(n15627), .IN2(n15628), .QN(g26814) );
  INVX0 U15679 ( .INP(n15629), .ZN(n15628) );
  NOR2X0 U15680 ( .IN1(g6712), .IN2(n9749), .QN(n15629) );
  NAND2X0 U15681 ( .IN1(n15592), .IN2(g6712), .QN(n15627) );
  NAND2X0 U15682 ( .IN1(n15630), .IN2(n15631), .QN(g26813) );
  NAND2X0 U15683 ( .IN1(n4381), .IN2(g1122), .QN(n15631) );
  NAND2X0 U15684 ( .IN1(n15632), .IN2(g1088), .QN(n15630) );
  NAND2X0 U15685 ( .IN1(n15633), .IN2(n15634), .QN(g26812) );
  NAND2X0 U15686 ( .IN1(n15635), .IN2(n4640), .QN(n15634) );
  INVX0 U15687 ( .INP(n15636), .ZN(n15633) );
  NOR2X0 U15688 ( .IN1(n13361), .IN2(n9774), .QN(n15636) );
  NAND2X0 U15689 ( .IN1(n15637), .IN2(n15638), .QN(g26811) );
  NAND2X0 U15690 ( .IN1(g5511), .IN2(n15588), .QN(n15638) );
  NAND2X0 U15691 ( .IN1(n15639), .IN2(n15640), .QN(n15588) );
  NAND2X0 U15692 ( .IN1(n14772), .IN2(g1690), .QN(n15640) );
  INVX0 U15693 ( .INP(n15622), .ZN(n14772) );
  NAND2X0 U15694 ( .IN1(n14060), .IN2(n15641), .QN(n15622) );
  NAND2X0 U15695 ( .IN1(n15642), .IN2(n15643), .QN(n15641) );
  NAND2X0 U15696 ( .IN1(n9903), .IN2(g6782), .QN(n15643) );
  NOR2X0 U15697 ( .IN1(n15644), .IN2(n15645), .QN(n15642) );
  NOR2X0 U15698 ( .IN1(n4368), .IN2(g1559), .QN(n15645) );
  NOR2X0 U15699 ( .IN1(n4317), .IN2(g1560), .QN(n15644) );
  INVX0 U15700 ( .INP(n15646), .ZN(n14060) );
  NAND2X0 U15701 ( .IN1(n4386), .IN2(n14776), .QN(n15639) );
  NAND2X0 U15702 ( .IN1(n15647), .IN2(n15648), .QN(n14776) );
  NAND2X0 U15703 ( .IN1(g5511), .IN2(g1810), .QN(n15648) );
  NOR2X0 U15704 ( .IN1(n15649), .IN2(n15650), .QN(n15647) );
  NOR2X0 U15705 ( .IN1(n9746), .IN2(n13179), .QN(n15650) );
  NOR2X0 U15706 ( .IN1(n9760), .IN2(n14055), .QN(n15649) );
  NAND2X0 U15707 ( .IN1(n4518), .IN2(g1810), .QN(n15637) );
  NAND2X0 U15708 ( .IN1(n15651), .IN2(n15652), .QN(g26810) );
  INVX0 U15709 ( .INP(n15653), .ZN(n15652) );
  NOR2X0 U15710 ( .IN1(g5472), .IN2(n9767), .QN(n15653) );
  NAND2X0 U15711 ( .IN1(n15592), .IN2(g5472), .QN(n15651) );
  NOR2X0 U15712 ( .IN1(n15654), .IN2(n15655), .QN(n15592) );
  NOR2X0 U15713 ( .IN1(n14799), .IN2(n15656), .QN(n15655) );
  INVX0 U15714 ( .INP(n15657), .ZN(n15654) );
  NAND2X0 U15715 ( .IN1(n15656), .IN2(n14799), .QN(n15657) );
  NOR2X0 U15716 ( .IN1(n14789), .IN2(n15658), .QN(n15656) );
  NOR2X0 U15717 ( .IN1(n14792), .IN2(n15659), .QN(n15658) );
  NOR2X0 U15718 ( .IN1(g1136), .IN2(n4364), .QN(n15659) );
  NAND2X0 U15719 ( .IN1(n15660), .IN2(n15661), .QN(n14792) );
  NAND2X0 U15720 ( .IN1(n9998), .IN2(g5472), .QN(n15661) );
  NAND2X0 U15721 ( .IN1(n9997), .IN2(g1088), .QN(n15660) );
  NAND2X0 U15722 ( .IN1(n15662), .IN2(g996), .QN(n14789) );
  NOR2X0 U15723 ( .IN1(n15663), .IN2(n15664), .QN(n15662) );
  NOR2X0 U15724 ( .IN1(n14796), .IN2(n14799), .QN(n15664) );
  NOR2X0 U15725 ( .IN1(n15665), .IN2(n15666), .QN(n14796) );
  INVX0 U15726 ( .INP(n14802), .ZN(n15665) );
  NOR2X0 U15727 ( .IN1(n14801), .IN2(n15667), .QN(n15663) );
  NOR2X0 U15728 ( .IN1(n14798), .IN2(n14802), .QN(n15667) );
  INVX0 U15729 ( .INP(n14799), .ZN(n14801) );
  NAND2X0 U15730 ( .IN1(n15668), .IN2(n15669), .QN(g26809) );
  NAND2X0 U15731 ( .IN1(n15632), .IN2(g6712), .QN(n15669) );
  NAND2X0 U15732 ( .IN1(n4364), .IN2(test_so38), .QN(n15668) );
  NAND2X0 U15733 ( .IN1(n15670), .IN2(n15671), .QN(g26808) );
  NAND2X0 U15734 ( .IN1(n15635), .IN2(g6447), .QN(n15671) );
  INVX0 U15735 ( .INP(n15672), .ZN(n15670) );
  NOR2X0 U15736 ( .IN1(n13382), .IN2(n9775), .QN(n15672) );
  NAND2X0 U15737 ( .IN1(n15673), .IN2(n15674), .QN(g26807) );
  NAND2X0 U15738 ( .IN1(n4640), .IN2(n15675), .QN(n15674) );
  INVX0 U15739 ( .INP(n15676), .ZN(n15673) );
  NOR2X0 U15740 ( .IN1(n13361), .IN2(n9777), .QN(n15676) );
  NAND2X0 U15741 ( .IN1(n15677), .IN2(n15678), .QN(g26806) );
  INVX0 U15742 ( .INP(n15679), .ZN(n15678) );
  NOR2X0 U15743 ( .IN1(g5472), .IN2(n9769), .QN(n15679) );
  NAND2X0 U15744 ( .IN1(n15632), .IN2(g5472), .QN(n15677) );
  NAND2X0 U15745 ( .IN1(n15680), .IN2(n15681), .QN(n15632) );
  NAND2X0 U15746 ( .IN1(n14798), .IN2(g996), .QN(n15681) );
  INVX0 U15747 ( .INP(n15666), .ZN(n14798) );
  NAND2X0 U15748 ( .IN1(n14100), .IN2(n15682), .QN(n15666) );
  NAND2X0 U15749 ( .IN1(n15683), .IN2(n15684), .QN(n15682) );
  NAND2X0 U15750 ( .IN1(n9913), .IN2(test_so31), .QN(n15684) );
  NOR2X0 U15751 ( .IN1(n15685), .IN2(n15686), .QN(n15683) );
  NOR2X0 U15752 ( .IN1(n4323), .IN2(g866), .QN(n15686) );
  NOR2X0 U15753 ( .IN1(n4312), .IN2(g867), .QN(n15685) );
  INVX0 U15754 ( .INP(n15687), .ZN(n14100) );
  NAND2X0 U15755 ( .IN1(n4387), .IN2(n14802), .QN(n15680) );
  NAND2X0 U15756 ( .IN1(n15688), .IN2(n15689), .QN(n14802) );
  NAND2X0 U15757 ( .IN1(g1088), .IN2(g1122), .QN(n15689) );
  NOR2X0 U15758 ( .IN1(n15690), .IN2(n15691), .QN(n15688) );
  INVX0 U15759 ( .INP(n15692), .ZN(n15691) );
  NAND2X0 U15760 ( .IN1(g6712), .IN2(test_so38), .QN(n15692) );
  NOR2X0 U15761 ( .IN1(n9769), .IN2(n4363), .QN(n15690) );
  NAND2X0 U15762 ( .IN1(n15693), .IN2(n15694), .QN(g26805) );
  NAND2X0 U15763 ( .IN1(n15635), .IN2(g5437), .QN(n15694) );
  NOR2X0 U15764 ( .IN1(n15695), .IN2(n15696), .QN(n15635) );
  NOR2X0 U15765 ( .IN1(n14820), .IN2(n15697), .QN(n15696) );
  INVX0 U15766 ( .INP(n15698), .ZN(n15695) );
  NAND2X0 U15767 ( .IN1(n15697), .IN2(n14820), .QN(n15698) );
  NOR2X0 U15768 ( .IN1(n14810), .IN2(n15699), .QN(n15697) );
  NOR2X0 U15769 ( .IN1(n14813), .IN2(n15700), .QN(n15699) );
  NOR2X0 U15770 ( .IN1(g447), .IN2(n4506), .QN(n15700) );
  NAND2X0 U15771 ( .IN1(n15701), .IN2(n15702), .QN(n14813) );
  NAND2X0 U15772 ( .IN1(n10005), .IN2(n13382), .QN(n15702) );
  NAND2X0 U15773 ( .IN1(n10006), .IN2(n12042), .QN(n15701) );
  NAND2X0 U15774 ( .IN1(n15703), .IN2(g309), .QN(n14810) );
  NOR2X0 U15775 ( .IN1(n15704), .IN2(n15705), .QN(n15703) );
  NOR2X0 U15776 ( .IN1(n14817), .IN2(n14820), .QN(n15705) );
  NOR2X0 U15777 ( .IN1(n15706), .IN2(n15707), .QN(n14817) );
  INVX0 U15778 ( .INP(n14823), .ZN(n15706) );
  NOR2X0 U15779 ( .IN1(n14822), .IN2(n15708), .QN(n15704) );
  NOR2X0 U15780 ( .IN1(n14819), .IN2(n14823), .QN(n15708) );
  INVX0 U15781 ( .INP(n14820), .ZN(n14822) );
  NAND2X0 U15782 ( .IN1(n4520), .IN2(g438), .QN(n15693) );
  NAND2X0 U15783 ( .IN1(n15709), .IN2(n15710), .QN(g26804) );
  NAND2X0 U15784 ( .IN1(g6447), .IN2(n15675), .QN(n15710) );
  INVX0 U15785 ( .INP(n15711), .ZN(n15709) );
  NOR2X0 U15786 ( .IN1(n13382), .IN2(n9778), .QN(n15711) );
  NAND2X0 U15787 ( .IN1(n15712), .IN2(n15713), .QN(g26803) );
  NAND2X0 U15788 ( .IN1(g5437), .IN2(n15675), .QN(n15713) );
  NAND2X0 U15789 ( .IN1(n15714), .IN2(n15715), .QN(n15675) );
  NAND2X0 U15790 ( .IN1(n14819), .IN2(g309), .QN(n15715) );
  INVX0 U15791 ( .INP(n15707), .ZN(n14819) );
  NAND2X0 U15792 ( .IN1(n14136), .IN2(n15716), .QN(n15707) );
  NAND2X0 U15793 ( .IN1(n15717), .IN2(n15718), .QN(n15716) );
  NAND2X0 U15794 ( .IN1(n9925), .IN2(g6313), .QN(n15718) );
  NOR2X0 U15795 ( .IN1(n15719), .IN2(n15720), .QN(n15717) );
  NOR2X0 U15796 ( .IN1(n4369), .IN2(g177), .QN(n15720) );
  NOR2X0 U15797 ( .IN1(n4318), .IN2(g178), .QN(n15719) );
  INVX0 U15798 ( .INP(n15721), .ZN(n14136) );
  NAND2X0 U15799 ( .IN1(n4388), .IN2(n14823), .QN(n15714) );
  NAND2X0 U15800 ( .IN1(n15722), .IN2(n15723), .QN(n14823) );
  NAND2X0 U15801 ( .IN1(g5437), .IN2(g429), .QN(n15723) );
  NOR2X0 U15802 ( .IN1(n15724), .IN2(n15725), .QN(n15722) );
  NOR2X0 U15803 ( .IN1(n9778), .IN2(n14129), .QN(n15725) );
  NOR2X0 U15804 ( .IN1(n9777), .IN2(n14130), .QN(n15724) );
  NAND2X0 U15805 ( .IN1(n4520), .IN2(g429), .QN(n15712) );
  NOR2X0 U15806 ( .IN1(n10998), .IN2(n15726), .QN(g26798) );
  NAND2X0 U15807 ( .IN1(n15727), .IN2(n15728), .QN(n15726) );
  NAND2X0 U15808 ( .IN1(n4355), .IN2(n15729), .QN(n15728) );
  NAND2X0 U15809 ( .IN1(n15730), .IN2(g2908), .QN(n15727) );
  NOR2X0 U15810 ( .IN1(n14690), .IN2(n15731), .QN(g26795) );
  NOR2X0 U15811 ( .IN1(n15732), .IN2(n15733), .QN(n15731) );
  NOR2X0 U15812 ( .IN1(test_so92), .IN2(n15538), .QN(n15733) );
  INVX0 U15813 ( .INP(n15734), .ZN(n15732) );
  NAND2X0 U15814 ( .IN1(n15538), .IN2(test_so92), .QN(n15734) );
  NOR2X0 U15815 ( .IN1(n15735), .IN2(n15736), .QN(g26789) );
  NAND2X0 U15816 ( .IN1(n15737), .IN2(n15738), .QN(n15736) );
  NAND2X0 U15817 ( .IN1(n4468), .IN2(n14842), .QN(n15738) );
  NAND2X0 U15818 ( .IN1(n14840), .IN2(g2046), .QN(n15737) );
  INVX0 U15819 ( .INP(n14842), .ZN(n14840) );
  NOR2X0 U15820 ( .IN1(n15739), .IN2(n15740), .QN(g26786) );
  NOR2X0 U15821 ( .IN1(n15741), .IN2(n15742), .QN(n15739) );
  INVX0 U15822 ( .INP(n15743), .ZN(n15742) );
  NAND2X0 U15823 ( .IN1(g3024), .IN2(n3741), .QN(n15743) );
  NOR2X0 U15824 ( .IN1(n3741), .IN2(g3024), .QN(n15741) );
  NOR2X0 U15825 ( .IN1(n14704), .IN2(n15744), .QN(g26781) );
  NAND2X0 U15826 ( .IN1(n15745), .IN2(n15746), .QN(n15744) );
  NAND2X0 U15827 ( .IN1(n4469), .IN2(n14848), .QN(n15746) );
  NAND2X0 U15828 ( .IN1(n14846), .IN2(g1352), .QN(n15745) );
  INVX0 U15829 ( .INP(n14848), .ZN(n14846) );
  NOR2X0 U15830 ( .IN1(n14141), .IN2(n15747), .QN(g26776) );
  NOR2X0 U15831 ( .IN1(n15748), .IN2(n15749), .QN(n15747) );
  NOR2X0 U15832 ( .IN1(test_so28), .IN2(n14852), .QN(n15749) );
  INVX0 U15833 ( .INP(n15750), .ZN(n15748) );
  NAND2X0 U15834 ( .IN1(n14852), .IN2(test_so28), .QN(n15750) );
  NOR2X0 U15835 ( .IN1(n15751), .IN2(n15752), .QN(g26677) );
  NAND2X0 U15836 ( .IN1(n15538), .IN2(n14826), .QN(n15752) );
  NAND2X0 U15837 ( .IN1(n15753), .IN2(n15754), .QN(n15538) );
  NOR2X0 U15838 ( .IN1(n4407), .IN2(n4397), .QN(n15753) );
  NOR2X0 U15839 ( .IN1(n15755), .IN2(g2746), .QN(n15751) );
  NOR2X0 U15840 ( .IN1(n4397), .IN2(n15756), .QN(n15755) );
  NAND2X0 U15841 ( .IN1(n15757), .IN2(n15758), .QN(g26676) );
  NAND2X0 U15842 ( .IN1(n15759), .IN2(g2479), .QN(n15758) );
  NAND2X0 U15843 ( .IN1(n15760), .IN2(n11937), .QN(n15759) );
  NAND2X0 U15844 ( .IN1(n15761), .IN2(n11937), .QN(n15757) );
  NAND2X0 U15845 ( .IN1(n15762), .IN2(n15763), .QN(g26675) );
  NAND2X0 U15846 ( .IN1(n15764), .IN2(g1783), .QN(n15763) );
  NAND2X0 U15847 ( .IN1(n11720), .IN2(n13315), .QN(n15764) );
  NAND2X0 U15848 ( .IN1(n15765), .IN2(n13315), .QN(n15762) );
  INVX0 U15849 ( .INP(n4511), .ZN(n13315) );
  NAND2X0 U15850 ( .IN1(n15766), .IN2(n15767), .QN(g26672) );
  NAND2X0 U15851 ( .IN1(n15768), .IN2(g2478), .QN(n15767) );
  NAND2X0 U15852 ( .IN1(n15760), .IN2(n13416), .QN(n15768) );
  NAND2X0 U15853 ( .IN1(n15761), .IN2(n13416), .QN(n15766) );
  INVX0 U15854 ( .INP(n4516), .ZN(n13416) );
  NOR2X0 U15855 ( .IN1(n15769), .IN2(n15770), .QN(g26671) );
  NAND2X0 U15856 ( .IN1(n14842), .IN2(n14703), .QN(n15770) );
  NAND2X0 U15857 ( .IN1(n15771), .IN2(n15772), .QN(n14842) );
  NOR2X0 U15858 ( .IN1(n4409), .IN2(n4399), .QN(n15771) );
  NOR2X0 U15859 ( .IN1(n15773), .IN2(g2052), .QN(n15769) );
  NOR2X0 U15860 ( .IN1(n4399), .IN2(n15774), .QN(n15773) );
  NAND2X0 U15861 ( .IN1(n15775), .IN2(n15776), .QN(g26670) );
  NAND2X0 U15862 ( .IN1(n15777), .IN2(g1785), .QN(n15776) );
  NAND2X0 U15863 ( .IN1(n11720), .IN2(n11946), .QN(n15777) );
  NAND2X0 U15864 ( .IN1(n15765), .IN2(n11946), .QN(n15775) );
  NAND2X0 U15865 ( .IN1(n15778), .IN2(n15779), .QN(g26669) );
  NAND2X0 U15866 ( .IN1(n15780), .IN2(g1089), .QN(n15779) );
  NAND2X0 U15867 ( .IN1(n11719), .IN2(g1088), .QN(n15780) );
  NAND2X0 U15868 ( .IN1(n15781), .IN2(g1088), .QN(n15778) );
  NAND2X0 U15869 ( .IN1(n15782), .IN2(n15783), .QN(g26667) );
  NAND2X0 U15870 ( .IN1(test_so60), .IN2(n15784), .QN(n15783) );
  NAND2X0 U15871 ( .IN1(n11720), .IN2(n13555), .QN(n15784) );
  NAND2X0 U15872 ( .IN1(n15765), .IN2(n13555), .QN(n15782) );
  INVX0 U15873 ( .INP(n4518), .ZN(n13555) );
  NOR2X0 U15874 ( .IN1(n11720), .IN2(n4386), .QN(n15765) );
  NOR2X0 U15875 ( .IN1(n15785), .IN2(n13230), .QN(n11720) );
  NAND2X0 U15876 ( .IN1(n15786), .IN2(n15787), .QN(n13230) );
  NAND2X0 U15877 ( .IN1(n9980), .IN2(n11946), .QN(n15787) );
  NOR2X0 U15878 ( .IN1(n15788), .IN2(n15789), .QN(n15786) );
  NOR2X0 U15879 ( .IN1(test_so60), .IN2(n4518), .QN(n15789) );
  NOR2X0 U15880 ( .IN1(n4511), .IN2(g1783), .QN(n15788) );
  NAND2X0 U15881 ( .IN1(g1690), .IN2(n13229), .QN(n15785) );
  INVX0 U15882 ( .INP(n13001), .ZN(n13229) );
  NAND2X0 U15883 ( .IN1(n15790), .IN2(n15791), .QN(n13001) );
  NOR2X0 U15884 ( .IN1(n15792), .IN2(n15793), .QN(n15791) );
  NAND2X0 U15885 ( .IN1(n15794), .IN2(n15795), .QN(n15793) );
  NOR2X0 U15886 ( .IN1(n15796), .IN2(n15797), .QN(n15795) );
  NOR2X0 U15887 ( .IN1(n12365), .IN2(n15798), .QN(n15797) );
  INVX0 U15888 ( .INP(n15799), .ZN(n15796) );
  NAND2X0 U15889 ( .IN1(n15798), .IN2(n12365), .QN(n15799) );
  NAND2X0 U15890 ( .IN1(n15800), .IN2(n15801), .QN(n15798) );
  NAND2X0 U15891 ( .IN1(n9829), .IN2(g6782), .QN(n15801) );
  NOR2X0 U15892 ( .IN1(n15802), .IN2(n15803), .QN(n15800) );
  NOR2X0 U15893 ( .IN1(n4368), .IN2(g1541), .QN(n15803) );
  NOR2X0 U15894 ( .IN1(n4317), .IN2(g1542), .QN(n15802) );
  NOR2X0 U15895 ( .IN1(n15804), .IN2(n15805), .QN(n15794) );
  NAND2X0 U15896 ( .IN1(n15806), .IN2(n15807), .QN(n15805) );
  NAND2X0 U15897 ( .IN1(n12132), .IN2(n15808), .QN(n15807) );
  INVX0 U15898 ( .INP(n15809), .ZN(n15806) );
  NOR2X0 U15899 ( .IN1(n15808), .IN2(n12132), .QN(n15809) );
  NAND2X0 U15900 ( .IN1(n15810), .IN2(n15811), .QN(n15808) );
  NAND2X0 U15901 ( .IN1(n9845), .IN2(g6782), .QN(n15811) );
  NOR2X0 U15902 ( .IN1(n15812), .IN2(n15813), .QN(n15810) );
  NOR2X0 U15903 ( .IN1(n4368), .IN2(g1544), .QN(n15813) );
  NOR2X0 U15904 ( .IN1(n4317), .IN2(g1545), .QN(n15812) );
  NAND2X0 U15905 ( .IN1(n15814), .IN2(n15815), .QN(n15804) );
  NAND2X0 U15906 ( .IN1(n4320), .IN2(n15816), .QN(n15815) );
  INVX0 U15907 ( .INP(n15817), .ZN(n15814) );
  NOR2X0 U15908 ( .IN1(n15816), .IN2(n4320), .QN(n15817) );
  NAND2X0 U15909 ( .IN1(n15818), .IN2(n15819), .QN(n15816) );
  NAND2X0 U15910 ( .IN1(n9852), .IN2(g1547), .QN(n15819) );
  NOR2X0 U15911 ( .IN1(n15820), .IN2(n15821), .QN(n15818) );
  NOR2X0 U15912 ( .IN1(n4317), .IN2(g1524), .QN(n15821) );
  NOR2X0 U15913 ( .IN1(n4515), .IN2(g1525), .QN(n15820) );
  NAND2X0 U15914 ( .IN1(n15822), .IN2(n15823), .QN(n15792) );
  NOR2X0 U15915 ( .IN1(n15824), .IN2(n15825), .QN(n15823) );
  NOR2X0 U15916 ( .IN1(n4374), .IN2(n15826), .QN(n15825) );
  INVX0 U15917 ( .INP(n15827), .ZN(n15824) );
  NAND2X0 U15918 ( .IN1(n15826), .IN2(n4374), .QN(n15827) );
  NAND2X0 U15919 ( .IN1(n15828), .IN2(n15829), .QN(n15826) );
  NAND2X0 U15920 ( .IN1(n9853), .IN2(g1547), .QN(n15829) );
  NOR2X0 U15921 ( .IN1(n15830), .IN2(n15831), .QN(n15828) );
  NOR2X0 U15922 ( .IN1(test_so52), .IN2(n4317), .QN(n15831) );
  NOR2X0 U15923 ( .IN1(n4515), .IN2(g1516), .QN(n15830) );
  NOR2X0 U15924 ( .IN1(n13613), .IN2(n15832), .QN(n15822) );
  NAND2X0 U15925 ( .IN1(n15833), .IN2(n15834), .QN(n15832) );
  NAND2X0 U15926 ( .IN1(n4378), .IN2(n15835), .QN(n15834) );
  INVX0 U15927 ( .INP(n15836), .ZN(n15833) );
  NOR2X0 U15928 ( .IN1(n15835), .IN2(n4378), .QN(n15836) );
  NAND2X0 U15929 ( .IN1(n15837), .IN2(n15838), .QN(n15835) );
  NAND2X0 U15930 ( .IN1(n9854), .IN2(g1547), .QN(n15838) );
  NOR2X0 U15931 ( .IN1(n15839), .IN2(n15840), .QN(n15837) );
  NOR2X0 U15932 ( .IN1(n4317), .IN2(g1512), .QN(n15840) );
  NOR2X0 U15933 ( .IN1(n4515), .IN2(g1513), .QN(n15839) );
  INVX0 U15934 ( .INP(n3070), .ZN(n13613) );
  NOR2X0 U15935 ( .IN1(n15841), .IN2(n15842), .QN(n15790) );
  NAND2X0 U15936 ( .IN1(n15843), .IN2(n15844), .QN(n15842) );
  NOR2X0 U15937 ( .IN1(n15845), .IN2(n15846), .QN(n15844) );
  INVX0 U15938 ( .INP(n15847), .ZN(n15846) );
  NAND2X0 U15939 ( .IN1(g1501), .IN2(n15848), .QN(n15847) );
  NOR2X0 U15940 ( .IN1(n15848), .IN2(g1501), .QN(n15845) );
  NOR2X0 U15941 ( .IN1(n15849), .IN2(n15850), .QN(n15848) );
  NOR2X0 U15942 ( .IN1(n4515), .IN2(test_so53), .QN(n15850) );
  INVX0 U15943 ( .INP(n15851), .ZN(n15849) );
  NOR2X0 U15944 ( .IN1(n15852), .IN2(n15853), .QN(n15851) );
  NOR2X0 U15945 ( .IN1(n4368), .IN2(g1535), .QN(n15853) );
  NOR2X0 U15946 ( .IN1(n4317), .IN2(g1536), .QN(n15852) );
  NOR2X0 U15947 ( .IN1(n15854), .IN2(n15855), .QN(n15843) );
  NOR2X0 U15948 ( .IN1(n4390), .IN2(n15856), .QN(n15855) );
  INVX0 U15949 ( .INP(n15857), .ZN(n15854) );
  NAND2X0 U15950 ( .IN1(n15856), .IN2(n4390), .QN(n15857) );
  NAND2X0 U15951 ( .IN1(n15858), .IN2(n15859), .QN(n15856) );
  NAND2X0 U15952 ( .IN1(n9851), .IN2(g1547), .QN(n15859) );
  NOR2X0 U15953 ( .IN1(n15860), .IN2(n15861), .QN(n15858) );
  NOR2X0 U15954 ( .IN1(n4317), .IN2(g1527), .QN(n15861) );
  NOR2X0 U15955 ( .IN1(n4515), .IN2(g1528), .QN(n15860) );
  NAND2X0 U15956 ( .IN1(n15862), .IN2(n15863), .QN(n15841) );
  NOR2X0 U15957 ( .IN1(n15864), .IN2(n15865), .QN(n15863) );
  NOR2X0 U15958 ( .IN1(n4326), .IN2(n15866), .QN(n15865) );
  INVX0 U15959 ( .INP(n15867), .ZN(n15864) );
  NAND2X0 U15960 ( .IN1(n15866), .IN2(n4326), .QN(n15867) );
  NAND2X0 U15961 ( .IN1(n15868), .IN2(n15869), .QN(n15866) );
  NAND2X0 U15962 ( .IN1(n9850), .IN2(g1547), .QN(n15869) );
  NOR2X0 U15963 ( .IN1(n15870), .IN2(n15871), .QN(n15868) );
  NOR2X0 U15964 ( .IN1(n4317), .IN2(g1530), .QN(n15871) );
  NOR2X0 U15965 ( .IN1(n4515), .IN2(g1531), .QN(n15870) );
  NOR2X0 U15966 ( .IN1(n15872), .IN2(n15873), .QN(n15862) );
  NAND2X0 U15967 ( .IN1(n15874), .IN2(n15875), .QN(n15873) );
  NAND2X0 U15968 ( .IN1(n4288), .IN2(n15876), .QN(n15875) );
  INVX0 U15969 ( .INP(n15877), .ZN(n15874) );
  NOR2X0 U15970 ( .IN1(n15876), .IN2(n4288), .QN(n15877) );
  NAND2X0 U15971 ( .IN1(n15878), .IN2(n15879), .QN(n15876) );
  NAND2X0 U15972 ( .IN1(n9847), .IN2(g1547), .QN(n15879) );
  NOR2X0 U15973 ( .IN1(n15880), .IN2(n15881), .QN(n15878) );
  NOR2X0 U15974 ( .IN1(n4317), .IN2(g1539), .QN(n15881) );
  NOR2X0 U15975 ( .IN1(n4515), .IN2(g1540), .QN(n15880) );
  NAND2X0 U15976 ( .IN1(n15882), .IN2(n15883), .QN(n15872) );
  NAND2X0 U15977 ( .IN1(n4557), .IN2(n15884), .QN(n15883) );
  INVX0 U15978 ( .INP(n15885), .ZN(n15882) );
  NOR2X0 U15979 ( .IN1(n15884), .IN2(n4557), .QN(n15885) );
  NAND2X0 U15980 ( .IN1(n15886), .IN2(n15887), .QN(n15884) );
  NAND2X0 U15981 ( .IN1(n9849), .IN2(g1547), .QN(n15887) );
  NOR2X0 U15982 ( .IN1(n15888), .IN2(n15889), .QN(n15886) );
  NOR2X0 U15983 ( .IN1(n4317), .IN2(g1533), .QN(n15889) );
  NOR2X0 U15984 ( .IN1(n4515), .IN2(g1534), .QN(n15888) );
  NOR2X0 U15985 ( .IN1(n15890), .IN2(n15891), .QN(g26666) );
  NAND2X0 U15986 ( .IN1(n14848), .IN2(n14834), .QN(n15891) );
  NAND2X0 U15987 ( .IN1(n15892), .IN2(n15893), .QN(n14848) );
  NOR2X0 U15988 ( .IN1(n4411), .IN2(n4401), .QN(n15892) );
  NOR2X0 U15989 ( .IN1(n15894), .IN2(g1358), .QN(n15890) );
  NOR2X0 U15990 ( .IN1(n4401), .IN2(n15895), .QN(n15894) );
  NAND2X0 U15991 ( .IN1(n15896), .IN2(n15897), .QN(g26665) );
  NAND2X0 U15992 ( .IN1(n15898), .IN2(g1091), .QN(n15897) );
  NAND2X0 U15993 ( .IN1(n11719), .IN2(g6712), .QN(n15898) );
  NAND2X0 U15994 ( .IN1(n15781), .IN2(g6712), .QN(n15896) );
  NAND2X0 U15995 ( .IN1(n15899), .IN2(n15900), .QN(g26664) );
  NAND2X0 U15996 ( .IN1(n15901), .IN2(g402), .QN(n15900) );
  NAND2X0 U15997 ( .IN1(n11718), .IN2(n13361), .QN(n15901) );
  NAND2X0 U15998 ( .IN1(n15902), .IN2(n13361), .QN(n15899) );
  INVX0 U15999 ( .INP(n4506), .ZN(n13361) );
  NAND2X0 U16000 ( .IN1(n15903), .IN2(n15904), .QN(g26661) );
  NAND2X0 U16001 ( .IN1(n15905), .IN2(g1090), .QN(n15904) );
  NAND2X0 U16002 ( .IN1(n11719), .IN2(g5472), .QN(n15905) );
  NAND2X0 U16003 ( .IN1(n15781), .IN2(g5472), .QN(n15903) );
  NOR2X0 U16004 ( .IN1(n11719), .IN2(n4387), .QN(n15781) );
  NOR2X0 U16005 ( .IN1(n15906), .IN2(n13245), .QN(n11719) );
  NAND2X0 U16006 ( .IN1(n15907), .IN2(n15908), .QN(n13245) );
  NAND2X0 U16007 ( .IN1(n9995), .IN2(g1088), .QN(n15908) );
  NOR2X0 U16008 ( .IN1(n15909), .IN2(n15910), .QN(n15907) );
  NOR2X0 U16009 ( .IN1(n4364), .IN2(g1091), .QN(n15910) );
  NOR2X0 U16010 ( .IN1(n4363), .IN2(g1090), .QN(n15909) );
  NAND2X0 U16011 ( .IN1(g996), .IN2(n13067), .QN(n15906) );
  INVX0 U16012 ( .INP(n15911), .ZN(n13067) );
  NAND2X0 U16013 ( .IN1(n15912), .IN2(n15913), .QN(n15911) );
  NOR2X0 U16014 ( .IN1(n15914), .IN2(n15915), .QN(n15913) );
  NAND2X0 U16015 ( .IN1(n15916), .IN2(n15917), .QN(n15915) );
  NOR2X0 U16016 ( .IN1(n15918), .IN2(n15919), .QN(n15917) );
  NOR2X0 U16017 ( .IN1(n13804), .IN2(n15920), .QN(n15919) );
  INVX0 U16018 ( .INP(n15921), .ZN(n15918) );
  NAND2X0 U16019 ( .IN1(n15920), .IN2(n13804), .QN(n15921) );
  NAND2X0 U16020 ( .IN1(n15922), .IN2(n15923), .QN(n15920) );
  NAND2X0 U16021 ( .IN1(n9858), .IN2(test_so31), .QN(n15923) );
  NOR2X0 U16022 ( .IN1(n15924), .IN2(n15925), .QN(n15922) );
  NOR2X0 U16023 ( .IN1(n4323), .IN2(g848), .QN(n15925) );
  NOR2X0 U16024 ( .IN1(n4312), .IN2(g849), .QN(n15924) );
  NOR2X0 U16025 ( .IN1(n15926), .IN2(n15927), .QN(n15916) );
  NAND2X0 U16026 ( .IN1(n15928), .IN2(n15929), .QN(n15927) );
  NAND2X0 U16027 ( .IN1(n12178), .IN2(n15930), .QN(n15929) );
  INVX0 U16028 ( .INP(n15931), .ZN(n15928) );
  NOR2X0 U16029 ( .IN1(n15930), .IN2(n12178), .QN(n15931) );
  NAND2X0 U16030 ( .IN1(n15932), .IN2(n15933), .QN(n15930) );
  NAND2X0 U16031 ( .IN1(n9855), .IN2(test_so31), .QN(n15933) );
  NOR2X0 U16032 ( .IN1(n15934), .IN2(n15935), .QN(n15932) );
  NOR2X0 U16033 ( .IN1(n4323), .IN2(g851), .QN(n15935) );
  NOR2X0 U16034 ( .IN1(n4312), .IN2(g852), .QN(n15934) );
  NAND2X0 U16035 ( .IN1(n15936), .IN2(n15937), .QN(n15926) );
  NAND2X0 U16036 ( .IN1(n4321), .IN2(n15938), .QN(n15937) );
  INVX0 U16037 ( .INP(n15939), .ZN(n15936) );
  NOR2X0 U16038 ( .IN1(n15938), .IN2(n4321), .QN(n15939) );
  NAND2X0 U16039 ( .IN1(n15940), .IN2(n15941), .QN(n15938) );
  NAND2X0 U16040 ( .IN1(n9866), .IN2(test_so31), .QN(n15941) );
  NOR2X0 U16041 ( .IN1(n15942), .IN2(n15943), .QN(n15940) );
  NOR2X0 U16042 ( .IN1(n4323), .IN2(g830), .QN(n15943) );
  NOR2X0 U16043 ( .IN1(n4312), .IN2(g831), .QN(n15942) );
  NAND2X0 U16044 ( .IN1(n15944), .IN2(n15945), .QN(n15914) );
  NOR2X0 U16045 ( .IN1(n15946), .IN2(n15947), .QN(n15945) );
  NOR2X0 U16046 ( .IN1(n4375), .IN2(n15948), .QN(n15947) );
  INVX0 U16047 ( .INP(n15949), .ZN(n15946) );
  NAND2X0 U16048 ( .IN1(n15948), .IN2(n4375), .QN(n15949) );
  NAND2X0 U16049 ( .IN1(n15950), .IN2(n15951), .QN(n15948) );
  NAND2X0 U16050 ( .IN1(n9867), .IN2(test_so31), .QN(n15951) );
  NOR2X0 U16051 ( .IN1(n15952), .IN2(n15953), .QN(n15950) );
  NOR2X0 U16052 ( .IN1(n4323), .IN2(g821), .QN(n15953) );
  NOR2X0 U16053 ( .IN1(n4312), .IN2(g822), .QN(n15952) );
  NOR2X0 U16054 ( .IN1(n11799), .IN2(n15954), .QN(n15944) );
  NAND2X0 U16055 ( .IN1(n15955), .IN2(n15956), .QN(n15954) );
  NAND2X0 U16056 ( .IN1(n4379), .IN2(n15957), .QN(n15956) );
  INVX0 U16057 ( .INP(n15958), .ZN(n15955) );
  NOR2X0 U16058 ( .IN1(n15957), .IN2(n4379), .QN(n15958) );
  NAND2X0 U16059 ( .IN1(n15959), .IN2(n15960), .QN(n15957) );
  NAND2X0 U16060 ( .IN1(n9868), .IN2(test_so31), .QN(n15960) );
  NOR2X0 U16061 ( .IN1(n15961), .IN2(n15962), .QN(n15959) );
  NOR2X0 U16062 ( .IN1(n4323), .IN2(g818), .QN(n15962) );
  NOR2X0 U16063 ( .IN1(n4312), .IN2(g819), .QN(n15961) );
  INVX0 U16064 ( .INP(n3102), .ZN(n11799) );
  NOR2X0 U16065 ( .IN1(n15963), .IN2(n15964), .QN(n15912) );
  NAND2X0 U16066 ( .IN1(n15965), .IN2(n15966), .QN(n15964) );
  NOR2X0 U16067 ( .IN1(n15967), .IN2(n15968), .QN(n15966) );
  NOR2X0 U16068 ( .IN1(n4567), .IN2(n15969), .QN(n15968) );
  INVX0 U16069 ( .INP(n15970), .ZN(n15967) );
  NAND2X0 U16070 ( .IN1(n15969), .IN2(n4567), .QN(n15970) );
  NAND2X0 U16071 ( .IN1(n15971), .IN2(n15972), .QN(n15969) );
  NAND2X0 U16072 ( .IN1(n9862), .IN2(test_so31), .QN(n15972) );
  NOR2X0 U16073 ( .IN1(n15973), .IN2(n15974), .QN(n15971) );
  NOR2X0 U16074 ( .IN1(n4323), .IN2(g842), .QN(n15974) );
  NOR2X0 U16075 ( .IN1(n4312), .IN2(g843), .QN(n15973) );
  NOR2X0 U16076 ( .IN1(n15975), .IN2(n15976), .QN(n15965) );
  NOR2X0 U16077 ( .IN1(n4391), .IN2(n15977), .QN(n15976) );
  INVX0 U16078 ( .INP(n15978), .ZN(n15975) );
  NAND2X0 U16079 ( .IN1(n15977), .IN2(n4391), .QN(n15978) );
  NAND2X0 U16080 ( .IN1(n15979), .IN2(n15980), .QN(n15977) );
  NAND2X0 U16081 ( .IN1(n9865), .IN2(test_so31), .QN(n15980) );
  NOR2X0 U16082 ( .IN1(n15981), .IN2(n15982), .QN(n15979) );
  NOR2X0 U16083 ( .IN1(n4323), .IN2(g833), .QN(n15982) );
  NOR2X0 U16084 ( .IN1(n4312), .IN2(g834), .QN(n15981) );
  NAND2X0 U16085 ( .IN1(n15983), .IN2(n15984), .QN(n15963) );
  NOR2X0 U16086 ( .IN1(n15985), .IN2(n15986), .QN(n15984) );
  NOR2X0 U16087 ( .IN1(n4327), .IN2(n15987), .QN(n15986) );
  INVX0 U16088 ( .INP(n15988), .ZN(n15985) );
  NAND2X0 U16089 ( .IN1(n15987), .IN2(n4327), .QN(n15988) );
  NAND2X0 U16090 ( .IN1(n15989), .IN2(n15990), .QN(n15987) );
  NAND2X0 U16091 ( .IN1(n9864), .IN2(test_so31), .QN(n15990) );
  NOR2X0 U16092 ( .IN1(n15991), .IN2(n15992), .QN(n15989) );
  NOR2X0 U16093 ( .IN1(n4323), .IN2(g836), .QN(n15992) );
  NOR2X0 U16094 ( .IN1(n4312), .IN2(g837), .QN(n15991) );
  NOR2X0 U16095 ( .IN1(n15993), .IN2(n15994), .QN(n15983) );
  NAND2X0 U16096 ( .IN1(n15995), .IN2(n15996), .QN(n15994) );
  NAND2X0 U16097 ( .IN1(n4289), .IN2(n15997), .QN(n15996) );
  INVX0 U16098 ( .INP(n15998), .ZN(n15995) );
  NOR2X0 U16099 ( .IN1(n15997), .IN2(n4289), .QN(n15998) );
  NAND2X0 U16100 ( .IN1(n15999), .IN2(n16000), .QN(n15997) );
  NAND2X0 U16101 ( .IN1(n9861), .IN2(test_so31), .QN(n16000) );
  NOR2X0 U16102 ( .IN1(n16001), .IN2(n16002), .QN(n15999) );
  NOR2X0 U16103 ( .IN1(n4323), .IN2(g845), .QN(n16002) );
  NOR2X0 U16104 ( .IN1(n4312), .IN2(g846), .QN(n16001) );
  NAND2X0 U16105 ( .IN1(n16003), .IN2(n16004), .QN(n15993) );
  NAND2X0 U16106 ( .IN1(n4559), .IN2(n16005), .QN(n16004) );
  INVX0 U16107 ( .INP(n16006), .ZN(n16003) );
  NOR2X0 U16108 ( .IN1(n16005), .IN2(n4559), .QN(n16006) );
  NAND2X0 U16109 ( .IN1(n16007), .IN2(n16008), .QN(n16005) );
  NAND2X0 U16110 ( .IN1(n9863), .IN2(test_so31), .QN(n16008) );
  NOR2X0 U16111 ( .IN1(n16009), .IN2(n16010), .QN(n16007) );
  NOR2X0 U16112 ( .IN1(test_so32), .IN2(n4323), .QN(n16010) );
  NOR2X0 U16113 ( .IN1(n4312), .IN2(g840), .QN(n16009) );
  NOR2X0 U16114 ( .IN1(n16011), .IN2(n16012), .QN(g26660) );
  NAND2X0 U16115 ( .IN1(n14852), .IN2(n14712), .QN(n16012) );
  NAND2X0 U16116 ( .IN1(n16013), .IN2(n16014), .QN(n14852) );
  NOR2X0 U16117 ( .IN1(n4413), .IN2(n4403), .QN(n16013) );
  NOR2X0 U16118 ( .IN1(n16015), .IN2(g672), .QN(n16011) );
  NOR2X0 U16119 ( .IN1(n4403), .IN2(n16016), .QN(n16015) );
  NAND2X0 U16120 ( .IN1(n16017), .IN2(n16018), .QN(g26659) );
  NAND2X0 U16121 ( .IN1(n16019), .IN2(g404), .QN(n16018) );
  NAND2X0 U16122 ( .IN1(n11718), .IN2(n13382), .QN(n16019) );
  NAND2X0 U16123 ( .IN1(n15902), .IN2(n13382), .QN(n16017) );
  INVX0 U16124 ( .INP(n4499), .ZN(n13382) );
  NAND2X0 U16125 ( .IN1(n16020), .IN2(n16021), .QN(g26655) );
  NAND2X0 U16126 ( .IN1(n16022), .IN2(g403), .QN(n16021) );
  NAND2X0 U16127 ( .IN1(n11718), .IN2(n12042), .QN(n16022) );
  NAND2X0 U16128 ( .IN1(n15902), .IN2(n12042), .QN(n16020) );
  NOR2X0 U16129 ( .IN1(n11718), .IN2(n4388), .QN(n15902) );
  NOR2X0 U16130 ( .IN1(n16023), .IN2(n13256), .QN(n11718) );
  NAND2X0 U16131 ( .IN1(n16024), .IN2(n16025), .QN(n13256) );
  NAND2X0 U16132 ( .IN1(n10003), .IN2(n12042), .QN(n16025) );
  NOR2X0 U16133 ( .IN1(n16026), .IN2(n16027), .QN(n16024) );
  NOR2X0 U16134 ( .IN1(n4499), .IN2(g404), .QN(n16027) );
  NOR2X0 U16135 ( .IN1(n4506), .IN2(g402), .QN(n16026) );
  NAND2X0 U16136 ( .IN1(g309), .IN2(n13255), .QN(n16023) );
  INVX0 U16137 ( .INP(n13136), .ZN(n13255) );
  NAND2X0 U16138 ( .IN1(n16028), .IN2(n16029), .QN(n13136) );
  NOR2X0 U16139 ( .IN1(n16030), .IN2(n16031), .QN(n16029) );
  NAND2X0 U16140 ( .IN1(n16032), .IN2(n16033), .QN(n16031) );
  NOR2X0 U16141 ( .IN1(n16034), .IN2(n16035), .QN(n16033) );
  NOR2X0 U16142 ( .IN1(n12454), .IN2(n16036), .QN(n16035) );
  INVX0 U16143 ( .INP(n16037), .ZN(n16034) );
  NAND2X0 U16144 ( .IN1(n16036), .IN2(n12454), .QN(n16037) );
  NAND2X0 U16145 ( .IN1(n16038), .IN2(n16039), .QN(n16036) );
  NAND2X0 U16146 ( .IN1(n9832), .IN2(g6313), .QN(n16039) );
  NOR2X0 U16147 ( .IN1(n16040), .IN2(n16041), .QN(n16038) );
  NOR2X0 U16148 ( .IN1(n4369), .IN2(g159), .QN(n16041) );
  NOR2X0 U16149 ( .IN1(n4318), .IN2(g160), .QN(n16040) );
  NOR2X0 U16150 ( .IN1(n16042), .IN2(n16043), .QN(n16032) );
  NAND2X0 U16151 ( .IN1(n16044), .IN2(n16045), .QN(n16043) );
  NAND2X0 U16152 ( .IN1(n12247), .IN2(n16046), .QN(n16045) );
  INVX0 U16153 ( .INP(n16047), .ZN(n16044) );
  NOR2X0 U16154 ( .IN1(n16046), .IN2(n12247), .QN(n16047) );
  NAND2X0 U16155 ( .IN1(n16048), .IN2(n16049), .QN(n16046) );
  NAND2X0 U16156 ( .IN1(n9870), .IN2(g6313), .QN(n16049) );
  NOR2X0 U16157 ( .IN1(n16050), .IN2(n16051), .QN(n16048) );
  NOR2X0 U16158 ( .IN1(n4369), .IN2(g162), .QN(n16051) );
  NOR2X0 U16159 ( .IN1(test_so12), .IN2(n4318), .QN(n16050) );
  NAND2X0 U16160 ( .IN1(n16052), .IN2(n16053), .QN(n16042) );
  NAND2X0 U16161 ( .IN1(n4322), .IN2(n16054), .QN(n16053) );
  INVX0 U16162 ( .INP(n16055), .ZN(n16052) );
  NOR2X0 U16163 ( .IN1(n16054), .IN2(n4322), .QN(n16055) );
  NAND2X0 U16164 ( .IN1(n16056), .IN2(n16057), .QN(n16054) );
  NAND2X0 U16165 ( .IN1(n9875), .IN2(g165), .QN(n16057) );
  NOR2X0 U16166 ( .IN1(n16058), .IN2(n16059), .QN(n16056) );
  NOR2X0 U16167 ( .IN1(n4318), .IN2(g142), .QN(n16059) );
  NOR2X0 U16168 ( .IN1(n4512), .IN2(g143), .QN(n16058) );
  NAND2X0 U16169 ( .IN1(n16060), .IN2(n16061), .QN(n16030) );
  NOR2X0 U16170 ( .IN1(n16062), .IN2(n16063), .QN(n16061) );
  NOR2X0 U16171 ( .IN1(n4376), .IN2(n16064), .QN(n16063) );
  INVX0 U16172 ( .INP(n16065), .ZN(n16062) );
  NAND2X0 U16173 ( .IN1(n16064), .IN2(n4376), .QN(n16065) );
  NAND2X0 U16174 ( .IN1(n16066), .IN2(n16067), .QN(n16064) );
  NAND2X0 U16175 ( .IN1(n9876), .IN2(g165), .QN(n16067) );
  NOR2X0 U16176 ( .IN1(n16068), .IN2(n16069), .QN(n16066) );
  NOR2X0 U16177 ( .IN1(n4318), .IN2(g133), .QN(n16069) );
  NOR2X0 U16178 ( .IN1(n4512), .IN2(g134), .QN(n16068) );
  NOR2X0 U16179 ( .IN1(n13884), .IN2(n16070), .QN(n16060) );
  NAND2X0 U16180 ( .IN1(n16071), .IN2(n16072), .QN(n16070) );
  NAND2X0 U16181 ( .IN1(n4380), .IN2(n16073), .QN(n16072) );
  INVX0 U16182 ( .INP(n16074), .ZN(n16071) );
  NOR2X0 U16183 ( .IN1(n16073), .IN2(n4380), .QN(n16074) );
  NAND2X0 U16184 ( .IN1(n16075), .IN2(n16076), .QN(n16073) );
  NAND2X0 U16185 ( .IN1(n9877), .IN2(g165), .QN(n16076) );
  NOR2X0 U16186 ( .IN1(n16077), .IN2(n16078), .QN(n16075) );
  NOR2X0 U16187 ( .IN1(n4318), .IN2(g130), .QN(n16078) );
  NOR2X0 U16188 ( .IN1(n4512), .IN2(g131), .QN(n16077) );
  INVX0 U16189 ( .INP(n3130), .ZN(n13884) );
  NOR2X0 U16190 ( .IN1(n16079), .IN2(n16080), .QN(n16028) );
  NAND2X0 U16191 ( .IN1(n16081), .IN2(n16082), .QN(n16080) );
  NOR2X0 U16192 ( .IN1(n16083), .IN2(n16084), .QN(n16082) );
  NOR2X0 U16193 ( .IN1(n4569), .IN2(n16085), .QN(n16084) );
  INVX0 U16194 ( .INP(n16086), .ZN(n16083) );
  NAND2X0 U16195 ( .IN1(n16085), .IN2(n4569), .QN(n16086) );
  NAND2X0 U16196 ( .IN1(n16087), .IN2(n16088), .QN(n16085) );
  NAND2X0 U16197 ( .IN1(n9872), .IN2(g165), .QN(n16088) );
  NOR2X0 U16198 ( .IN1(n16089), .IN2(n16090), .QN(n16087) );
  NOR2X0 U16199 ( .IN1(n4318), .IN2(g154), .QN(n16090) );
  NOR2X0 U16200 ( .IN1(n4512), .IN2(g155), .QN(n16089) );
  NOR2X0 U16201 ( .IN1(n16091), .IN2(n16092), .QN(n16081) );
  INVX0 U16202 ( .INP(n16093), .ZN(n16092) );
  NAND2X0 U16203 ( .IN1(g109), .IN2(n16094), .QN(n16093) );
  NOR2X0 U16204 ( .IN1(n16094), .IN2(g109), .QN(n16091) );
  NOR2X0 U16205 ( .IN1(n16095), .IN2(n16096), .QN(n16094) );
  NOR2X0 U16206 ( .IN1(n4369), .IN2(test_so11), .QN(n16096) );
  INVX0 U16207 ( .INP(n16097), .ZN(n16095) );
  NOR2X0 U16208 ( .IN1(n16098), .IN2(n16099), .QN(n16097) );
  NOR2X0 U16209 ( .IN1(n4318), .IN2(g145), .QN(n16099) );
  NOR2X0 U16210 ( .IN1(n4512), .IN2(g146), .QN(n16098) );
  NAND2X0 U16211 ( .IN1(n16100), .IN2(n16101), .QN(n16079) );
  NOR2X0 U16212 ( .IN1(n16102), .IN2(n16103), .QN(n16101) );
  NOR2X0 U16213 ( .IN1(n4328), .IN2(n16104), .QN(n16103) );
  INVX0 U16214 ( .INP(n16105), .ZN(n16102) );
  NAND2X0 U16215 ( .IN1(n16104), .IN2(n4328), .QN(n16105) );
  NAND2X0 U16216 ( .IN1(n16106), .IN2(n16107), .QN(n16104) );
  NAND2X0 U16217 ( .IN1(n9874), .IN2(g165), .QN(n16107) );
  NOR2X0 U16218 ( .IN1(n16108), .IN2(n16109), .QN(n16106) );
  NOR2X0 U16219 ( .IN1(n4318), .IN2(g148), .QN(n16109) );
  NOR2X0 U16220 ( .IN1(n4512), .IN2(g149), .QN(n16108) );
  NOR2X0 U16221 ( .IN1(n16110), .IN2(n16111), .QN(n16100) );
  NAND2X0 U16222 ( .IN1(n16112), .IN2(n16113), .QN(n16111) );
  NAND2X0 U16223 ( .IN1(n4290), .IN2(n16114), .QN(n16113) );
  INVX0 U16224 ( .INP(n16115), .ZN(n16112) );
  NOR2X0 U16225 ( .IN1(n16114), .IN2(n4290), .QN(n16115) );
  NAND2X0 U16226 ( .IN1(n16116), .IN2(n16117), .QN(n16114) );
  NAND2X0 U16227 ( .IN1(n9871), .IN2(g165), .QN(n16117) );
  NOR2X0 U16228 ( .IN1(n16118), .IN2(n16119), .QN(n16116) );
  NOR2X0 U16229 ( .IN1(n4318), .IN2(g157), .QN(n16119) );
  NOR2X0 U16230 ( .IN1(n4512), .IN2(g158), .QN(n16118) );
  NAND2X0 U16231 ( .IN1(n16120), .IN2(n16121), .QN(n16110) );
  NAND2X0 U16232 ( .IN1(n4561), .IN2(n16122), .QN(n16121) );
  INVX0 U16233 ( .INP(n16123), .ZN(n16120) );
  NOR2X0 U16234 ( .IN1(n16122), .IN2(n4561), .QN(n16123) );
  NAND2X0 U16235 ( .IN1(n16124), .IN2(n16125), .QN(n16122) );
  NAND2X0 U16236 ( .IN1(n9873), .IN2(g165), .QN(n16125) );
  NOR2X0 U16237 ( .IN1(n16126), .IN2(n16127), .QN(n16124) );
  NOR2X0 U16238 ( .IN1(n4318), .IN2(g151), .QN(n16127) );
  NOR2X0 U16239 ( .IN1(n4512), .IN2(g152), .QN(n16126) );
  NAND2X0 U16240 ( .IN1(n16128), .IN2(n16129), .QN(g26616) );
  INVX0 U16241 ( .INP(n16130), .ZN(n16129) );
  NOR2X0 U16242 ( .IN1(g2624), .IN2(n9788), .QN(n16130) );
  NAND2X0 U16243 ( .IN1(n16131), .IN2(g2624), .QN(n16128) );
  NAND2X0 U16244 ( .IN1(n16132), .IN2(n16133), .QN(g26596) );
  NAND2X0 U16245 ( .IN1(n4370), .IN2(g2568), .QN(n16133) );
  NAND2X0 U16246 ( .IN1(n16131), .IN2(g7390), .QN(n16132) );
  NAND2X0 U16247 ( .IN1(n16134), .IN2(n16135), .QN(g26592) );
  NAND2X0 U16248 ( .IN1(n4366), .IN2(g1877), .QN(n16135) );
  NAND2X0 U16249 ( .IN1(n16136), .IN2(g1930), .QN(n16134) );
  NAND2X0 U16250 ( .IN1(n16137), .IN2(n16138), .QN(g26575) );
  INVX0 U16251 ( .INP(n16139), .ZN(n16138) );
  NOR2X0 U16252 ( .IN1(n13147), .IN2(n9786), .QN(n16139) );
  NAND2X0 U16253 ( .IN1(n16131), .IN2(n13147), .QN(n16137) );
  NOR2X0 U16254 ( .IN1(n16140), .IN2(n16141), .QN(n16131) );
  NAND2X0 U16255 ( .IN1(g2584), .IN2(n11267), .QN(n16140) );
  NAND2X0 U16256 ( .IN1(n16142), .IN2(n16143), .QN(g26573) );
  INVX0 U16257 ( .INP(n16144), .ZN(n16143) );
  NOR2X0 U16258 ( .IN1(g7194), .IN2(n9793), .QN(n16144) );
  NAND2X0 U16259 ( .IN1(n16136), .IN2(g7194), .QN(n16142) );
  NAND2X0 U16260 ( .IN1(n16145), .IN2(n16146), .QN(g26569) );
  INVX0 U16261 ( .INP(n16147), .ZN(n16146) );
  NOR2X0 U16262 ( .IN1(g1236), .IN2(n9790), .QN(n16147) );
  NAND2X0 U16263 ( .IN1(n16148), .IN2(g1236), .QN(n16145) );
  NAND2X0 U16264 ( .IN1(n16149), .IN2(n16150), .QN(g26559) );
  NAND2X0 U16265 ( .IN1(n16136), .IN2(n14321), .QN(n16150) );
  NOR2X0 U16266 ( .IN1(n16151), .IN2(n16152), .QN(n16136) );
  NAND2X0 U16267 ( .IN1(g1890), .IN2(n11438), .QN(n16151) );
  NAND2X0 U16268 ( .IN1(test_so68), .IN2(n4296), .QN(n16149) );
  NAND2X0 U16269 ( .IN1(n16153), .IN2(n16154), .QN(g26557) );
  INVX0 U16270 ( .INP(n16155), .ZN(n16154) );
  NOR2X0 U16271 ( .IN1(g6944), .IN2(n9794), .QN(n16155) );
  NAND2X0 U16272 ( .IN1(n16148), .IN2(g6944), .QN(n16153) );
  NAND2X0 U16273 ( .IN1(n16156), .IN2(n16157), .QN(g26553) );
  INVX0 U16274 ( .INP(n16158), .ZN(n16157) );
  NOR2X0 U16275 ( .IN1(g550), .IN2(n9791), .QN(n16158) );
  NAND2X0 U16276 ( .IN1(n16159), .IN2(g550), .QN(n16156) );
  NAND2X0 U16277 ( .IN1(n16160), .IN2(n16161), .QN(g26547) );
  NAND2X0 U16278 ( .IN1(n16148), .IN2(n14180), .QN(n16161) );
  NOR2X0 U16279 ( .IN1(n16162), .IN2(n16163), .QN(n16148) );
  NAND2X0 U16280 ( .IN1(g1196), .IN2(n11614), .QN(n16162) );
  NAND2X0 U16281 ( .IN1(test_so47), .IN2(n4371), .QN(n16160) );
  NAND2X0 U16282 ( .IN1(n16164), .IN2(n16165), .QN(g26545) );
  NAND2X0 U16283 ( .IN1(n4372), .IN2(g493), .QN(n16165) );
  NAND2X0 U16284 ( .IN1(n16159), .IN2(g6642), .QN(n16164) );
  NAND2X0 U16285 ( .IN1(n16166), .IN2(n16167), .QN(g26541) );
  INVX0 U16286 ( .INP(n16168), .ZN(n16167) );
  NOR2X0 U16287 ( .IN1(n14574), .IN2(n9787), .QN(n16168) );
  NAND2X0 U16288 ( .IN1(n16159), .IN2(n14574), .QN(n16166) );
  NOR2X0 U16289 ( .IN1(n16169), .IN2(n16170), .QN(n16159) );
  NAND2X0 U16290 ( .IN1(n11130), .IN2(test_so22), .QN(n16169) );
  NOR2X0 U16291 ( .IN1(n13263), .IN2(n16171), .QN(g26532) );
  NOR2X0 U16292 ( .IN1(n16172), .IN2(n16173), .QN(n16171) );
  NOR2X0 U16293 ( .IN1(n4526), .IN2(g2151), .QN(n16173) );
  NOR2X0 U16294 ( .IN1(n10012), .IN2(n16174), .QN(n16172) );
  NOR2X0 U16295 ( .IN1(n13268), .IN2(n16175), .QN(g26531) );
  NOR2X0 U16296 ( .IN1(n16176), .IN2(n16177), .QN(n16175) );
  NOR2X0 U16297 ( .IN1(n4527), .IN2(g1457), .QN(n16177) );
  NOR2X0 U16298 ( .IN1(n10016), .IN2(n16178), .QN(n16176) );
  NAND2X0 U16299 ( .IN1(n16179), .IN2(n16180), .QN(g26530) );
  NAND2X0 U16300 ( .IN1(n16181), .IN2(g771), .QN(n16180) );
  INVX0 U16301 ( .INP(n16182), .ZN(n16181) );
  NAND2X0 U16302 ( .IN1(n16183), .IN2(n10020), .QN(n16179) );
  NOR2X0 U16303 ( .IN1(n13273), .IN2(n3690), .QN(n16183) );
  NOR2X0 U16304 ( .IN1(n13278), .IN2(n16184), .QN(g26529) );
  NOR2X0 U16305 ( .IN1(n16185), .IN2(n16186), .QN(n16184) );
  NOR2X0 U16306 ( .IN1(n4528), .IN2(g83), .QN(n16186) );
  NOR2X0 U16307 ( .IN1(n10024), .IN2(n16187), .QN(n16185) );
  NAND2X0 U16308 ( .IN1(n16188), .IN2(n16189), .QN(g26149) );
  NOR2X0 U16309 ( .IN1(n16190), .IN2(n16191), .QN(n16189) );
  NAND2X0 U16310 ( .IN1(n16192), .IN2(n16193), .QN(n16191) );
  NAND2X0 U16311 ( .IN1(n16194), .IN2(g3161), .QN(n16193) );
  NOR2X0 U16312 ( .IN1(n16195), .IN2(n16196), .QN(n16192) );
  NOR2X0 U16313 ( .IN1(n4338), .IN2(n16197), .QN(n16196) );
  NOR2X0 U16314 ( .IN1(n4441), .IN2(n16198), .QN(n16195) );
  NAND2X0 U16315 ( .IN1(n16199), .IN2(n16200), .QN(n16190) );
  NAND2X0 U16316 ( .IN1(n3936), .IN2(n16201), .QN(n16200) );
  NAND2X0 U16317 ( .IN1(n16202), .IN2(n16203), .QN(n16201) );
  NOR2X0 U16318 ( .IN1(n16204), .IN2(n16205), .QN(n16203) );
  NOR2X0 U16319 ( .IN1(n4339), .IN2(n16206), .QN(n16205) );
  NOR2X0 U16320 ( .IN1(n4341), .IN2(n16207), .QN(n16204) );
  NOR2X0 U16321 ( .IN1(n16208), .IN2(n16209), .QN(n16202) );
  NOR2X0 U16322 ( .IN1(n4453), .IN2(n16210), .QN(n16209) );
  NOR2X0 U16323 ( .IN1(n4436), .IN2(n16211), .QN(n16208) );
  NOR2X0 U16324 ( .IN1(n16212), .IN2(n16213), .QN(n16199) );
  NOR2X0 U16325 ( .IN1(n16214), .IN2(n16215), .QN(n16213) );
  NOR2X0 U16326 ( .IN1(n16216), .IN2(n16217), .QN(n16214) );
  NAND2X0 U16327 ( .IN1(n16218), .IN2(n16219), .QN(n16217) );
  NAND2X0 U16328 ( .IN1(test_so8), .IN2(n16220), .QN(n16219) );
  NAND2X0 U16329 ( .IN1(n16221), .IN2(g3155), .QN(n16218) );
  NOR2X0 U16330 ( .IN1(n4442), .IN2(n16222), .QN(n16216) );
  NOR2X0 U16331 ( .IN1(n4348), .IN2(n16223), .QN(n16212) );
  NOR2X0 U16332 ( .IN1(n16224), .IN2(n16225), .QN(n16188) );
  NAND2X0 U16333 ( .IN1(n3700), .IN2(n16226), .QN(n16225) );
  NAND2X0 U16334 ( .IN1(n14900), .IN2(n8086), .QN(n16226) );
  NAND2X0 U16335 ( .IN1(n16227), .IN2(n16228), .QN(n16224) );
  NAND2X0 U16336 ( .IN1(n16229), .IN2(n8080), .QN(n16228) );
  INVX0 U16337 ( .INP(n16230), .ZN(n16229) );
  NOR2X0 U16338 ( .IN1(n16231), .IN2(n16232), .QN(n16227) );
  NOR2X0 U16339 ( .IN1(n4450), .IN2(n16233), .QN(n16232) );
  NOR2X0 U16340 ( .IN1(n14899), .IN2(DFF_156_n1), .QN(n16231) );
  NAND2X0 U16341 ( .IN1(n16234), .IN2(n16235), .QN(g26135) );
  NOR2X0 U16342 ( .IN1(n16236), .IN2(n16237), .QN(n16235) );
  NAND2X0 U16343 ( .IN1(n16238), .IN2(n16239), .QN(n16237) );
  NAND2X0 U16344 ( .IN1(test_so7), .IN2(n16240), .QN(n16239) );
  NOR2X0 U16345 ( .IN1(n16241), .IN2(n16242), .QN(n16238) );
  NOR2X0 U16346 ( .IN1(n14884), .IN2(n10329), .QN(n16242) );
  NOR2X0 U16347 ( .IN1(n16243), .IN2(g3128), .QN(n16241) );
  NAND2X0 U16348 ( .IN1(n16244), .IN2(n16245), .QN(n16236) );
  NOR2X0 U16349 ( .IN1(n16246), .IN2(n16247), .QN(n16245) );
  NOR2X0 U16350 ( .IN1(n14899), .IN2(DFF_155_n1), .QN(n16247) );
  NOR2X0 U16351 ( .IN1(n4443), .IN2(n16248), .QN(n16246) );
  NOR2X0 U16352 ( .IN1(n16249), .IN2(n16250), .QN(n16244) );
  NOR2X0 U16353 ( .IN1(n18869), .IN2(n16230), .QN(n16250) );
  NOR2X0 U16354 ( .IN1(n4452), .IN2(n16233), .QN(n16249) );
  NOR2X0 U16355 ( .IN1(n16251), .IN2(n16252), .QN(n16234) );
  NAND2X0 U16356 ( .IN1(n16253), .IN2(n3700), .QN(n16252) );
  NOR2X0 U16357 ( .IN1(n16254), .IN2(n16255), .QN(n16253) );
  NOR2X0 U16358 ( .IN1(n4447), .IN2(n16197), .QN(n16255) );
  NOR2X0 U16359 ( .IN1(n4343), .IN2(n16198), .QN(n16254) );
  NAND2X0 U16360 ( .IN1(n16256), .IN2(n16257), .QN(n16251) );
  NAND2X0 U16361 ( .IN1(n3936), .IN2(n16258), .QN(n16257) );
  NAND2X0 U16362 ( .IN1(n16259), .IN2(n16260), .QN(n16258) );
  NOR2X0 U16363 ( .IN1(n16261), .IN2(n16262), .QN(n16260) );
  NOR2X0 U16364 ( .IN1(n4342), .IN2(n16206), .QN(n16262) );
  NOR2X0 U16365 ( .IN1(n4334), .IN2(n16207), .QN(n16261) );
  NOR2X0 U16366 ( .IN1(n16263), .IN2(n16264), .QN(n16259) );
  NOR2X0 U16367 ( .IN1(n4438), .IN2(n16210), .QN(n16264) );
  NOR2X0 U16368 ( .IN1(n4434), .IN2(n16211), .QN(n16263) );
  NOR2X0 U16369 ( .IN1(n16265), .IN2(n16266), .QN(n16256) );
  NOR2X0 U16370 ( .IN1(n16267), .IN2(n16215), .QN(n16266) );
  NOR2X0 U16371 ( .IN1(n16268), .IN2(n16269), .QN(n16267) );
  NAND2X0 U16372 ( .IN1(n16270), .IN2(n16271), .QN(n16269) );
  NAND2X0 U16373 ( .IN1(n16220), .IN2(g3105), .QN(n16271) );
  NAND2X0 U16374 ( .IN1(n16221), .IN2(g3097), .QN(n16270) );
  NOR2X0 U16375 ( .IN1(n4437), .IN2(n16222), .QN(n16268) );
  NOR2X0 U16376 ( .IN1(n14892), .IN2(n14886), .QN(n16265) );
  INVX0 U16377 ( .INP(n16272), .ZN(n14892) );
  NAND2X0 U16378 ( .IN1(n16273), .IN2(n16274), .QN(g26104) );
  NOR2X0 U16379 ( .IN1(n16275), .IN2(n16276), .QN(n16274) );
  NAND2X0 U16380 ( .IN1(n16277), .IN2(n16278), .QN(n16276) );
  NAND2X0 U16381 ( .IN1(n16279), .IN2(g3091), .QN(n16278) );
  INVX0 U16382 ( .INP(n16197), .ZN(n16279) );
  NAND2X0 U16383 ( .IN1(n16280), .IN2(n3933), .QN(n16197) );
  NOR2X0 U16384 ( .IN1(g3201), .IN2(n14882), .QN(n16280) );
  NOR2X0 U16385 ( .IN1(n16281), .IN2(n16282), .QN(n16277) );
  NOR2X0 U16386 ( .IN1(n4344), .IN2(n16198), .QN(n16282) );
  NAND2X0 U16387 ( .IN1(n16283), .IN2(n4329), .QN(n16198) );
  NOR2X0 U16388 ( .IN1(n16284), .IN2(n16285), .QN(n16281) );
  INVX0 U16389 ( .INP(n3936), .ZN(n16285) );
  NOR2X0 U16390 ( .IN1(n16286), .IN2(n16287), .QN(n16284) );
  NAND2X0 U16391 ( .IN1(n16288), .IN2(n16289), .QN(n16287) );
  NAND2X0 U16392 ( .IN1(n16290), .IN2(g3211), .QN(n16289) );
  NAND2X0 U16393 ( .IN1(n14877), .IN2(g3094), .QN(n16288) );
  INVX0 U16394 ( .INP(n16291), .ZN(n16286) );
  NOR2X0 U16395 ( .IN1(n16292), .IN2(n16293), .QN(n16291) );
  NOR2X0 U16396 ( .IN1(n16207), .IN2(n4336), .QN(n16293) );
  NAND2X0 U16397 ( .IN1(g3207), .IN2(g3201), .QN(n16207) );
  NOR2X0 U16398 ( .IN1(n16206), .IN2(n4340), .QN(n16292) );
  NAND2X0 U16399 ( .IN1(n4406), .IN2(g3207), .QN(n16206) );
  NAND2X0 U16400 ( .IN1(n16294), .IN2(n16295), .QN(n16275) );
  NOR2X0 U16401 ( .IN1(n16296), .IN2(n16297), .QN(n16295) );
  NOR2X0 U16402 ( .IN1(n4337), .IN2(n16223), .QN(n16297) );
  INVX0 U16403 ( .INP(n16240), .ZN(n16223) );
  NOR2X0 U16404 ( .IN1(n14882), .IN2(n16298), .QN(n16240) );
  NOR2X0 U16405 ( .IN1(n4301), .IN2(n14884), .QN(n16296) );
  NAND2X0 U16406 ( .IN1(n16299), .IN2(n4073), .QN(n14884) );
  NOR2X0 U16407 ( .IN1(n10296), .IN2(n16222), .QN(n16299) );
  NOR2X0 U16408 ( .IN1(n16300), .IN2(n16301), .QN(n16294) );
  NOR2X0 U16409 ( .IN1(n16302), .IN2(n16215), .QN(n16301) );
  NOR2X0 U16410 ( .IN1(n16303), .IN2(n16304), .QN(n16302) );
  NAND2X0 U16411 ( .IN1(n16305), .IN2(n16306), .QN(n16304) );
  NAND2X0 U16412 ( .IN1(n16220), .IN2(g3093), .QN(n16306) );
  NAND2X0 U16413 ( .IN1(test_so6), .IN2(n16221), .QN(n16305) );
  NOR2X0 U16414 ( .IN1(n4439), .IN2(n16222), .QN(n16303) );
  NOR2X0 U16415 ( .IN1(n14891), .IN2(n14886), .QN(n16300) );
  NAND2X0 U16416 ( .IN1(n3705), .IN2(n16221), .QN(n14886) );
  INVX0 U16417 ( .INP(n16307), .ZN(n14891) );
  NOR2X0 U16418 ( .IN1(n16308), .IN2(n16309), .QN(n16273) );
  NAND2X0 U16419 ( .IN1(n16310), .IN2(n3700), .QN(n16309) );
  NOR2X0 U16420 ( .IN1(n16311), .IN2(n16312), .QN(n16310) );
  NOR2X0 U16421 ( .IN1(n16243), .IN2(DFF_140_n1), .QN(n16312) );
  NOR2X0 U16422 ( .IN1(n18868), .IN2(n16230), .QN(n16311) );
  NAND2X0 U16423 ( .IN1(n16313), .IN2(n16314), .QN(n16308) );
  NAND2X0 U16424 ( .IN1(n16315), .IN2(g3092), .QN(n16314) );
  INVX0 U16425 ( .INP(n16233), .ZN(n16315) );
  NAND2X0 U16426 ( .IN1(n16283), .IN2(g3207), .QN(n16233) );
  NOR2X0 U16427 ( .IN1(n16316), .IN2(n14882), .QN(n16283) );
  INVX0 U16428 ( .INP(n16317), .ZN(n14882) );
  NOR2X0 U16429 ( .IN1(n11728), .IN2(n10296), .QN(n16317) );
  NAND2X0 U16430 ( .IN1(n307), .IN2(g3197), .QN(n11728) );
  INVX0 U16431 ( .INP(n16318), .ZN(n307) );
  NAND2X0 U16432 ( .IN1(n16319), .IN2(n18863), .QN(n16318) );
  NOR2X0 U16433 ( .IN1(n8088), .IN2(n8090), .QN(n16319) );
  NAND2X0 U16434 ( .IN1(g3188), .IN2(n4406), .QN(n16316) );
  NOR2X0 U16435 ( .IN1(n16320), .IN2(n16321), .QN(n16313) );
  NOR2X0 U16436 ( .IN1(n18871), .IN2(n14899), .QN(n16321) );
  NAND2X0 U16437 ( .IN1(n16322), .IN2(n4073), .QN(n14899) );
  NOR2X0 U16438 ( .IN1(n10296), .IN2(n14893), .QN(n16322) );
  INVX0 U16439 ( .INP(n16220), .ZN(n14893) );
  NOR2X0 U16440 ( .IN1(n16210), .IN2(g3188), .QN(n16220) );
  INVX0 U16441 ( .INP(n14877), .ZN(n16210) );
  NOR2X0 U16442 ( .IN1(g3207), .IN2(n4406), .QN(n14877) );
  NOR2X0 U16443 ( .IN1(n4445), .IN2(n16248), .QN(n16320) );
  INVX0 U16444 ( .INP(n16194), .ZN(n16248) );
  NOR2X0 U16445 ( .IN1(n16323), .IN2(n16215), .QN(n16194) );
  INVX0 U16446 ( .INP(n3939), .ZN(n16215) );
  NAND2X0 U16447 ( .IN1(n4406), .IN2(n3933), .QN(n16323) );
  NOR2X0 U16448 ( .IN1(g3188), .IN2(n4329), .QN(n3933) );
  NAND2X0 U16449 ( .IN1(n11062), .IN2(n16324), .QN(g26048) );
  NAND2X0 U16450 ( .IN1(n16325), .IN2(n16326), .QN(n16324) );
  NOR2X0 U16451 ( .IN1(n16327), .IN2(n16328), .QN(n16325) );
  NOR2X0 U16452 ( .IN1(n18873), .IN2(n16329), .QN(n16328) );
  INVX0 U16453 ( .INP(n16330), .ZN(n16329) );
  NOR2X0 U16454 ( .IN1(n16330), .IN2(n7909), .QN(n16327) );
  NOR2X0 U16455 ( .IN1(n10998), .IN2(n16331), .QN(g26037) );
  NAND2X0 U16456 ( .IN1(n16332), .IN2(n15729), .QN(n16331) );
  INVX0 U16457 ( .INP(n15730), .ZN(n15729) );
  NOR2X0 U16458 ( .IN1(n16333), .IN2(n4291), .QN(n15730) );
  NAND2X0 U16459 ( .IN1(n4291), .IN2(n16333), .QN(n16332) );
  NOR2X0 U16460 ( .IN1(n16334), .IN2(n15740), .QN(g26031) );
  NOR2X0 U16461 ( .IN1(n16335), .IN2(n16336), .QN(n16334) );
  NOR2X0 U16462 ( .IN1(test_so98), .IN2(n3742), .QN(n16336) );
  NOR2X0 U16463 ( .IN1(n16337), .IN2(n10327), .QN(n16335) );
  INVX0 U16464 ( .INP(n3742), .ZN(n16337) );
  NAND2X0 U16465 ( .IN1(n16338), .IN2(n16339), .QN(g26025) );
  NAND2X0 U16466 ( .IN1(test_so82), .IN2(n16340), .QN(n16339) );
  NAND2X0 U16467 ( .IN1(n15760), .IN2(n13307), .QN(n16340) );
  NAND2X0 U16468 ( .IN1(n15761), .IN2(n13307), .QN(n16338) );
  INVX0 U16469 ( .INP(n4509), .ZN(n13307) );
  NOR2X0 U16470 ( .IN1(n10322), .IN2(n15760), .QN(n15761) );
  INVX0 U16471 ( .INP(n3749), .ZN(n15760) );
  NAND2X0 U16472 ( .IN1(n16341), .IN2(test_so79), .QN(n3749) );
  NOR2X0 U16473 ( .IN1(n13423), .IN2(n13214), .QN(n16341) );
  NAND2X0 U16474 ( .IN1(n16342), .IN2(n16343), .QN(n13214) );
  NAND2X0 U16475 ( .IN1(n9977), .IN2(n11937), .QN(n16343) );
  NOR2X0 U16476 ( .IN1(n16344), .IN2(n16345), .QN(n16342) );
  NOR2X0 U16477 ( .IN1(n4516), .IN2(g2478), .QN(n16345) );
  NOR2X0 U16478 ( .IN1(test_so82), .IN2(n4509), .QN(n16344) );
  NAND2X0 U16479 ( .IN1(n16346), .IN2(n16347), .QN(n13423) );
  NOR2X0 U16480 ( .IN1(n16348), .IN2(n16349), .QN(n16347) );
  NAND2X0 U16481 ( .IN1(n16350), .IN2(n16351), .QN(n16349) );
  NOR2X0 U16482 ( .IN1(n16352), .IN2(n16353), .QN(n16351) );
  NOR2X0 U16483 ( .IN1(n13519), .IN2(n16354), .QN(n16353) );
  INVX0 U16484 ( .INP(n16355), .ZN(n16352) );
  NAND2X0 U16485 ( .IN1(n16354), .IN2(n13519), .QN(n16355) );
  NAND2X0 U16486 ( .IN1(n16356), .IN2(n16357), .QN(n16354) );
  NAND2X0 U16487 ( .IN1(n9826), .IN2(test_so73), .QN(n16357) );
  NOR2X0 U16488 ( .IN1(n16358), .IN2(n16359), .QN(n16356) );
  NOR2X0 U16489 ( .IN1(n4367), .IN2(g2235), .QN(n16359) );
  NOR2X0 U16490 ( .IN1(n4324), .IN2(g2236), .QN(n16358) );
  NOR2X0 U16491 ( .IN1(n16360), .IN2(n16361), .QN(n16350) );
  NAND2X0 U16492 ( .IN1(n16362), .IN2(n16363), .QN(n16361) );
  INVX0 U16493 ( .INP(n16364), .ZN(n16363) );
  NOR2X0 U16494 ( .IN1(n13485), .IN2(n16365), .QN(n16364) );
  NAND2X0 U16495 ( .IN1(n16365), .IN2(n13485), .QN(n16362) );
  NOR2X0 U16496 ( .IN1(n16366), .IN2(n16367), .QN(n16365) );
  NOR2X0 U16497 ( .IN1(n10320), .IN2(test_so75), .QN(n16367) );
  INVX0 U16498 ( .INP(n16368), .ZN(n16366) );
  NOR2X0 U16499 ( .IN1(n16369), .IN2(n16370), .QN(n16368) );
  NOR2X0 U16500 ( .IN1(n4367), .IN2(g2238), .QN(n16370) );
  NOR2X0 U16501 ( .IN1(n4324), .IN2(g2239), .QN(n16369) );
  NAND2X0 U16502 ( .IN1(n16371), .IN2(n16372), .QN(n16360) );
  NAND2X0 U16503 ( .IN1(n4319), .IN2(n16373), .QN(n16372) );
  INVX0 U16504 ( .INP(n16374), .ZN(n16371) );
  NOR2X0 U16505 ( .IN1(n16373), .IN2(n4319), .QN(n16374) );
  NAND2X0 U16506 ( .IN1(n16375), .IN2(n16376), .QN(n16373) );
  NAND2X0 U16507 ( .IN1(n9841), .IN2(g2241), .QN(n16376) );
  NOR2X0 U16508 ( .IN1(n16377), .IN2(n16378), .QN(n16375) );
  NOR2X0 U16509 ( .IN1(n4324), .IN2(g2218), .QN(n16378) );
  NOR2X0 U16510 ( .IN1(n10320), .IN2(g2219), .QN(n16377) );
  NAND2X0 U16511 ( .IN1(n16379), .IN2(n16380), .QN(n16348) );
  NOR2X0 U16512 ( .IN1(n16381), .IN2(n16382), .QN(n16380) );
  NOR2X0 U16513 ( .IN1(n4373), .IN2(n16383), .QN(n16382) );
  INVX0 U16514 ( .INP(n16384), .ZN(n16381) );
  NAND2X0 U16515 ( .IN1(n16383), .IN2(n4373), .QN(n16384) );
  NAND2X0 U16516 ( .IN1(n16385), .IN2(n16386), .QN(n16383) );
  NAND2X0 U16517 ( .IN1(n9842), .IN2(g2241), .QN(n16386) );
  NOR2X0 U16518 ( .IN1(n16387), .IN2(n16388), .QN(n16385) );
  NOR2X0 U16519 ( .IN1(n4324), .IN2(g2209), .QN(n16388) );
  NOR2X0 U16520 ( .IN1(n10320), .IN2(g2210), .QN(n16387) );
  NOR2X0 U16521 ( .IN1(n12566), .IN2(n16389), .QN(n16379) );
  NAND2X0 U16522 ( .IN1(n16390), .IN2(n16391), .QN(n16389) );
  NAND2X0 U16523 ( .IN1(n4377), .IN2(n16392), .QN(n16391) );
  INVX0 U16524 ( .INP(n16393), .ZN(n16390) );
  NOR2X0 U16525 ( .IN1(n16392), .IN2(n4377), .QN(n16393) );
  NAND2X0 U16526 ( .IN1(n16394), .IN2(n16395), .QN(n16392) );
  NAND2X0 U16527 ( .IN1(n9843), .IN2(g2241), .QN(n16395) );
  NOR2X0 U16528 ( .IN1(n16396), .IN2(n16397), .QN(n16394) );
  NOR2X0 U16529 ( .IN1(n4324), .IN2(g2206), .QN(n16397) );
  NOR2X0 U16530 ( .IN1(n10320), .IN2(g2207), .QN(n16396) );
  INVX0 U16531 ( .INP(n3038), .ZN(n12566) );
  NOR2X0 U16532 ( .IN1(n16398), .IN2(n16399), .QN(n16346) );
  NAND2X0 U16533 ( .IN1(n16400), .IN2(n16401), .QN(n16399) );
  NOR2X0 U16534 ( .IN1(n16402), .IN2(n16403), .QN(n16401) );
  NOR2X0 U16535 ( .IN1(n4563), .IN2(n16404), .QN(n16403) );
  INVX0 U16536 ( .INP(n16405), .ZN(n16402) );
  NAND2X0 U16537 ( .IN1(n16404), .IN2(n4563), .QN(n16405) );
  NAND2X0 U16538 ( .IN1(n16406), .IN2(n16407), .QN(n16404) );
  NAND2X0 U16539 ( .IN1(n9837), .IN2(g2241), .QN(n16407) );
  NOR2X0 U16540 ( .IN1(n16408), .IN2(n16409), .QN(n16406) );
  NOR2X0 U16541 ( .IN1(n4324), .IN2(g2230), .QN(n16409) );
  NOR2X0 U16542 ( .IN1(n10320), .IN2(g2231), .QN(n16408) );
  NOR2X0 U16543 ( .IN1(n16410), .IN2(n16411), .QN(n16400) );
  NOR2X0 U16544 ( .IN1(n4389), .IN2(n16412), .QN(n16411) );
  INVX0 U16545 ( .INP(n16413), .ZN(n16410) );
  NAND2X0 U16546 ( .IN1(n16412), .IN2(n4389), .QN(n16413) );
  NAND2X0 U16547 ( .IN1(n16414), .IN2(n16415), .QN(n16412) );
  NAND2X0 U16548 ( .IN1(n9840), .IN2(g2241), .QN(n16415) );
  NOR2X0 U16549 ( .IN1(n16416), .IN2(n16417), .QN(n16414) );
  NOR2X0 U16550 ( .IN1(n4324), .IN2(g2221), .QN(n16417) );
  NOR2X0 U16551 ( .IN1(n10320), .IN2(g2222), .QN(n16416) );
  NAND2X0 U16552 ( .IN1(n16418), .IN2(n16419), .QN(n16398) );
  NOR2X0 U16553 ( .IN1(n16420), .IN2(n16421), .QN(n16419) );
  INVX0 U16554 ( .INP(n16422), .ZN(n16421) );
  NAND2X0 U16555 ( .IN1(g2185), .IN2(n16423), .QN(n16422) );
  NOR2X0 U16556 ( .IN1(n16423), .IN2(g2185), .QN(n16420) );
  NOR2X0 U16557 ( .IN1(n16424), .IN2(n16425), .QN(n16423) );
  NOR2X0 U16558 ( .IN1(n10320), .IN2(test_so74), .QN(n16425) );
  INVX0 U16559 ( .INP(n16426), .ZN(n16424) );
  NOR2X0 U16560 ( .IN1(n16427), .IN2(n16428), .QN(n16426) );
  NOR2X0 U16561 ( .IN1(n4367), .IN2(g2223), .QN(n16428) );
  NOR2X0 U16562 ( .IN1(n4324), .IN2(g2224), .QN(n16427) );
  NOR2X0 U16563 ( .IN1(n16429), .IN2(n16430), .QN(n16418) );
  NAND2X0 U16564 ( .IN1(n16431), .IN2(n16432), .QN(n16430) );
  NAND2X0 U16565 ( .IN1(n4287), .IN2(n16433), .QN(n16432) );
  INVX0 U16566 ( .INP(n16434), .ZN(n16431) );
  NOR2X0 U16567 ( .IN1(n16433), .IN2(n4287), .QN(n16434) );
  NAND2X0 U16568 ( .IN1(n16435), .IN2(n16436), .QN(n16433) );
  NAND2X0 U16569 ( .IN1(n9836), .IN2(g2241), .QN(n16436) );
  NOR2X0 U16570 ( .IN1(n16437), .IN2(n16438), .QN(n16435) );
  NOR2X0 U16571 ( .IN1(n4324), .IN2(g2233), .QN(n16438) );
  NOR2X0 U16572 ( .IN1(n10320), .IN2(g2234), .QN(n16437) );
  NAND2X0 U16573 ( .IN1(n16439), .IN2(n16440), .QN(n16429) );
  NAND2X0 U16574 ( .IN1(n4555), .IN2(n16441), .QN(n16440) );
  INVX0 U16575 ( .INP(n16442), .ZN(n16439) );
  NOR2X0 U16576 ( .IN1(n16441), .IN2(n4555), .QN(n16442) );
  NAND2X0 U16577 ( .IN1(n16443), .IN2(n16444), .QN(n16441) );
  NAND2X0 U16578 ( .IN1(n9838), .IN2(g2241), .QN(n16444) );
  NOR2X0 U16579 ( .IN1(n16445), .IN2(n16446), .QN(n16443) );
  NOR2X0 U16580 ( .IN1(n4324), .IN2(g2227), .QN(n16446) );
  NOR2X0 U16581 ( .IN1(n10320), .IN2(g2228), .QN(n16445) );
  NOR2X0 U16582 ( .IN1(n16174), .IN2(n16447), .QN(g25940) );
  NAND2X0 U16583 ( .IN1(n16448), .IN2(n13952), .QN(n16447) );
  INVX0 U16584 ( .INP(n13263), .ZN(n13952) );
  INVX0 U16585 ( .INP(n16449), .ZN(n16448) );
  NOR2X0 U16586 ( .IN1(test_so78), .IN2(n3887), .QN(n16449) );
  INVX0 U16587 ( .INP(n4526), .ZN(n16174) );
  NOR2X0 U16588 ( .IN1(n16178), .IN2(n16450), .QN(g25938) );
  NAND2X0 U16589 ( .IN1(n16451), .IN2(n13954), .QN(n16450) );
  INVX0 U16590 ( .INP(n13268), .ZN(n13954) );
  INVX0 U16591 ( .INP(n16452), .ZN(n16451) );
  NOR2X0 U16592 ( .IN1(g1462), .IN2(n3890), .QN(n16452) );
  INVX0 U16593 ( .INP(n4527), .ZN(n16178) );
  NOR2X0 U16594 ( .IN1(n16453), .IN2(n16182), .QN(g25935) );
  NAND2X0 U16595 ( .IN1(n3690), .IN2(n13956), .QN(n16182) );
  NAND2X0 U16596 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NOR2X0 U16597 ( .IN1(n3893), .IN2(g776), .QN(n16453) );
  NOR2X0 U16598 ( .IN1(n16187), .IN2(n16454), .QN(g25932) );
  NAND2X0 U16599 ( .IN1(n16455), .IN2(n13958), .QN(n16454) );
  INVX0 U16600 ( .INP(n13278), .ZN(n13958) );
  INVX0 U16601 ( .INP(n16456), .ZN(n16455) );
  NOR2X0 U16602 ( .IN1(g88), .IN2(n3896), .QN(n16456) );
  INVX0 U16603 ( .INP(n4528), .ZN(n16187) );
  NAND2X0 U16604 ( .IN1(n16457), .IN2(n16458), .QN(g25489) );
  NAND2X0 U16605 ( .IN1(n16459), .IN2(n16460), .QN(n16458) );
  NOR2X0 U16606 ( .IN1(n4433), .IN2(n4424), .QN(n16460) );
  NOR2X0 U16607 ( .IN1(n4301), .IN2(n16461), .QN(n16459) );
  NAND2X0 U16608 ( .IN1(n16462), .IN2(n10329), .QN(n16457) );
  NAND2X0 U16609 ( .IN1(n16461), .IN2(n16463), .QN(n16462) );
  NAND2X0 U16610 ( .IN1(n4301), .IN2(n16307), .QN(n16463) );
  NAND2X0 U16611 ( .IN1(DFF_15_n1), .IN2(DFF_16_n1), .QN(n16307) );
  NOR2X0 U16612 ( .IN1(test_so10), .IN2(n16464), .QN(n16461) );
  INVX0 U16613 ( .INP(n16465), .ZN(n16464) );
  NAND2X0 U16614 ( .IN1(n4424), .IN2(n16466), .QN(n16465) );
  INVX0 U16615 ( .INP(n16467), .ZN(n16466) );
  NOR2X0 U16616 ( .IN1(n16272), .IN2(n4301), .QN(n16467) );
  NAND2X0 U16617 ( .IN1(n9739), .IN2(n9738), .QN(n16272) );
  NAND2X0 U16618 ( .IN1(n16468), .IN2(n16469), .QN(g25452) );
  INVX0 U16619 ( .INP(n16470), .ZN(n16469) );
  NOR2X0 U16620 ( .IN1(g3109), .IN2(n4443), .QN(n16470) );
  NAND2X0 U16621 ( .IN1(g21851), .IN2(g3109), .QN(n16468) );
  NAND2X0 U16622 ( .IN1(n16471), .IN2(n16472), .QN(g25451) );
  INVX0 U16623 ( .INP(n16473), .ZN(n16472) );
  NOR2X0 U16624 ( .IN1(g8030), .IN2(n4434), .QN(n16473) );
  NAND2X0 U16625 ( .IN1(g21851), .IN2(g8030), .QN(n16471) );
  NAND2X0 U16626 ( .IN1(n16474), .IN2(n16475), .QN(g25450) );
  NAND2X0 U16627 ( .IN1(n4382), .IN2(g3097), .QN(n16475) );
  NAND2X0 U16628 ( .IN1(g21851), .IN2(g8106), .QN(n16474) );
  NAND2X0 U16629 ( .IN1(n16476), .IN2(n3700), .QN(g25442) );
  NOR2X0 U16630 ( .IN1(n16477), .IN2(n16478), .QN(n16476) );
  NOR2X0 U16631 ( .IN1(n9638), .IN2(n16243), .QN(n16478) );
  NOR2X0 U16632 ( .IN1(n9639), .IN2(n16230), .QN(n16477) );
  NAND2X0 U16633 ( .IN1(n16479), .IN2(n3700), .QN(g25435) );
  NOR2X0 U16634 ( .IN1(n16480), .IN2(n16481), .QN(n16479) );
  NOR2X0 U16635 ( .IN1(n16243), .IN2(n8084), .QN(n16481) );
  NOR2X0 U16636 ( .IN1(n9604), .IN2(n16230), .QN(n16480) );
  NAND2X0 U16637 ( .IN1(n16482), .IN2(n3700), .QN(g25420) );
  NOR2X0 U16638 ( .IN1(n16483), .IN2(n16484), .QN(n16482) );
  NOR2X0 U16639 ( .IN1(n16243), .IN2(n9636), .QN(n16484) );
  INVX0 U16640 ( .INP(n14900), .ZN(n16243) );
  NOR2X0 U16641 ( .IN1(n9637), .IN2(n16230), .QN(n16483) );
  NAND2X0 U16642 ( .IN1(n16485), .IN2(n4073), .QN(n16230) );
  NOR2X0 U16643 ( .IN1(n10296), .IN2(n16298), .QN(n16485) );
  INVX0 U16644 ( .INP(n16221), .ZN(n16298) );
  NOR2X0 U16645 ( .IN1(g3188), .IN2(n16211), .QN(n16221) );
  INVX0 U16646 ( .INP(n16290), .ZN(n16211) );
  NOR2X0 U16647 ( .IN1(g3201), .IN2(g3207), .QN(n16290) );
  NAND2X0 U16648 ( .IN1(n16486), .IN2(n16487), .QN(g25288) );
  NAND2X0 U16649 ( .IN1(n16488), .IN2(g2808), .QN(n16487) );
  NAND2X0 U16650 ( .IN1(n16489), .IN2(n16490), .QN(n16486) );
  NAND2X0 U16651 ( .IN1(n16491), .IN2(n16492), .QN(g25280) );
  NAND2X0 U16652 ( .IN1(n16493), .IN2(g2810), .QN(n16492) );
  NAND2X0 U16653 ( .IN1(n16494), .IN2(n16489), .QN(n16491) );
  NAND2X0 U16654 ( .IN1(n16495), .IN2(n16496), .QN(g25279) );
  NAND2X0 U16655 ( .IN1(n16497), .IN2(g2114), .QN(n16496) );
  NAND2X0 U16656 ( .IN1(n16498), .IN2(n16499), .QN(n16495) );
  NAND2X0 U16657 ( .IN1(n16500), .IN2(n16501), .QN(g25272) );
  NAND2X0 U16658 ( .IN1(n16502), .IN2(g2809), .QN(n16501) );
  NAND2X0 U16659 ( .IN1(n16503), .IN2(n16489), .QN(n16500) );
  INVX0 U16660 ( .INP(n16504), .ZN(n16489) );
  NAND2X0 U16661 ( .IN1(n16505), .IN2(n16506), .QN(n16504) );
  NOR2X0 U16662 ( .IN1(n16507), .IN2(n16508), .QN(n16506) );
  NAND2X0 U16663 ( .IN1(n16509), .IN2(n16510), .QN(n16508) );
  NAND2X0 U16664 ( .IN1(n16511), .IN2(n16512), .QN(n16510) );
  NOR2X0 U16665 ( .IN1(n16513), .IN2(n16514), .QN(n16512) );
  NAND2X0 U16666 ( .IN1(n16515), .IN2(n16516), .QN(n16514) );
  NOR2X0 U16667 ( .IN1(n16517), .IN2(n16518), .QN(n16516) );
  NOR2X0 U16668 ( .IN1(n4408), .IN2(n11338), .QN(n16518) );
  NOR2X0 U16669 ( .IN1(n11337), .IN2(g2720), .QN(n16517) );
  INVX0 U16670 ( .INP(n11338), .ZN(n11337) );
  NAND2X0 U16671 ( .IN1(n16519), .IN2(n16520), .QN(n11338) );
  NAND2X0 U16672 ( .IN1(g2703), .IN2(n10334), .QN(n16520) );
  NOR2X0 U16673 ( .IN1(n16521), .IN2(n16522), .QN(n16519) );
  NOR2X0 U16674 ( .IN1(n4306), .IN2(g2782), .QN(n16522) );
  NOR2X0 U16675 ( .IN1(n4356), .IN2(g2783), .QN(n16521) );
  NOR2X0 U16676 ( .IN1(n16523), .IN2(n16524), .QN(n16515) );
  NOR2X0 U16677 ( .IN1(n4407), .IN2(n11345), .QN(n16524) );
  NOR2X0 U16678 ( .IN1(n11343), .IN2(g2746), .QN(n16523) );
  INVX0 U16679 ( .INP(n11345), .ZN(n11343) );
  NAND2X0 U16680 ( .IN1(n16525), .IN2(n16526), .QN(n11345) );
  NAND2X0 U16681 ( .IN1(n10158), .IN2(g2703), .QN(n16526) );
  NOR2X0 U16682 ( .IN1(n16527), .IN2(n16528), .QN(n16525) );
  NOR2X0 U16683 ( .IN1(n4306), .IN2(g2788), .QN(n16528) );
  NOR2X0 U16684 ( .IN1(n4356), .IN2(g2789), .QN(n16527) );
  NAND2X0 U16685 ( .IN1(n16529), .IN2(n16530), .QN(n16513) );
  NOR2X0 U16686 ( .IN1(n16531), .IN2(n16532), .QN(n16530) );
  NOR2X0 U16687 ( .IN1(n4415), .IN2(n11276), .QN(n16532) );
  NOR2X0 U16688 ( .IN1(n11273), .IN2(g2766), .QN(n16531) );
  INVX0 U16689 ( .INP(n11276), .ZN(n11273) );
  NAND2X0 U16690 ( .IN1(n16533), .IN2(n16534), .QN(n11276) );
  NAND2X0 U16691 ( .IN1(n10155), .IN2(g2703), .QN(n16534) );
  NOR2X0 U16692 ( .IN1(n16535), .IN2(n16536), .QN(n16533) );
  NOR2X0 U16693 ( .IN1(n4306), .IN2(g2800), .QN(n16536) );
  NOR2X0 U16694 ( .IN1(n4356), .IN2(g2801), .QN(n16535) );
  NOR2X0 U16695 ( .IN1(n16537), .IN2(n16538), .QN(n16529) );
  NAND2X0 U16696 ( .IN1(n16539), .IN2(n16540), .QN(n16538) );
  NAND2X0 U16697 ( .IN1(n4393), .IN2(n11268), .QN(n16540) );
  NAND2X0 U16698 ( .IN1(n11265), .IN2(g2760), .QN(n16539) );
  INVX0 U16699 ( .INP(n11268), .ZN(n11265) );
  NAND2X0 U16700 ( .IN1(n16541), .IN2(n16542), .QN(n11268) );
  NAND2X0 U16701 ( .IN1(g2703), .IN2(n10335), .QN(n16542) );
  NOR2X0 U16702 ( .IN1(n16543), .IN2(n16544), .QN(n16541) );
  NOR2X0 U16703 ( .IN1(n4306), .IN2(g2797), .QN(n16544) );
  NOR2X0 U16704 ( .IN1(n4356), .IN2(g2798), .QN(n16543) );
  NOR2X0 U16705 ( .IN1(n16545), .IN2(n16546), .QN(n16537) );
  NOR2X0 U16706 ( .IN1(test_so92), .IN2(n11295), .QN(n16546) );
  NOR2X0 U16707 ( .IN1(n11294), .IN2(n10324), .QN(n16545) );
  INVX0 U16708 ( .INP(n11295), .ZN(n11294) );
  NAND2X0 U16709 ( .IN1(n16547), .IN2(n16548), .QN(n11295) );
  NAND2X0 U16710 ( .IN1(n10157), .IN2(g2703), .QN(n16548) );
  NOR2X0 U16711 ( .IN1(n16549), .IN2(n16550), .QN(n16547) );
  NOR2X0 U16712 ( .IN1(n4306), .IN2(g2791), .QN(n16550) );
  NOR2X0 U16713 ( .IN1(n4356), .IN2(g2792), .QN(n16549) );
  NOR2X0 U16714 ( .IN1(n16551), .IN2(n16552), .QN(n16511) );
  NAND2X0 U16715 ( .IN1(n16553), .IN2(n16554), .QN(n16552) );
  NOR2X0 U16716 ( .IN1(n16555), .IN2(n16556), .QN(n16554) );
  NOR2X0 U16717 ( .IN1(n4419), .IN2(n11358), .QN(n16556) );
  NOR2X0 U16718 ( .IN1(n11357), .IN2(g2727), .QN(n16555) );
  INVX0 U16719 ( .INP(n11358), .ZN(n11357) );
  NAND2X0 U16720 ( .IN1(n16557), .IN2(n16558), .QN(n11358) );
  NAND2X0 U16721 ( .IN1(n10160), .IN2(g2703), .QN(n16558) );
  NOR2X0 U16722 ( .IN1(n16559), .IN2(n16560), .QN(n16557) );
  NOR2X0 U16723 ( .IN1(n4306), .IN2(g2779), .QN(n16560) );
  NOR2X0 U16724 ( .IN1(n4356), .IN2(g2780), .QN(n16559) );
  NOR2X0 U16725 ( .IN1(n16561), .IN2(n16562), .QN(n16553) );
  NOR2X0 U16726 ( .IN1(n4472), .IN2(n11325), .QN(n16562) );
  NOR2X0 U16727 ( .IN1(n11324), .IN2(g2707), .QN(n16561) );
  INVX0 U16728 ( .INP(n11325), .ZN(n11324) );
  NAND2X0 U16729 ( .IN1(n16563), .IN2(n16564), .QN(n11325) );
  NAND2X0 U16730 ( .IN1(n10161), .IN2(g2703), .QN(n16564) );
  NOR2X0 U16731 ( .IN1(n16565), .IN2(n16566), .QN(n16563) );
  NOR2X0 U16732 ( .IN1(n4306), .IN2(g2776), .QN(n16566) );
  NOR2X0 U16733 ( .IN1(n4356), .IN2(g2777), .QN(n16565) );
  NAND2X0 U16734 ( .IN1(n16567), .IN2(n16568), .QN(n16551) );
  NOR2X0 U16735 ( .IN1(n16569), .IN2(n16570), .QN(n16568) );
  NOR2X0 U16736 ( .IN1(n4471), .IN2(n11332), .QN(n16570) );
  NOR2X0 U16737 ( .IN1(n11331), .IN2(g2753), .QN(n16569) );
  INVX0 U16738 ( .INP(n11332), .ZN(n11331) );
  NAND2X0 U16739 ( .IN1(n16571), .IN2(n16572), .QN(n11332) );
  NAND2X0 U16740 ( .IN1(n10156), .IN2(g2703), .QN(n16572) );
  NOR2X0 U16741 ( .IN1(n16573), .IN2(n16574), .QN(n16571) );
  NOR2X0 U16742 ( .IN1(n4306), .IN2(g2794), .QN(n16574) );
  NOR2X0 U16743 ( .IN1(n4356), .IN2(g2795), .QN(n16573) );
  NOR2X0 U16744 ( .IN1(n16575), .IN2(n16576), .QN(n16567) );
  NAND2X0 U16745 ( .IN1(n16577), .IN2(n16578), .QN(n16576) );
  NAND2X0 U16746 ( .IN1(n4398), .IN2(n11320), .QN(n16578) );
  NAND2X0 U16747 ( .IN1(n11319), .IN2(g2714), .QN(n16577) );
  INVX0 U16748 ( .INP(n11320), .ZN(n11319) );
  NAND2X0 U16749 ( .IN1(n16579), .IN2(n16580), .QN(n11320) );
  NAND2X0 U16750 ( .IN1(n10162), .IN2(g2703), .QN(n16580) );
  NOR2X0 U16751 ( .IN1(n16581), .IN2(n16582), .QN(n16579) );
  NOR2X0 U16752 ( .IN1(n4306), .IN2(g2773), .QN(n16582) );
  NOR2X0 U16753 ( .IN1(n4356), .IN2(g2774), .QN(n16581) );
  NAND2X0 U16754 ( .IN1(n16583), .IN2(n16584), .QN(n16575) );
  NAND2X0 U16755 ( .IN1(n4397), .IN2(n11363), .QN(n16584) );
  NAND2X0 U16756 ( .IN1(n11362), .IN2(g2734), .QN(n16583) );
  INVX0 U16757 ( .INP(n11363), .ZN(n11362) );
  NAND2X0 U16758 ( .IN1(n16585), .IN2(n16586), .QN(n11363) );
  NAND2X0 U16759 ( .IN1(n10159), .IN2(g2703), .QN(n16586) );
  NOR2X0 U16760 ( .IN1(n16587), .IN2(n16588), .QN(n16585) );
  NOR2X0 U16761 ( .IN1(n4306), .IN2(g2785), .QN(n16588) );
  NOR2X0 U16762 ( .IN1(n4356), .IN2(g2786), .QN(n16587) );
  NAND2X0 U16763 ( .IN1(n10300), .IN2(g7425), .QN(n16509) );
  NOR2X0 U16764 ( .IN1(n4292), .IN2(g2802), .QN(n16507) );
  NOR2X0 U16765 ( .IN1(n16589), .IN2(n11854), .QN(n16505) );
  NAND2X0 U16766 ( .IN1(n16590), .IN2(n16591), .QN(n11854) );
  NAND2X0 U16767 ( .IN1(n9878), .IN2(g7487), .QN(n16591) );
  NOR2X0 U16768 ( .IN1(n16592), .IN2(n16593), .QN(n16590) );
  NOR2X0 U16769 ( .IN1(n4306), .IN2(g2806), .QN(n16593) );
  NOR2X0 U16770 ( .IN1(n4292), .IN2(g2805), .QN(n16592) );
  NOR2X0 U16771 ( .IN1(n4356), .IN2(g2804), .QN(n16589) );
  NAND2X0 U16772 ( .IN1(n16594), .IN2(n16595), .QN(g25271) );
  NAND2X0 U16773 ( .IN1(n16596), .IN2(n16498), .QN(n16595) );
  NAND2X0 U16774 ( .IN1(n16597), .IN2(g2116), .QN(n16594) );
  NAND2X0 U16775 ( .IN1(n16598), .IN2(n16599), .QN(g25270) );
  NAND2X0 U16776 ( .IN1(n16600), .IN2(g1420), .QN(n16599) );
  NAND2X0 U16777 ( .IN1(n16601), .IN2(n16602), .QN(n16598) );
  NAND2X0 U16778 ( .IN1(n16603), .IN2(n16604), .QN(g25268) );
  NAND2X0 U16779 ( .IN1(n16605), .IN2(n16498), .QN(n16604) );
  INVX0 U16780 ( .INP(n16606), .ZN(n16498) );
  NAND2X0 U16781 ( .IN1(n16607), .IN2(n16608), .QN(n16606) );
  NOR2X0 U16782 ( .IN1(n16609), .IN2(n16610), .QN(n16608) );
  NAND2X0 U16783 ( .IN1(n16611), .IN2(n16612), .QN(n16610) );
  NAND2X0 U16784 ( .IN1(n16613), .IN2(n16614), .QN(n16612) );
  NOR2X0 U16785 ( .IN1(n16615), .IN2(n16616), .QN(n16614) );
  NAND2X0 U16786 ( .IN1(n16617), .IN2(n16618), .QN(n16616) );
  NOR2X0 U16787 ( .IN1(n16619), .IN2(n16620), .QN(n16618) );
  NOR2X0 U16788 ( .IN1(n4400), .IN2(n11491), .QN(n16620) );
  NOR2X0 U16789 ( .IN1(n11490), .IN2(g2020), .QN(n16619) );
  INVX0 U16790 ( .INP(n11491), .ZN(n11490) );
  NAND2X0 U16791 ( .IN1(n16621), .IN2(n16622), .QN(n11491) );
  NAND2X0 U16792 ( .IN1(n10172), .IN2(g2009), .QN(n16622) );
  NOR2X0 U16793 ( .IN1(n16623), .IN2(n16624), .QN(n16621) );
  NOR2X0 U16794 ( .IN1(n4307), .IN2(g2079), .QN(n16624) );
  NOR2X0 U16795 ( .IN1(n4357), .IN2(g2080), .QN(n16623) );
  NOR2X0 U16796 ( .IN1(n16625), .IN2(n16626), .QN(n16617) );
  NOR2X0 U16797 ( .IN1(n4410), .IN2(n11512), .QN(n16626) );
  NOR2X0 U16798 ( .IN1(n11511), .IN2(g2026), .QN(n16625) );
  INVX0 U16799 ( .INP(n11512), .ZN(n11511) );
  NAND2X0 U16800 ( .IN1(n16627), .IN2(n16628), .QN(n11512) );
  NAND2X0 U16801 ( .IN1(n10169), .IN2(g2009), .QN(n16628) );
  NOR2X0 U16802 ( .IN1(n16629), .IN2(n16630), .QN(n16627) );
  NOR2X0 U16803 ( .IN1(n4307), .IN2(g2088), .QN(n16630) );
  NOR2X0 U16804 ( .IN1(n4357), .IN2(g2089), .QN(n16629) );
  NAND2X0 U16805 ( .IN1(n16631), .IN2(n16632), .QN(n16615) );
  NOR2X0 U16806 ( .IN1(n16633), .IN2(n16634), .QN(n16632) );
  NOR2X0 U16807 ( .IN1(n4416), .IN2(n11447), .QN(n16634) );
  NOR2X0 U16808 ( .IN1(n11444), .IN2(g2072), .QN(n16633) );
  INVX0 U16809 ( .INP(n11447), .ZN(n11444) );
  NAND2X0 U16810 ( .IN1(n16635), .IN2(n16636), .QN(n11447) );
  NAND2X0 U16811 ( .IN1(g7357), .IN2(n10336), .QN(n16636) );
  NOR2X0 U16812 ( .IN1(n16637), .IN2(n16638), .QN(n16635) );
  NOR2X0 U16813 ( .IN1(n4293), .IN2(g2105), .QN(n16638) );
  NOR2X0 U16814 ( .IN1(n4307), .IN2(g2106), .QN(n16637) );
  NOR2X0 U16815 ( .IN1(n16639), .IN2(n16640), .QN(n16631) );
  NAND2X0 U16816 ( .IN1(n16641), .IN2(n16642), .QN(n16640) );
  NAND2X0 U16817 ( .IN1(n4409), .IN2(n11519), .QN(n16642) );
  NAND2X0 U16818 ( .IN1(n11517), .IN2(g2052), .QN(n16641) );
  INVX0 U16819 ( .INP(n11519), .ZN(n11517) );
  NAND2X0 U16820 ( .IN1(n16643), .IN2(n16644), .QN(n11519) );
  NAND2X0 U16821 ( .IN1(n10167), .IN2(g2009), .QN(n16644) );
  NOR2X0 U16822 ( .IN1(n16645), .IN2(n16646), .QN(n16643) );
  NOR2X0 U16823 ( .IN1(n4307), .IN2(g2094), .QN(n16646) );
  NOR2X0 U16824 ( .IN1(n4357), .IN2(g2095), .QN(n16645) );
  NOR2X0 U16825 ( .IN1(n16647), .IN2(n16648), .QN(n16639) );
  NOR2X0 U16826 ( .IN1(test_so70), .IN2(n11439), .QN(n16648) );
  NOR2X0 U16827 ( .IN1(n11436), .IN2(n10323), .QN(n16647) );
  INVX0 U16828 ( .INP(n11439), .ZN(n11436) );
  NAND2X0 U16829 ( .IN1(n16649), .IN2(n16650), .QN(n11439) );
  NAND2X0 U16830 ( .IN1(n10164), .IN2(g2009), .QN(n16650) );
  NOR2X0 U16831 ( .IN1(n16651), .IN2(n16652), .QN(n16649) );
  NOR2X0 U16832 ( .IN1(n4307), .IN2(g2103), .QN(n16652) );
  NOR2X0 U16833 ( .IN1(n4357), .IN2(g2104), .QN(n16651) );
  NOR2X0 U16834 ( .IN1(n16653), .IN2(n16654), .QN(n16613) );
  NAND2X0 U16835 ( .IN1(n16655), .IN2(n16656), .QN(n16654) );
  NOR2X0 U16836 ( .IN1(n16657), .IN2(n16658), .QN(n16656) );
  NOR2X0 U16837 ( .IN1(n4420), .IN2(n11531), .QN(n16658) );
  NOR2X0 U16838 ( .IN1(n11530), .IN2(g2033), .QN(n16657) );
  INVX0 U16839 ( .INP(n11531), .ZN(n11530) );
  NAND2X0 U16840 ( .IN1(n16659), .IN2(n16660), .QN(n11531) );
  NAND2X0 U16841 ( .IN1(n10170), .IN2(g2009), .QN(n16660) );
  NOR2X0 U16842 ( .IN1(n16661), .IN2(n16662), .QN(n16659) );
  NOR2X0 U16843 ( .IN1(n4307), .IN2(g2085), .QN(n16662) );
  NOR2X0 U16844 ( .IN1(n4357), .IN2(g2086), .QN(n16661) );
  NOR2X0 U16845 ( .IN1(n16663), .IN2(n16664), .QN(n16655) );
  NOR2X0 U16846 ( .IN1(n4474), .IN2(n11496), .QN(n16664) );
  NOR2X0 U16847 ( .IN1(n11495), .IN2(g2013), .QN(n16663) );
  INVX0 U16848 ( .INP(n11496), .ZN(n11495) );
  NAND2X0 U16849 ( .IN1(n16665), .IN2(n16666), .QN(n11496) );
  NAND2X0 U16850 ( .IN1(n10171), .IN2(g2009), .QN(n16666) );
  NOR2X0 U16851 ( .IN1(n16667), .IN2(n16668), .QN(n16665) );
  NOR2X0 U16852 ( .IN1(n4307), .IN2(g2082), .QN(n16668) );
  NOR2X0 U16853 ( .IN1(n4357), .IN2(g2083), .QN(n16667) );
  NAND2X0 U16854 ( .IN1(n16669), .IN2(n16670), .QN(n16653) );
  NOR2X0 U16855 ( .IN1(n16671), .IN2(n16672), .QN(n16670) );
  NOR2X0 U16856 ( .IN1(n4399), .IN2(n11536), .QN(n16672) );
  INVX0 U16857 ( .INP(n11535), .ZN(n11536) );
  NOR2X0 U16858 ( .IN1(n11535), .IN2(g2040), .QN(n16671) );
  NOR2X0 U16859 ( .IN1(n16673), .IN2(n16674), .QN(n11535) );
  NOR2X0 U16860 ( .IN1(n4357), .IN2(test_so71), .QN(n16674) );
  INVX0 U16861 ( .INP(n16675), .ZN(n16673) );
  NOR2X0 U16862 ( .IN1(n16676), .IN2(n16677), .QN(n16675) );
  NOR2X0 U16863 ( .IN1(n4293), .IN2(g2090), .QN(n16677) );
  NOR2X0 U16864 ( .IN1(n4307), .IN2(g2091), .QN(n16676) );
  NOR2X0 U16865 ( .IN1(n16678), .IN2(n16679), .QN(n16669) );
  NAND2X0 U16866 ( .IN1(n16680), .IN2(n16681), .QN(n16679) );
  NAND2X0 U16867 ( .IN1(n4473), .IN2(n11503), .QN(n16681) );
  NAND2X0 U16868 ( .IN1(n11502), .IN2(g2059), .QN(n16680) );
  INVX0 U16869 ( .INP(n11503), .ZN(n11502) );
  NAND2X0 U16870 ( .IN1(n16682), .IN2(n16683), .QN(n11503) );
  NAND2X0 U16871 ( .IN1(n10165), .IN2(g2009), .QN(n16683) );
  NOR2X0 U16872 ( .IN1(n16684), .IN2(n16685), .QN(n16682) );
  NOR2X0 U16873 ( .IN1(n4307), .IN2(g2100), .QN(n16685) );
  NOR2X0 U16874 ( .IN1(n4357), .IN2(g2101), .QN(n16684) );
  NAND2X0 U16875 ( .IN1(n16686), .IN2(n16687), .QN(n16678) );
  NAND2X0 U16876 ( .IN1(n4468), .IN2(n11466), .QN(n16687) );
  NAND2X0 U16877 ( .IN1(n11465), .IN2(g2046), .QN(n16686) );
  INVX0 U16878 ( .INP(n11466), .ZN(n11465) );
  NAND2X0 U16879 ( .IN1(n16688), .IN2(n16689), .QN(n11466) );
  NAND2X0 U16880 ( .IN1(n10166), .IN2(g2009), .QN(n16689) );
  NOR2X0 U16881 ( .IN1(n16690), .IN2(n16691), .QN(n16688) );
  NOR2X0 U16882 ( .IN1(n4307), .IN2(g2097), .QN(n16691) );
  NOR2X0 U16883 ( .IN1(n4357), .IN2(g2098), .QN(n16690) );
  NAND2X0 U16884 ( .IN1(n10299), .IN2(g7229), .QN(n16611) );
  NOR2X0 U16885 ( .IN1(n4293), .IN2(g2108), .QN(n16609) );
  NOR2X0 U16886 ( .IN1(n16692), .IN2(n11876), .QN(n16607) );
  NAND2X0 U16887 ( .IN1(n16693), .IN2(n16694), .QN(n11876) );
  NAND2X0 U16888 ( .IN1(n9880), .IN2(g7357), .QN(n16694) );
  NOR2X0 U16889 ( .IN1(n16695), .IN2(n16696), .QN(n16693) );
  INVX0 U16890 ( .INP(n16697), .ZN(n16696) );
  NAND2X0 U16891 ( .IN1(g7229), .IN2(n9887), .QN(n16697) );
  NOR2X0 U16892 ( .IN1(n4293), .IN2(g2111), .QN(n16695) );
  NOR2X0 U16893 ( .IN1(n4357), .IN2(g2110), .QN(n16692) );
  NAND2X0 U16894 ( .IN1(n16698), .IN2(g2115), .QN(n16603) );
  NAND2X0 U16895 ( .IN1(n16699), .IN2(n16700), .QN(g25267) );
  NAND2X0 U16896 ( .IN1(n16701), .IN2(g1422), .QN(n16700) );
  NAND2X0 U16897 ( .IN1(n16702), .IN2(n16601), .QN(n16699) );
  NAND2X0 U16898 ( .IN1(n16703), .IN2(n16704), .QN(g25266) );
  NAND2X0 U16899 ( .IN1(n16705), .IN2(g734), .QN(n16704) );
  NAND2X0 U16900 ( .IN1(n16706), .IN2(n16707), .QN(n16703) );
  NAND2X0 U16901 ( .IN1(n16708), .IN2(n16709), .QN(g25265) );
  NAND2X0 U16902 ( .IN1(n15740), .IN2(n11062), .QN(n16709) );
  NAND2X0 U16903 ( .IN1(n16710), .IN2(n16326), .QN(n16708) );
  INVX0 U16904 ( .INP(n15740), .ZN(n16326) );
  NAND2X0 U16905 ( .IN1(n16711), .IN2(n16712), .QN(n16710) );
  INVX0 U16906 ( .INP(n16713), .ZN(n16712) );
  NOR2X0 U16907 ( .IN1(g2993), .IN2(n10302), .QN(n16713) );
  NAND2X0 U16908 ( .IN1(n10302), .IN2(g2993), .QN(n16711) );
  NAND2X0 U16909 ( .IN1(n16714), .IN2(n16715), .QN(g25263) );
  NAND2X0 U16910 ( .IN1(n16716), .IN2(g1421), .QN(n16715) );
  NAND2X0 U16911 ( .IN1(n16717), .IN2(n16601), .QN(n16714) );
  INVX0 U16912 ( .INP(n16718), .ZN(n16601) );
  NAND2X0 U16913 ( .IN1(n16719), .IN2(n16720), .QN(n16718) );
  NOR2X0 U16914 ( .IN1(n16721), .IN2(n16722), .QN(n16720) );
  NAND2X0 U16915 ( .IN1(n16723), .IN2(n16724), .QN(n16722) );
  NAND2X0 U16916 ( .IN1(n16725), .IN2(n16726), .QN(n16724) );
  NOR2X0 U16917 ( .IN1(n16727), .IN2(n16728), .QN(n16726) );
  NAND2X0 U16918 ( .IN1(n16729), .IN2(n16730), .QN(n16728) );
  NOR2X0 U16919 ( .IN1(n16731), .IN2(n16732), .QN(n16730) );
  NOR2X0 U16920 ( .IN1(n4402), .IN2(n11667), .QN(n16732) );
  NOR2X0 U16921 ( .IN1(n11666), .IN2(g1326), .QN(n16731) );
  INVX0 U16922 ( .INP(n11667), .ZN(n11666) );
  NAND2X0 U16923 ( .IN1(n16733), .IN2(n16734), .QN(n11667) );
  NAND2X0 U16924 ( .IN1(g6979), .IN2(n10337), .QN(n16734) );
  NOR2X0 U16925 ( .IN1(n16735), .IN2(n16736), .QN(n16733) );
  NOR2X0 U16926 ( .IN1(n4294), .IN2(g1384), .QN(n16736) );
  NOR2X0 U16927 ( .IN1(n4358), .IN2(g1386), .QN(n16735) );
  NOR2X0 U16928 ( .IN1(n16737), .IN2(n16738), .QN(n16729) );
  NOR2X0 U16929 ( .IN1(n4412), .IN2(n11688), .QN(n16738) );
  NOR2X0 U16930 ( .IN1(n11687), .IN2(g1332), .QN(n16737) );
  INVX0 U16931 ( .INP(n11688), .ZN(n11687) );
  NAND2X0 U16932 ( .IN1(n16739), .IN2(n16740), .QN(n11688) );
  NAND2X0 U16933 ( .IN1(n10179), .IN2(g1315), .QN(n16740) );
  NOR2X0 U16934 ( .IN1(n16741), .IN2(n16742), .QN(n16739) );
  NOR2X0 U16935 ( .IN1(n4308), .IN2(g1394), .QN(n16742) );
  NOR2X0 U16936 ( .IN1(n4358), .IN2(g1395), .QN(n16741) );
  NAND2X0 U16937 ( .IN1(n16743), .IN2(n16744), .QN(n16727) );
  NOR2X0 U16938 ( .IN1(n16745), .IN2(n16746), .QN(n16744) );
  NOR2X0 U16939 ( .IN1(n4395), .IN2(n11615), .QN(n16746) );
  NOR2X0 U16940 ( .IN1(n11612), .IN2(g1372), .QN(n16745) );
  INVX0 U16941 ( .INP(n11615), .ZN(n11612) );
  NAND2X0 U16942 ( .IN1(n16747), .IN2(n16748), .QN(n11615) );
  NAND2X0 U16943 ( .IN1(n10174), .IN2(g1315), .QN(n16748) );
  NOR2X0 U16944 ( .IN1(n16749), .IN2(n16750), .QN(n16747) );
  NOR2X0 U16945 ( .IN1(n4308), .IN2(g1409), .QN(n16750) );
  NOR2X0 U16946 ( .IN1(n4358), .IN2(g1410), .QN(n16749) );
  NOR2X0 U16947 ( .IN1(n16751), .IN2(n16752), .QN(n16743) );
  NAND2X0 U16948 ( .IN1(n16753), .IN2(n16754), .QN(n16752) );
  NAND2X0 U16949 ( .IN1(n4417), .IN2(n11623), .QN(n16754) );
  NAND2X0 U16950 ( .IN1(n11620), .IN2(g1378), .QN(n16753) );
  INVX0 U16951 ( .INP(n11623), .ZN(n11620) );
  NAND2X0 U16952 ( .IN1(n16755), .IN2(n16756), .QN(n11623) );
  NAND2X0 U16953 ( .IN1(n10173), .IN2(g1315), .QN(n16756) );
  NOR2X0 U16954 ( .IN1(n16757), .IN2(n16758), .QN(n16755) );
  NOR2X0 U16955 ( .IN1(n4308), .IN2(g1412), .QN(n16758) );
  NOR2X0 U16956 ( .IN1(n4358), .IN2(g1413), .QN(n16757) );
  NAND2X0 U16957 ( .IN1(n16759), .IN2(n16760), .QN(n16751) );
  NAND2X0 U16958 ( .IN1(n4411), .IN2(n11695), .QN(n16760) );
  INVX0 U16959 ( .INP(n11693), .ZN(n11695) );
  NAND2X0 U16960 ( .IN1(n11693), .IN2(g1358), .QN(n16759) );
  NOR2X0 U16961 ( .IN1(n16761), .IN2(n16762), .QN(n11693) );
  NOR2X0 U16962 ( .IN1(n4358), .IN2(test_so50), .QN(n16762) );
  INVX0 U16963 ( .INP(n16763), .ZN(n16761) );
  NOR2X0 U16964 ( .IN1(n16764), .IN2(n16765), .QN(n16763) );
  NOR2X0 U16965 ( .IN1(n4294), .IN2(g1399), .QN(n16765) );
  NOR2X0 U16966 ( .IN1(n4308), .IN2(g1400), .QN(n16764) );
  NOR2X0 U16967 ( .IN1(n16766), .IN2(n16767), .QN(n16725) );
  NAND2X0 U16968 ( .IN1(n16768), .IN2(n16769), .QN(n16767) );
  NOR2X0 U16969 ( .IN1(n16770), .IN2(n16771), .QN(n16769) );
  NOR2X0 U16970 ( .IN1(n4421), .IN2(n11707), .QN(n16771) );
  NOR2X0 U16971 ( .IN1(n11706), .IN2(g1339), .QN(n16770) );
  INVX0 U16972 ( .INP(n11707), .ZN(n11706) );
  NAND2X0 U16973 ( .IN1(n16772), .IN2(n16773), .QN(n11707) );
  NAND2X0 U16974 ( .IN1(n10180), .IN2(g1315), .QN(n16773) );
  NOR2X0 U16975 ( .IN1(n16774), .IN2(n16775), .QN(n16772) );
  NOR2X0 U16976 ( .IN1(n4308), .IN2(g1391), .QN(n16775) );
  NOR2X0 U16977 ( .IN1(n4358), .IN2(g1392), .QN(n16774) );
  NOR2X0 U16978 ( .IN1(n16776), .IN2(n16777), .QN(n16768) );
  NOR2X0 U16979 ( .IN1(n4476), .IN2(n11672), .QN(n16777) );
  NOR2X0 U16980 ( .IN1(n11671), .IN2(g1319), .QN(n16776) );
  INVX0 U16981 ( .INP(n11672), .ZN(n11671) );
  NAND2X0 U16982 ( .IN1(n16778), .IN2(n16779), .QN(n11672) );
  NAND2X0 U16983 ( .IN1(n10181), .IN2(g1315), .QN(n16779) );
  NOR2X0 U16984 ( .IN1(n16780), .IN2(n16781), .QN(n16778) );
  NOR2X0 U16985 ( .IN1(n4308), .IN2(g1388), .QN(n16781) );
  NOR2X0 U16986 ( .IN1(n4358), .IN2(g1389), .QN(n16780) );
  NAND2X0 U16987 ( .IN1(n16782), .IN2(n16783), .QN(n16766) );
  NOR2X0 U16988 ( .IN1(n16784), .IN2(n16785), .QN(n16783) );
  NOR2X0 U16989 ( .IN1(n4401), .IN2(n11712), .QN(n16785) );
  NOR2X0 U16990 ( .IN1(n11711), .IN2(g1346), .QN(n16784) );
  INVX0 U16991 ( .INP(n11712), .ZN(n11711) );
  NAND2X0 U16992 ( .IN1(n16786), .IN2(n16787), .QN(n11712) );
  NAND2X0 U16993 ( .IN1(n10178), .IN2(g1315), .QN(n16787) );
  NOR2X0 U16994 ( .IN1(n16788), .IN2(n16789), .QN(n16786) );
  NOR2X0 U16995 ( .IN1(n4308), .IN2(g1397), .QN(n16789) );
  NOR2X0 U16996 ( .IN1(n4358), .IN2(g1398), .QN(n16788) );
  NOR2X0 U16997 ( .IN1(n16790), .IN2(n16791), .QN(n16782) );
  NAND2X0 U16998 ( .IN1(n16792), .IN2(n16793), .QN(n16791) );
  NAND2X0 U16999 ( .IN1(n4475), .IN2(n11679), .QN(n16793) );
  NAND2X0 U17000 ( .IN1(n11678), .IN2(g1365), .QN(n16792) );
  INVX0 U17001 ( .INP(n11679), .ZN(n11678) );
  NAND2X0 U17002 ( .IN1(n16794), .IN2(n16795), .QN(n11679) );
  NAND2X0 U17003 ( .IN1(n10175), .IN2(g1315), .QN(n16795) );
  NOR2X0 U17004 ( .IN1(n16796), .IN2(n16797), .QN(n16794) );
  NOR2X0 U17005 ( .IN1(n4308), .IN2(g1406), .QN(n16797) );
  NOR2X0 U17006 ( .IN1(n4358), .IN2(g1407), .QN(n16796) );
  NAND2X0 U17007 ( .IN1(n16798), .IN2(n16799), .QN(n16790) );
  NAND2X0 U17008 ( .IN1(n4469), .IN2(n11642), .QN(n16799) );
  NAND2X0 U17009 ( .IN1(n11641), .IN2(g1352), .QN(n16798) );
  INVX0 U17010 ( .INP(n11642), .ZN(n11641) );
  NAND2X0 U17011 ( .IN1(n16800), .IN2(n16801), .QN(n11642) );
  NAND2X0 U17012 ( .IN1(n10176), .IN2(g1315), .QN(n16801) );
  NOR2X0 U17013 ( .IN1(n16802), .IN2(n16803), .QN(n16800) );
  NOR2X0 U17014 ( .IN1(n4308), .IN2(g1403), .QN(n16803) );
  NOR2X0 U17015 ( .IN1(n4358), .IN2(g1404), .QN(n16802) );
  NAND2X0 U17016 ( .IN1(n10298), .IN2(g6979), .QN(n16723) );
  NOR2X0 U17017 ( .IN1(test_so51), .IN2(n4294), .QN(n16721) );
  NOR2X0 U17018 ( .IN1(n16804), .IN2(n11901), .QN(n16719) );
  NAND2X0 U17019 ( .IN1(n16805), .IN2(n16806), .QN(n11901) );
  NAND2X0 U17020 ( .IN1(n9882), .IN2(g7161), .QN(n16806) );
  NOR2X0 U17021 ( .IN1(n16807), .IN2(n16808), .QN(n16805) );
  INVX0 U17022 ( .INP(n16809), .ZN(n16808) );
  NAND2X0 U17023 ( .IN1(g6979), .IN2(n9888), .QN(n16809) );
  NOR2X0 U17024 ( .IN1(n4294), .IN2(g1417), .QN(n16807) );
  NOR2X0 U17025 ( .IN1(n4358), .IN2(g1416), .QN(n16804) );
  NAND2X0 U17026 ( .IN1(n16810), .IN2(n16811), .QN(g25262) );
  NAND2X0 U17027 ( .IN1(n16812), .IN2(g736), .QN(n16811) );
  NAND2X0 U17028 ( .IN1(n16813), .IN2(n16706), .QN(n16810) );
  NAND2X0 U17029 ( .IN1(n16814), .IN2(n16815), .QN(g25260) );
  NAND2X0 U17030 ( .IN1(n16816), .IN2(g735), .QN(n16815) );
  NAND2X0 U17031 ( .IN1(n16817), .IN2(n16706), .QN(n16814) );
  INVX0 U17032 ( .INP(n16818), .ZN(n16706) );
  NAND2X0 U17033 ( .IN1(n16819), .IN2(n16820), .QN(n16818) );
  NOR2X0 U17034 ( .IN1(n16821), .IN2(n16822), .QN(n16820) );
  NAND2X0 U17035 ( .IN1(n16823), .IN2(n16824), .QN(n16822) );
  NAND2X0 U17036 ( .IN1(n16825), .IN2(n16826), .QN(n16824) );
  NOR2X0 U17037 ( .IN1(n16827), .IN2(n16828), .QN(n16826) );
  NAND2X0 U17038 ( .IN1(n16829), .IN2(n16830), .QN(n16828) );
  NOR2X0 U17039 ( .IN1(n16831), .IN2(n16832), .QN(n16830) );
  NOR2X0 U17040 ( .IN1(n4414), .IN2(n11163), .QN(n16832) );
  NOR2X0 U17041 ( .IN1(n11162), .IN2(g646), .QN(n16831) );
  INVX0 U17042 ( .INP(n11163), .ZN(n11162) );
  NAND2X0 U17043 ( .IN1(n16833), .IN2(n16834), .QN(n11163) );
  NAND2X0 U17044 ( .IN1(n10189), .IN2(g629), .QN(n16834) );
  NOR2X0 U17045 ( .IN1(n16835), .IN2(n16836), .QN(n16833) );
  NOR2X0 U17046 ( .IN1(n4309), .IN2(g708), .QN(n16836) );
  NOR2X0 U17047 ( .IN1(n4359), .IN2(g709), .QN(n16835) );
  NOR2X0 U17048 ( .IN1(n16837), .IN2(n16838), .QN(n16829) );
  NOR2X0 U17049 ( .IN1(n4413), .IN2(n11108), .QN(n16838) );
  NOR2X0 U17050 ( .IN1(n11107), .IN2(g672), .QN(n16837) );
  INVX0 U17051 ( .INP(n11108), .ZN(n11107) );
  NAND2X0 U17052 ( .IN1(n16839), .IN2(n16840), .QN(n11108) );
  NAND2X0 U17053 ( .IN1(n10187), .IN2(g629), .QN(n16840) );
  NOR2X0 U17054 ( .IN1(n16841), .IN2(n16842), .QN(n16839) );
  NOR2X0 U17055 ( .IN1(n4309), .IN2(g714), .QN(n16842) );
  NOR2X0 U17056 ( .IN1(n4359), .IN2(g715), .QN(n16841) );
  NAND2X0 U17057 ( .IN1(n16843), .IN2(n16844), .QN(n16827) );
  NOR2X0 U17058 ( .IN1(n16845), .IN2(n16846), .QN(n16844) );
  NOR2X0 U17059 ( .IN1(n4418), .IN2(n11179), .QN(n16846) );
  NOR2X0 U17060 ( .IN1(n11177), .IN2(g692), .QN(n16845) );
  INVX0 U17061 ( .INP(n11179), .ZN(n11177) );
  NAND2X0 U17062 ( .IN1(n16847), .IN2(n16848), .QN(n11179) );
  INVX0 U17063 ( .INP(n16849), .ZN(n16848) );
  NOR2X0 U17064 ( .IN1(n4359), .IN2(test_so30), .QN(n16849) );
  NOR2X0 U17065 ( .IN1(n16850), .IN2(n16851), .QN(n16847) );
  NOR2X0 U17066 ( .IN1(n4295), .IN2(g725), .QN(n16851) );
  NOR2X0 U17067 ( .IN1(n4309), .IN2(g726), .QN(n16850) );
  NOR2X0 U17068 ( .IN1(n16852), .IN2(n16853), .QN(n16843) );
  NAND2X0 U17069 ( .IN1(n16854), .IN2(n16855), .QN(n16853) );
  NAND2X0 U17070 ( .IN1(n4396), .IN2(n11187), .QN(n16855) );
  NAND2X0 U17071 ( .IN1(n11186), .IN2(g686), .QN(n16854) );
  INVX0 U17072 ( .INP(n11187), .ZN(n11186) );
  NAND2X0 U17073 ( .IN1(n16856), .IN2(n16857), .QN(n11187) );
  NAND2X0 U17074 ( .IN1(n10184), .IN2(g629), .QN(n16857) );
  NOR2X0 U17075 ( .IN1(n16858), .IN2(n16859), .QN(n16856) );
  NOR2X0 U17076 ( .IN1(n4309), .IN2(g723), .QN(n16859) );
  NOR2X0 U17077 ( .IN1(n4359), .IN2(g724), .QN(n16858) );
  NOR2X0 U17078 ( .IN1(n16860), .IN2(n16861), .QN(n16852) );
  NOR2X0 U17079 ( .IN1(test_so28), .IN2(n11131), .QN(n16861) );
  NOR2X0 U17080 ( .IN1(n11128), .IN2(n10325), .QN(n16860) );
  INVX0 U17081 ( .INP(n11131), .ZN(n11128) );
  NAND2X0 U17082 ( .IN1(n16862), .IN2(n16863), .QN(n11131) );
  NAND2X0 U17083 ( .IN1(n10186), .IN2(g629), .QN(n16863) );
  NOR2X0 U17084 ( .IN1(n16864), .IN2(n16865), .QN(n16862) );
  NOR2X0 U17085 ( .IN1(n4309), .IN2(g717), .QN(n16865) );
  NOR2X0 U17086 ( .IN1(n4359), .IN2(g718), .QN(n16864) );
  NOR2X0 U17087 ( .IN1(n16866), .IN2(n16867), .QN(n16825) );
  NAND2X0 U17088 ( .IN1(n16868), .IN2(n16869), .QN(n16867) );
  NOR2X0 U17089 ( .IN1(n16870), .IN2(n16871), .QN(n16869) );
  NOR2X0 U17090 ( .IN1(n4422), .IN2(n11144), .QN(n16871) );
  NOR2X0 U17091 ( .IN1(n11143), .IN2(g653), .QN(n16870) );
  INVX0 U17092 ( .INP(n11144), .ZN(n11143) );
  NAND2X0 U17093 ( .IN1(n16872), .IN2(n16873), .QN(n11144) );
  NAND2X0 U17094 ( .IN1(n10190), .IN2(g629), .QN(n16873) );
  NOR2X0 U17095 ( .IN1(n16874), .IN2(n16875), .QN(n16872) );
  NOR2X0 U17096 ( .IN1(n4309), .IN2(g705), .QN(n16875) );
  NOR2X0 U17097 ( .IN1(n4359), .IN2(g706), .QN(n16874) );
  NOR2X0 U17098 ( .IN1(n16876), .IN2(n16877), .QN(n16868) );
  NOR2X0 U17099 ( .IN1(n4478), .IN2(n11097), .QN(n16877) );
  NOR2X0 U17100 ( .IN1(n11094), .IN2(g633), .QN(n16876) );
  INVX0 U17101 ( .INP(n11097), .ZN(n11094) );
  NAND2X0 U17102 ( .IN1(n16878), .IN2(n16879), .QN(n11097) );
  NAND2X0 U17103 ( .IN1(n10191), .IN2(g629), .QN(n16879) );
  NOR2X0 U17104 ( .IN1(n16880), .IN2(n16881), .QN(n16878) );
  NOR2X0 U17105 ( .IN1(n4309), .IN2(g702), .QN(n16881) );
  NOR2X0 U17106 ( .IN1(n4359), .IN2(g703), .QN(n16880) );
  NAND2X0 U17107 ( .IN1(n16882), .IN2(n16883), .QN(n16866) );
  NOR2X0 U17108 ( .IN1(n16884), .IN2(n16885), .QN(n16883) );
  NOR2X0 U17109 ( .IN1(n4477), .IN2(n11149), .QN(n16885) );
  NOR2X0 U17110 ( .IN1(n11148), .IN2(g679), .QN(n16884) );
  INVX0 U17111 ( .INP(n11149), .ZN(n11148) );
  NAND2X0 U17112 ( .IN1(n16886), .IN2(n16887), .QN(n11149) );
  NAND2X0 U17113 ( .IN1(n10185), .IN2(g629), .QN(n16887) );
  NOR2X0 U17114 ( .IN1(n16888), .IN2(n16889), .QN(n16886) );
  NOR2X0 U17115 ( .IN1(n4309), .IN2(g720), .QN(n16889) );
  NOR2X0 U17116 ( .IN1(n4359), .IN2(g721), .QN(n16888) );
  NOR2X0 U17117 ( .IN1(n16890), .IN2(n16891), .QN(n16882) );
  NAND2X0 U17118 ( .IN1(n16892), .IN2(n16893), .QN(n16891) );
  NAND2X0 U17119 ( .IN1(n4404), .IN2(n11158), .QN(n16893) );
  NAND2X0 U17120 ( .IN1(n11157), .IN2(g640), .QN(n16892) );
  INVX0 U17121 ( .INP(n11158), .ZN(n11157) );
  NAND2X0 U17122 ( .IN1(n16894), .IN2(n16895), .QN(n11158) );
  NAND2X0 U17123 ( .IN1(n10192), .IN2(g629), .QN(n16895) );
  NOR2X0 U17124 ( .IN1(n16896), .IN2(n16897), .QN(n16894) );
  NOR2X0 U17125 ( .IN1(n4309), .IN2(g699), .QN(n16897) );
  NOR2X0 U17126 ( .IN1(n4359), .IN2(g700), .QN(n16896) );
  NAND2X0 U17127 ( .IN1(n16898), .IN2(n16899), .QN(n16890) );
  NAND2X0 U17128 ( .IN1(n4403), .IN2(n11136), .QN(n16899) );
  NAND2X0 U17129 ( .IN1(n11135), .IN2(g660), .QN(n16898) );
  INVX0 U17130 ( .INP(n11136), .ZN(n11135) );
  NAND2X0 U17131 ( .IN1(n16900), .IN2(n16901), .QN(n11136) );
  NAND2X0 U17132 ( .IN1(g6677), .IN2(n10338), .QN(n16901) );
  NOR2X0 U17133 ( .IN1(n16902), .IN2(n16903), .QN(n16900) );
  NOR2X0 U17134 ( .IN1(n4295), .IN2(g710), .QN(n16903) );
  NOR2X0 U17135 ( .IN1(n4359), .IN2(g712), .QN(n16902) );
  NAND2X0 U17136 ( .IN1(n10297), .IN2(g6677), .QN(n16823) );
  NOR2X0 U17137 ( .IN1(n4295), .IN2(g728), .QN(n16821) );
  NOR2X0 U17138 ( .IN1(n16904), .IN2(n11826), .QN(n16819) );
  NAND2X0 U17139 ( .IN1(n16905), .IN2(n16906), .QN(n11826) );
  NAND2X0 U17140 ( .IN1(n9884), .IN2(g6911), .QN(n16906) );
  NOR2X0 U17141 ( .IN1(n16907), .IN2(n16908), .QN(n16905) );
  INVX0 U17142 ( .INP(n16909), .ZN(n16908) );
  NAND2X0 U17143 ( .IN1(g6677), .IN2(n9889), .QN(n16909) );
  NOR2X0 U17144 ( .IN1(n4295), .IN2(g731), .QN(n16907) );
  NOR2X0 U17145 ( .IN1(n4359), .IN2(g730), .QN(n16904) );
  NAND2X0 U17146 ( .IN1(n16910), .IN2(n16911), .QN(g25259) );
  NAND2X0 U17147 ( .IN1(n16912), .IN2(n15602), .QN(n16911) );
  NAND2X0 U17148 ( .IN1(n16913), .IN2(g2253), .QN(n16910) );
  NAND2X0 U17149 ( .IN1(n16914), .IN2(n16915), .QN(g25257) );
  NAND2X0 U17150 ( .IN1(n16916), .IN2(n15602), .QN(n16915) );
  INVX0 U17151 ( .INP(n16917), .ZN(n16914) );
  NOR2X0 U17152 ( .IN1(n16916), .IN2(n9891), .QN(n16917) );
  NAND2X0 U17153 ( .IN1(n16918), .IN2(n16919), .QN(g25256) );
  NAND2X0 U17154 ( .IN1(n16912), .IN2(n4377), .QN(n16919) );
  NAND2X0 U17155 ( .IN1(n16913), .IN2(g2250), .QN(n16918) );
  NAND2X0 U17156 ( .IN1(n16920), .IN2(n16921), .QN(g25255) );
  NAND2X0 U17157 ( .IN1(n16922), .IN2(n15646), .QN(n16921) );
  NAND2X0 U17158 ( .IN1(n16923), .IN2(g1559), .QN(n16920) );
  NAND2X0 U17159 ( .IN1(n16924), .IN2(n16925), .QN(g25253) );
  NAND2X0 U17160 ( .IN1(n16926), .IN2(n15602), .QN(n16925) );
  NAND2X0 U17161 ( .IN1(n16927), .IN2(n16928), .QN(n15602) );
  NOR2X0 U17162 ( .IN1(n16929), .IN2(n16930), .QN(n16928) );
  NAND2X0 U17163 ( .IN1(g2165), .IN2(g2180), .QN(n16930) );
  NAND2X0 U17164 ( .IN1(g2190), .IN2(g2195), .QN(n16929) );
  NOR2X0 U17165 ( .IN1(n16931), .IN2(n16932), .QN(n16927) );
  NAND2X0 U17166 ( .IN1(g2200), .IN2(g2175), .QN(n16932) );
  NAND2X0 U17167 ( .IN1(g2185), .IN2(g2170), .QN(n16931) );
  NAND2X0 U17168 ( .IN1(n16933), .IN2(g2254), .QN(n16924) );
  NAND2X0 U17169 ( .IN1(n16934), .IN2(n16935), .QN(g25252) );
  NAND2X0 U17170 ( .IN1(n16916), .IN2(n4377), .QN(n16935) );
  INVX0 U17171 ( .INP(n16936), .ZN(n16934) );
  NOR2X0 U17172 ( .IN1(n16916), .IN2(n9894), .QN(n16936) );
  NAND2X0 U17173 ( .IN1(n16937), .IN2(n16938), .QN(g25251) );
  NAND2X0 U17174 ( .IN1(n16912), .IN2(n4373), .QN(n16938) );
  NAND2X0 U17175 ( .IN1(n16913), .IN2(g2247), .QN(n16937) );
  NAND2X0 U17176 ( .IN1(n16939), .IN2(n16940), .QN(g25250) );
  NAND2X0 U17177 ( .IN1(n16941), .IN2(n15646), .QN(n16940) );
  INVX0 U17178 ( .INP(n16942), .ZN(n16939) );
  NOR2X0 U17179 ( .IN1(n16941), .IN2(n9903), .QN(n16942) );
  NAND2X0 U17180 ( .IN1(n16943), .IN2(n16944), .QN(g25249) );
  NAND2X0 U17181 ( .IN1(n16922), .IN2(n4378), .QN(n16944) );
  NAND2X0 U17182 ( .IN1(n16923), .IN2(g1556), .QN(n16943) );
  NAND2X0 U17183 ( .IN1(n16945), .IN2(n16946), .QN(g25248) );
  NAND2X0 U17184 ( .IN1(n16947), .IN2(n15687), .QN(n16946) );
  INVX0 U17185 ( .INP(n16948), .ZN(n16945) );
  NOR2X0 U17186 ( .IN1(n16947), .IN2(n9913), .QN(n16948) );
  NAND2X0 U17187 ( .IN1(n16949), .IN2(n16950), .QN(g25247) );
  NAND2X0 U17188 ( .IN1(n16926), .IN2(n4377), .QN(n16950) );
  NAND2X0 U17189 ( .IN1(n16933), .IN2(g2251), .QN(n16949) );
  NAND2X0 U17190 ( .IN1(n16951), .IN2(n16952), .QN(g25246) );
  NAND2X0 U17191 ( .IN1(n16916), .IN2(n4373), .QN(n16952) );
  INVX0 U17192 ( .INP(n16953), .ZN(n16951) );
  NOR2X0 U17193 ( .IN1(n16916), .IN2(n9897), .QN(n16953) );
  NAND2X0 U17194 ( .IN1(n16954), .IN2(n16955), .QN(g25245) );
  NAND2X0 U17195 ( .IN1(n16913), .IN2(g2244), .QN(n16955) );
  INVX0 U17196 ( .INP(n16912), .ZN(n16913) );
  NAND2X0 U17197 ( .IN1(n16956), .IN2(n16912), .QN(n16954) );
  NOR2X0 U17198 ( .IN1(n11722), .IN2(n4367), .QN(n16912) );
  NAND2X0 U17199 ( .IN1(n16957), .IN2(n16958), .QN(g25244) );
  NAND2X0 U17200 ( .IN1(n16959), .IN2(n15646), .QN(n16958) );
  NAND2X0 U17201 ( .IN1(n16960), .IN2(n16961), .QN(n15646) );
  NOR2X0 U17202 ( .IN1(n16962), .IN2(n16963), .QN(n16961) );
  NAND2X0 U17203 ( .IN1(g1471), .IN2(g1486), .QN(n16963) );
  NAND2X0 U17204 ( .IN1(g1496), .IN2(g1501), .QN(n16962) );
  NOR2X0 U17205 ( .IN1(n16964), .IN2(n16965), .QN(n16960) );
  NAND2X0 U17206 ( .IN1(g1506), .IN2(g1481), .QN(n16965) );
  NAND2X0 U17207 ( .IN1(g1491), .IN2(g1476), .QN(n16964) );
  NAND2X0 U17208 ( .IN1(n16966), .IN2(g1560), .QN(n16957) );
  NAND2X0 U17209 ( .IN1(n16967), .IN2(n16968), .QN(g25243) );
  NAND2X0 U17210 ( .IN1(n16941), .IN2(n4378), .QN(n16968) );
  INVX0 U17211 ( .INP(n16969), .ZN(n16967) );
  NOR2X0 U17212 ( .IN1(n16941), .IN2(n9906), .QN(n16969) );
  NAND2X0 U17213 ( .IN1(n16970), .IN2(n16971), .QN(g25242) );
  NAND2X0 U17214 ( .IN1(test_so54), .IN2(n16923), .QN(n16971) );
  NAND2X0 U17215 ( .IN1(n16922), .IN2(n4374), .QN(n16970) );
  NAND2X0 U17216 ( .IN1(n16972), .IN2(n16973), .QN(g25241) );
  NAND2X0 U17217 ( .IN1(n16974), .IN2(n15687), .QN(n16973) );
  NAND2X0 U17218 ( .IN1(n16975), .IN2(g867), .QN(n16972) );
  NAND2X0 U17219 ( .IN1(n16976), .IN2(n16977), .QN(g25240) );
  NAND2X0 U17220 ( .IN1(n16947), .IN2(n4379), .QN(n16977) );
  INVX0 U17221 ( .INP(n16978), .ZN(n16976) );
  NOR2X0 U17222 ( .IN1(n16947), .IN2(n9916), .QN(n16978) );
  NAND2X0 U17223 ( .IN1(n16979), .IN2(n16980), .QN(g25239) );
  NAND2X0 U17224 ( .IN1(n16981), .IN2(n15721), .QN(n16980) );
  NAND2X0 U17225 ( .IN1(n16982), .IN2(g177), .QN(n16979) );
  NAND2X0 U17226 ( .IN1(n16983), .IN2(n16984), .QN(g25237) );
  NAND2X0 U17227 ( .IN1(n16926), .IN2(n4373), .QN(n16984) );
  NAND2X0 U17228 ( .IN1(n16933), .IN2(g2248), .QN(n16983) );
  NAND2X0 U17229 ( .IN1(n16985), .IN2(n16986), .QN(g25236) );
  INVX0 U17230 ( .INP(n16987), .ZN(n16986) );
  NOR2X0 U17231 ( .IN1(n16916), .IN2(n9900), .QN(n16987) );
  NAND2X0 U17232 ( .IN1(n16956), .IN2(n16916), .QN(n16985) );
  NOR2X0 U17233 ( .IN1(n11722), .IN2(n10320), .QN(n16916) );
  NAND2X0 U17234 ( .IN1(n16988), .IN2(n16989), .QN(g25235) );
  NAND2X0 U17235 ( .IN1(n16959), .IN2(n4378), .QN(n16989) );
  NAND2X0 U17236 ( .IN1(n16966), .IN2(g1557), .QN(n16988) );
  NAND2X0 U17237 ( .IN1(n16990), .IN2(n16991), .QN(g25234) );
  NAND2X0 U17238 ( .IN1(n16941), .IN2(n4374), .QN(n16991) );
  INVX0 U17239 ( .INP(n16992), .ZN(n16990) );
  NOR2X0 U17240 ( .IN1(n16941), .IN2(n9908), .QN(n16992) );
  NAND2X0 U17241 ( .IN1(n16993), .IN2(n16994), .QN(g25233) );
  NAND2X0 U17242 ( .IN1(n16923), .IN2(g1550), .QN(n16994) );
  INVX0 U17243 ( .INP(n16922), .ZN(n16923) );
  NAND2X0 U17244 ( .IN1(n16995), .IN2(n16922), .QN(n16993) );
  NOR2X0 U17245 ( .IN1(n11722), .IN2(n4368), .QN(n16922) );
  NAND2X0 U17246 ( .IN1(n16996), .IN2(n16997), .QN(g25232) );
  NAND2X0 U17247 ( .IN1(n16998), .IN2(n15687), .QN(n16997) );
  NAND2X0 U17248 ( .IN1(n16999), .IN2(n17000), .QN(n15687) );
  NOR2X0 U17249 ( .IN1(n17001), .IN2(n17002), .QN(n17000) );
  NAND2X0 U17250 ( .IN1(g785), .IN2(g797), .QN(n17002) );
  NAND2X0 U17251 ( .IN1(g805), .IN2(g809), .QN(n17001) );
  NOR2X0 U17252 ( .IN1(n17003), .IN2(n17004), .QN(n16999) );
  NAND2X0 U17253 ( .IN1(g813), .IN2(g793), .QN(n17004) );
  NAND2X0 U17254 ( .IN1(g801), .IN2(g789), .QN(n17003) );
  NAND2X0 U17255 ( .IN1(n17005), .IN2(g866), .QN(n16996) );
  NAND2X0 U17256 ( .IN1(n17006), .IN2(n17007), .QN(g25231) );
  NAND2X0 U17257 ( .IN1(n16974), .IN2(n4379), .QN(n17007) );
  NAND2X0 U17258 ( .IN1(n16975), .IN2(g864), .QN(n17006) );
  NAND2X0 U17259 ( .IN1(n17008), .IN2(n17009), .QN(g25230) );
  NAND2X0 U17260 ( .IN1(n16947), .IN2(n4375), .QN(n17009) );
  INVX0 U17261 ( .INP(n17010), .ZN(n17008) );
  NOR2X0 U17262 ( .IN1(n16947), .IN2(n9919), .QN(n17010) );
  NAND2X0 U17263 ( .IN1(n17011), .IN2(n17012), .QN(g25229) );
  NAND2X0 U17264 ( .IN1(n17013), .IN2(n15721), .QN(n17012) );
  INVX0 U17265 ( .INP(n17014), .ZN(n17011) );
  NOR2X0 U17266 ( .IN1(n17013), .IN2(n9925), .QN(n17014) );
  NAND2X0 U17267 ( .IN1(n17015), .IN2(n17016), .QN(g25228) );
  NAND2X0 U17268 ( .IN1(n16981), .IN2(n4380), .QN(n17016) );
  NAND2X0 U17269 ( .IN1(n16982), .IN2(g174), .QN(n17015) );
  NAND2X0 U17270 ( .IN1(n17017), .IN2(n17018), .QN(g25227) );
  NAND2X0 U17271 ( .IN1(n16933), .IN2(g2245), .QN(n17018) );
  INVX0 U17272 ( .INP(n16926), .ZN(n16933) );
  NAND2X0 U17273 ( .IN1(n16956), .IN2(n16926), .QN(n17017) );
  NOR2X0 U17274 ( .IN1(n11722), .IN2(n4324), .QN(n16926) );
  INVX0 U17275 ( .INP(n17019), .ZN(n16956) );
  NAND2X0 U17276 ( .IN1(n17020), .IN2(n17021), .QN(n17019) );
  NOR2X0 U17277 ( .IN1(n4325), .IN2(n4287), .QN(n17021) );
  NOR2X0 U17278 ( .IN1(g2190), .IN2(g2195), .QN(n17020) );
  NAND2X0 U17279 ( .IN1(n17022), .IN2(n17023), .QN(g25225) );
  NAND2X0 U17280 ( .IN1(n16959), .IN2(n4374), .QN(n17023) );
  NAND2X0 U17281 ( .IN1(n16966), .IN2(g1554), .QN(n17022) );
  NAND2X0 U17282 ( .IN1(n17024), .IN2(n17025), .QN(g25224) );
  INVX0 U17283 ( .INP(n17026), .ZN(n17025) );
  NOR2X0 U17284 ( .IN1(n16941), .IN2(n9911), .QN(n17026) );
  NAND2X0 U17285 ( .IN1(n16995), .IN2(n16941), .QN(n17024) );
  NOR2X0 U17286 ( .IN1(n11722), .IN2(n4515), .QN(n16941) );
  NAND2X0 U17287 ( .IN1(n17027), .IN2(n17028), .QN(g25223) );
  NAND2X0 U17288 ( .IN1(n16998), .IN2(n4379), .QN(n17028) );
  NAND2X0 U17289 ( .IN1(n17005), .IN2(g863), .QN(n17027) );
  NAND2X0 U17290 ( .IN1(n17029), .IN2(n17030), .QN(g25222) );
  NAND2X0 U17291 ( .IN1(n16974), .IN2(n4375), .QN(n17030) );
  NAND2X0 U17292 ( .IN1(n16975), .IN2(g861), .QN(n17029) );
  NAND2X0 U17293 ( .IN1(n17031), .IN2(n17032), .QN(g25221) );
  INVX0 U17294 ( .INP(n17033), .ZN(n17032) );
  NOR2X0 U17295 ( .IN1(n16947), .IN2(n9922), .QN(n17033) );
  NAND2X0 U17296 ( .IN1(n17034), .IN2(n16947), .QN(n17031) );
  NOR2X0 U17297 ( .IN1(n11722), .IN2(n10321), .QN(n16947) );
  NAND2X0 U17298 ( .IN1(n17035), .IN2(n17036), .QN(g25220) );
  NAND2X0 U17299 ( .IN1(n17037), .IN2(n15721), .QN(n17036) );
  NAND2X0 U17300 ( .IN1(n17038), .IN2(n17039), .QN(n15721) );
  NOR2X0 U17301 ( .IN1(n17040), .IN2(n17041), .QN(n17039) );
  NAND2X0 U17302 ( .IN1(g97), .IN2(g109), .QN(n17041) );
  NAND2X0 U17303 ( .IN1(g117), .IN2(g121), .QN(n17040) );
  NOR2X0 U17304 ( .IN1(n17042), .IN2(n17043), .QN(n17038) );
  NAND2X0 U17305 ( .IN1(g125), .IN2(g105), .QN(n17043) );
  NAND2X0 U17306 ( .IN1(g113), .IN2(g101), .QN(n17042) );
  NAND2X0 U17307 ( .IN1(n17044), .IN2(g178), .QN(n17035) );
  NAND2X0 U17308 ( .IN1(n17045), .IN2(n17046), .QN(g25219) );
  NAND2X0 U17309 ( .IN1(n17013), .IN2(n4380), .QN(n17046) );
  INVX0 U17310 ( .INP(n17047), .ZN(n17045) );
  NOR2X0 U17311 ( .IN1(n17013), .IN2(n9928), .QN(n17047) );
  NAND2X0 U17312 ( .IN1(n17048), .IN2(n17049), .QN(g25218) );
  NAND2X0 U17313 ( .IN1(n16981), .IN2(n4376), .QN(n17049) );
  NAND2X0 U17314 ( .IN1(n16982), .IN2(g171), .QN(n17048) );
  NAND2X0 U17315 ( .IN1(n17050), .IN2(n17051), .QN(g25217) );
  NAND2X0 U17316 ( .IN1(n16966), .IN2(g1551), .QN(n17051) );
  INVX0 U17317 ( .INP(n16959), .ZN(n16966) );
  NAND2X0 U17318 ( .IN1(n16995), .IN2(n16959), .QN(n17050) );
  NOR2X0 U17319 ( .IN1(n11722), .IN2(n4317), .QN(n16959) );
  INVX0 U17320 ( .INP(n17052), .ZN(n16995) );
  NAND2X0 U17321 ( .IN1(n17053), .IN2(n17054), .QN(n17052) );
  NOR2X0 U17322 ( .IN1(n4326), .IN2(n4288), .QN(n17054) );
  NOR2X0 U17323 ( .IN1(g1496), .IN2(g1501), .QN(n17053) );
  NAND2X0 U17324 ( .IN1(n17055), .IN2(n17056), .QN(g25215) );
  NAND2X0 U17325 ( .IN1(n16998), .IN2(n4375), .QN(n17056) );
  NAND2X0 U17326 ( .IN1(n17005), .IN2(g860), .QN(n17055) );
  NAND2X0 U17327 ( .IN1(n17057), .IN2(n17058), .QN(g25214) );
  NAND2X0 U17328 ( .IN1(test_so33), .IN2(n16975), .QN(n17058) );
  INVX0 U17329 ( .INP(n16974), .ZN(n16975) );
  NAND2X0 U17330 ( .IN1(n17034), .IN2(n16974), .QN(n17057) );
  NOR2X0 U17331 ( .IN1(n11722), .IN2(n4312), .QN(n16974) );
  NAND2X0 U17332 ( .IN1(n17059), .IN2(n17060), .QN(g25213) );
  NAND2X0 U17333 ( .IN1(n17037), .IN2(n4380), .QN(n17060) );
  NAND2X0 U17334 ( .IN1(n17044), .IN2(g175), .QN(n17059) );
  NAND2X0 U17335 ( .IN1(n17061), .IN2(n17062), .QN(g25212) );
  NAND2X0 U17336 ( .IN1(n17013), .IN2(n4376), .QN(n17062) );
  INVX0 U17337 ( .INP(n17063), .ZN(n17061) );
  NOR2X0 U17338 ( .IN1(n17013), .IN2(n9931), .QN(n17063) );
  NAND2X0 U17339 ( .IN1(n17064), .IN2(n17065), .QN(g25211) );
  NAND2X0 U17340 ( .IN1(n16982), .IN2(g168), .QN(n17065) );
  INVX0 U17341 ( .INP(n16981), .ZN(n16982) );
  NAND2X0 U17342 ( .IN1(n17066), .IN2(n16981), .QN(n17064) );
  NOR2X0 U17343 ( .IN1(n11722), .IN2(n4369), .QN(n16981) );
  NAND2X0 U17344 ( .IN1(n17067), .IN2(n17068), .QN(g25209) );
  NAND2X0 U17345 ( .IN1(n17005), .IN2(g857), .QN(n17068) );
  INVX0 U17346 ( .INP(n16998), .ZN(n17005) );
  NAND2X0 U17347 ( .IN1(n17034), .IN2(n16998), .QN(n17067) );
  NOR2X0 U17348 ( .IN1(n11722), .IN2(n4323), .QN(n16998) );
  INVX0 U17349 ( .INP(n17069), .ZN(n17034) );
  NAND2X0 U17350 ( .IN1(n17070), .IN2(n17071), .QN(n17069) );
  NOR2X0 U17351 ( .IN1(n4327), .IN2(n4289), .QN(n17071) );
  NOR2X0 U17352 ( .IN1(g805), .IN2(g809), .QN(n17070) );
  NAND2X0 U17353 ( .IN1(n17072), .IN2(n17073), .QN(g25207) );
  NAND2X0 U17354 ( .IN1(n17037), .IN2(n4376), .QN(n17073) );
  NAND2X0 U17355 ( .IN1(n17044), .IN2(g172), .QN(n17072) );
  NAND2X0 U17356 ( .IN1(n17074), .IN2(n17075), .QN(g25206) );
  INVX0 U17357 ( .INP(n17076), .ZN(n17075) );
  NOR2X0 U17358 ( .IN1(n17013), .IN2(n9934), .QN(n17076) );
  NAND2X0 U17359 ( .IN1(n17066), .IN2(n17013), .QN(n17074) );
  NOR2X0 U17360 ( .IN1(n11722), .IN2(n4512), .QN(n17013) );
  NAND2X0 U17361 ( .IN1(n17077), .IN2(n17078), .QN(g25204) );
  NAND2X0 U17362 ( .IN1(n17044), .IN2(g169), .QN(n17078) );
  INVX0 U17363 ( .INP(n17037), .ZN(n17044) );
  NAND2X0 U17364 ( .IN1(n17066), .IN2(n17037), .QN(n17077) );
  NOR2X0 U17365 ( .IN1(n11722), .IN2(n4318), .QN(n17037) );
  NAND2X0 U17366 ( .IN1(n17079), .IN2(n17080), .QN(n11722) );
  NOR2X0 U17367 ( .IN1(n17081), .IN2(n17082), .QN(n17080) );
  NAND2X0 U17368 ( .IN1(n4479), .IN2(n4482), .QN(n17082) );
  NAND2X0 U17369 ( .IN1(g2883), .IN2(g2924), .QN(n17081) );
  NOR2X0 U17370 ( .IN1(g2888), .IN2(n17083), .QN(n17079) );
  NAND2X0 U17371 ( .IN1(n10026), .IN2(n15466), .QN(n17083) );
  INVX0 U17372 ( .INP(n17084), .ZN(n17066) );
  NAND2X0 U17373 ( .IN1(n17085), .IN2(n17086), .QN(n17084) );
  NOR2X0 U17374 ( .IN1(n4328), .IN2(n4290), .QN(n17086) );
  NOR2X0 U17375 ( .IN1(g117), .IN2(g121), .QN(n17085) );
  NOR2X0 U17376 ( .IN1(n17087), .IN2(n17088), .QN(g25202) );
  NAND2X0 U17377 ( .IN1(n17089), .IN2(n17090), .QN(n17088) );
  NAND2X0 U17378 ( .IN1(n9736), .IN2(n17091), .QN(n17090) );
  NAND2X0 U17379 ( .IN1(n17092), .IN2(g3032), .QN(n17089) );
  NOR2X0 U17380 ( .IN1(n10998), .IN2(n17093), .QN(g25201) );
  NAND2X0 U17381 ( .IN1(n17094), .IN2(n16333), .QN(n17093) );
  INVX0 U17382 ( .INP(n17095), .ZN(n16333) );
  NOR2X0 U17383 ( .IN1(n18), .IN2(n4305), .QN(n17095) );
  INVX0 U17384 ( .INP(n4057), .ZN(n17094) );
  NAND2X0 U17385 ( .IN1(n17096), .IN2(n17097), .QN(g25199) );
  INVX0 U17386 ( .INP(n17098), .ZN(n17097) );
  NOR2X0 U17387 ( .IN1(n17099), .IN2(n10026), .QN(n17098) );
  NAND2X0 U17388 ( .IN1(n17100), .IN2(n10026), .QN(n17096) );
  NOR2X0 U17389 ( .IN1(n17101), .IN2(n17102), .QN(n17100) );
  NOR2X0 U17390 ( .IN1(n14690), .IN2(n17103), .QN(g25197) );
  NAND2X0 U17391 ( .IN1(n17104), .IN2(n17105), .QN(n17103) );
  NAND2X0 U17392 ( .IN1(n4397), .IN2(n15756), .QN(n17105) );
  NAND2X0 U17393 ( .IN1(n15754), .IN2(g2734), .QN(n17104) );
  INVX0 U17394 ( .INP(n15756), .ZN(n15754) );
  NOR2X0 U17395 ( .IN1(n15735), .IN2(n17106), .QN(g25194) );
  NAND2X0 U17396 ( .IN1(n17107), .IN2(n17108), .QN(n17106) );
  NAND2X0 U17397 ( .IN1(n4399), .IN2(n15774), .QN(n17108) );
  NAND2X0 U17398 ( .IN1(n15772), .IN2(g2040), .QN(n17107) );
  INVX0 U17399 ( .INP(n15774), .ZN(n15772) );
  NOR2X0 U17400 ( .IN1(n15740), .IN2(n17109), .QN(g25191) );
  NAND2X0 U17401 ( .IN1(n17110), .IN2(n3742), .QN(n17109) );
  NAND2X0 U17402 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  NAND2X0 U17403 ( .IN1(n10311), .IN2(n17111), .QN(n17110) );
  INVX0 U17404 ( .INP(n4065), .ZN(n17111) );
  NOR2X0 U17405 ( .IN1(n14704), .IN2(n17112), .QN(g25189) );
  NAND2X0 U17406 ( .IN1(n17113), .IN2(n17114), .QN(n17112) );
  NAND2X0 U17407 ( .IN1(n4401), .IN2(n15895), .QN(n17114) );
  NAND2X0 U17408 ( .IN1(n15893), .IN2(g1346), .QN(n17113) );
  INVX0 U17409 ( .INP(n15895), .ZN(n15893) );
  NOR2X0 U17410 ( .IN1(n14141), .IN2(n17115), .QN(g25185) );
  NAND2X0 U17411 ( .IN1(n17116), .IN2(n17117), .QN(n17115) );
  NAND2X0 U17412 ( .IN1(n4403), .IN2(n16016), .QN(n17117) );
  NAND2X0 U17413 ( .IN1(n16014), .IN2(g660), .QN(n17116) );
  INVX0 U17414 ( .INP(n16016), .ZN(n16014) );
  NOR2X0 U17415 ( .IN1(n13263), .IN2(n17118), .QN(g25067) );
  NAND2X0 U17416 ( .IN1(n17119), .IN2(n17120), .QN(n17118) );
  NAND2X0 U17417 ( .IN1(n10013), .IN2(n3888), .QN(n17120) );
  INVX0 U17418 ( .INP(n17121), .ZN(n3888) );
  NAND2X0 U17419 ( .IN1(n17121), .IN2(g2160), .QN(n17119) );
  NOR2X0 U17420 ( .IN1(n4367), .IN2(n15466), .QN(n17121) );
  NOR2X0 U17421 ( .IN1(n17122), .IN2(n10780), .QN(n13263) );
  NOR2X0 U17422 ( .IN1(n13268), .IN2(n17123), .QN(g25056) );
  NAND2X0 U17423 ( .IN1(n17124), .IN2(n17125), .QN(n17123) );
  NAND2X0 U17424 ( .IN1(n10017), .IN2(n3891), .QN(n17125) );
  INVX0 U17425 ( .INP(n17126), .ZN(n3891) );
  NAND2X0 U17426 ( .IN1(n17126), .IN2(g1466), .QN(n17124) );
  NOR2X0 U17427 ( .IN1(n4368), .IN2(n15466), .QN(n17126) );
  NOR2X0 U17428 ( .IN1(n17127), .IN2(n10780), .QN(n13268) );
  NOR2X0 U17429 ( .IN1(n13273), .IN2(n17128), .QN(g25042) );
  NAND2X0 U17430 ( .IN1(n17129), .IN2(n17130), .QN(n17128) );
  NAND2X0 U17431 ( .IN1(n10021), .IN2(n3894), .QN(n17130) );
  INVX0 U17432 ( .INP(n17131), .ZN(n3894) );
  NAND2X0 U17433 ( .IN1(n17131), .IN2(g780), .QN(n17129) );
  NOR2X0 U17434 ( .IN1(n10321), .IN2(n15466), .QN(n17131) );
  INVX0 U17435 ( .INP(n13956), .ZN(n13273) );
  NAND2X0 U17436 ( .IN1(n17132), .IN2(n15466), .QN(n13956) );
  NOR2X0 U17437 ( .IN1(n13278), .IN2(n17133), .QN(g25027) );
  NAND2X0 U17438 ( .IN1(n17134), .IN2(n17135), .QN(n17133) );
  NAND2X0 U17439 ( .IN1(n10025), .IN2(n3897), .QN(n17135) );
  INVX0 U17440 ( .INP(n17136), .ZN(n3897) );
  NAND2X0 U17441 ( .IN1(n17136), .IN2(g92), .QN(n17134) );
  NOR2X0 U17442 ( .IN1(n4369), .IN2(n15466), .QN(n17136) );
  NOR2X0 U17443 ( .IN1(n17137), .IN2(n10780), .QN(n13278) );
  INVX0 U17444 ( .INP(n15466), .ZN(n10780) );
  NOR2X0 U17445 ( .IN1(n17138), .IN2(n17139), .QN(n15466) );
  NAND2X0 U17446 ( .IN1(n4305), .IN2(n17140), .QN(n17139) );
  NOR2X0 U17447 ( .IN1(g2900), .IN2(g2892), .QN(n17140) );
  NAND2X0 U17448 ( .IN1(n4355), .IN2(n4431), .QN(n17138) );
  NAND2X0 U17449 ( .IN1(n3700), .IN2(n17141), .QN(g24734) );
  NAND2X0 U17450 ( .IN1(n14900), .IN2(DFF_146_n1), .QN(n17141) );
  NOR2X0 U17451 ( .IN1(n16222), .IN2(n14879), .QN(n14900) );
  INVX0 U17452 ( .INP(n3705), .ZN(n14879) );
  INVX0 U17453 ( .INP(n3940), .ZN(n16222) );
  NAND2X0 U17454 ( .IN1(n17142), .IN2(n17143), .QN(g24557) );
  NAND2X0 U17455 ( .IN1(n11916), .IN2(n11726), .QN(n17143) );
  INVX0 U17456 ( .INP(n17144), .ZN(n17142) );
  NOR2X0 U17457 ( .IN1(g2624), .IN2(n9689), .QN(n17144) );
  NAND2X0 U17458 ( .IN1(n17145), .IN2(n17146), .QN(g24548) );
  INVX0 U17459 ( .INP(n17147), .ZN(n17146) );
  NOR2X0 U17460 ( .IN1(g7390), .IN2(n9690), .QN(n17147) );
  NAND2X0 U17461 ( .IN1(n17148), .IN2(g7390), .QN(n17145) );
  NAND2X0 U17462 ( .IN1(n17149), .IN2(n17150), .QN(g24547) );
  NAND2X0 U17463 ( .IN1(n11916), .IN2(n14267), .QN(n17150) );
  NOR2X0 U17464 ( .IN1(n14200), .IN2(n4299), .QN(n11916) );
  INVX0 U17465 ( .INP(n17151), .ZN(n17149) );
  NOR2X0 U17466 ( .IN1(g2624), .IN2(n9702), .QN(n17151) );
  NAND2X0 U17467 ( .IN1(n17152), .IN2(n17153), .QN(g24545) );
  NAND2X0 U17468 ( .IN1(n11921), .IN2(n14330), .QN(n17153) );
  INVX0 U17469 ( .INP(n17154), .ZN(n17152) );
  NOR2X0 U17470 ( .IN1(g1930), .IN2(n9692), .QN(n17154) );
  NAND2X0 U17471 ( .IN1(n17155), .IN2(n17156), .QN(g24538) );
  NAND2X0 U17472 ( .IN1(n17148), .IN2(g7302), .QN(n17156) );
  NOR2X0 U17473 ( .IN1(n14200), .IN2(n17157), .QN(n17148) );
  INVX0 U17474 ( .INP(n11726), .ZN(n17157) );
  NAND2X0 U17475 ( .IN1(n17158), .IN2(n17159), .QN(n11726) );
  NOR2X0 U17476 ( .IN1(n17160), .IN2(n17161), .QN(n17159) );
  NOR2X0 U17477 ( .IN1(n9689), .IN2(n4299), .QN(n17161) );
  NOR2X0 U17478 ( .IN1(n9688), .IN2(n17162), .QN(n17160) );
  NAND2X0 U17479 ( .IN1(n11918), .IN2(g185), .QN(n17162) );
  NAND2X0 U17480 ( .IN1(n17163), .IN2(n17164), .QN(n11918) );
  NAND2X0 U17481 ( .IN1(g7390), .IN2(g2641), .QN(n17164) );
  NOR2X0 U17482 ( .IN1(n17165), .IN2(n17166), .QN(n17163) );
  NOR2X0 U17483 ( .IN1(n9809), .IN2(n4314), .QN(n17166) );
  NOR2X0 U17484 ( .IN1(n9810), .IN2(n4299), .QN(n17165) );
  NOR2X0 U17485 ( .IN1(n17167), .IN2(n17168), .QN(n17158) );
  NOR2X0 U17486 ( .IN1(n9690), .IN2(n4370), .QN(n17168) );
  NOR2X0 U17487 ( .IN1(n9687), .IN2(n4314), .QN(n17167) );
  INVX0 U17488 ( .INP(n17169), .ZN(n17155) );
  NOR2X0 U17489 ( .IN1(n13147), .IN2(n9687), .QN(n17169) );
  NAND2X0 U17490 ( .IN1(n17170), .IN2(n17171), .QN(g24537) );
  INVX0 U17491 ( .INP(n17172), .ZN(n17171) );
  NOR2X0 U17492 ( .IN1(g7390), .IN2(n9703), .QN(n17172) );
  NAND2X0 U17493 ( .IN1(n17173), .IN2(g7390), .QN(n17170) );
  NAND2X0 U17494 ( .IN1(n17174), .IN2(n17175), .QN(g24535) );
  INVX0 U17495 ( .INP(n17176), .ZN(n17175) );
  NOR2X0 U17496 ( .IN1(g7194), .IN2(n9693), .QN(n17176) );
  NAND2X0 U17497 ( .IN1(n17177), .IN2(g7194), .QN(n17174) );
  NAND2X0 U17498 ( .IN1(n17178), .IN2(n17179), .QN(g24534) );
  NAND2X0 U17499 ( .IN1(n11921), .IN2(n14399), .QN(n17179) );
  NOR2X0 U17500 ( .IN1(n14200), .IN2(n4366), .QN(n11921) );
  INVX0 U17501 ( .INP(n17180), .ZN(n17178) );
  NOR2X0 U17502 ( .IN1(g1930), .IN2(n9705), .QN(n17180) );
  NAND2X0 U17503 ( .IN1(n17181), .IN2(n17182), .QN(g24532) );
  NAND2X0 U17504 ( .IN1(n10715), .IN2(n14458), .QN(n17182) );
  INVX0 U17505 ( .INP(n17183), .ZN(n17181) );
  NOR2X0 U17506 ( .IN1(g1236), .IN2(n9696), .QN(n17183) );
  NAND2X0 U17507 ( .IN1(n17184), .IN2(n17185), .QN(g24527) );
  INVX0 U17508 ( .INP(n17186), .ZN(n17185) );
  NOR2X0 U17509 ( .IN1(n13147), .IN2(n9701), .QN(n17186) );
  NAND2X0 U17510 ( .IN1(n17173), .IN2(n13147), .QN(n17184) );
  NOR2X0 U17511 ( .IN1(n14200), .IN2(n14268), .QN(n17173) );
  INVX0 U17512 ( .INP(n14267), .ZN(n14268) );
  NAND2X0 U17513 ( .IN1(n17187), .IN2(n17188), .QN(n14267) );
  NOR2X0 U17514 ( .IN1(n17189), .IN2(n17190), .QN(n17188) );
  NOR2X0 U17515 ( .IN1(n9701), .IN2(n13148), .QN(n17190) );
  NOR2X0 U17516 ( .IN1(n1684), .IN2(n17191), .QN(n17189) );
  NAND2X0 U17517 ( .IN1(g185), .IN2(g2598), .QN(n17191) );
  INVX0 U17518 ( .INP(n17192), .ZN(n1684) );
  NAND2X0 U17519 ( .IN1(n17193), .IN2(n17194), .QN(n17192) );
  NAND2X0 U17520 ( .IN1(g7390), .IN2(g2645), .QN(n17194) );
  NOR2X0 U17521 ( .IN1(n17195), .IN2(n17196), .QN(n17193) );
  NOR2X0 U17522 ( .IN1(n9812), .IN2(n4299), .QN(n17196) );
  NOR2X0 U17523 ( .IN1(n9811), .IN2(n13148), .QN(n17195) );
  NOR2X0 U17524 ( .IN1(n17197), .IN2(n17198), .QN(n17187) );
  NOR2X0 U17525 ( .IN1(n9703), .IN2(n4370), .QN(n17198) );
  NOR2X0 U17526 ( .IN1(n9702), .IN2(n4299), .QN(n17197) );
  NAND2X0 U17527 ( .IN1(n17199), .IN2(n17200), .QN(g24525) );
  NAND2X0 U17528 ( .IN1(n17177), .IN2(g7052), .QN(n17200) );
  NOR2X0 U17529 ( .IN1(n14200), .IN2(n17201), .QN(n17177) );
  INVX0 U17530 ( .INP(n14330), .ZN(n17201) );
  NAND2X0 U17531 ( .IN1(n17202), .IN2(n17203), .QN(n14330) );
  NOR2X0 U17532 ( .IN1(n17204), .IN2(n17205), .QN(n17203) );
  NOR2X0 U17533 ( .IN1(n9691), .IN2(n4296), .QN(n17205) );
  NOR2X0 U17534 ( .IN1(n1330), .IN2(n17206), .QN(n17204) );
  NAND2X0 U17535 ( .IN1(g185), .IN2(g1922), .QN(n17206) );
  INVX0 U17536 ( .INP(n17207), .ZN(n1330) );
  NAND2X0 U17537 ( .IN1(n17208), .IN2(n17209), .QN(n17207) );
  NAND2X0 U17538 ( .IN1(g1930), .IN2(g1870), .QN(n17209) );
  NOR2X0 U17539 ( .IN1(n17210), .IN2(n17211), .QN(n17208) );
  NOR2X0 U17540 ( .IN1(n18866), .IN2(n4315), .QN(n17211) );
  NOR2X0 U17541 ( .IN1(n9813), .IN2(n4296), .QN(n17210) );
  NOR2X0 U17542 ( .IN1(n17212), .IN2(n17213), .QN(n17202) );
  NOR2X0 U17543 ( .IN1(n9692), .IN2(n4366), .QN(n17213) );
  NOR2X0 U17544 ( .IN1(n9693), .IN2(n4315), .QN(n17212) );
  INVX0 U17545 ( .INP(n17214), .ZN(n17199) );
  NOR2X0 U17546 ( .IN1(n14321), .IN2(n9691), .QN(n17214) );
  NAND2X0 U17547 ( .IN1(n17215), .IN2(n17216), .QN(g24524) );
  INVX0 U17548 ( .INP(n17217), .ZN(n17216) );
  NOR2X0 U17549 ( .IN1(g7194), .IN2(n9706), .QN(n17217) );
  NAND2X0 U17550 ( .IN1(n17218), .IN2(g7194), .QN(n17215) );
  NAND2X0 U17551 ( .IN1(n17219), .IN2(n17220), .QN(g24522) );
  INVX0 U17552 ( .INP(n17221), .ZN(n17220) );
  NOR2X0 U17553 ( .IN1(g6944), .IN2(n9697), .QN(n17221) );
  NAND2X0 U17554 ( .IN1(n17222), .IN2(g6944), .QN(n17219) );
  NAND2X0 U17555 ( .IN1(n17223), .IN2(n17224), .QN(g24521) );
  NAND2X0 U17556 ( .IN1(n10715), .IN2(n14522), .QN(n17224) );
  NOR2X0 U17557 ( .IN1(n14200), .IN2(n4300), .QN(n10715) );
  INVX0 U17558 ( .INP(n17225), .ZN(n17223) );
  NOR2X0 U17559 ( .IN1(g1236), .IN2(n9708), .QN(n17225) );
  NAND2X0 U17560 ( .IN1(n17226), .IN2(n17227), .QN(g24519) );
  NAND2X0 U17561 ( .IN1(n10720), .IN2(n14583), .QN(n17227) );
  INVX0 U17562 ( .INP(n17228), .ZN(n17226) );
  NOR2X0 U17563 ( .IN1(g550), .IN2(n9699), .QN(n17228) );
  NAND2X0 U17564 ( .IN1(n17229), .IN2(n17230), .QN(g24513) );
  INVX0 U17565 ( .INP(n17231), .ZN(n17230) );
  NOR2X0 U17566 ( .IN1(n14321), .IN2(n9704), .QN(n17231) );
  NAND2X0 U17567 ( .IN1(n17218), .IN2(n14321), .QN(n17229) );
  NOR2X0 U17568 ( .IN1(n14200), .IN2(n17232), .QN(n17218) );
  INVX0 U17569 ( .INP(n14399), .ZN(n17232) );
  NAND2X0 U17570 ( .IN1(n17233), .IN2(n17234), .QN(n14399) );
  NOR2X0 U17571 ( .IN1(n17235), .IN2(n17236), .QN(n17234) );
  NOR2X0 U17572 ( .IN1(n9704), .IN2(n17237), .QN(n17236) );
  NOR2X0 U17573 ( .IN1(n1333), .IN2(n17238), .QN(n17235) );
  NAND2X0 U17574 ( .IN1(g185), .IN2(g1904), .QN(n17238) );
  INVX0 U17575 ( .INP(n17239), .ZN(n1333) );
  NAND2X0 U17576 ( .IN1(n17240), .IN2(n17241), .QN(n17239) );
  NAND2X0 U17577 ( .IN1(g1930), .IN2(g1953), .QN(n17241) );
  NOR2X0 U17578 ( .IN1(n17242), .IN2(n17243), .QN(n17240) );
  NOR2X0 U17579 ( .IN1(n18864), .IN2(n4315), .QN(n17243) );
  NOR2X0 U17580 ( .IN1(n9815), .IN2(n17237), .QN(n17242) );
  NOR2X0 U17581 ( .IN1(n17244), .IN2(n17245), .QN(n17233) );
  NOR2X0 U17582 ( .IN1(n9705), .IN2(n4366), .QN(n17245) );
  NOR2X0 U17583 ( .IN1(n9706), .IN2(n4315), .QN(n17244) );
  NAND2X0 U17584 ( .IN1(n17246), .IN2(n17247), .QN(g24511) );
  NAND2X0 U17585 ( .IN1(n17222), .IN2(g6750), .QN(n17247) );
  NOR2X0 U17586 ( .IN1(n14200), .IN2(n17248), .QN(n17222) );
  INVX0 U17587 ( .INP(n14458), .ZN(n17248) );
  NAND2X0 U17588 ( .IN1(n17249), .IN2(n17250), .QN(n14458) );
  NOR2X0 U17589 ( .IN1(n17251), .IN2(n17252), .QN(n17250) );
  NOR2X0 U17590 ( .IN1(n9696), .IN2(n4300), .QN(n17252) );
  NOR2X0 U17591 ( .IN1(n9695), .IN2(n17253), .QN(n17251) );
  NAND2X0 U17592 ( .IN1(n10717), .IN2(g185), .QN(n17253) );
  NAND2X0 U17593 ( .IN1(n17254), .IN2(n17255), .QN(n10717) );
  NAND2X0 U17594 ( .IN1(g6944), .IN2(g1253), .QN(n17255) );
  NOR2X0 U17595 ( .IN1(n17256), .IN2(n17257), .QN(n17254) );
  NOR2X0 U17596 ( .IN1(n9818), .IN2(n4300), .QN(n17257) );
  NOR2X0 U17597 ( .IN1(n9817), .IN2(n17258), .QN(n17256) );
  NOR2X0 U17598 ( .IN1(n17259), .IN2(n17260), .QN(n17249) );
  NOR2X0 U17599 ( .IN1(n9694), .IN2(n4371), .QN(n17260) );
  NOR2X0 U17600 ( .IN1(n9697), .IN2(n4316), .QN(n17259) );
  INVX0 U17601 ( .INP(n17261), .ZN(n17246) );
  NOR2X0 U17602 ( .IN1(n14180), .IN2(n9694), .QN(n17261) );
  NAND2X0 U17603 ( .IN1(n17262), .IN2(n17263), .QN(g24510) );
  INVX0 U17604 ( .INP(n17264), .ZN(n17263) );
  NOR2X0 U17605 ( .IN1(g6944), .IN2(n9709), .QN(n17264) );
  NAND2X0 U17606 ( .IN1(n17265), .IN2(g6944), .QN(n17262) );
  NAND2X0 U17607 ( .IN1(n17266), .IN2(n17267), .QN(g24508) );
  INVX0 U17608 ( .INP(n17268), .ZN(n17267) );
  NOR2X0 U17609 ( .IN1(g6642), .IN2(n9700), .QN(n17268) );
  NAND2X0 U17610 ( .IN1(n17269), .IN2(g6642), .QN(n17266) );
  NAND2X0 U17611 ( .IN1(n17270), .IN2(n17271), .QN(g24507) );
  NAND2X0 U17612 ( .IN1(n10720), .IN2(n14641), .QN(n17271) );
  NOR2X0 U17613 ( .IN1(n14200), .IN2(n4313), .QN(n10720) );
  INVX0 U17614 ( .INP(n17272), .ZN(n17270) );
  NOR2X0 U17615 ( .IN1(g550), .IN2(n9711), .QN(n17272) );
  NAND2X0 U17616 ( .IN1(n17273), .IN2(n17274), .QN(g24501) );
  INVX0 U17617 ( .INP(n17275), .ZN(n17274) );
  NOR2X0 U17618 ( .IN1(n14180), .IN2(n9707), .QN(n17275) );
  NAND2X0 U17619 ( .IN1(n17265), .IN2(n14180), .QN(n17273) );
  NOR2X0 U17620 ( .IN1(n14200), .IN2(n17276), .QN(n17265) );
  INVX0 U17621 ( .INP(n14522), .ZN(n17276) );
  NAND2X0 U17622 ( .IN1(n17277), .IN2(n17278), .QN(n14522) );
  NOR2X0 U17623 ( .IN1(n17279), .IN2(n17280), .QN(n17278) );
  NOR2X0 U17624 ( .IN1(n9707), .IN2(n17258), .QN(n17280) );
  NOR2X0 U17625 ( .IN1(n982), .IN2(n17281), .QN(n17279) );
  NAND2X0 U17626 ( .IN1(g185), .IN2(g1210), .QN(n17281) );
  INVX0 U17627 ( .INP(n17282), .ZN(n982) );
  NAND2X0 U17628 ( .IN1(n17283), .IN2(n17284), .QN(n17282) );
  NAND2X0 U17629 ( .IN1(n14180), .IN2(g1255), .QN(n17284) );
  NOR2X0 U17630 ( .IN1(n17285), .IN2(n17286), .QN(n17283) );
  NOR2X0 U17631 ( .IN1(n18865), .IN2(n4316), .QN(n17286) );
  NOR2X0 U17632 ( .IN1(n9820), .IN2(n4300), .QN(n17285) );
  NOR2X0 U17633 ( .IN1(n17287), .IN2(n17288), .QN(n17277) );
  NOR2X0 U17634 ( .IN1(n9709), .IN2(n4316), .QN(n17288) );
  NOR2X0 U17635 ( .IN1(n9708), .IN2(n4300), .QN(n17287) );
  NAND2X0 U17636 ( .IN1(n17289), .IN2(n17290), .QN(g24499) );
  NAND2X0 U17637 ( .IN1(n17269), .IN2(g6485), .QN(n17290) );
  NOR2X0 U17638 ( .IN1(n14200), .IN2(n17291), .QN(n17269) );
  INVX0 U17639 ( .INP(n14583), .ZN(n17291) );
  NAND2X0 U17640 ( .IN1(n17292), .IN2(n17293), .QN(n14583) );
  NOR2X0 U17641 ( .IN1(n17294), .IN2(n17295), .QN(n17293) );
  NOR2X0 U17642 ( .IN1(n9698), .IN2(n17296), .QN(n17295) );
  NOR2X0 U17643 ( .IN1(n621), .IN2(n17297), .QN(n17294) );
  NAND2X0 U17644 ( .IN1(g185), .IN2(g542), .QN(n17297) );
  INVX0 U17645 ( .INP(n17298), .ZN(n621) );
  NAND2X0 U17646 ( .IN1(n17299), .IN2(n17300), .QN(n17298) );
  NAND2X0 U17647 ( .IN1(g6642), .IN2(g567), .QN(n17300) );
  NOR2X0 U17648 ( .IN1(n17301), .IN2(n17302), .QN(n17299) );
  NOR2X0 U17649 ( .IN1(n9806), .IN2(n4313), .QN(n17302) );
  NOR2X0 U17650 ( .IN1(n9805), .IN2(n4298), .QN(n17301) );
  NOR2X0 U17651 ( .IN1(n17303), .IN2(n17304), .QN(n17292) );
  NOR2X0 U17652 ( .IN1(n9700), .IN2(n4372), .QN(n17304) );
  NOR2X0 U17653 ( .IN1(n9699), .IN2(n4313), .QN(n17303) );
  INVX0 U17654 ( .INP(n17305), .ZN(n17289) );
  NOR2X0 U17655 ( .IN1(n14574), .IN2(n9698), .QN(n17305) );
  NAND2X0 U17656 ( .IN1(n17306), .IN2(n17307), .QN(g24498) );
  INVX0 U17657 ( .INP(n17308), .ZN(n17307) );
  NOR2X0 U17658 ( .IN1(g6642), .IN2(n9712), .QN(n17308) );
  NAND2X0 U17659 ( .IN1(n17309), .IN2(g6642), .QN(n17306) );
  NAND2X0 U17660 ( .IN1(n17310), .IN2(n17311), .QN(g24491) );
  INVX0 U17661 ( .INP(n17312), .ZN(n17311) );
  NOR2X0 U17662 ( .IN1(n14574), .IN2(n9710), .QN(n17312) );
  NAND2X0 U17663 ( .IN1(n17309), .IN2(n14574), .QN(n17310) );
  NOR2X0 U17664 ( .IN1(n14200), .IN2(n17313), .QN(n17309) );
  INVX0 U17665 ( .INP(n14641), .ZN(n17313) );
  NAND2X0 U17666 ( .IN1(n17314), .IN2(n17315), .QN(n14641) );
  NOR2X0 U17667 ( .IN1(n17316), .IN2(n17317), .QN(n17315) );
  NOR2X0 U17668 ( .IN1(n9710), .IN2(n4298), .QN(n17317) );
  NOR2X0 U17669 ( .IN1(n622), .IN2(n17318), .QN(n17316) );
  NAND2X0 U17670 ( .IN1(g185), .IN2(g524), .QN(n17318) );
  INVX0 U17671 ( .INP(n17319), .ZN(n622) );
  NAND2X0 U17672 ( .IN1(n17320), .IN2(n17321), .QN(n17319) );
  NAND2X0 U17673 ( .IN1(g6642), .IN2(g571), .QN(n17321) );
  NOR2X0 U17674 ( .IN1(n17322), .IN2(n17323), .QN(n17320) );
  NOR2X0 U17675 ( .IN1(n9808), .IN2(n4313), .QN(n17323) );
  NOR2X0 U17676 ( .IN1(n9807), .IN2(n17296), .QN(n17322) );
  NOR2X0 U17677 ( .IN1(n17324), .IN2(n17325), .QN(n17314) );
  NOR2X0 U17678 ( .IN1(n9712), .IN2(n4372), .QN(n17325) );
  NOR2X0 U17679 ( .IN1(n9711), .IN2(n4313), .QN(n17324) );
  INVX0 U17680 ( .INP(n14201), .ZN(n14200) );
  NAND2X0 U17681 ( .IN1(n17326), .IN2(n17327), .QN(n14201) );
  NOR2X0 U17682 ( .IN1(n17328), .IN2(n17329), .QN(n17327) );
  NAND2X0 U17683 ( .IN1(g3028), .IN2(g3018), .QN(n17329) );
  NOR2X0 U17684 ( .IN1(g3036), .IN2(g3032), .QN(n17326) );
  NOR2X0 U17685 ( .IN1(n17330), .IN2(n17099), .QN(g24476) );
  NAND2X0 U17686 ( .IN1(n11001), .IN2(n17102), .QN(n17099) );
  NAND2X0 U17687 ( .IN1(n17331), .IN2(n17332), .QN(n17102) );
  NOR2X0 U17688 ( .IN1(n4479), .IN2(n4349), .QN(n17331) );
  NOR2X0 U17689 ( .IN1(n17333), .IN2(g2924), .QN(n17330) );
  NOR2X0 U17690 ( .IN1(n4479), .IN2(n11004), .QN(n17333) );
  NOR2X0 U17691 ( .IN1(n10998), .IN2(n17334), .QN(g24473) );
  NAND2X0 U17692 ( .IN1(n18), .IN2(n17335), .QN(n17334) );
  NAND2X0 U17693 ( .IN1(n10079), .IN2(n17336), .QN(n17335) );
  INVX0 U17694 ( .INP(n17337), .ZN(n17336) );
  NAND2X0 U17695 ( .IN1(n17337), .IN2(g2892), .QN(n18) );
  NOR2X0 U17696 ( .IN1(n17087), .IN2(n17338), .QN(g24446) );
  NAND2X0 U17697 ( .IN1(n17091), .IN2(n17339), .QN(n17338) );
  INVX0 U17698 ( .INP(n4101), .ZN(n17339) );
  INVX0 U17699 ( .INP(n17092), .ZN(n17091) );
  NOR2X0 U17700 ( .IN1(n4102), .IN2(n4480), .QN(n17092) );
  NOR2X0 U17701 ( .IN1(n15740), .IN2(n17340), .QN(g24445) );
  NAND2X0 U17702 ( .IN1(n17341), .IN2(n17342), .QN(n17340) );
  NAND2X0 U17703 ( .IN1(n10304), .IN2(n4066), .QN(n17342) );
  INVX0 U17704 ( .INP(n17343), .ZN(n17341) );
  NOR2X0 U17705 ( .IN1(n4066), .IN2(n10304), .QN(n17343) );
  NOR2X0 U17706 ( .IN1(n17344), .IN2(n17345), .QN(g24438) );
  NAND2X0 U17707 ( .IN1(n15756), .IN2(n14826), .QN(n17345) );
  NAND2X0 U17708 ( .IN1(n17346), .IN2(n17347), .QN(n15756) );
  NOR2X0 U17709 ( .IN1(n4419), .IN2(n4408), .QN(n17346) );
  NOR2X0 U17710 ( .IN1(n17348), .IN2(g2720), .QN(n17344) );
  NOR2X0 U17711 ( .IN1(n4419), .IN2(n17349), .QN(n17348) );
  NOR2X0 U17712 ( .IN1(n17350), .IN2(n17351), .QN(g24434) );
  NAND2X0 U17713 ( .IN1(n15774), .IN2(n14703), .QN(n17351) );
  NAND2X0 U17714 ( .IN1(n17352), .IN2(n17353), .QN(n15774) );
  NOR2X0 U17715 ( .IN1(n4420), .IN2(n4410), .QN(n17352) );
  NOR2X0 U17716 ( .IN1(n17354), .IN2(g2026), .QN(n17350) );
  NOR2X0 U17717 ( .IN1(n4420), .IN2(n17355), .QN(n17354) );
  NOR2X0 U17718 ( .IN1(n17356), .IN2(n17357), .QN(g24430) );
  NAND2X0 U17719 ( .IN1(n15895), .IN2(n14834), .QN(n17357) );
  NAND2X0 U17720 ( .IN1(n17358), .IN2(n17359), .QN(n15895) );
  NOR2X0 U17721 ( .IN1(n4421), .IN2(n4412), .QN(n17358) );
  NOR2X0 U17722 ( .IN1(n17360), .IN2(g1332), .QN(n17356) );
  NOR2X0 U17723 ( .IN1(n4421), .IN2(n17361), .QN(n17360) );
  NOR2X0 U17724 ( .IN1(n17362), .IN2(n17363), .QN(g24426) );
  NAND2X0 U17725 ( .IN1(n16016), .IN2(n14712), .QN(n17363) );
  NAND2X0 U17726 ( .IN1(n17364), .IN2(n17365), .QN(n16016) );
  NOR2X0 U17727 ( .IN1(n4422), .IN2(n4414), .QN(n17364) );
  NOR2X0 U17728 ( .IN1(n17366), .IN2(g646), .QN(n17362) );
  NOR2X0 U17729 ( .IN1(n4422), .IN2(n17367), .QN(n17366) );
  NAND2X0 U17730 ( .IN1(n17368), .IN2(n17369), .QN(g24250) );
  NAND2X0 U17731 ( .IN1(n4463), .IN2(g2546), .QN(n17369) );
  NAND2X0 U17732 ( .IN1(n12926), .IN2(g2560), .QN(n17368) );
  NAND2X0 U17733 ( .IN1(n17370), .IN2(n17371), .QN(g24243) );
  NAND2X0 U17734 ( .IN1(n4464), .IN2(g1852), .QN(n17371) );
  NAND2X0 U17735 ( .IN1(n12975), .IN2(g1866), .QN(n17370) );
  NAND2X0 U17736 ( .IN1(n17372), .IN2(n17373), .QN(g24238) );
  INVX0 U17737 ( .INP(n17374), .ZN(n17373) );
  NOR2X0 U17738 ( .IN1(g2560), .IN2(n10043), .QN(n17374) );
  NAND2X0 U17739 ( .IN1(n12932), .IN2(g2560), .QN(n17372) );
  NAND2X0 U17740 ( .IN1(n17375), .IN2(n17376), .QN(g24237) );
  NAND2X0 U17741 ( .IN1(n4455), .IN2(g2543), .QN(n17376) );
  NAND2X0 U17742 ( .IN1(n12926), .IN2(g8167), .QN(n17375) );
  NAND2X0 U17743 ( .IN1(n17377), .IN2(n17378), .QN(g24235) );
  NAND2X0 U17744 ( .IN1(n4465), .IN2(g1158), .QN(n17378) );
  NAND2X0 U17745 ( .IN1(n13036), .IN2(g1172), .QN(n17377) );
  NAND2X0 U17746 ( .IN1(n17379), .IN2(n17380), .QN(g24231) );
  INVX0 U17747 ( .INP(n17381), .ZN(n17380) );
  NOR2X0 U17748 ( .IN1(g1866), .IN2(n10052), .QN(n17381) );
  NAND2X0 U17749 ( .IN1(n13234), .IN2(g1866), .QN(n17379) );
  NAND2X0 U17750 ( .IN1(n17382), .IN2(n17383), .QN(g24230) );
  NAND2X0 U17751 ( .IN1(n4457), .IN2(g1849), .QN(n17383) );
  NAND2X0 U17752 ( .IN1(n12975), .IN2(g8082), .QN(n17382) );
  NAND2X0 U17753 ( .IN1(n17384), .IN2(n17385), .QN(g24228) );
  NAND2X0 U17754 ( .IN1(n4466), .IN2(g471), .QN(n17385) );
  NAND2X0 U17755 ( .IN1(n13109), .IN2(g485), .QN(n17384) );
  NAND2X0 U17756 ( .IN1(n17386), .IN2(n17387), .QN(g24226) );
  NAND2X0 U17757 ( .IN1(n4455), .IN2(g2553), .QN(n17387) );
  NAND2X0 U17758 ( .IN1(n12932), .IN2(g8167), .QN(n17386) );
  NAND2X0 U17759 ( .IN1(n17388), .IN2(n17389), .QN(g24225) );
  NAND2X0 U17760 ( .IN1(n4456), .IN2(g2540), .QN(n17389) );
  NAND2X0 U17761 ( .IN1(n12926), .IN2(g8087), .QN(n17388) );
  NOR2X0 U17762 ( .IN1(n12476), .IN2(n12478), .QN(n12926) );
  NAND2X0 U17763 ( .IN1(n12491), .IN2(n12498), .QN(n12476) );
  NAND2X0 U17764 ( .IN1(n17390), .IN2(n17391), .QN(g24223) );
  INVX0 U17765 ( .INP(n17392), .ZN(n17391) );
  NOR2X0 U17766 ( .IN1(g1172), .IN2(n10060), .QN(n17392) );
  NAND2X0 U17767 ( .IN1(n13065), .IN2(g1172), .QN(n17390) );
  NAND2X0 U17768 ( .IN1(n17393), .IN2(n17394), .QN(g24222) );
  NAND2X0 U17769 ( .IN1(n4459), .IN2(g1155), .QN(n17394) );
  NAND2X0 U17770 ( .IN1(n13036), .IN2(g8007), .QN(n17393) );
  NAND2X0 U17771 ( .IN1(n17395), .IN2(n17396), .QN(g24219) );
  NAND2X0 U17772 ( .IN1(n4457), .IN2(g1859), .QN(n17396) );
  NAND2X0 U17773 ( .IN1(n13234), .IN2(g8082), .QN(n17395) );
  NAND2X0 U17774 ( .IN1(n17397), .IN2(n17398), .QN(g24218) );
  NAND2X0 U17775 ( .IN1(n4458), .IN2(g1846), .QN(n17398) );
  NAND2X0 U17776 ( .IN1(n12975), .IN2(g8012), .QN(n17397) );
  NOR2X0 U17777 ( .IN1(n11962), .IN2(n11964), .QN(n12975) );
  NAND2X0 U17778 ( .IN1(n11978), .IN2(n11985), .QN(n11962) );
  NAND2X0 U17779 ( .IN1(n17399), .IN2(n17400), .QN(g24216) );
  INVX0 U17780 ( .INP(n17401), .ZN(n17400) );
  NOR2X0 U17781 ( .IN1(g485), .IN2(n10069), .QN(n17401) );
  NAND2X0 U17782 ( .IN1(n13260), .IN2(g485), .QN(n17399) );
  NAND2X0 U17783 ( .IN1(n17402), .IN2(n17403), .QN(g24215) );
  NAND2X0 U17784 ( .IN1(n13109), .IN2(g7956), .QN(n17403) );
  NAND2X0 U17785 ( .IN1(test_so24), .IN2(n4461), .QN(n17402) );
  NAND2X0 U17786 ( .IN1(n17404), .IN2(n17405), .QN(g24214) );
  INVX0 U17787 ( .INP(n17406), .ZN(n17405) );
  NOR2X0 U17788 ( .IN1(g8087), .IN2(n10042), .QN(n17406) );
  NAND2X0 U17789 ( .IN1(n12932), .IN2(g8087), .QN(n17404) );
  NOR2X0 U17790 ( .IN1(n17407), .IN2(n12470), .QN(n12932) );
  NAND2X0 U17791 ( .IN1(n12487), .IN2(n12478), .QN(n17407) );
  NAND2X0 U17792 ( .IN1(n17408), .IN2(n17409), .QN(g24213) );
  NAND2X0 U17793 ( .IN1(n4459), .IN2(g1165), .QN(n17409) );
  NAND2X0 U17794 ( .IN1(n13065), .IN2(g8007), .QN(n17408) );
  NAND2X0 U17795 ( .IN1(n17410), .IN2(n17411), .QN(g24212) );
  NAND2X0 U17796 ( .IN1(n4460), .IN2(g1152), .QN(n17411) );
  NAND2X0 U17797 ( .IN1(n13036), .IN2(g7961), .QN(n17410) );
  INVX0 U17798 ( .INP(n10804), .ZN(n13036) );
  NAND2X0 U17799 ( .IN1(n17412), .IN2(n11766), .QN(n10804) );
  NOR2X0 U17800 ( .IN1(n11759), .IN2(n11753), .QN(n17412) );
  NAND2X0 U17801 ( .IN1(n17413), .IN2(n17414), .QN(g24209) );
  NAND2X0 U17802 ( .IN1(n4463), .IN2(g2536), .QN(n17414) );
  NAND2X0 U17803 ( .IN1(n15268), .IN2(g2560), .QN(n17413) );
  NAND2X0 U17804 ( .IN1(n17415), .IN2(n17416), .QN(g24208) );
  INVX0 U17805 ( .INP(n17417), .ZN(n17416) );
  NOR2X0 U17806 ( .IN1(g8012), .IN2(n10051), .QN(n17417) );
  NAND2X0 U17807 ( .IN1(n13234), .IN2(g8012), .QN(n17415) );
  INVX0 U17808 ( .INP(n13609), .ZN(n13234) );
  NAND2X0 U17809 ( .IN1(n17418), .IN2(n11978), .QN(n13609) );
  NOR2X0 U17810 ( .IN1(n11985), .IN2(n11961), .QN(n17418) );
  NAND2X0 U17811 ( .IN1(n17419), .IN2(n17420), .QN(g24207) );
  NAND2X0 U17812 ( .IN1(n4461), .IN2(g478), .QN(n17420) );
  NAND2X0 U17813 ( .IN1(n13260), .IN2(g7956), .QN(n17419) );
  NAND2X0 U17814 ( .IN1(n17421), .IN2(n17422), .QN(g24206) );
  NAND2X0 U17815 ( .IN1(g465), .IN2(n10328), .QN(n17422) );
  NAND2X0 U17816 ( .IN1(test_so23), .IN2(n13109), .QN(n17421) );
  NOR2X0 U17817 ( .IN1(n12012), .IN2(n12014), .QN(n13109) );
  NAND2X0 U17818 ( .IN1(n12028), .IN2(n12035), .QN(n12012) );
  NAND2X0 U17819 ( .IN1(n17423), .IN2(n17424), .QN(g24182) );
  NAND2X0 U17820 ( .IN1(n4464), .IN2(g1842), .QN(n17424) );
  NAND2X0 U17821 ( .IN1(n15378), .IN2(g1866), .QN(n17423) );
  NAND2X0 U17822 ( .IN1(n17425), .IN2(n17426), .QN(g24181) );
  INVX0 U17823 ( .INP(n17427), .ZN(n17426) );
  NOR2X0 U17824 ( .IN1(g7961), .IN2(n10059), .QN(n17427) );
  NAND2X0 U17825 ( .IN1(n13065), .IN2(g7961), .QN(n17425) );
  INVX0 U17826 ( .INP(n13749), .ZN(n13065) );
  NAND2X0 U17827 ( .IN1(n17428), .IN2(n11766), .QN(n13749) );
  NOR2X0 U17828 ( .IN1(n11756), .IN2(n11787), .QN(n17428) );
  NAND2X0 U17829 ( .IN1(n17429), .IN2(n17430), .QN(g24179) );
  NAND2X0 U17830 ( .IN1(n4465), .IN2(g1148), .QN(n17430) );
  NAND2X0 U17831 ( .IN1(n17431), .IN2(g1172), .QN(n17429) );
  NAND2X0 U17832 ( .IN1(n17432), .IN2(n17433), .QN(g24178) );
  INVX0 U17833 ( .INP(n17434), .ZN(n17433) );
  NOR2X0 U17834 ( .IN1(n10068), .IN2(test_so23), .QN(n17434) );
  NAND2X0 U17835 ( .IN1(test_so23), .IN2(n13260), .QN(n17432) );
  INVX0 U17836 ( .INP(n13880), .ZN(n13260) );
  NAND2X0 U17837 ( .IN1(n17435), .IN2(n12028), .QN(n13880) );
  NOR2X0 U17838 ( .IN1(n12035), .IN2(n12011), .QN(n17435) );
  NAND2X0 U17839 ( .IN1(n17436), .IN2(n17437), .QN(g24174) );
  NAND2X0 U17840 ( .IN1(n4466), .IN2(g461), .QN(n17437) );
  NAND2X0 U17841 ( .IN1(n15508), .IN2(g485), .QN(n17436) );
  NAND2X0 U17842 ( .IN1(n17438), .IN2(n17439), .QN(g24092) );
  NAND2X0 U17843 ( .IN1(g3229), .IN2(n4483), .QN(n17439) );
  NAND2X0 U17844 ( .IN1(n11195), .IN2(g2380), .QN(n17438) );
  INVX0 U17845 ( .INP(g3229), .ZN(n11195) );
  NAND2X0 U17846 ( .IN1(n17440), .IN2(n17441), .QN(g24083) );
  NAND2X0 U17847 ( .IN1(g3229), .IN2(n4484), .QN(n17441) );
  INVX0 U17848 ( .INP(n17442), .ZN(n17440) );
  NOR2X0 U17849 ( .IN1(g3229), .IN2(n10027), .QN(n17442) );
  NAND2X0 U17850 ( .IN1(n17443), .IN2(n17444), .QN(g24072) );
  NAND2X0 U17851 ( .IN1(g3229), .IN2(n4486), .QN(n17444) );
  INVX0 U17852 ( .INP(n17445), .ZN(n17443) );
  NOR2X0 U17853 ( .IN1(g3229), .IN2(n10028), .QN(n17445) );
  NAND2X0 U17854 ( .IN1(n17446), .IN2(n17447), .QN(g24059) );
  NAND2X0 U17855 ( .IN1(g3229), .IN2(n4485), .QN(n17447) );
  INVX0 U17856 ( .INP(n17448), .ZN(n17446) );
  NOR2X0 U17857 ( .IN1(g3229), .IN2(n9740), .QN(n17448) );
  NAND2X0 U17858 ( .IN1(n17449), .IN2(n17450), .QN(g23418) );
  NAND2X0 U17859 ( .IN1(n4455), .IN2(g2533), .QN(n17450) );
  NAND2X0 U17860 ( .IN1(n15268), .IN2(g8167), .QN(n17449) );
  NAND2X0 U17861 ( .IN1(n17451), .IN2(n17452), .QN(g23413) );
  NAND2X0 U17862 ( .IN1(n15378), .IN2(g8082), .QN(n17452) );
  NAND2X0 U17863 ( .IN1(test_so65), .IN2(n4457), .QN(n17451) );
  NAND2X0 U17864 ( .IN1(n17453), .IN2(n17454), .QN(g23407) );
  NAND2X0 U17865 ( .IN1(n4456), .IN2(g2530), .QN(n17454) );
  NAND2X0 U17866 ( .IN1(n15268), .IN2(g8087), .QN(n17453) );
  INVX0 U17867 ( .INP(n10975), .ZN(n15268) );
  NAND2X0 U17868 ( .IN1(n17455), .IN2(n12475), .QN(n10975) );
  INVX0 U17869 ( .INP(n12478), .ZN(n12475) );
  NAND2X0 U17870 ( .IN1(n17456), .IN2(n17457), .QN(n12478) );
  NAND2X0 U17871 ( .IN1(n9536), .IN2(n11937), .QN(n17457) );
  NOR2X0 U17872 ( .IN1(n17458), .IN2(n17459), .QN(n17456) );
  NOR2X0 U17873 ( .IN1(n4516), .IN2(g2387), .QN(n17459) );
  NOR2X0 U17874 ( .IN1(n4509), .IN2(g2389), .QN(n17458) );
  NOR2X0 U17875 ( .IN1(n12491), .IN2(n12498), .QN(n17455) );
  INVX0 U17876 ( .INP(n12487), .ZN(n12498) );
  NAND2X0 U17877 ( .IN1(n17460), .IN2(n17461), .QN(n12487) );
  NAND2X0 U17878 ( .IN1(n9534), .IN2(n11937), .QN(n17461) );
  NOR2X0 U17879 ( .IN1(n17462), .IN2(n17463), .QN(n17460) );
  NOR2X0 U17880 ( .IN1(n4516), .IN2(g2393), .QN(n17463) );
  NOR2X0 U17881 ( .IN1(n4509), .IN2(g2395), .QN(n17462) );
  INVX0 U17882 ( .INP(n12470), .ZN(n12491) );
  NAND2X0 U17883 ( .IN1(n17464), .IN2(n17465), .QN(n12470) );
  NAND2X0 U17884 ( .IN1(n9535), .IN2(n11937), .QN(n17465) );
  INVX0 U17885 ( .INP(n4524), .ZN(n11937) );
  NOR2X0 U17886 ( .IN1(n17466), .IN2(n17467), .QN(n17464) );
  NOR2X0 U17887 ( .IN1(n4516), .IN2(g2390), .QN(n17467) );
  NOR2X0 U17888 ( .IN1(n4509), .IN2(g2392), .QN(n17466) );
  NAND2X0 U17889 ( .IN1(n17468), .IN2(n17469), .QN(g23406) );
  NAND2X0 U17890 ( .IN1(n4459), .IN2(g1145), .QN(n17469) );
  NAND2X0 U17891 ( .IN1(n17431), .IN2(g8007), .QN(n17468) );
  NAND2X0 U17892 ( .IN1(n17470), .IN2(n17471), .QN(g23400) );
  NAND2X0 U17893 ( .IN1(n4458), .IN2(g1836), .QN(n17471) );
  NAND2X0 U17894 ( .IN1(n15378), .IN2(g8012), .QN(n17470) );
  INVX0 U17895 ( .INP(n10910), .ZN(n15378) );
  NAND2X0 U17896 ( .IN1(n17472), .IN2(n11961), .QN(n10910) );
  INVX0 U17897 ( .INP(n11964), .ZN(n11961) );
  NAND2X0 U17898 ( .IN1(n17473), .IN2(n17474), .QN(n11964) );
  NAND2X0 U17899 ( .IN1(n9539), .IN2(n11946), .QN(n17474) );
  NOR2X0 U17900 ( .IN1(n17475), .IN2(n17476), .QN(n17473) );
  NOR2X0 U17901 ( .IN1(n4518), .IN2(g1693), .QN(n17476) );
  NOR2X0 U17902 ( .IN1(n4511), .IN2(g1695), .QN(n17475) );
  NOR2X0 U17903 ( .IN1(n11978), .IN2(n11985), .QN(n17472) );
  INVX0 U17904 ( .INP(n11975), .ZN(n11985) );
  NAND2X0 U17905 ( .IN1(n17477), .IN2(n17478), .QN(n11975) );
  NAND2X0 U17906 ( .IN1(n9537), .IN2(n11946), .QN(n17478) );
  NOR2X0 U17907 ( .IN1(n17479), .IN2(n17480), .QN(n17477) );
  NOR2X0 U17908 ( .IN1(n4518), .IN2(g1699), .QN(n17480) );
  NOR2X0 U17909 ( .IN1(n4511), .IN2(g1701), .QN(n17479) );
  INVX0 U17910 ( .INP(n11956), .ZN(n11978) );
  NAND2X0 U17911 ( .IN1(n17481), .IN2(n17482), .QN(n11956) );
  NAND2X0 U17912 ( .IN1(n9538), .IN2(n11946), .QN(n17482) );
  INVX0 U17913 ( .INP(n4525), .ZN(n11946) );
  NOR2X0 U17914 ( .IN1(n17483), .IN2(n17484), .QN(n17481) );
  NOR2X0 U17915 ( .IN1(n4518), .IN2(g1696), .QN(n17484) );
  NOR2X0 U17916 ( .IN1(n4511), .IN2(g1698), .QN(n17483) );
  NAND2X0 U17917 ( .IN1(n17485), .IN2(n17486), .QN(g23399) );
  NAND2X0 U17918 ( .IN1(n4461), .IN2(g458), .QN(n17486) );
  NAND2X0 U17919 ( .IN1(n15508), .IN2(g7956), .QN(n17485) );
  NAND2X0 U17920 ( .IN1(n17487), .IN2(n17488), .QN(g23392) );
  NAND2X0 U17921 ( .IN1(n4460), .IN2(g1142), .QN(n17488) );
  NAND2X0 U17922 ( .IN1(n17431), .IN2(g7961), .QN(n17487) );
  INVX0 U17923 ( .INP(n10845), .ZN(n17431) );
  NAND2X0 U17924 ( .IN1(n17489), .IN2(n11787), .QN(n10845) );
  INVX0 U17925 ( .INP(n11759), .ZN(n11787) );
  NAND2X0 U17926 ( .IN1(n17490), .IN2(n17491), .QN(n11759) );
  NAND2X0 U17927 ( .IN1(n9558), .IN2(g1088), .QN(n17491) );
  NOR2X0 U17928 ( .IN1(n17492), .IN2(n17493), .QN(n17490) );
  NOR2X0 U17929 ( .IN1(n4364), .IN2(g1000), .QN(n17493) );
  NOR2X0 U17930 ( .IN1(n4363), .IN2(g999), .QN(n17492) );
  NOR2X0 U17931 ( .IN1(n11766), .IN2(n11756), .QN(n17489) );
  INVX0 U17932 ( .INP(n11753), .ZN(n11756) );
  NAND2X0 U17933 ( .IN1(n17494), .IN2(n17495), .QN(n11753) );
  NAND2X0 U17934 ( .IN1(g1088), .IN2(n10339), .QN(n17495) );
  NOR2X0 U17935 ( .IN1(n17496), .IN2(n17497), .QN(n17494) );
  NOR2X0 U17936 ( .IN1(n4364), .IN2(g1006), .QN(n17497) );
  NOR2X0 U17937 ( .IN1(n4363), .IN2(g1005), .QN(n17496) );
  INVX0 U17938 ( .INP(n11762), .ZN(n11766) );
  NAND2X0 U17939 ( .IN1(n17498), .IN2(n17499), .QN(n11762) );
  NAND2X0 U17940 ( .IN1(n9556), .IN2(g1088), .QN(n17499) );
  NOR2X0 U17941 ( .IN1(n17500), .IN2(n17501), .QN(n17498) );
  NOR2X0 U17942 ( .IN1(n4364), .IN2(g1003), .QN(n17501) );
  NOR2X0 U17943 ( .IN1(n4363), .IN2(g1002), .QN(n17500) );
  NAND2X0 U17944 ( .IN1(n17502), .IN2(n17503), .QN(g23385) );
  NAND2X0 U17945 ( .IN1(g455), .IN2(n10328), .QN(n17503) );
  NAND2X0 U17946 ( .IN1(n15508), .IN2(test_so23), .QN(n17502) );
  INVX0 U17947 ( .INP(n10781), .ZN(n15508) );
  NAND2X0 U17948 ( .IN1(n17504), .IN2(n12011), .QN(n10781) );
  INVX0 U17949 ( .INP(n12014), .ZN(n12011) );
  NAND2X0 U17950 ( .IN1(n17505), .IN2(n17506), .QN(n12014) );
  NAND2X0 U17951 ( .IN1(n9567), .IN2(n12042), .QN(n17506) );
  NOR2X0 U17952 ( .IN1(n17507), .IN2(n17508), .QN(n17505) );
  NOR2X0 U17953 ( .IN1(n4506), .IN2(g314), .QN(n17508) );
  NOR2X0 U17954 ( .IN1(n4499), .IN2(g313), .QN(n17507) );
  NOR2X0 U17955 ( .IN1(n12028), .IN2(n12035), .QN(n17504) );
  INVX0 U17956 ( .INP(n12025), .ZN(n12035) );
  NAND2X0 U17957 ( .IN1(n17509), .IN2(n17510), .QN(n12025) );
  NAND2X0 U17958 ( .IN1(n9562), .IN2(n12042), .QN(n17510) );
  NOR2X0 U17959 ( .IN1(n17511), .IN2(n17512), .QN(n17509) );
  NOR2X0 U17960 ( .IN1(n4506), .IN2(g320), .QN(n17512) );
  NOR2X0 U17961 ( .IN1(n4499), .IN2(g319), .QN(n17511) );
  INVX0 U17962 ( .INP(n12006), .ZN(n12028) );
  NAND2X0 U17963 ( .IN1(n17513), .IN2(n17514), .QN(n12006) );
  NAND2X0 U17964 ( .IN1(n9564), .IN2(n12042), .QN(n17514) );
  INVX0 U17965 ( .INP(n4520), .ZN(n12042) );
  NOR2X0 U17966 ( .IN1(n17515), .IN2(n17516), .QN(n17513) );
  NOR2X0 U17967 ( .IN1(n4506), .IN2(g317), .QN(n17516) );
  NOR2X0 U17968 ( .IN1(test_so18), .IN2(n4499), .QN(n17515) );
  NOR2X0 U17969 ( .IN1(n17087), .IN2(n17517), .QN(g23359) );
  NAND2X0 U17970 ( .IN1(n4102), .IN2(n17518), .QN(n17517) );
  NAND2X0 U17971 ( .IN1(n4350), .IN2(n11065), .QN(n17518) );
  NAND2X0 U17972 ( .IN1(n17519), .IN2(g3028), .QN(n4102) );
  INVX0 U17973 ( .INP(n11065), .ZN(n17519) );
  NAND2X0 U17974 ( .IN1(n17520), .IN2(g3018), .QN(n11065) );
  INVX0 U17975 ( .INP(n11064), .ZN(n17087) );
  NAND2X0 U17976 ( .IN1(n15740), .IN2(n17521), .QN(n11064) );
  NAND2X0 U17977 ( .IN1(n17522), .IN2(n11062), .QN(n17521) );
  NAND2X0 U17978 ( .IN1(n17523), .IN2(n17524), .QN(n17522) );
  NOR2X0 U17979 ( .IN1(n9736), .IN2(n4481), .QN(n17524) );
  NOR2X0 U17980 ( .IN1(g3036), .IN2(g3028), .QN(n17523) );
  NOR2X0 U17981 ( .IN1(n10998), .IN2(n17525), .QN(g23358) );
  INVX0 U17982 ( .INP(n17526), .ZN(n17525) );
  NOR2X0 U17983 ( .IN1(n4122), .IN2(n17337), .QN(n17526) );
  NOR2X0 U17984 ( .IN1(n4123), .IN2(n4431), .QN(n17337) );
  NOR2X0 U17985 ( .IN1(n17101), .IN2(n17527), .QN(g23357) );
  NAND2X0 U17986 ( .IN1(n17528), .IN2(n17529), .QN(n17527) );
  NAND2X0 U17987 ( .IN1(n4479), .IN2(n11004), .QN(n17529) );
  INVX0 U17988 ( .INP(n17332), .ZN(n11004) );
  NAND2X0 U17989 ( .IN1(n17332), .IN2(g2917), .QN(n17528) );
  NOR2X0 U17990 ( .IN1(n11005), .IN2(n4482), .QN(n17332) );
  INVX0 U17991 ( .INP(n11001), .ZN(n17101) );
  NAND2X0 U17992 ( .IN1(n10998), .IN2(n17530), .QN(n11001) );
  NAND2X0 U17993 ( .IN1(n18867), .IN2(n17531), .QN(n17530) );
  NAND2X0 U17994 ( .IN1(n17532), .IN2(n17533), .QN(n17531) );
  NOR2X0 U17995 ( .IN1(n4482), .IN2(n10026), .QN(n17533) );
  NOR2X0 U17996 ( .IN1(g2924), .IN2(g2917), .QN(n17532) );
  NOR2X0 U17997 ( .IN1(n14690), .IN2(n17534), .QN(g23348) );
  NAND2X0 U17998 ( .IN1(n17535), .IN2(n17536), .QN(n17534) );
  NAND2X0 U17999 ( .IN1(n4419), .IN2(n17349), .QN(n17536) );
  NAND2X0 U18000 ( .IN1(n17347), .IN2(g2727), .QN(n17535) );
  INVX0 U18001 ( .INP(n17349), .ZN(n17347) );
  NOR2X0 U18002 ( .IN1(n15735), .IN2(n17537), .QN(g23339) );
  NAND2X0 U18003 ( .IN1(n17538), .IN2(n17539), .QN(n17537) );
  NAND2X0 U18004 ( .IN1(n4420), .IN2(n17355), .QN(n17539) );
  NAND2X0 U18005 ( .IN1(n17353), .IN2(g2033), .QN(n17538) );
  INVX0 U18006 ( .INP(n17355), .ZN(n17353) );
  NOR2X0 U18007 ( .IN1(n15740), .IN2(n17540), .QN(g23330) );
  NAND2X0 U18008 ( .IN1(n17541), .IN2(n4066), .QN(n17540) );
  NAND2X0 U18009 ( .IN1(n17542), .IN2(n16330), .QN(n4066) );
  NOR2X0 U18010 ( .IN1(n18873), .IN2(n10305), .QN(n17542) );
  NAND2X0 U18011 ( .IN1(n10305), .IN2(n17543), .QN(n17541) );
  NAND2X0 U18012 ( .IN1(n16330), .IN2(n7909), .QN(n17543) );
  NOR2X0 U18013 ( .IN1(n10303), .IN2(n10302), .QN(n16330) );
  NAND2X0 U18014 ( .IN1(n11062), .IN2(n11067), .QN(n15740) );
  INVX0 U18015 ( .INP(n17520), .ZN(n11067) );
  NOR2X0 U18016 ( .IN1(n17328), .IN2(n10302), .QN(n17520) );
  NAND2X0 U18017 ( .IN1(n17544), .IN2(n17545), .QN(n17328) );
  NOR2X0 U18018 ( .IN1(n17546), .IN2(n17547), .QN(n17545) );
  NAND2X0 U18019 ( .IN1(g3013), .IN2(g3024), .QN(n17547) );
  NAND2X0 U18020 ( .IN1(n7909), .IN2(n10327), .QN(n17546) );
  NOR2X0 U18021 ( .IN1(g3006), .IN2(n17548), .QN(n17544) );
  NAND2X0 U18022 ( .IN1(n10303), .IN2(g3002), .QN(n17548) );
  INVX0 U18023 ( .INP(g3234), .ZN(n11062) );
  NOR2X0 U18024 ( .IN1(n14704), .IN2(n17549), .QN(g23329) );
  NAND2X0 U18025 ( .IN1(n17550), .IN2(n17551), .QN(n17549) );
  NAND2X0 U18026 ( .IN1(n4421), .IN2(n17361), .QN(n17551) );
  NAND2X0 U18027 ( .IN1(n17359), .IN2(g1339), .QN(n17550) );
  INVX0 U18028 ( .INP(n17361), .ZN(n17359) );
  NOR2X0 U18029 ( .IN1(n14141), .IN2(n17552), .QN(g23324) );
  NAND2X0 U18030 ( .IN1(n17553), .IN2(n17554), .QN(n17552) );
  NAND2X0 U18031 ( .IN1(n4422), .IN2(n17367), .QN(n17554) );
  NAND2X0 U18032 ( .IN1(n17365), .IN2(g653), .QN(n17553) );
  INVX0 U18033 ( .INP(n17367), .ZN(n17365) );
  NAND2X0 U18034 ( .IN1(n17555), .IN2(n17556), .QN(g23137) );
  INVX0 U18035 ( .INP(n17557), .ZN(n17556) );
  NOR2X0 U18036 ( .IN1(g1866), .IN2(n10046), .QN(n17557) );
  NAND2X0 U18037 ( .IN1(n14773), .IN2(g1866), .QN(n17555) );
  NOR2X0 U18038 ( .IN1(n17558), .IN2(n17559), .QN(g23136) );
  NAND2X0 U18039 ( .IN1(n17367), .IN2(n14712), .QN(n17559) );
  NAND2X0 U18040 ( .IN1(n17560), .IN2(n17561), .QN(n17367) );
  NOR2X0 U18041 ( .IN1(n4478), .IN2(n4404), .QN(n17560) );
  NOR2X0 U18042 ( .IN1(n17562), .IN2(g633), .QN(n17558) );
  NOR2X0 U18043 ( .IN1(n4404), .IN2(n17563), .QN(n17562) );
  NAND2X0 U18044 ( .IN1(n17564), .IN2(n17565), .QN(g23133) );
  NAND2X0 U18045 ( .IN1(n4455), .IN2(g2562), .QN(n17565) );
  NAND2X0 U18046 ( .IN1(n14747), .IN2(g8167), .QN(n17564) );
  NAND2X0 U18047 ( .IN1(n17566), .IN2(n17567), .QN(g23132) );
  INVX0 U18048 ( .INP(n17568), .ZN(n17567) );
  NOR2X0 U18049 ( .IN1(g8087), .IN2(n10039), .QN(n17568) );
  NAND2X0 U18050 ( .IN1(n13322), .IN2(g8087), .QN(n17566) );
  NAND2X0 U18051 ( .IN1(n17569), .IN2(n17570), .QN(g23126) );
  NAND2X0 U18052 ( .IN1(n4465), .IN2(g1175), .QN(n17570) );
  NAND2X0 U18053 ( .IN1(n14799), .IN2(g1172), .QN(n17569) );
  NAND2X0 U18054 ( .IN1(n17571), .IN2(n17572), .QN(g23124) );
  NAND2X0 U18055 ( .IN1(n4457), .IN2(g1868), .QN(n17572) );
  NAND2X0 U18056 ( .IN1(n14773), .IN2(g8082), .QN(n17571) );
  NAND2X0 U18057 ( .IN1(n17573), .IN2(n17574), .QN(g23123) );
  INVX0 U18058 ( .INP(n17575), .ZN(n17574) );
  NOR2X0 U18059 ( .IN1(g8012), .IN2(n10048), .QN(n17575) );
  NAND2X0 U18060 ( .IN1(n13344), .IN2(g8012), .QN(n17573) );
  NAND2X0 U18061 ( .IN1(n17576), .IN2(n17577), .QN(g23117) );
  INVX0 U18062 ( .INP(n17578), .ZN(n17577) );
  NOR2X0 U18063 ( .IN1(g485), .IN2(n10063), .QN(n17578) );
  NAND2X0 U18064 ( .IN1(n14820), .IN2(g485), .QN(n17576) );
  NAND2X0 U18065 ( .IN1(n17579), .IN2(n17580), .QN(g23114) );
  INVX0 U18066 ( .INP(n17581), .ZN(n17580) );
  NOR2X0 U18067 ( .IN1(g8087), .IN2(n10037), .QN(n17581) );
  NAND2X0 U18068 ( .IN1(n14747), .IN2(g8087), .QN(n17579) );
  NAND2X0 U18069 ( .IN1(n17582), .IN2(n17583), .QN(g23111) );
  NAND2X0 U18070 ( .IN1(test_so44), .IN2(n4459), .QN(n17583) );
  NAND2X0 U18071 ( .IN1(n14799), .IN2(g8007), .QN(n17582) );
  NAND2X0 U18072 ( .IN1(n17584), .IN2(n17585), .QN(g23110) );
  INVX0 U18073 ( .INP(n17586), .ZN(n17585) );
  NOR2X0 U18074 ( .IN1(g7961), .IN2(n10056), .QN(n17586) );
  NAND2X0 U18075 ( .IN1(n13369), .IN2(g7961), .QN(n17584) );
  NAND2X0 U18076 ( .IN1(n17587), .IN2(n17588), .QN(g23097) );
  INVX0 U18077 ( .INP(n17589), .ZN(n17588) );
  NOR2X0 U18078 ( .IN1(g8012), .IN2(n10045), .QN(n17589) );
  NAND2X0 U18079 ( .IN1(n14773), .IN2(g8012), .QN(n17587) );
  NAND2X0 U18080 ( .IN1(n17590), .IN2(n17591), .QN(n14773) );
  NAND2X0 U18081 ( .IN1(g5511), .IN2(g1819), .QN(n17591) );
  NOR2X0 U18082 ( .IN1(n17592), .IN2(n17593), .QN(n17590) );
  NOR2X0 U18083 ( .IN1(n9745), .IN2(n13179), .QN(n17593) );
  INVX0 U18084 ( .INP(n17594), .ZN(n17592) );
  NAND2X0 U18085 ( .IN1(n4618), .IN2(test_so59), .QN(n17594) );
  NAND2X0 U18086 ( .IN1(n17595), .IN2(n17596), .QN(g23093) );
  NAND2X0 U18087 ( .IN1(n4461), .IN2(g487), .QN(n17596) );
  NAND2X0 U18088 ( .IN1(n14820), .IN2(g7956), .QN(n17595) );
  NAND2X0 U18089 ( .IN1(n17597), .IN2(n17598), .QN(g23092) );
  INVX0 U18090 ( .INP(n17599), .ZN(n17598) );
  NOR2X0 U18091 ( .IN1(n10065), .IN2(test_so23), .QN(n17599) );
  NAND2X0 U18092 ( .IN1(test_so23), .IN2(n13389), .QN(n17597) );
  NAND2X0 U18093 ( .IN1(n17600), .IN2(n17601), .QN(g23081) );
  INVX0 U18094 ( .INP(n17602), .ZN(n17601) );
  NOR2X0 U18095 ( .IN1(g7961), .IN2(n10054), .QN(n17602) );
  NAND2X0 U18096 ( .IN1(n14799), .IN2(g7961), .QN(n17600) );
  NAND2X0 U18097 ( .IN1(n17603), .IN2(n17604), .QN(n14799) );
  NAND2X0 U18098 ( .IN1(g1088), .IN2(g1131), .QN(n17604) );
  NOR2X0 U18099 ( .IN1(n17605), .IN2(n17606), .QN(n17603) );
  NOR2X0 U18100 ( .IN1(n9749), .IN2(n4364), .QN(n17606) );
  NOR2X0 U18101 ( .IN1(n9767), .IN2(n4363), .QN(n17605) );
  NAND2X0 U18102 ( .IN1(n17607), .IN2(n17608), .QN(g23076) );
  INVX0 U18103 ( .INP(n17609), .ZN(n17608) );
  NOR2X0 U18104 ( .IN1(g2560), .IN2(n10040), .QN(n17609) );
  NAND2X0 U18105 ( .IN1(n13322), .IN2(g2560), .QN(n17607) );
  NAND2X0 U18106 ( .IN1(n17610), .IN2(n17611), .QN(g23067) );
  INVX0 U18107 ( .INP(n17612), .ZN(n17611) );
  NOR2X0 U18108 ( .IN1(n10062), .IN2(test_so23), .QN(n17612) );
  NAND2X0 U18109 ( .IN1(test_so23), .IN2(n14820), .QN(n17610) );
  NAND2X0 U18110 ( .IN1(n17613), .IN2(n17614), .QN(n14820) );
  NAND2X0 U18111 ( .IN1(g5437), .IN2(g438), .QN(n17614) );
  NOR2X0 U18112 ( .IN1(n17615), .IN2(n17616), .QN(n17613) );
  NOR2X0 U18113 ( .IN1(n9775), .IN2(n14129), .QN(n17616) );
  NOR2X0 U18114 ( .IN1(n9774), .IN2(n14130), .QN(n17615) );
  NAND2X0 U18115 ( .IN1(n17617), .IN2(n17618), .QN(g23058) );
  INVX0 U18116 ( .INP(n17619), .ZN(n17618) );
  NOR2X0 U18117 ( .IN1(g1866), .IN2(n10049), .QN(n17619) );
  NAND2X0 U18118 ( .IN1(n13344), .IN2(g1866), .QN(n17617) );
  NAND2X0 U18119 ( .IN1(n17620), .IN2(n17621), .QN(g23047) );
  NAND2X0 U18120 ( .IN1(n4455), .IN2(g2559), .QN(n17621) );
  NAND2X0 U18121 ( .IN1(n13322), .IN2(g8167), .QN(n17620) );
  INVX0 U18122 ( .INP(n4285), .ZN(n13322) );
  NAND2X0 U18123 ( .IN1(n17622), .IN2(n17623), .QN(n4285) );
  NAND2X0 U18124 ( .IN1(g5555), .IN2(g2492), .QN(n17623) );
  NOR2X0 U18125 ( .IN1(n17624), .IN2(n17625), .QN(n17622) );
  NOR2X0 U18126 ( .IN1(n9743), .IN2(n14010), .QN(n17625) );
  NOR2X0 U18127 ( .IN1(n9756), .IN2(n15607), .QN(n17624) );
  NAND2X0 U18128 ( .IN1(n17626), .IN2(n17627), .QN(g23039) );
  INVX0 U18129 ( .INP(n17628), .ZN(n17627) );
  NOR2X0 U18130 ( .IN1(g1172), .IN2(n10057), .QN(n17628) );
  NAND2X0 U18131 ( .IN1(n13369), .IN2(g1172), .QN(n17626) );
  NAND2X0 U18132 ( .IN1(n17629), .IN2(n17630), .QN(g23030) );
  NAND2X0 U18133 ( .IN1(n4457), .IN2(g1865), .QN(n17630) );
  NAND2X0 U18134 ( .IN1(n13344), .IN2(g8082), .QN(n17629) );
  INVX0 U18135 ( .INP(n4284), .ZN(n13344) );
  NAND2X0 U18136 ( .IN1(n17631), .IN2(n17632), .QN(n4284) );
  NAND2X0 U18137 ( .IN1(g5511), .IN2(g1798), .QN(n17632) );
  NOR2X0 U18138 ( .IN1(n17633), .IN2(n17634), .QN(n17631) );
  NOR2X0 U18139 ( .IN1(n9747), .IN2(n13179), .QN(n17634) );
  INVX0 U18140 ( .INP(g7014), .ZN(n13179) );
  NOR2X0 U18141 ( .IN1(n9762), .IN2(n14055), .QN(n17633) );
  INVX0 U18142 ( .INP(n4618), .ZN(n14055) );
  NAND2X0 U18143 ( .IN1(n17635), .IN2(n17636), .QN(g23022) );
  INVX0 U18144 ( .INP(n17637), .ZN(n17636) );
  NOR2X0 U18145 ( .IN1(g485), .IN2(n10066), .QN(n17637) );
  NAND2X0 U18146 ( .IN1(n13389), .IN2(g485), .QN(n17635) );
  NAND2X0 U18147 ( .IN1(n17638), .IN2(n17639), .QN(g23014) );
  NAND2X0 U18148 ( .IN1(n4459), .IN2(g1171), .QN(n17639) );
  NAND2X0 U18149 ( .IN1(n13369), .IN2(g8007), .QN(n17638) );
  INVX0 U18150 ( .INP(n4283), .ZN(n13369) );
  NAND2X0 U18151 ( .IN1(n17640), .IN2(n17641), .QN(n4283) );
  NAND2X0 U18152 ( .IN1(g1088), .IN2(g1110), .QN(n17641) );
  NOR2X0 U18153 ( .IN1(n17642), .IN2(n17643), .QN(n17640) );
  NOR2X0 U18154 ( .IN1(n9750), .IN2(n4364), .QN(n17643) );
  NOR2X0 U18155 ( .IN1(n9771), .IN2(n4363), .QN(n17642) );
  NAND2X0 U18156 ( .IN1(n17644), .IN2(n17645), .QN(g23000) );
  NAND2X0 U18157 ( .IN1(n4461), .IN2(g484), .QN(n17645) );
  NAND2X0 U18158 ( .IN1(n13389), .IN2(g7956), .QN(n17644) );
  INVX0 U18159 ( .INP(n4282), .ZN(n13389) );
  NAND2X0 U18160 ( .IN1(n17646), .IN2(n17647), .QN(n4282) );
  NAND2X0 U18161 ( .IN1(g5437), .IN2(g417), .QN(n17647) );
  NOR2X0 U18162 ( .IN1(n17648), .IN2(n17649), .QN(n17646) );
  NOR2X0 U18163 ( .IN1(n9781), .IN2(n14129), .QN(n17649) );
  INVX0 U18164 ( .INP(g6447), .ZN(n14129) );
  NOR2X0 U18165 ( .IN1(n9780), .IN2(n14130), .QN(n17648) );
  INVX0 U18166 ( .INP(n4640), .ZN(n14130) );
  NAND2X0 U18167 ( .IN1(n17650), .IN2(n17651), .QN(g22687) );
  NAND2X0 U18168 ( .IN1(n17652), .IN2(n17653), .QN(n17651) );
  INVX0 U18169 ( .INP(n16141), .ZN(n17653) );
  NOR2X0 U18170 ( .IN1(n4303), .IN2(n11267), .QN(n17652) );
  NAND2X0 U18171 ( .IN1(n17654), .IN2(n17655), .QN(n17650) );
  NAND2X0 U18172 ( .IN1(n11846), .IN2(n16141), .QN(n17654) );
  NAND2X0 U18173 ( .IN1(n17656), .IN2(n17657), .QN(n16141) );
  NAND2X0 U18174 ( .IN1(g7390), .IN2(g2568), .QN(n17657) );
  NOR2X0 U18175 ( .IN1(n17658), .IN2(n17659), .QN(n17656) );
  NOR2X0 U18176 ( .IN1(n9786), .IN2(n4314), .QN(n17659) );
  NOR2X0 U18177 ( .IN1(n9788), .IN2(n4299), .QN(n17658) );
  NAND2X0 U18178 ( .IN1(n17660), .IN2(n17661), .QN(g22651) );
  NAND2X0 U18179 ( .IN1(n17662), .IN2(n17663), .QN(n17661) );
  INVX0 U18180 ( .INP(n16152), .ZN(n17663) );
  NOR2X0 U18181 ( .IN1(n4297), .IN2(n11438), .QN(n17662) );
  NAND2X0 U18182 ( .IN1(n17664), .IN2(n17655), .QN(n17660) );
  NAND2X0 U18183 ( .IN1(n11508), .IN2(n16152), .QN(n17664) );
  NAND2X0 U18184 ( .IN1(n17665), .IN2(n17666), .QN(n16152) );
  NAND2X0 U18185 ( .IN1(g1930), .IN2(g1877), .QN(n17666) );
  NOR2X0 U18186 ( .IN1(n17667), .IN2(n17668), .QN(n17665) );
  NOR2X0 U18187 ( .IN1(n9793), .IN2(n4315), .QN(n17668) );
  INVX0 U18188 ( .INP(n17669), .ZN(n17667) );
  NAND2X0 U18189 ( .IN1(n14321), .IN2(test_so68), .QN(n17669) );
  NAND2X0 U18190 ( .IN1(n17670), .IN2(n17671), .QN(g22615) );
  NAND2X0 U18191 ( .IN1(n17672), .IN2(n17673), .QN(n17671) );
  INVX0 U18192 ( .INP(n16163), .ZN(n17673) );
  NOR2X0 U18193 ( .IN1(n4304), .IN2(n11614), .QN(n17672) );
  NAND2X0 U18194 ( .IN1(n17674), .IN2(n17655), .QN(n17670) );
  NAND2X0 U18195 ( .IN1(n11684), .IN2(n16163), .QN(n17674) );
  NAND2X0 U18196 ( .IN1(n17675), .IN2(n17676), .QN(n16163) );
  NAND2X0 U18197 ( .IN1(test_so47), .IN2(n14180), .QN(n17676) );
  NOR2X0 U18198 ( .IN1(n17677), .IN2(n17678), .QN(n17675) );
  NOR2X0 U18199 ( .IN1(n9794), .IN2(n4316), .QN(n17678) );
  NOR2X0 U18200 ( .IN1(n9790), .IN2(n4300), .QN(n17677) );
  NAND2X0 U18201 ( .IN1(n17679), .IN2(n17680), .QN(g22578) );
  NAND2X0 U18202 ( .IN1(n17681), .IN2(n17682), .QN(n17680) );
  INVX0 U18203 ( .INP(n16170), .ZN(n17682) );
  NOR2X0 U18204 ( .IN1(n11130), .IN2(n10326), .QN(n17681) );
  NAND2X0 U18205 ( .IN1(n17683), .IN2(n17655), .QN(n17679) );
  NAND2X0 U18206 ( .IN1(n11174), .IN2(n16170), .QN(n17683) );
  NAND2X0 U18207 ( .IN1(n17684), .IN2(n17685), .QN(n16170) );
  NAND2X0 U18208 ( .IN1(g6642), .IN2(g493), .QN(n17685) );
  NOR2X0 U18209 ( .IN1(n17686), .IN2(n17687), .QN(n17684) );
  NOR2X0 U18210 ( .IN1(n9791), .IN2(n4313), .QN(n17687) );
  NOR2X0 U18211 ( .IN1(n9787), .IN2(n17296), .QN(n17686) );
  NOR2X0 U18212 ( .IN1(n17688), .IN2(n17689), .QN(g22299) );
  NOR2X0 U18213 ( .IN1(n16490), .IN2(test_so95), .QN(n17689) );
  NOR2X0 U18214 ( .IN1(n14690), .IN2(n17690), .QN(g22284) );
  NOR2X0 U18215 ( .IN1(n16494), .IN2(g2813), .QN(n17690) );
  NOR2X0 U18216 ( .IN1(n17691), .IN2(n17692), .QN(g22280) );
  NOR2X0 U18217 ( .IN1(n16499), .IN2(g2117), .QN(n17692) );
  INVX0 U18218 ( .INP(n17693), .ZN(g22269) );
  NAND2X0 U18219 ( .IN1(n17694), .IN2(n17695), .QN(n17693) );
  NAND2X0 U18220 ( .IN1(n16502), .IN2(n10193), .QN(n17695) );
  NOR2X0 U18221 ( .IN1(n15735), .IN2(n17696), .QN(g22267) );
  NOR2X0 U18222 ( .IN1(n16596), .IN2(g2119), .QN(n17696) );
  NOR2X0 U18223 ( .IN1(n17697), .IN2(n17698), .QN(g22263) );
  NOR2X0 U18224 ( .IN1(n16602), .IN2(g1423), .QN(n17698) );
  NOR2X0 U18225 ( .IN1(n17699), .IN2(n17700), .QN(g22249) );
  INVX0 U18226 ( .INP(n17701), .ZN(n17700) );
  NAND2X0 U18227 ( .IN1(n16698), .IN2(n10194), .QN(n17701) );
  NOR2X0 U18228 ( .IN1(n14704), .IN2(n17702), .QN(g22247) );
  NOR2X0 U18229 ( .IN1(n16702), .IN2(g1425), .QN(n17702) );
  NOR2X0 U18230 ( .IN1(n17703), .IN2(n17704), .QN(g22242) );
  NOR2X0 U18231 ( .IN1(n16707), .IN2(g737), .QN(n17704) );
  NOR2X0 U18232 ( .IN1(n17705), .IN2(n17706), .QN(g22234) );
  INVX0 U18233 ( .INP(n17707), .ZN(n17706) );
  NAND2X0 U18234 ( .IN1(n16716), .IN2(n10195), .QN(n17707) );
  NOR2X0 U18235 ( .IN1(n14141), .IN2(n17708), .QN(g22231) );
  NOR2X0 U18236 ( .IN1(n16813), .IN2(g739), .QN(n17708) );
  NOR2X0 U18237 ( .IN1(n17709), .IN2(n17710), .QN(g22218) );
  INVX0 U18238 ( .INP(n17711), .ZN(n17710) );
  NAND2X0 U18239 ( .IN1(n16816), .IN2(n10196), .QN(n17711) );
  NAND2X0 U18240 ( .IN1(n17712), .IN2(n17713), .QN(g22200) );
  NAND2X0 U18241 ( .IN1(n17714), .IN2(n4373), .QN(n17713) );
  INVX0 U18242 ( .INP(n17715), .ZN(n17712) );
  NOR2X0 U18243 ( .IN1(n17714), .IN2(n9842), .QN(n17715) );
  NAND2X0 U18244 ( .IN1(n17716), .IN2(n17717), .QN(g22194) );
  NAND2X0 U18245 ( .IN1(n17122), .IN2(g2238), .QN(n17717) );
  NAND2X0 U18246 ( .IN1(n17714), .IN2(n12088), .QN(n17716) );
  NAND2X0 U18247 ( .IN1(n17718), .IN2(n17719), .QN(g22193) );
  NAND2X0 U18248 ( .IN1(n17720), .IN2(n4373), .QN(n17719) );
  NAND2X0 U18249 ( .IN1(n17721), .IN2(g2210), .QN(n17718) );
  NAND2X0 U18250 ( .IN1(n17722), .IN2(n17723), .QN(g22192) );
  NAND2X0 U18251 ( .IN1(n17714), .IN2(n4377), .QN(n17723) );
  INVX0 U18252 ( .INP(n17724), .ZN(n17722) );
  NOR2X0 U18253 ( .IN1(n17714), .IN2(n9843), .QN(n17724) );
  NAND2X0 U18254 ( .IN1(n17725), .IN2(n17726), .QN(g22191) );
  NAND2X0 U18255 ( .IN1(n17727), .IN2(n4374), .QN(n17726) );
  INVX0 U18256 ( .INP(n17728), .ZN(n17725) );
  NOR2X0 U18257 ( .IN1(n17727), .IN2(n9853), .QN(n17728) );
  NAND2X0 U18258 ( .IN1(n17729), .IN2(n17730), .QN(g22185) );
  NAND2X0 U18259 ( .IN1(test_so75), .IN2(n17721), .QN(n17730) );
  NAND2X0 U18260 ( .IN1(n17720), .IN2(n12088), .QN(n17729) );
  NAND2X0 U18261 ( .IN1(n17731), .IN2(n17732), .QN(g22184) );
  NAND2X0 U18262 ( .IN1(n17122), .IN2(g2235), .QN(n17732) );
  NAND2X0 U18263 ( .IN1(n13519), .IN2(n17714), .QN(n17731) );
  NAND2X0 U18264 ( .IN1(n17733), .IN2(n17734), .QN(g22183) );
  NAND2X0 U18265 ( .IN1(n17735), .IN2(n4373), .QN(n17734) );
  NAND2X0 U18266 ( .IN1(n17736), .IN2(g2209), .QN(n17733) );
  NAND2X0 U18267 ( .IN1(n17737), .IN2(n17738), .QN(g22182) );
  NAND2X0 U18268 ( .IN1(n17720), .IN2(n4377), .QN(n17738) );
  NAND2X0 U18269 ( .IN1(n17721), .IN2(g2207), .QN(n17737) );
  NAND2X0 U18270 ( .IN1(n17739), .IN2(n17740), .QN(g22180) );
  NAND2X0 U18271 ( .IN1(n17127), .IN2(g1544), .QN(n17740) );
  NAND2X0 U18272 ( .IN1(n17727), .IN2(n12132), .QN(n17739) );
  NAND2X0 U18273 ( .IN1(n17741), .IN2(n17742), .QN(g22179) );
  NAND2X0 U18274 ( .IN1(n17743), .IN2(n4374), .QN(n17742) );
  NAND2X0 U18275 ( .IN1(n17744), .IN2(g1516), .QN(n17741) );
  NAND2X0 U18276 ( .IN1(n17745), .IN2(n17746), .QN(g22178) );
  NAND2X0 U18277 ( .IN1(n17727), .IN2(n4378), .QN(n17746) );
  INVX0 U18278 ( .INP(n17747), .ZN(n17745) );
  NOR2X0 U18279 ( .IN1(n17727), .IN2(n9854), .QN(n17747) );
  NAND2X0 U18280 ( .IN1(n17748), .IN2(n17749), .QN(g22177) );
  NAND2X0 U18281 ( .IN1(n17132), .IN2(n4375), .QN(n17749) );
  INVX0 U18282 ( .INP(n17750), .ZN(n17748) );
  NOR2X0 U18283 ( .IN1(n17132), .IN2(n9867), .QN(n17750) );
  NAND2X0 U18284 ( .IN1(n17751), .IN2(n17752), .QN(g22173) );
  NAND2X0 U18285 ( .IN1(n17736), .IN2(g2239), .QN(n17752) );
  NAND2X0 U18286 ( .IN1(n17735), .IN2(n12088), .QN(n17751) );
  INVX0 U18287 ( .INP(n13485), .ZN(n12088) );
  NAND2X0 U18288 ( .IN1(n17753), .IN2(n17754), .QN(n13485) );
  NAND2X0 U18289 ( .IN1(n9897), .IN2(test_so73), .QN(n17754) );
  NOR2X0 U18290 ( .IN1(n17755), .IN2(n17756), .QN(n17753) );
  NOR2X0 U18291 ( .IN1(n4367), .IN2(g2247), .QN(n17756) );
  NOR2X0 U18292 ( .IN1(n4324), .IN2(g2248), .QN(n17755) );
  NAND2X0 U18293 ( .IN1(n17757), .IN2(n17758), .QN(g22172) );
  INVX0 U18294 ( .INP(n17759), .ZN(n17758) );
  NOR2X0 U18295 ( .IN1(n17720), .IN2(n9826), .QN(n17759) );
  NAND2X0 U18296 ( .IN1(n17720), .IN2(n13519), .QN(n17757) );
  NAND2X0 U18297 ( .IN1(n17760), .IN2(n17761), .QN(g22171) );
  NAND2X0 U18298 ( .IN1(n17714), .IN2(n4287), .QN(n17761) );
  INVX0 U18299 ( .INP(n17762), .ZN(n17760) );
  NOR2X0 U18300 ( .IN1(n17714), .IN2(n9836), .QN(n17762) );
  NAND2X0 U18301 ( .IN1(n17763), .IN2(n17764), .QN(g22170) );
  NAND2X0 U18302 ( .IN1(n17735), .IN2(n4377), .QN(n17764) );
  NAND2X0 U18303 ( .IN1(n17736), .IN2(g2206), .QN(n17763) );
  NAND2X0 U18304 ( .IN1(n17765), .IN2(n17766), .QN(g22169) );
  INVX0 U18305 ( .INP(n17767), .ZN(n17766) );
  NOR2X0 U18306 ( .IN1(n17743), .IN2(n9845), .QN(n17767) );
  NAND2X0 U18307 ( .IN1(n17743), .IN2(n12132), .QN(n17765) );
  NAND2X0 U18308 ( .IN1(n17768), .IN2(n17769), .QN(g22168) );
  NAND2X0 U18309 ( .IN1(n17127), .IN2(g1541), .QN(n17769) );
  NAND2X0 U18310 ( .IN1(n12365), .IN2(n17727), .QN(n17768) );
  NAND2X0 U18311 ( .IN1(n17770), .IN2(n17771), .QN(g22167) );
  NAND2X0 U18312 ( .IN1(test_so52), .IN2(n17772), .QN(n17771) );
  NAND2X0 U18313 ( .IN1(n17773), .IN2(n4374), .QN(n17770) );
  NAND2X0 U18314 ( .IN1(n17774), .IN2(n17775), .QN(g22166) );
  NAND2X0 U18315 ( .IN1(n17743), .IN2(n4378), .QN(n17775) );
  NAND2X0 U18316 ( .IN1(n17744), .IN2(g1513), .QN(n17774) );
  NAND2X0 U18317 ( .IN1(n17776), .IN2(n17777), .QN(g22164) );
  INVX0 U18318 ( .INP(n17778), .ZN(n17777) );
  NOR2X0 U18319 ( .IN1(n17132), .IN2(n9855), .QN(n17778) );
  NAND2X0 U18320 ( .IN1(n17132), .IN2(n12178), .QN(n17776) );
  NAND2X0 U18321 ( .IN1(n17779), .IN2(n17780), .QN(g22163) );
  NAND2X0 U18322 ( .IN1(n17781), .IN2(n4375), .QN(n17780) );
  NAND2X0 U18323 ( .IN1(n17782), .IN2(g822), .QN(n17779) );
  NAND2X0 U18324 ( .IN1(n17783), .IN2(n17784), .QN(g22162) );
  NAND2X0 U18325 ( .IN1(n4379), .IN2(n17132), .QN(n17784) );
  INVX0 U18326 ( .INP(n17785), .ZN(n17783) );
  NOR2X0 U18327 ( .IN1(n17132), .IN2(n9868), .QN(n17785) );
  NAND2X0 U18328 ( .IN1(n17786), .IN2(n17787), .QN(g22161) );
  NAND2X0 U18329 ( .IN1(n17788), .IN2(n4376), .QN(n17787) );
  INVX0 U18330 ( .INP(n17789), .ZN(n17786) );
  NOR2X0 U18331 ( .IN1(n17788), .IN2(n9876), .QN(n17789) );
  NAND2X0 U18332 ( .IN1(n17790), .IN2(n17791), .QN(g22155) );
  NAND2X0 U18333 ( .IN1(n17736), .IN2(g2236), .QN(n17791) );
  NAND2X0 U18334 ( .IN1(n17735), .IN2(n13519), .QN(n17790) );
  INVX0 U18335 ( .INP(n12307), .ZN(n13519) );
  NAND2X0 U18336 ( .IN1(n17792), .IN2(n17793), .QN(n12307) );
  NAND2X0 U18337 ( .IN1(n9894), .IN2(test_so73), .QN(n17793) );
  NOR2X0 U18338 ( .IN1(n17794), .IN2(n17795), .QN(n17792) );
  NOR2X0 U18339 ( .IN1(n4367), .IN2(g2250), .QN(n17795) );
  NOR2X0 U18340 ( .IN1(n4324), .IN2(g2251), .QN(n17794) );
  NAND2X0 U18341 ( .IN1(n17796), .IN2(n17797), .QN(g22154) );
  NAND2X0 U18342 ( .IN1(n17720), .IN2(n4287), .QN(n17797) );
  NAND2X0 U18343 ( .IN1(n17721), .IN2(g2234), .QN(n17796) );
  NAND2X0 U18344 ( .IN1(n17798), .IN2(n17799), .QN(g22153) );
  NAND2X0 U18345 ( .IN1(n17714), .IN2(n4563), .QN(n17799) );
  INVX0 U18346 ( .INP(n17800), .ZN(n17798) );
  NOR2X0 U18347 ( .IN1(n17714), .IN2(n9837), .QN(n17800) );
  NAND2X0 U18348 ( .IN1(n17801), .IN2(n17802), .QN(g22152) );
  NAND2X0 U18349 ( .IN1(n17772), .IN2(g1545), .QN(n17802) );
  NAND2X0 U18350 ( .IN1(n17773), .IN2(n12132), .QN(n17801) );
  INVX0 U18351 ( .INP(n13626), .ZN(n12132) );
  NAND2X0 U18352 ( .IN1(n17803), .IN2(n17804), .QN(n13626) );
  NAND2X0 U18353 ( .IN1(n9908), .IN2(g6782), .QN(n17804) );
  NOR2X0 U18354 ( .IN1(n17805), .IN2(n17806), .QN(n17803) );
  NOR2X0 U18355 ( .IN1(test_so54), .IN2(n4368), .QN(n17806) );
  NOR2X0 U18356 ( .IN1(n4317), .IN2(g1554), .QN(n17805) );
  NAND2X0 U18357 ( .IN1(n17807), .IN2(n17808), .QN(g22151) );
  INVX0 U18358 ( .INP(n17809), .ZN(n17808) );
  NOR2X0 U18359 ( .IN1(n17743), .IN2(n9829), .QN(n17809) );
  NAND2X0 U18360 ( .IN1(n17743), .IN2(n12365), .QN(n17807) );
  NAND2X0 U18361 ( .IN1(n17810), .IN2(n17811), .QN(g22150) );
  NAND2X0 U18362 ( .IN1(n17727), .IN2(n4288), .QN(n17811) );
  INVX0 U18363 ( .INP(n17812), .ZN(n17810) );
  NOR2X0 U18364 ( .IN1(n17727), .IN2(n9847), .QN(n17812) );
  NAND2X0 U18365 ( .IN1(n17813), .IN2(n17814), .QN(g22149) );
  NAND2X0 U18366 ( .IN1(n17773), .IN2(n4378), .QN(n17814) );
  NAND2X0 U18367 ( .IN1(n17772), .IN2(g1512), .QN(n17813) );
  NAND2X0 U18368 ( .IN1(n17815), .IN2(n17816), .QN(g22148) );
  NAND2X0 U18369 ( .IN1(n17782), .IN2(g852), .QN(n17816) );
  NAND2X0 U18370 ( .IN1(n17781), .IN2(n12178), .QN(n17815) );
  NAND2X0 U18371 ( .IN1(n17817), .IN2(n17818), .QN(g22147) );
  INVX0 U18372 ( .INP(n17819), .ZN(n17818) );
  NOR2X0 U18373 ( .IN1(n17132), .IN2(n9858), .QN(n17819) );
  NAND2X0 U18374 ( .IN1(n13804), .IN2(n17132), .QN(n17817) );
  NAND2X0 U18375 ( .IN1(n17820), .IN2(n17821), .QN(g22146) );
  NAND2X0 U18376 ( .IN1(n17822), .IN2(n4375), .QN(n17821) );
  NAND2X0 U18377 ( .IN1(n17823), .IN2(g821), .QN(n17820) );
  NAND2X0 U18378 ( .IN1(n17824), .IN2(n17825), .QN(g22145) );
  NAND2X0 U18379 ( .IN1(n17781), .IN2(n4379), .QN(n17825) );
  NAND2X0 U18380 ( .IN1(n17782), .IN2(g819), .QN(n17824) );
  NAND2X0 U18381 ( .IN1(n17826), .IN2(n17827), .QN(g22143) );
  NAND2X0 U18382 ( .IN1(n17137), .IN2(g162), .QN(n17827) );
  NAND2X0 U18383 ( .IN1(n17788), .IN2(n12247), .QN(n17826) );
  NAND2X0 U18384 ( .IN1(n17828), .IN2(n17829), .QN(g22142) );
  NAND2X0 U18385 ( .IN1(n17830), .IN2(n4376), .QN(n17829) );
  NAND2X0 U18386 ( .IN1(n17831), .IN2(g134), .QN(n17828) );
  NAND2X0 U18387 ( .IN1(n17832), .IN2(n17833), .QN(g22141) );
  NAND2X0 U18388 ( .IN1(n4380), .IN2(n17788), .QN(n17833) );
  INVX0 U18389 ( .INP(n17834), .ZN(n17832) );
  NOR2X0 U18390 ( .IN1(n17788), .IN2(n9877), .QN(n17834) );
  NAND2X0 U18391 ( .IN1(n17835), .IN2(n17836), .QN(g22140) );
  NAND2X0 U18392 ( .IN1(n17735), .IN2(n4287), .QN(n17836) );
  NAND2X0 U18393 ( .IN1(n17736), .IN2(g2233), .QN(n17835) );
  NAND2X0 U18394 ( .IN1(n17837), .IN2(n17838), .QN(g22139) );
  NAND2X0 U18395 ( .IN1(n17720), .IN2(n4563), .QN(n17838) );
  NAND2X0 U18396 ( .IN1(n17721), .IN2(g2231), .QN(n17837) );
  NAND2X0 U18397 ( .IN1(n17839), .IN2(n17840), .QN(g22138) );
  NAND2X0 U18398 ( .IN1(n17714), .IN2(n4555), .QN(n17840) );
  INVX0 U18399 ( .INP(n17841), .ZN(n17839) );
  NOR2X0 U18400 ( .IN1(n17714), .IN2(n9838), .QN(n17841) );
  NAND2X0 U18401 ( .IN1(n17842), .IN2(n17843), .QN(g22132) );
  NAND2X0 U18402 ( .IN1(n17772), .IN2(g1542), .QN(n17843) );
  NAND2X0 U18403 ( .IN1(n17773), .IN2(n12365), .QN(n17842) );
  INVX0 U18404 ( .INP(n13660), .ZN(n12365) );
  NAND2X0 U18405 ( .IN1(n17844), .IN2(n17845), .QN(n13660) );
  NAND2X0 U18406 ( .IN1(n9906), .IN2(g6782), .QN(n17845) );
  NOR2X0 U18407 ( .IN1(n17846), .IN2(n17847), .QN(n17844) );
  NOR2X0 U18408 ( .IN1(n4368), .IN2(g1556), .QN(n17847) );
  NOR2X0 U18409 ( .IN1(n4317), .IN2(g1557), .QN(n17846) );
  NAND2X0 U18410 ( .IN1(n17848), .IN2(n17849), .QN(g22131) );
  NAND2X0 U18411 ( .IN1(n17743), .IN2(n4288), .QN(n17849) );
  NAND2X0 U18412 ( .IN1(n17744), .IN2(g1540), .QN(n17848) );
  NAND2X0 U18413 ( .IN1(n17850), .IN2(n17851), .QN(g22130) );
  NAND2X0 U18414 ( .IN1(n17727), .IN2(n4565), .QN(n17851) );
  NAND2X0 U18415 ( .IN1(n17127), .IN2(g1535), .QN(n17850) );
  INVX0 U18416 ( .INP(n17727), .ZN(n17127) );
  NAND2X0 U18417 ( .IN1(n17852), .IN2(n17853), .QN(g22129) );
  NAND2X0 U18418 ( .IN1(n17823), .IN2(g851), .QN(n17853) );
  NAND2X0 U18419 ( .IN1(n17822), .IN2(n12178), .QN(n17852) );
  INVX0 U18420 ( .INP(n13796), .ZN(n12178) );
  NAND2X0 U18421 ( .IN1(n17854), .IN2(n17855), .QN(n13796) );
  NAND2X0 U18422 ( .IN1(n9919), .IN2(test_so31), .QN(n17855) );
  NOR2X0 U18423 ( .IN1(n17856), .IN2(n17857), .QN(n17854) );
  NOR2X0 U18424 ( .IN1(n4323), .IN2(g860), .QN(n17857) );
  NOR2X0 U18425 ( .IN1(n4312), .IN2(g861), .QN(n17856) );
  NAND2X0 U18426 ( .IN1(n17858), .IN2(n17859), .QN(g22128) );
  NAND2X0 U18427 ( .IN1(n17782), .IN2(g849), .QN(n17859) );
  NAND2X0 U18428 ( .IN1(n17781), .IN2(n13804), .QN(n17858) );
  NAND2X0 U18429 ( .IN1(n17860), .IN2(n17861), .QN(g22127) );
  NAND2X0 U18430 ( .IN1(n4289), .IN2(n17132), .QN(n17861) );
  INVX0 U18431 ( .INP(n17862), .ZN(n17860) );
  NOR2X0 U18432 ( .IN1(n17132), .IN2(n9861), .QN(n17862) );
  NAND2X0 U18433 ( .IN1(n17863), .IN2(n17864), .QN(g22126) );
  NAND2X0 U18434 ( .IN1(n17822), .IN2(n4379), .QN(n17864) );
  NAND2X0 U18435 ( .IN1(n17823), .IN2(g818), .QN(n17863) );
  NAND2X0 U18436 ( .IN1(n17865), .IN2(n17866), .QN(g22125) );
  INVX0 U18437 ( .INP(n17867), .ZN(n17866) );
  NOR2X0 U18438 ( .IN1(n17830), .IN2(n9870), .QN(n17867) );
  NAND2X0 U18439 ( .IN1(n17830), .IN2(n12247), .QN(n17865) );
  NAND2X0 U18440 ( .IN1(n17868), .IN2(n17869), .QN(g22124) );
  NAND2X0 U18441 ( .IN1(n17137), .IN2(g159), .QN(n17869) );
  NAND2X0 U18442 ( .IN1(n12454), .IN2(n17788), .QN(n17868) );
  NAND2X0 U18443 ( .IN1(n17870), .IN2(n17871), .QN(g22123) );
  NAND2X0 U18444 ( .IN1(n17872), .IN2(n4376), .QN(n17871) );
  NAND2X0 U18445 ( .IN1(n17873), .IN2(g133), .QN(n17870) );
  NAND2X0 U18446 ( .IN1(n17874), .IN2(n17875), .QN(g22122) );
  NAND2X0 U18447 ( .IN1(n17830), .IN2(n4380), .QN(n17875) );
  NAND2X0 U18448 ( .IN1(n17831), .IN2(g131), .QN(n17874) );
  NAND2X0 U18449 ( .IN1(n17876), .IN2(n17877), .QN(g22117) );
  NAND2X0 U18450 ( .IN1(n17735), .IN2(n4563), .QN(n17877) );
  NAND2X0 U18451 ( .IN1(n17736), .IN2(g2230), .QN(n17876) );
  NAND2X0 U18452 ( .IN1(n17878), .IN2(n17879), .QN(g22116) );
  NAND2X0 U18453 ( .IN1(n17720), .IN2(n4555), .QN(n17879) );
  NAND2X0 U18454 ( .IN1(n17721), .IN2(g2228), .QN(n17878) );
  NAND2X0 U18455 ( .IN1(n17880), .IN2(n17881), .QN(g22115) );
  NAND2X0 U18456 ( .IN1(n17714), .IN2(n4325), .QN(n17881) );
  NAND2X0 U18457 ( .IN1(n17122), .IN2(g2223), .QN(n17880) );
  INVX0 U18458 ( .INP(n17714), .ZN(n17122) );
  NAND2X0 U18459 ( .IN1(n17882), .IN2(n17883), .QN(g22114) );
  NAND2X0 U18460 ( .IN1(n17773), .IN2(n4288), .QN(n17883) );
  NAND2X0 U18461 ( .IN1(n17772), .IN2(g1539), .QN(n17882) );
  NAND2X0 U18462 ( .IN1(n17884), .IN2(n17885), .QN(g22113) );
  NAND2X0 U18463 ( .IN1(test_so53), .IN2(n17744), .QN(n17885) );
  NAND2X0 U18464 ( .IN1(n17743), .IN2(n4565), .QN(n17884) );
  NAND2X0 U18465 ( .IN1(n17886), .IN2(n17887), .QN(g22112) );
  NAND2X0 U18466 ( .IN1(n17727), .IN2(n4557), .QN(n17887) );
  INVX0 U18467 ( .INP(n17888), .ZN(n17886) );
  NOR2X0 U18468 ( .IN1(n17727), .IN2(n9849), .QN(n17888) );
  NAND2X0 U18469 ( .IN1(n17889), .IN2(n17890), .QN(g22106) );
  NAND2X0 U18470 ( .IN1(n17823), .IN2(g848), .QN(n17890) );
  NAND2X0 U18471 ( .IN1(n17822), .IN2(n13804), .QN(n17889) );
  INVX0 U18472 ( .INP(n12419), .ZN(n13804) );
  NAND2X0 U18473 ( .IN1(n17891), .IN2(n17892), .QN(n12419) );
  NAND2X0 U18474 ( .IN1(n9916), .IN2(test_so31), .QN(n17892) );
  NOR2X0 U18475 ( .IN1(n17893), .IN2(n17894), .QN(n17891) );
  NOR2X0 U18476 ( .IN1(n4323), .IN2(g863), .QN(n17894) );
  NOR2X0 U18477 ( .IN1(n4312), .IN2(g864), .QN(n17893) );
  NAND2X0 U18478 ( .IN1(n17895), .IN2(n17896), .QN(g22105) );
  NAND2X0 U18479 ( .IN1(n17781), .IN2(n4289), .QN(n17896) );
  NAND2X0 U18480 ( .IN1(n17782), .IN2(g846), .QN(n17895) );
  NAND2X0 U18481 ( .IN1(n17897), .IN2(n17898), .QN(g22104) );
  NAND2X0 U18482 ( .IN1(n17132), .IN2(n4567), .QN(n17898) );
  INVX0 U18483 ( .INP(n17899), .ZN(n17897) );
  NOR2X0 U18484 ( .IN1(n17132), .IN2(n9862), .QN(n17899) );
  NAND2X0 U18485 ( .IN1(n17900), .IN2(n17901), .QN(g22103) );
  NAND2X0 U18486 ( .IN1(test_so12), .IN2(n17873), .QN(n17901) );
  NAND2X0 U18487 ( .IN1(n17872), .IN2(n12247), .QN(n17900) );
  INVX0 U18488 ( .INP(n13898), .ZN(n12247) );
  NAND2X0 U18489 ( .IN1(n17902), .IN2(n17903), .QN(n13898) );
  NAND2X0 U18490 ( .IN1(n9931), .IN2(g6313), .QN(n17903) );
  NOR2X0 U18491 ( .IN1(n17904), .IN2(n17905), .QN(n17902) );
  NOR2X0 U18492 ( .IN1(n4369), .IN2(g171), .QN(n17905) );
  NOR2X0 U18493 ( .IN1(n4318), .IN2(g172), .QN(n17904) );
  NAND2X0 U18494 ( .IN1(n17906), .IN2(n17907), .QN(g22102) );
  INVX0 U18495 ( .INP(n17908), .ZN(n17907) );
  NOR2X0 U18496 ( .IN1(n17830), .IN2(n9832), .QN(n17908) );
  NAND2X0 U18497 ( .IN1(n17830), .IN2(n12454), .QN(n17906) );
  NAND2X0 U18498 ( .IN1(n17909), .IN2(n17910), .QN(g22101) );
  NAND2X0 U18499 ( .IN1(n4290), .IN2(n17788), .QN(n17910) );
  INVX0 U18500 ( .INP(n17911), .ZN(n17909) );
  NOR2X0 U18501 ( .IN1(n17788), .IN2(n9871), .QN(n17911) );
  NAND2X0 U18502 ( .IN1(n17912), .IN2(n17913), .QN(g22100) );
  NAND2X0 U18503 ( .IN1(n17872), .IN2(n4380), .QN(n17913) );
  NAND2X0 U18504 ( .IN1(n17873), .IN2(g130), .QN(n17912) );
  NAND2X0 U18505 ( .IN1(n17914), .IN2(n17915), .QN(g22099) );
  NAND2X0 U18506 ( .IN1(n17735), .IN2(n4555), .QN(n17915) );
  NAND2X0 U18507 ( .IN1(n17736), .IN2(g2227), .QN(n17914) );
  NAND2X0 U18508 ( .IN1(n17916), .IN2(n17917), .QN(g22098) );
  NAND2X0 U18509 ( .IN1(test_so74), .IN2(n17721), .QN(n17917) );
  NAND2X0 U18510 ( .IN1(n17720), .IN2(n4325), .QN(n17916) );
  NAND2X0 U18511 ( .IN1(n17918), .IN2(n17919), .QN(g22097) );
  NAND2X0 U18512 ( .IN1(n17714), .IN2(n4389), .QN(n17919) );
  INVX0 U18513 ( .INP(n17920), .ZN(n17918) );
  NOR2X0 U18514 ( .IN1(n17714), .IN2(n9840), .QN(n17920) );
  NAND2X0 U18515 ( .IN1(n17921), .IN2(n17922), .QN(g22092) );
  NAND2X0 U18516 ( .IN1(n17773), .IN2(n4565), .QN(n17922) );
  NAND2X0 U18517 ( .IN1(n17772), .IN2(g1536), .QN(n17921) );
  NAND2X0 U18518 ( .IN1(n17923), .IN2(n17924), .QN(g22091) );
  NAND2X0 U18519 ( .IN1(n17743), .IN2(n4557), .QN(n17924) );
  NAND2X0 U18520 ( .IN1(n17744), .IN2(g1534), .QN(n17923) );
  NAND2X0 U18521 ( .IN1(n17925), .IN2(n17926), .QN(g22090) );
  NAND2X0 U18522 ( .IN1(n17727), .IN2(n4326), .QN(n17926) );
  INVX0 U18523 ( .INP(n17927), .ZN(n17925) );
  NOR2X0 U18524 ( .IN1(n17727), .IN2(n9850), .QN(n17927) );
  NAND2X0 U18525 ( .IN1(n17928), .IN2(n17929), .QN(g22089) );
  NAND2X0 U18526 ( .IN1(n17822), .IN2(n4289), .QN(n17929) );
  NAND2X0 U18527 ( .IN1(n17823), .IN2(g845), .QN(n17928) );
  NAND2X0 U18528 ( .IN1(n17930), .IN2(n17931), .QN(g22088) );
  NAND2X0 U18529 ( .IN1(n17781), .IN2(n4567), .QN(n17931) );
  NAND2X0 U18530 ( .IN1(n17782), .IN2(g843), .QN(n17930) );
  NAND2X0 U18531 ( .IN1(n17932), .IN2(n17933), .QN(g22087) );
  NAND2X0 U18532 ( .IN1(n17132), .IN2(n4559), .QN(n17933) );
  INVX0 U18533 ( .INP(n17934), .ZN(n17932) );
  NOR2X0 U18534 ( .IN1(n17132), .IN2(n9863), .QN(n17934) );
  NAND2X0 U18535 ( .IN1(n17935), .IN2(n17936), .QN(g22081) );
  NAND2X0 U18536 ( .IN1(n17873), .IN2(g160), .QN(n17936) );
  NAND2X0 U18537 ( .IN1(n17872), .IN2(n12454), .QN(n17935) );
  INVX0 U18538 ( .INP(n13931), .ZN(n12454) );
  NAND2X0 U18539 ( .IN1(n17937), .IN2(n17938), .QN(n13931) );
  NAND2X0 U18540 ( .IN1(n9928), .IN2(g6313), .QN(n17938) );
  NOR2X0 U18541 ( .IN1(n17939), .IN2(n17940), .QN(n17937) );
  NOR2X0 U18542 ( .IN1(n4369), .IN2(g174), .QN(n17940) );
  NOR2X0 U18543 ( .IN1(n4318), .IN2(g175), .QN(n17939) );
  NAND2X0 U18544 ( .IN1(n17941), .IN2(n17942), .QN(g22080) );
  NAND2X0 U18545 ( .IN1(n17830), .IN2(n4290), .QN(n17942) );
  NAND2X0 U18546 ( .IN1(n17831), .IN2(g158), .QN(n17941) );
  NAND2X0 U18547 ( .IN1(n17943), .IN2(n17944), .QN(g22079) );
  NAND2X0 U18548 ( .IN1(n17788), .IN2(n4569), .QN(n17944) );
  INVX0 U18549 ( .INP(n17945), .ZN(n17943) );
  NOR2X0 U18550 ( .IN1(n17788), .IN2(n9872), .QN(n17945) );
  NAND2X0 U18551 ( .IN1(n17946), .IN2(n17947), .QN(g22078) );
  NAND2X0 U18552 ( .IN1(n17735), .IN2(n4325), .QN(n17947) );
  NAND2X0 U18553 ( .IN1(n17736), .IN2(g2224), .QN(n17946) );
  NAND2X0 U18554 ( .IN1(n17948), .IN2(n17949), .QN(g22077) );
  NAND2X0 U18555 ( .IN1(n17720), .IN2(n4389), .QN(n17949) );
  NAND2X0 U18556 ( .IN1(n17721), .IN2(g2222), .QN(n17948) );
  NAND2X0 U18557 ( .IN1(n17950), .IN2(n17951), .QN(g22076) );
  NAND2X0 U18558 ( .IN1(n17714), .IN2(n4319), .QN(n17951) );
  INVX0 U18559 ( .INP(n17952), .ZN(n17950) );
  NOR2X0 U18560 ( .IN1(n17714), .IN2(n9841), .QN(n17952) );
  NOR2X0 U18561 ( .IN1(n10029), .IN2(n4367), .QN(n17714) );
  NAND2X0 U18562 ( .IN1(n17953), .IN2(n17954), .QN(g22075) );
  NAND2X0 U18563 ( .IN1(n17773), .IN2(n4557), .QN(n17954) );
  NAND2X0 U18564 ( .IN1(n17772), .IN2(g1533), .QN(n17953) );
  NAND2X0 U18565 ( .IN1(n17955), .IN2(n17956), .QN(g22074) );
  NAND2X0 U18566 ( .IN1(n17743), .IN2(n4326), .QN(n17956) );
  NAND2X0 U18567 ( .IN1(n17744), .IN2(g1531), .QN(n17955) );
  NAND2X0 U18568 ( .IN1(n17957), .IN2(n17958), .QN(g22073) );
  NAND2X0 U18569 ( .IN1(n17727), .IN2(n4390), .QN(n17958) );
  INVX0 U18570 ( .INP(n17959), .ZN(n17957) );
  NOR2X0 U18571 ( .IN1(n17727), .IN2(n9851), .QN(n17959) );
  NAND2X0 U18572 ( .IN1(n17960), .IN2(n17961), .QN(g22068) );
  NAND2X0 U18573 ( .IN1(n17822), .IN2(n4567), .QN(n17961) );
  NAND2X0 U18574 ( .IN1(n17823), .IN2(g842), .QN(n17960) );
  NAND2X0 U18575 ( .IN1(n17962), .IN2(n17963), .QN(g22067) );
  NAND2X0 U18576 ( .IN1(n17781), .IN2(n4559), .QN(n17963) );
  NAND2X0 U18577 ( .IN1(n17782), .IN2(g840), .QN(n17962) );
  NAND2X0 U18578 ( .IN1(n17964), .IN2(n17965), .QN(g22066) );
  NAND2X0 U18579 ( .IN1(n4327), .IN2(n17132), .QN(n17965) );
  INVX0 U18580 ( .INP(n17966), .ZN(n17964) );
  NOR2X0 U18581 ( .IN1(n17132), .IN2(n9864), .QN(n17966) );
  NAND2X0 U18582 ( .IN1(n17967), .IN2(n17968), .QN(g22065) );
  NAND2X0 U18583 ( .IN1(n17872), .IN2(n4290), .QN(n17968) );
  NAND2X0 U18584 ( .IN1(n17873), .IN2(g157), .QN(n17967) );
  NAND2X0 U18585 ( .IN1(n17969), .IN2(n17970), .QN(g22064) );
  NAND2X0 U18586 ( .IN1(n17830), .IN2(n4569), .QN(n17970) );
  NAND2X0 U18587 ( .IN1(n17831), .IN2(g155), .QN(n17969) );
  NAND2X0 U18588 ( .IN1(n17971), .IN2(n17972), .QN(g22063) );
  NAND2X0 U18589 ( .IN1(n17788), .IN2(n4561), .QN(n17972) );
  INVX0 U18590 ( .INP(n17973), .ZN(n17971) );
  NOR2X0 U18591 ( .IN1(n17788), .IN2(n9873), .QN(n17973) );
  NAND2X0 U18592 ( .IN1(n17974), .IN2(n17975), .QN(g22061) );
  NAND2X0 U18593 ( .IN1(n17735), .IN2(n4389), .QN(n17975) );
  NAND2X0 U18594 ( .IN1(n17736), .IN2(g2221), .QN(n17974) );
  NAND2X0 U18595 ( .IN1(n17976), .IN2(n17977), .QN(g22060) );
  NAND2X0 U18596 ( .IN1(n17720), .IN2(n4319), .QN(n17977) );
  NAND2X0 U18597 ( .IN1(n17721), .IN2(g2219), .QN(n17976) );
  INVX0 U18598 ( .INP(n17720), .ZN(n17721) );
  NOR2X0 U18599 ( .IN1(n10320), .IN2(n10029), .QN(n17720) );
  NAND2X0 U18600 ( .IN1(n17978), .IN2(n17979), .QN(g22059) );
  NAND2X0 U18601 ( .IN1(n17773), .IN2(n4326), .QN(n17979) );
  NAND2X0 U18602 ( .IN1(n17772), .IN2(g1530), .QN(n17978) );
  NAND2X0 U18603 ( .IN1(n17980), .IN2(n17981), .QN(g22058) );
  NAND2X0 U18604 ( .IN1(n17743), .IN2(n4390), .QN(n17981) );
  NAND2X0 U18605 ( .IN1(n17744), .IN2(g1528), .QN(n17980) );
  NAND2X0 U18606 ( .IN1(n17982), .IN2(n17983), .QN(g22057) );
  NAND2X0 U18607 ( .IN1(n17727), .IN2(n4320), .QN(n17983) );
  INVX0 U18608 ( .INP(n17984), .ZN(n17982) );
  NOR2X0 U18609 ( .IN1(n17727), .IN2(n9852), .QN(n17984) );
  NOR2X0 U18610 ( .IN1(n10030), .IN2(n4368), .QN(n17727) );
  NAND2X0 U18611 ( .IN1(n17985), .IN2(n17986), .QN(g22056) );
  NAND2X0 U18612 ( .IN1(test_so32), .IN2(n17823), .QN(n17986) );
  NAND2X0 U18613 ( .IN1(n17822), .IN2(n4559), .QN(n17985) );
  NAND2X0 U18614 ( .IN1(n17987), .IN2(n17988), .QN(g22055) );
  NAND2X0 U18615 ( .IN1(n17781), .IN2(n4327), .QN(n17988) );
  NAND2X0 U18616 ( .IN1(n17782), .IN2(g837), .QN(n17987) );
  NAND2X0 U18617 ( .IN1(n17989), .IN2(n17990), .QN(g22054) );
  NAND2X0 U18618 ( .IN1(n17132), .IN2(n4391), .QN(n17990) );
  INVX0 U18619 ( .INP(n17991), .ZN(n17989) );
  NOR2X0 U18620 ( .IN1(n17132), .IN2(n9865), .QN(n17991) );
  NAND2X0 U18621 ( .IN1(n17992), .IN2(n17993), .QN(g22049) );
  NAND2X0 U18622 ( .IN1(n17872), .IN2(n4569), .QN(n17993) );
  NAND2X0 U18623 ( .IN1(n17873), .IN2(g154), .QN(n17992) );
  NAND2X0 U18624 ( .IN1(n17994), .IN2(n17995), .QN(g22048) );
  NAND2X0 U18625 ( .IN1(n17830), .IN2(n4561), .QN(n17995) );
  NAND2X0 U18626 ( .IN1(n17831), .IN2(g152), .QN(n17994) );
  NAND2X0 U18627 ( .IN1(n17996), .IN2(n17997), .QN(g22047) );
  NAND2X0 U18628 ( .IN1(n4328), .IN2(n17788), .QN(n17997) );
  INVX0 U18629 ( .INP(n17998), .ZN(n17996) );
  NOR2X0 U18630 ( .IN1(n17788), .IN2(n9874), .QN(n17998) );
  NAND2X0 U18631 ( .IN1(n17999), .IN2(n18000), .QN(g22045) );
  NAND2X0 U18632 ( .IN1(n17735), .IN2(n4319), .QN(n18000) );
  NAND2X0 U18633 ( .IN1(n17736), .IN2(g2218), .QN(n17999) );
  INVX0 U18634 ( .INP(n17735), .ZN(n17736) );
  NOR2X0 U18635 ( .IN1(n10029), .IN2(n4324), .QN(n17735) );
  NAND2X0 U18636 ( .IN1(n18001), .IN2(n18002), .QN(g22044) );
  NAND2X0 U18637 ( .IN1(n17773), .IN2(n4390), .QN(n18002) );
  NAND2X0 U18638 ( .IN1(n17772), .IN2(g1527), .QN(n18001) );
  NAND2X0 U18639 ( .IN1(n18003), .IN2(n18004), .QN(g22043) );
  NAND2X0 U18640 ( .IN1(n17743), .IN2(n4320), .QN(n18004) );
  NAND2X0 U18641 ( .IN1(n17744), .IN2(g1525), .QN(n18003) );
  INVX0 U18642 ( .INP(n17743), .ZN(n17744) );
  NOR2X0 U18643 ( .IN1(n10030), .IN2(n4515), .QN(n17743) );
  NAND2X0 U18644 ( .IN1(n18005), .IN2(n18006), .QN(g22042) );
  NAND2X0 U18645 ( .IN1(n17822), .IN2(n4327), .QN(n18006) );
  NAND2X0 U18646 ( .IN1(n17823), .IN2(g836), .QN(n18005) );
  NAND2X0 U18647 ( .IN1(n18007), .IN2(n18008), .QN(g22041) );
  NAND2X0 U18648 ( .IN1(n17781), .IN2(n4391), .QN(n18008) );
  NAND2X0 U18649 ( .IN1(n17782), .IN2(g834), .QN(n18007) );
  NAND2X0 U18650 ( .IN1(n18009), .IN2(n18010), .QN(g22040) );
  NAND2X0 U18651 ( .IN1(n4321), .IN2(n17132), .QN(n18010) );
  INVX0 U18652 ( .INP(n18011), .ZN(n18009) );
  NOR2X0 U18653 ( .IN1(n17132), .IN2(n9866), .QN(n18011) );
  NOR2X0 U18654 ( .IN1(n10321), .IN2(n10031), .QN(n17132) );
  NAND2X0 U18655 ( .IN1(n18012), .IN2(n18013), .QN(g22039) );
  NAND2X0 U18656 ( .IN1(n17872), .IN2(n4561), .QN(n18013) );
  NAND2X0 U18657 ( .IN1(n17873), .IN2(g151), .QN(n18012) );
  NAND2X0 U18658 ( .IN1(n18014), .IN2(n18015), .QN(g22038) );
  NAND2X0 U18659 ( .IN1(n17830), .IN2(n4328), .QN(n18015) );
  NAND2X0 U18660 ( .IN1(n17831), .IN2(g149), .QN(n18014) );
  NAND2X0 U18661 ( .IN1(n18016), .IN2(n18017), .QN(g22037) );
  NAND2X0 U18662 ( .IN1(test_so11), .IN2(n17137), .QN(n18017) );
  INVX0 U18663 ( .INP(n17788), .ZN(n17137) );
  NAND2X0 U18664 ( .IN1(n17788), .IN2(n4392), .QN(n18016) );
  NAND2X0 U18665 ( .IN1(n18018), .IN2(n18019), .QN(g22035) );
  NAND2X0 U18666 ( .IN1(n17773), .IN2(n4320), .QN(n18019) );
  NAND2X0 U18667 ( .IN1(n17772), .IN2(g1524), .QN(n18018) );
  INVX0 U18668 ( .INP(n17773), .ZN(n17772) );
  NOR2X0 U18669 ( .IN1(n10030), .IN2(n4317), .QN(n17773) );
  NAND2X0 U18670 ( .IN1(n18020), .IN2(n18021), .QN(g22034) );
  NAND2X0 U18671 ( .IN1(n17822), .IN2(n4391), .QN(n18021) );
  NAND2X0 U18672 ( .IN1(n17823), .IN2(g833), .QN(n18020) );
  NAND2X0 U18673 ( .IN1(n18022), .IN2(n18023), .QN(g22033) );
  NAND2X0 U18674 ( .IN1(n17781), .IN2(n4321), .QN(n18023) );
  NAND2X0 U18675 ( .IN1(n17782), .IN2(g831), .QN(n18022) );
  INVX0 U18676 ( .INP(n17781), .ZN(n17782) );
  NOR2X0 U18677 ( .IN1(n10031), .IN2(n4312), .QN(n17781) );
  NAND2X0 U18678 ( .IN1(n18024), .IN2(n18025), .QN(g22032) );
  NAND2X0 U18679 ( .IN1(n17872), .IN2(n4328), .QN(n18025) );
  NAND2X0 U18680 ( .IN1(n17873), .IN2(g148), .QN(n18024) );
  NAND2X0 U18681 ( .IN1(n18026), .IN2(n18027), .QN(g22031) );
  NAND2X0 U18682 ( .IN1(n17830), .IN2(n4392), .QN(n18027) );
  NAND2X0 U18683 ( .IN1(n17831), .IN2(g146), .QN(n18026) );
  NAND2X0 U18684 ( .IN1(n18028), .IN2(n18029), .QN(g22030) );
  NAND2X0 U18685 ( .IN1(n4322), .IN2(n17788), .QN(n18029) );
  INVX0 U18686 ( .INP(n18030), .ZN(n18028) );
  NOR2X0 U18687 ( .IN1(n17788), .IN2(n9875), .QN(n18030) );
  NOR2X0 U18688 ( .IN1(n10032), .IN2(n4369), .QN(n17788) );
  NAND2X0 U18689 ( .IN1(n18031), .IN2(n18032), .QN(g22029) );
  NAND2X0 U18690 ( .IN1(n17822), .IN2(n4321), .QN(n18032) );
  NAND2X0 U18691 ( .IN1(n17823), .IN2(g830), .QN(n18031) );
  INVX0 U18692 ( .INP(n17822), .ZN(n17823) );
  NOR2X0 U18693 ( .IN1(n10031), .IN2(n4323), .QN(n17822) );
  NAND2X0 U18694 ( .IN1(n18033), .IN2(n18034), .QN(g22028) );
  NAND2X0 U18695 ( .IN1(n17872), .IN2(n4392), .QN(n18034) );
  NAND2X0 U18696 ( .IN1(n17873), .IN2(g145), .QN(n18033) );
  NAND2X0 U18697 ( .IN1(n18035), .IN2(n18036), .QN(g22027) );
  NAND2X0 U18698 ( .IN1(n17830), .IN2(n4322), .QN(n18036) );
  NAND2X0 U18699 ( .IN1(n17831), .IN2(g143), .QN(n18035) );
  INVX0 U18700 ( .INP(n17830), .ZN(n17831) );
  NOR2X0 U18701 ( .IN1(n10032), .IN2(n4512), .QN(n17830) );
  NOR2X0 U18702 ( .IN1(n10998), .IN2(n18037), .QN(g22026) );
  NAND2X0 U18703 ( .IN1(n4123), .IN2(n18038), .QN(n18037) );
  INVX0 U18704 ( .INP(n18039), .ZN(n18038) );
  NOR2X0 U18705 ( .IN1(g2888), .IN2(n18040), .QN(n18039) );
  NAND2X0 U18706 ( .IN1(n18040), .IN2(g2888), .QN(n4123) );
  NOR2X0 U18707 ( .IN1(n4423), .IN2(n4330), .QN(n18040) );
  NAND2X0 U18708 ( .IN1(n18867), .IN2(n11005), .QN(n10998) );
  NAND2X0 U18709 ( .IN1(n18041), .IN2(n18042), .QN(n11005) );
  NOR2X0 U18710 ( .IN1(n18043), .IN2(n18044), .QN(n18042) );
  NAND2X0 U18711 ( .IN1(n4291), .IN2(g2888), .QN(n18044) );
  NAND2X0 U18712 ( .IN1(g2908), .IN2(g2950), .QN(n18043) );
  NOR2X0 U18713 ( .IN1(g2883), .IN2(n18045), .QN(n18041) );
  NAND2X0 U18714 ( .IN1(n4182), .IN2(n4431), .QN(n18045) );
  NAND2X0 U18715 ( .IN1(n18046), .IN2(n18047), .QN(g22025) );
  NAND2X0 U18716 ( .IN1(n17872), .IN2(n4322), .QN(n18047) );
  NAND2X0 U18717 ( .IN1(n17873), .IN2(g142), .QN(n18046) );
  INVX0 U18718 ( .INP(n17872), .ZN(n17873) );
  NOR2X0 U18719 ( .IN1(n10032), .IN2(n4318), .QN(n17872) );
  NOR2X0 U18720 ( .IN1(n18048), .IN2(n18049), .QN(g21974) );
  NAND2X0 U18721 ( .IN1(n17349), .IN2(n14826), .QN(n18049) );
  NAND2X0 U18722 ( .IN1(n18050), .IN2(n18051), .QN(n17349) );
  NOR2X0 U18723 ( .IN1(n4472), .IN2(n4398), .QN(n18050) );
  NOR2X0 U18724 ( .IN1(n18052), .IN2(g2707), .QN(n18048) );
  NOR2X0 U18725 ( .IN1(n4398), .IN2(n18053), .QN(n18052) );
  NOR2X0 U18726 ( .IN1(n18054), .IN2(n18055), .QN(g21972) );
  NAND2X0 U18727 ( .IN1(n17355), .IN2(n14703), .QN(n18055) );
  NAND2X0 U18728 ( .IN1(n18056), .IN2(n18057), .QN(n17355) );
  NOR2X0 U18729 ( .IN1(n4474), .IN2(n4400), .QN(n18056) );
  NOR2X0 U18730 ( .IN1(n18058), .IN2(g2013), .QN(n18054) );
  NOR2X0 U18731 ( .IN1(n4400), .IN2(n18059), .QN(n18058) );
  NAND2X0 U18732 ( .IN1(n18060), .IN2(n18061), .QN(g21970) );
  NAND2X0 U18733 ( .IN1(test_so87), .IN2(n4463), .QN(n18061) );
  NAND2X0 U18734 ( .IN1(n14747), .IN2(g2560), .QN(n18060) );
  NAND2X0 U18735 ( .IN1(n18062), .IN2(n18063), .QN(n14747) );
  NAND2X0 U18736 ( .IN1(g5555), .IN2(g2513), .QN(n18063) );
  NOR2X0 U18737 ( .IN1(n18064), .IN2(n18065), .QN(n18062) );
  NOR2X0 U18738 ( .IN1(n9741), .IN2(n14010), .QN(n18065) );
  INVX0 U18739 ( .INP(g7264), .ZN(n14010) );
  NOR2X0 U18740 ( .IN1(n9752), .IN2(n15607), .QN(n18064) );
  INVX0 U18741 ( .INP(n4606), .ZN(n15607) );
  NOR2X0 U18742 ( .IN1(n18066), .IN2(n18067), .QN(g21969) );
  NAND2X0 U18743 ( .IN1(n17361), .IN2(n14834), .QN(n18067) );
  NAND2X0 U18744 ( .IN1(n18068), .IN2(n18069), .QN(n17361) );
  NOR2X0 U18745 ( .IN1(n4476), .IN2(n4402), .QN(n18068) );
  NOR2X0 U18746 ( .IN1(n18070), .IN2(g1319), .QN(n18066) );
  NOR2X0 U18747 ( .IN1(n4402), .IN2(n18071), .QN(n18070) );
  NAND2X0 U18748 ( .IN1(n18072), .IN2(n18073), .QN(g21882) );
  NAND2X0 U18749 ( .IN1(n4351), .IN2(g2878), .QN(n18073) );
  NAND2X0 U18750 ( .IN1(n18074), .IN2(g2879), .QN(n18072) );
  NAND2X0 U18751 ( .IN1(n18075), .IN2(n18076), .QN(g21880) );
  NAND2X0 U18752 ( .IN1(n4351), .IN2(g2877), .QN(n18076) );
  NAND2X0 U18753 ( .IN1(n18077), .IN2(g2879), .QN(n18075) );
  NAND2X0 U18754 ( .IN1(n18078), .IN2(n18079), .QN(g21878) );
  NAND2X0 U18755 ( .IN1(test_so4), .IN2(g2879), .QN(n18079) );
  NAND2X0 U18756 ( .IN1(n4351), .IN2(n18074), .QN(n18078) );
  NAND2X0 U18757 ( .IN1(n18080), .IN2(n18081), .QN(n18074) );
  NAND2X0 U18758 ( .IN1(n18082), .IN2(n10729), .QN(n18081) );
  INVX0 U18759 ( .INP(n18083), .ZN(n18080) );
  NOR2X0 U18760 ( .IN1(n10729), .IN2(n18082), .QN(n18083) );
  NOR2X0 U18761 ( .IN1(n18084), .IN2(n18085), .QN(n10729) );
  INVX0 U18762 ( .INP(n18086), .ZN(n18085) );
  NAND2X0 U18763 ( .IN1(n18087), .IN2(n18088), .QN(n18086) );
  NOR2X0 U18764 ( .IN1(n18088), .IN2(n18087), .QN(n18084) );
  NAND2X0 U18765 ( .IN1(n18089), .IN2(n18090), .QN(n18087) );
  INVX0 U18766 ( .INP(n18091), .ZN(n18090) );
  NOR2X0 U18767 ( .IN1(n18092), .IN2(n18093), .QN(n18091) );
  NAND2X0 U18768 ( .IN1(n18093), .IN2(n18092), .QN(n18089) );
  NOR2X0 U18769 ( .IN1(n18094), .IN2(n18095), .QN(n18092) );
  INVX0 U18770 ( .INP(n18096), .ZN(n18095) );
  NAND2X0 U18771 ( .IN1(test_so2), .IN2(g2981), .QN(n18096) );
  NOR2X0 U18772 ( .IN1(g2981), .IN2(test_so2), .QN(n18094) );
  NAND2X0 U18773 ( .IN1(n18097), .IN2(n18098), .QN(n18093) );
  NAND2X0 U18774 ( .IN1(n10286), .IN2(g2975), .QN(n18098) );
  NAND2X0 U18775 ( .IN1(n10285), .IN2(g2969), .QN(n18097) );
  NOR2X0 U18776 ( .IN1(n18099), .IN2(n18100), .QN(n18088) );
  NOR2X0 U18777 ( .IN1(n18101), .IN2(n18102), .QN(n18100) );
  INVX0 U18778 ( .INP(n18103), .ZN(n18099) );
  NAND2X0 U18779 ( .IN1(n18102), .IN2(n18101), .QN(n18103) );
  INVX0 U18780 ( .INP(n18104), .ZN(n18101) );
  NAND2X0 U18781 ( .IN1(n18105), .IN2(n18106), .QN(n18104) );
  NAND2X0 U18782 ( .IN1(n10284), .IN2(g2963), .QN(n18106) );
  NAND2X0 U18783 ( .IN1(n10283), .IN2(g2972), .QN(n18105) );
  NAND2X0 U18784 ( .IN1(n18107), .IN2(n18108), .QN(n18102) );
  NAND2X0 U18785 ( .IN1(n10282), .IN2(g2978), .QN(n18108) );
  NAND2X0 U18786 ( .IN1(n10281), .IN2(g2874), .QN(n18107) );
  NAND2X0 U18787 ( .IN1(n18109), .IN2(n18110), .QN(g21851) );
  NAND2X0 U18788 ( .IN1(g499), .IN2(g544), .QN(n18110) );
  NAND2X0 U18789 ( .IN1(n18111), .IN2(n4541), .QN(n18109) );
  NOR2X0 U18790 ( .IN1(n9416), .IN2(n14574), .QN(n18111) );
  NAND2X0 U18791 ( .IN1(n18112), .IN2(n18113), .QN(g21346) );
  NAND2X0 U18792 ( .IN1(n18872), .IN2(DFF_328_n1), .QN(n18113) );
  NAND2X0 U18793 ( .IN1(n18114), .IN2(n8056), .QN(n18112) );
  NOR2X0 U18794 ( .IN1(n9740), .IN2(g6447), .QN(n18114) );
  NAND2X0 U18795 ( .IN1(n18115), .IN2(n18116), .QN(g21094) );
  NAND2X0 U18796 ( .IN1(test_so94), .IN2(n16488), .QN(n18116) );
  NAND2X0 U18797 ( .IN1(n16490), .IN2(n4393), .QN(n18115) );
  NAND2X0 U18798 ( .IN1(n18117), .IN2(n18118), .QN(g21082) );
  NAND2X0 U18799 ( .IN1(n16494), .IN2(n4393), .QN(n18118) );
  NAND2X0 U18800 ( .IN1(n16493), .IN2(g2798), .QN(n18117) );
  NAND2X0 U18801 ( .IN1(n18119), .IN2(n18120), .QN(g21081) );
  NAND2X0 U18802 ( .IN1(n16490), .IN2(n4471), .QN(n18120) );
  INVX0 U18803 ( .INP(n18121), .ZN(n18119) );
  NOR2X0 U18804 ( .IN1(n16490), .IN2(n10156), .QN(n18121) );
  NAND2X0 U18805 ( .IN1(n18122), .IN2(n18123), .QN(g21080) );
  NAND2X0 U18806 ( .IN1(n16499), .IN2(n10323), .QN(n18123) );
  INVX0 U18807 ( .INP(n18124), .ZN(n18122) );
  NOR2X0 U18808 ( .IN1(n16499), .IN2(n10164), .QN(n18124) );
  NAND2X0 U18809 ( .IN1(n18125), .IN2(n18126), .QN(g21075) );
  NAND2X0 U18810 ( .IN1(n16503), .IN2(n4393), .QN(n18126) );
  NAND2X0 U18811 ( .IN1(n16502), .IN2(g2797), .QN(n18125) );
  NAND2X0 U18812 ( .IN1(n18127), .IN2(n18128), .QN(g21074) );
  NAND2X0 U18813 ( .IN1(n16494), .IN2(n4471), .QN(n18128) );
  NAND2X0 U18814 ( .IN1(n16493), .IN2(g2795), .QN(n18127) );
  NAND2X0 U18815 ( .IN1(n18129), .IN2(n18130), .QN(g21073) );
  NAND2X0 U18816 ( .IN1(n16490), .IN2(n10324), .QN(n18130) );
  INVX0 U18817 ( .INP(n18131), .ZN(n18129) );
  NOR2X0 U18818 ( .IN1(n16490), .IN2(n10157), .QN(n18131) );
  NAND2X0 U18819 ( .IN1(n18132), .IN2(n18133), .QN(g21072) );
  NAND2X0 U18820 ( .IN1(n16596), .IN2(n10323), .QN(n18133) );
  NAND2X0 U18821 ( .IN1(n16597), .IN2(g2104), .QN(n18132) );
  NAND2X0 U18822 ( .IN1(n18134), .IN2(n18135), .QN(g21071) );
  NAND2X0 U18823 ( .IN1(n16499), .IN2(n4473), .QN(n18135) );
  INVX0 U18824 ( .INP(n18136), .ZN(n18134) );
  NOR2X0 U18825 ( .IN1(n16499), .IN2(n10165), .QN(n18136) );
  NAND2X0 U18826 ( .IN1(n18137), .IN2(n18138), .QN(g21070) );
  NAND2X0 U18827 ( .IN1(n16602), .IN2(n4395), .QN(n18138) );
  INVX0 U18828 ( .INP(n18139), .ZN(n18137) );
  NOR2X0 U18829 ( .IN1(n16602), .IN2(n10174), .QN(n18139) );
  NAND2X0 U18830 ( .IN1(n18140), .IN2(n18141), .QN(g21063) );
  NAND2X0 U18831 ( .IN1(n18142), .IN2(g2805), .QN(n18141) );
  NAND2X0 U18832 ( .IN1(n17688), .IN2(n11275), .QN(n18140) );
  NAND2X0 U18833 ( .IN1(n18143), .IN2(n18144), .QN(g21062) );
  NAND2X0 U18834 ( .IN1(n16503), .IN2(n4471), .QN(n18144) );
  NAND2X0 U18835 ( .IN1(n16502), .IN2(g2794), .QN(n18143) );
  NAND2X0 U18836 ( .IN1(n18145), .IN2(n18146), .QN(g21061) );
  NAND2X0 U18837 ( .IN1(n16494), .IN2(n10324), .QN(n18146) );
  NAND2X0 U18838 ( .IN1(n16493), .IN2(g2792), .QN(n18145) );
  NAND2X0 U18839 ( .IN1(n18147), .IN2(n18148), .QN(g21060) );
  NAND2X0 U18840 ( .IN1(n16490), .IN2(n4407), .QN(n18148) );
  INVX0 U18841 ( .INP(n18149), .ZN(n18147) );
  NOR2X0 U18842 ( .IN1(n16490), .IN2(n10158), .QN(n18149) );
  NAND2X0 U18843 ( .IN1(n18150), .IN2(n18151), .QN(g21056) );
  NAND2X0 U18844 ( .IN1(n16605), .IN2(n10323), .QN(n18151) );
  NAND2X0 U18845 ( .IN1(n16698), .IN2(g2103), .QN(n18150) );
  NAND2X0 U18846 ( .IN1(n18152), .IN2(n18153), .QN(g21055) );
  NAND2X0 U18847 ( .IN1(n16596), .IN2(n4473), .QN(n18153) );
  NAND2X0 U18848 ( .IN1(n16597), .IN2(g2101), .QN(n18152) );
  NAND2X0 U18849 ( .IN1(n18154), .IN2(n18155), .QN(g21054) );
  NAND2X0 U18850 ( .IN1(n16499), .IN2(n4468), .QN(n18155) );
  INVX0 U18851 ( .INP(n18156), .ZN(n18154) );
  NOR2X0 U18852 ( .IN1(n16499), .IN2(n10166), .QN(n18156) );
  NAND2X0 U18853 ( .IN1(n18157), .IN2(n18158), .QN(g21053) );
  NAND2X0 U18854 ( .IN1(n16702), .IN2(n4395), .QN(n18158) );
  NAND2X0 U18855 ( .IN1(n16701), .IN2(g1410), .QN(n18157) );
  NAND2X0 U18856 ( .IN1(n18159), .IN2(n18160), .QN(g21052) );
  NAND2X0 U18857 ( .IN1(n16602), .IN2(n4475), .QN(n18160) );
  INVX0 U18858 ( .INP(n18161), .ZN(n18159) );
  NOR2X0 U18859 ( .IN1(n16602), .IN2(n10175), .QN(n18161) );
  NAND2X0 U18860 ( .IN1(n18162), .IN2(n18163), .QN(g21051) );
  NAND2X0 U18861 ( .IN1(n16707), .IN2(n4396), .QN(n18163) );
  INVX0 U18862 ( .INP(n18164), .ZN(n18162) );
  NOR2X0 U18863 ( .IN1(n16707), .IN2(n10184), .QN(n18164) );
  NAND2X0 U18864 ( .IN1(n18165), .IN2(n18166), .QN(g21047) );
  INVX0 U18865 ( .INP(n18167), .ZN(n18166) );
  NOR2X0 U18866 ( .IN1(n14690), .IN2(n9878), .QN(n18167) );
  NAND2X0 U18867 ( .IN1(n14690), .IN2(n11275), .QN(n18165) );
  NAND2X0 U18868 ( .IN1(n18168), .IN2(n18169), .QN(g21046) );
  NAND2X0 U18869 ( .IN1(n18142), .IN2(g2802), .QN(n18169) );
  INVX0 U18870 ( .INP(n17688), .ZN(n18142) );
  NAND2X0 U18871 ( .IN1(n17688), .IN2(n11267), .QN(n18168) );
  NOR2X0 U18872 ( .IN1(n10072), .IN2(n4292), .QN(n17688) );
  NAND2X0 U18873 ( .IN1(n18170), .IN2(n18171), .QN(g21045) );
  NAND2X0 U18874 ( .IN1(n16503), .IN2(n10324), .QN(n18171) );
  NAND2X0 U18875 ( .IN1(n16502), .IN2(g2791), .QN(n18170) );
  NAND2X0 U18876 ( .IN1(n18172), .IN2(n18173), .QN(g21044) );
  NAND2X0 U18877 ( .IN1(n16494), .IN2(n4407), .QN(n18173) );
  NAND2X0 U18878 ( .IN1(n16493), .IN2(g2789), .QN(n18172) );
  NAND2X0 U18879 ( .IN1(n18174), .IN2(n18175), .QN(g21043) );
  NAND2X0 U18880 ( .IN1(n16490), .IN2(n4397), .QN(n18175) );
  INVX0 U18881 ( .INP(n18176), .ZN(n18174) );
  NOR2X0 U18882 ( .IN1(n16490), .IN2(n10159), .QN(n18176) );
  NAND2X0 U18883 ( .IN1(n18177), .IN2(n18178), .QN(g21042) );
  NAND2X0 U18884 ( .IN1(n18179), .IN2(g2111), .QN(n18178) );
  NAND2X0 U18885 ( .IN1(n17691), .IN2(n11446), .QN(n18177) );
  NAND2X0 U18886 ( .IN1(n18180), .IN2(n18181), .QN(g21041) );
  NAND2X0 U18887 ( .IN1(n16605), .IN2(n4473), .QN(n18181) );
  NAND2X0 U18888 ( .IN1(n16698), .IN2(g2100), .QN(n18180) );
  NAND2X0 U18889 ( .IN1(n18182), .IN2(n18183), .QN(g21040) );
  NAND2X0 U18890 ( .IN1(n16596), .IN2(n4468), .QN(n18183) );
  NAND2X0 U18891 ( .IN1(n16597), .IN2(g2098), .QN(n18182) );
  NAND2X0 U18892 ( .IN1(n18184), .IN2(n18185), .QN(g21039) );
  NAND2X0 U18893 ( .IN1(n16499), .IN2(n4409), .QN(n18185) );
  INVX0 U18894 ( .INP(n18186), .ZN(n18184) );
  NOR2X0 U18895 ( .IN1(n16499), .IN2(n10167), .QN(n18186) );
  NAND2X0 U18896 ( .IN1(n18187), .IN2(n18188), .QN(g21035) );
  NAND2X0 U18897 ( .IN1(n16717), .IN2(n4395), .QN(n18188) );
  NAND2X0 U18898 ( .IN1(n16716), .IN2(g1409), .QN(n18187) );
  NAND2X0 U18899 ( .IN1(n18189), .IN2(n18190), .QN(g21034) );
  NAND2X0 U18900 ( .IN1(n16702), .IN2(n4475), .QN(n18190) );
  NAND2X0 U18901 ( .IN1(n16701), .IN2(g1407), .QN(n18189) );
  NAND2X0 U18902 ( .IN1(n18191), .IN2(n18192), .QN(g21033) );
  NAND2X0 U18903 ( .IN1(n16602), .IN2(n4469), .QN(n18192) );
  INVX0 U18904 ( .INP(n18193), .ZN(n18191) );
  NOR2X0 U18905 ( .IN1(n16602), .IN2(n10176), .QN(n18193) );
  NAND2X0 U18906 ( .IN1(n18194), .IN2(n18195), .QN(g21032) );
  NAND2X0 U18907 ( .IN1(n16813), .IN2(n4396), .QN(n18195) );
  NAND2X0 U18908 ( .IN1(n16812), .IN2(g724), .QN(n18194) );
  NAND2X0 U18909 ( .IN1(n18196), .IN2(n18197), .QN(g21031) );
  NAND2X0 U18910 ( .IN1(n16707), .IN2(n4477), .QN(n18197) );
  INVX0 U18911 ( .INP(n18198), .ZN(n18196) );
  NOR2X0 U18912 ( .IN1(n16707), .IN2(n10185), .QN(n18198) );
  NAND2X0 U18913 ( .IN1(n18199), .IN2(n18200), .QN(g21029) );
  NAND2X0 U18914 ( .IN1(n18201), .IN2(n11275), .QN(n18200) );
  INVX0 U18915 ( .INP(n11846), .ZN(n11275) );
  NAND2X0 U18916 ( .IN1(n18202), .IN2(n18203), .QN(n11846) );
  NAND2X0 U18917 ( .IN1(test_so90), .IN2(g7390), .QN(n18203) );
  NOR2X0 U18918 ( .IN1(n18204), .IN2(n18205), .QN(n18202) );
  NOR2X0 U18919 ( .IN1(n9729), .IN2(n4299), .QN(n18205) );
  NOR2X0 U18920 ( .IN1(n9728), .IN2(n13148), .QN(n18204) );
  INVX0 U18921 ( .INP(g7302), .ZN(n13148) );
  NAND2X0 U18922 ( .IN1(n17694), .IN2(g2806), .QN(n18199) );
  INVX0 U18923 ( .INP(n18201), .ZN(n17694) );
  NAND2X0 U18924 ( .IN1(n18206), .IN2(n18207), .QN(g21028) );
  NAND2X0 U18925 ( .IN1(n14826), .IN2(g2804), .QN(n18207) );
  INVX0 U18926 ( .INP(n14690), .ZN(n14826) );
  NAND2X0 U18927 ( .IN1(n14690), .IN2(n11267), .QN(n18206) );
  NAND2X0 U18928 ( .IN1(n18208), .IN2(n18209), .QN(g21027) );
  NAND2X0 U18929 ( .IN1(n16503), .IN2(n4407), .QN(n18209) );
  NAND2X0 U18930 ( .IN1(n16502), .IN2(g2788), .QN(n18208) );
  NAND2X0 U18931 ( .IN1(n18210), .IN2(n18211), .QN(g21026) );
  NAND2X0 U18932 ( .IN1(n16494), .IN2(n4397), .QN(n18211) );
  NAND2X0 U18933 ( .IN1(n16493), .IN2(g2786), .QN(n18210) );
  NAND2X0 U18934 ( .IN1(n18212), .IN2(n18213), .QN(g21025) );
  NAND2X0 U18935 ( .IN1(test_so93), .IN2(n16488), .QN(n18213) );
  NAND2X0 U18936 ( .IN1(n16490), .IN2(n4408), .QN(n18212) );
  NAND2X0 U18937 ( .IN1(n18214), .IN2(n18215), .QN(g21023) );
  NAND2X0 U18938 ( .IN1(n14703), .IN2(g2113), .QN(n18215) );
  NAND2X0 U18939 ( .IN1(n15735), .IN2(n11446), .QN(n18214) );
  NAND2X0 U18940 ( .IN1(n18216), .IN2(n18217), .QN(g21022) );
  NAND2X0 U18941 ( .IN1(n18179), .IN2(g2108), .QN(n18217) );
  NAND2X0 U18942 ( .IN1(n17691), .IN2(n11438), .QN(n18216) );
  INVX0 U18943 ( .INP(n18179), .ZN(n17691) );
  NAND2X0 U18944 ( .IN1(g2010), .IN2(g2009), .QN(n18179) );
  NAND2X0 U18945 ( .IN1(n18218), .IN2(n18219), .QN(g21021) );
  NAND2X0 U18946 ( .IN1(n16605), .IN2(n4468), .QN(n18219) );
  NAND2X0 U18947 ( .IN1(n16698), .IN2(g2097), .QN(n18218) );
  NAND2X0 U18948 ( .IN1(n18220), .IN2(n18221), .QN(g21020) );
  NAND2X0 U18949 ( .IN1(n16596), .IN2(n4409), .QN(n18221) );
  NAND2X0 U18950 ( .IN1(n16597), .IN2(g2095), .QN(n18220) );
  NAND2X0 U18951 ( .IN1(n18222), .IN2(n18223), .QN(g21019) );
  NAND2X0 U18952 ( .IN1(n16499), .IN2(n4399), .QN(n18223) );
  NAND2X0 U18953 ( .IN1(n16497), .IN2(g2090), .QN(n18222) );
  NAND2X0 U18954 ( .IN1(n18224), .IN2(n18225), .QN(g21018) );
  NAND2X0 U18955 ( .IN1(n18226), .IN2(g1417), .QN(n18225) );
  NAND2X0 U18956 ( .IN1(n17697), .IN2(n11622), .QN(n18224) );
  NAND2X0 U18957 ( .IN1(n18227), .IN2(n18228), .QN(g21017) );
  NAND2X0 U18958 ( .IN1(n16717), .IN2(n4475), .QN(n18228) );
  NAND2X0 U18959 ( .IN1(n16716), .IN2(g1406), .QN(n18227) );
  NAND2X0 U18960 ( .IN1(n18229), .IN2(n18230), .QN(g21016) );
  NAND2X0 U18961 ( .IN1(n16702), .IN2(n4469), .QN(n18230) );
  NAND2X0 U18962 ( .IN1(n16701), .IN2(g1404), .QN(n18229) );
  NAND2X0 U18963 ( .IN1(n18231), .IN2(n18232), .QN(g21015) );
  NAND2X0 U18964 ( .IN1(n16602), .IN2(n4411), .QN(n18232) );
  NAND2X0 U18965 ( .IN1(n16600), .IN2(g1399), .QN(n18231) );
  NAND2X0 U18966 ( .IN1(n18233), .IN2(n18234), .QN(g21011) );
  NAND2X0 U18967 ( .IN1(n16817), .IN2(n4396), .QN(n18234) );
  NAND2X0 U18968 ( .IN1(n16816), .IN2(g723), .QN(n18233) );
  NAND2X0 U18969 ( .IN1(n18235), .IN2(n18236), .QN(g21010) );
  NAND2X0 U18970 ( .IN1(n16813), .IN2(n4477), .QN(n18236) );
  NAND2X0 U18971 ( .IN1(n16812), .IN2(g721), .QN(n18235) );
  NAND2X0 U18972 ( .IN1(n18237), .IN2(n18238), .QN(g21009) );
  NAND2X0 U18973 ( .IN1(n16707), .IN2(n10325), .QN(n18238) );
  INVX0 U18974 ( .INP(n18239), .ZN(n18237) );
  NOR2X0 U18975 ( .IN1(n16707), .IN2(n10186), .QN(n18239) );
  NAND2X0 U18976 ( .IN1(n18240), .IN2(n18241), .QN(g21007) );
  NAND2X0 U18977 ( .IN1(n18201), .IN2(n11267), .QN(n18241) );
  INVX0 U18978 ( .INP(n11354), .ZN(n11267) );
  NAND2X0 U18979 ( .IN1(n18242), .IN2(n18243), .QN(n11354) );
  NAND2X0 U18980 ( .IN1(g7390), .IN2(g2691), .QN(n18243) );
  NOR2X0 U18981 ( .IN1(n18244), .IN2(n18245), .QN(n18242) );
  NOR2X0 U18982 ( .IN1(n9719), .IN2(n4314), .QN(n18245) );
  NOR2X0 U18983 ( .IN1(n9720), .IN2(n4299), .QN(n18244) );
  INVX0 U18984 ( .INP(n18246), .ZN(n18240) );
  NOR2X0 U18985 ( .IN1(n18201), .IN2(n10300), .QN(n18246) );
  NOR2X0 U18986 ( .IN1(n4306), .IN2(n10072), .QN(n18201) );
  NAND2X0 U18987 ( .IN1(n18247), .IN2(n18248), .QN(g21006) );
  NAND2X0 U18988 ( .IN1(n16503), .IN2(n4397), .QN(n18248) );
  NAND2X0 U18989 ( .IN1(n16502), .IN2(g2785), .QN(n18247) );
  NAND2X0 U18990 ( .IN1(n18249), .IN2(n18250), .QN(g21005) );
  NAND2X0 U18991 ( .IN1(n16494), .IN2(n4408), .QN(n18250) );
  NAND2X0 U18992 ( .IN1(n16493), .IN2(g2783), .QN(n18249) );
  NAND2X0 U18993 ( .IN1(n18251), .IN2(n18252), .QN(g21004) );
  NAND2X0 U18994 ( .IN1(n16490), .IN2(n4419), .QN(n18252) );
  INVX0 U18995 ( .INP(n18253), .ZN(n18251) );
  NOR2X0 U18996 ( .IN1(n16490), .IN2(n10160), .QN(n18253) );
  NAND2X0 U18997 ( .IN1(n18254), .IN2(n18255), .QN(g21003) );
  INVX0 U18998 ( .INP(n18256), .ZN(n18255) );
  NOR2X0 U18999 ( .IN1(n17699), .IN2(n9887), .QN(n18256) );
  NAND2X0 U19000 ( .IN1(n17699), .IN2(n11446), .QN(n18254) );
  INVX0 U19001 ( .INP(n11508), .ZN(n11446) );
  NAND2X0 U19002 ( .IN1(n18257), .IN2(n18258), .QN(n11508) );
  NAND2X0 U19003 ( .IN1(g1930), .IN2(g1991), .QN(n18258) );
  NOR2X0 U19004 ( .IN1(n18259), .IN2(n18260), .QN(n18257) );
  NOR2X0 U19005 ( .IN1(n9732), .IN2(n4315), .QN(n18260) );
  NOR2X0 U19006 ( .IN1(n9730), .IN2(n17237), .QN(n18259) );
  INVX0 U19007 ( .INP(g7052), .ZN(n17237) );
  NAND2X0 U19008 ( .IN1(n18261), .IN2(n18262), .QN(g21002) );
  NAND2X0 U19009 ( .IN1(n14703), .IN2(g2110), .QN(n18262) );
  NAND2X0 U19010 ( .IN1(n15735), .IN2(n11438), .QN(n18261) );
  NAND2X0 U19011 ( .IN1(n18263), .IN2(n18264), .QN(g21001) );
  NAND2X0 U19012 ( .IN1(n16605), .IN2(n4409), .QN(n18264) );
  NAND2X0 U19013 ( .IN1(n16698), .IN2(g2094), .QN(n18263) );
  NAND2X0 U19014 ( .IN1(n18265), .IN2(n18266), .QN(g21000) );
  NAND2X0 U19015 ( .IN1(test_so71), .IN2(n16597), .QN(n18266) );
  NAND2X0 U19016 ( .IN1(n16596), .IN2(n4399), .QN(n18265) );
  NAND2X0 U19017 ( .IN1(n18267), .IN2(n18268), .QN(g20999) );
  NAND2X0 U19018 ( .IN1(n16499), .IN2(n4410), .QN(n18268) );
  INVX0 U19019 ( .INP(n18269), .ZN(n18267) );
  NOR2X0 U19020 ( .IN1(n16499), .IN2(n10169), .QN(n18269) );
  NAND2X0 U19021 ( .IN1(n18270), .IN2(n18271), .QN(g20997) );
  NAND2X0 U19022 ( .IN1(n14834), .IN2(g1419), .QN(n18271) );
  NAND2X0 U19023 ( .IN1(n14704), .IN2(n11622), .QN(n18270) );
  NAND2X0 U19024 ( .IN1(n18272), .IN2(n18273), .QN(g20996) );
  NAND2X0 U19025 ( .IN1(test_so51), .IN2(n18226), .QN(n18273) );
  NAND2X0 U19026 ( .IN1(n17697), .IN2(n11614), .QN(n18272) );
  INVX0 U19027 ( .INP(n18226), .ZN(n17697) );
  NAND2X0 U19028 ( .IN1(g1316), .IN2(g1315), .QN(n18226) );
  NAND2X0 U19029 ( .IN1(n18274), .IN2(n18275), .QN(g20995) );
  NAND2X0 U19030 ( .IN1(n16717), .IN2(n4469), .QN(n18275) );
  NAND2X0 U19031 ( .IN1(n16716), .IN2(g1403), .QN(n18274) );
  NAND2X0 U19032 ( .IN1(n18276), .IN2(n18277), .QN(g20994) );
  NAND2X0 U19033 ( .IN1(test_so50), .IN2(n16701), .QN(n18277) );
  NAND2X0 U19034 ( .IN1(n16702), .IN2(n4411), .QN(n18276) );
  NAND2X0 U19035 ( .IN1(n18278), .IN2(n18279), .QN(g20993) );
  NAND2X0 U19036 ( .IN1(n16602), .IN2(n4401), .QN(n18279) );
  INVX0 U19037 ( .INP(n18280), .ZN(n18278) );
  NOR2X0 U19038 ( .IN1(n16602), .IN2(n10178), .QN(n18280) );
  NAND2X0 U19039 ( .IN1(n18281), .IN2(n18282), .QN(g20992) );
  NAND2X0 U19040 ( .IN1(n18283), .IN2(g731), .QN(n18282) );
  NAND2X0 U19041 ( .IN1(n17703), .IN2(n11096), .QN(n18281) );
  NAND2X0 U19042 ( .IN1(n18284), .IN2(n18285), .QN(g20991) );
  NAND2X0 U19043 ( .IN1(n16817), .IN2(n4477), .QN(n18285) );
  NAND2X0 U19044 ( .IN1(n16816), .IN2(g720), .QN(n18284) );
  NAND2X0 U19045 ( .IN1(n18286), .IN2(n18287), .QN(g20990) );
  NAND2X0 U19046 ( .IN1(n16813), .IN2(n10325), .QN(n18287) );
  NAND2X0 U19047 ( .IN1(n16812), .IN2(g718), .QN(n18286) );
  NAND2X0 U19048 ( .IN1(n18288), .IN2(n18289), .QN(g20989) );
  NAND2X0 U19049 ( .IN1(n16707), .IN2(n4413), .QN(n18289) );
  INVX0 U19050 ( .INP(n18290), .ZN(n18288) );
  NOR2X0 U19051 ( .IN1(n16707), .IN2(n10187), .QN(n18290) );
  NAND2X0 U19052 ( .IN1(n18291), .IN2(n18292), .QN(g20983) );
  NAND2X0 U19053 ( .IN1(n16503), .IN2(n4408), .QN(n18292) );
  NAND2X0 U19054 ( .IN1(n16502), .IN2(g2782), .QN(n18291) );
  NAND2X0 U19055 ( .IN1(n18293), .IN2(n18294), .QN(g20982) );
  NAND2X0 U19056 ( .IN1(n16494), .IN2(n4419), .QN(n18294) );
  NAND2X0 U19057 ( .IN1(n16493), .IN2(g2780), .QN(n18293) );
  NAND2X0 U19058 ( .IN1(n18295), .IN2(n18296), .QN(g20981) );
  NAND2X0 U19059 ( .IN1(n16490), .IN2(n4472), .QN(n18296) );
  INVX0 U19060 ( .INP(n18297), .ZN(n18295) );
  NOR2X0 U19061 ( .IN1(n16490), .IN2(n10161), .QN(n18297) );
  NAND2X0 U19062 ( .IN1(n18298), .IN2(n18299), .QN(g20980) );
  INVX0 U19063 ( .INP(n18300), .ZN(n18299) );
  NOR2X0 U19064 ( .IN1(n17699), .IN2(n10299), .QN(n18300) );
  NAND2X0 U19065 ( .IN1(n17699), .IN2(n11438), .QN(n18298) );
  INVX0 U19066 ( .INP(n11527), .ZN(n11438) );
  NAND2X0 U19067 ( .IN1(n18301), .IN2(n18302), .QN(n11527) );
  NAND2X0 U19068 ( .IN1(g1930), .IN2(g2000), .QN(n18302) );
  NOR2X0 U19069 ( .IN1(n18303), .IN2(n18304), .QN(n18301) );
  NOR2X0 U19070 ( .IN1(n9724), .IN2(n4315), .QN(n18304) );
  NOR2X0 U19071 ( .IN1(n9722), .IN2(n4296), .QN(n18303) );
  NOR2X0 U19072 ( .IN1(n10073), .IN2(n4307), .QN(n17699) );
  NAND2X0 U19073 ( .IN1(n18305), .IN2(n18306), .QN(g20979) );
  NAND2X0 U19074 ( .IN1(n16605), .IN2(n4399), .QN(n18306) );
  NAND2X0 U19075 ( .IN1(n16698), .IN2(g2091), .QN(n18305) );
  NAND2X0 U19076 ( .IN1(n18307), .IN2(n18308), .QN(g20978) );
  NAND2X0 U19077 ( .IN1(n16596), .IN2(n4410), .QN(n18308) );
  NAND2X0 U19078 ( .IN1(n16597), .IN2(g2089), .QN(n18307) );
  NAND2X0 U19079 ( .IN1(n18309), .IN2(n18310), .QN(g20977) );
  NAND2X0 U19080 ( .IN1(n16499), .IN2(n4420), .QN(n18310) );
  INVX0 U19081 ( .INP(n18311), .ZN(n18309) );
  NOR2X0 U19082 ( .IN1(n16499), .IN2(n10170), .QN(n18311) );
  NAND2X0 U19083 ( .IN1(n18312), .IN2(n18313), .QN(g20976) );
  INVX0 U19084 ( .INP(n18314), .ZN(n18313) );
  NOR2X0 U19085 ( .IN1(n17705), .IN2(n9888), .QN(n18314) );
  NAND2X0 U19086 ( .IN1(n17705), .IN2(n11622), .QN(n18312) );
  INVX0 U19087 ( .INP(n11684), .ZN(n11622) );
  NAND2X0 U19088 ( .IN1(n18315), .IN2(n18316), .QN(n11684) );
  NAND2X0 U19089 ( .IN1(g6944), .IN2(g1294), .QN(n18316) );
  NOR2X0 U19090 ( .IN1(n18317), .IN2(n18318), .QN(n18315) );
  NOR2X0 U19091 ( .IN1(n9734), .IN2(n4300), .QN(n18318) );
  NOR2X0 U19092 ( .IN1(n9733), .IN2(n17258), .QN(n18317) );
  INVX0 U19093 ( .INP(g6750), .ZN(n17258) );
  NAND2X0 U19094 ( .IN1(n18319), .IN2(n18320), .QN(g20975) );
  NAND2X0 U19095 ( .IN1(n14834), .IN2(g1416), .QN(n18320) );
  NAND2X0 U19096 ( .IN1(n14704), .IN2(n11614), .QN(n18319) );
  NAND2X0 U19097 ( .IN1(n18321), .IN2(n18322), .QN(g20974) );
  NAND2X0 U19098 ( .IN1(n16717), .IN2(n4411), .QN(n18322) );
  NAND2X0 U19099 ( .IN1(n16716), .IN2(g1400), .QN(n18321) );
  NAND2X0 U19100 ( .IN1(n18323), .IN2(n18324), .QN(g20973) );
  NAND2X0 U19101 ( .IN1(n16702), .IN2(n4401), .QN(n18324) );
  NAND2X0 U19102 ( .IN1(n16701), .IN2(g1398), .QN(n18323) );
  NAND2X0 U19103 ( .IN1(n18325), .IN2(n18326), .QN(g20972) );
  NAND2X0 U19104 ( .IN1(n16602), .IN2(n4412), .QN(n18326) );
  INVX0 U19105 ( .INP(n18327), .ZN(n18325) );
  NOR2X0 U19106 ( .IN1(n16602), .IN2(n10179), .QN(n18327) );
  NAND2X0 U19107 ( .IN1(n18328), .IN2(n18329), .QN(g20970) );
  INVX0 U19108 ( .INP(n18330), .ZN(n18329) );
  NOR2X0 U19109 ( .IN1(n14141), .IN2(n9884), .QN(n18330) );
  NAND2X0 U19110 ( .IN1(n14141), .IN2(n11096), .QN(n18328) );
  NAND2X0 U19111 ( .IN1(n18331), .IN2(n18332), .QN(g20969) );
  NAND2X0 U19112 ( .IN1(n18283), .IN2(g728), .QN(n18332) );
  INVX0 U19113 ( .INP(n17703), .ZN(n18283) );
  NAND2X0 U19114 ( .IN1(n17703), .IN2(n11130), .QN(n18331) );
  NOR2X0 U19115 ( .IN1(n10075), .IN2(n4295), .QN(n17703) );
  NAND2X0 U19116 ( .IN1(n18333), .IN2(n18334), .QN(g20968) );
  NAND2X0 U19117 ( .IN1(n16817), .IN2(n10325), .QN(n18334) );
  NAND2X0 U19118 ( .IN1(n16816), .IN2(g717), .QN(n18333) );
  NAND2X0 U19119 ( .IN1(n18335), .IN2(n18336), .QN(g20967) );
  NAND2X0 U19120 ( .IN1(n16813), .IN2(n4413), .QN(n18336) );
  NAND2X0 U19121 ( .IN1(n16812), .IN2(g715), .QN(n18335) );
  NAND2X0 U19122 ( .IN1(n18337), .IN2(n18338), .QN(g20966) );
  NAND2X0 U19123 ( .IN1(n16707), .IN2(n4403), .QN(n18338) );
  NAND2X0 U19124 ( .IN1(n16705), .IN2(g710), .QN(n18337) );
  NAND2X0 U19125 ( .IN1(n18339), .IN2(n18340), .QN(g20965) );
  NAND2X0 U19126 ( .IN1(n16490), .IN2(n4415), .QN(n18340) );
  INVX0 U19127 ( .INP(n18341), .ZN(n18339) );
  NOR2X0 U19128 ( .IN1(n16490), .IN2(n10155), .QN(n18341) );
  NAND2X0 U19129 ( .IN1(n18342), .IN2(n18343), .QN(g20964) );
  NAND2X0 U19130 ( .IN1(n16503), .IN2(n4419), .QN(n18343) );
  NAND2X0 U19131 ( .IN1(n16502), .IN2(g2779), .QN(n18342) );
  NAND2X0 U19132 ( .IN1(n18344), .IN2(n18345), .QN(g20963) );
  NAND2X0 U19133 ( .IN1(n16494), .IN2(n4472), .QN(n18345) );
  NAND2X0 U19134 ( .IN1(n16493), .IN2(g2777), .QN(n18344) );
  NAND2X0 U19135 ( .IN1(n18346), .IN2(n18347), .QN(g20962) );
  NAND2X0 U19136 ( .IN1(n16490), .IN2(n4398), .QN(n18347) );
  INVX0 U19137 ( .INP(n18348), .ZN(n18346) );
  NOR2X0 U19138 ( .IN1(n16490), .IN2(n10162), .QN(n18348) );
  INVX0 U19139 ( .INP(n16488), .ZN(n16490) );
  NAND2X0 U19140 ( .IN1(n18349), .IN2(n18051), .QN(n16488) );
  NAND2X0 U19141 ( .IN1(n18350), .IN2(n18351), .QN(g20955) );
  NAND2X0 U19142 ( .IN1(n16605), .IN2(n4410), .QN(n18351) );
  NAND2X0 U19143 ( .IN1(n16698), .IN2(g2088), .QN(n18350) );
  NAND2X0 U19144 ( .IN1(n18352), .IN2(n18353), .QN(g20954) );
  NAND2X0 U19145 ( .IN1(n16596), .IN2(n4420), .QN(n18353) );
  NAND2X0 U19146 ( .IN1(n16597), .IN2(g2086), .QN(n18352) );
  NAND2X0 U19147 ( .IN1(n18354), .IN2(n18355), .QN(g20953) );
  NAND2X0 U19148 ( .IN1(n16499), .IN2(n4474), .QN(n18355) );
  INVX0 U19149 ( .INP(n18356), .ZN(n18354) );
  NOR2X0 U19150 ( .IN1(n16499), .IN2(n10171), .QN(n18356) );
  NAND2X0 U19151 ( .IN1(n18357), .IN2(n18358), .QN(g20952) );
  INVX0 U19152 ( .INP(n18359), .ZN(n18358) );
  NOR2X0 U19153 ( .IN1(n17705), .IN2(n10298), .QN(n18359) );
  NAND2X0 U19154 ( .IN1(n17705), .IN2(n11614), .QN(n18357) );
  INVX0 U19155 ( .INP(n11703), .ZN(n11614) );
  NAND2X0 U19156 ( .IN1(n18360), .IN2(n18361), .QN(n11703) );
  NAND2X0 U19157 ( .IN1(n14180), .IN2(g1300), .QN(n18361) );
  NOR2X0 U19158 ( .IN1(n18362), .IN2(n18363), .QN(n18360) );
  NOR2X0 U19159 ( .IN1(n9727), .IN2(n4316), .QN(n18363) );
  NOR2X0 U19160 ( .IN1(n9726), .IN2(n4300), .QN(n18362) );
  NOR2X0 U19161 ( .IN1(n10074), .IN2(n4308), .QN(n17705) );
  NAND2X0 U19162 ( .IN1(n18364), .IN2(n18365), .QN(g20951) );
  NAND2X0 U19163 ( .IN1(n16717), .IN2(n4401), .QN(n18365) );
  NAND2X0 U19164 ( .IN1(n16716), .IN2(g1397), .QN(n18364) );
  NAND2X0 U19165 ( .IN1(n18366), .IN2(n18367), .QN(g20950) );
  NAND2X0 U19166 ( .IN1(n16702), .IN2(n4412), .QN(n18367) );
  NAND2X0 U19167 ( .IN1(n16701), .IN2(g1395), .QN(n18366) );
  NAND2X0 U19168 ( .IN1(n18368), .IN2(n18369), .QN(g20949) );
  NAND2X0 U19169 ( .IN1(n16602), .IN2(n4421), .QN(n18369) );
  INVX0 U19170 ( .INP(n18370), .ZN(n18368) );
  NOR2X0 U19171 ( .IN1(n16602), .IN2(n10180), .QN(n18370) );
  NAND2X0 U19172 ( .IN1(n18371), .IN2(n18372), .QN(g20948) );
  NAND2X0 U19173 ( .IN1(n17709), .IN2(n11096), .QN(n18372) );
  INVX0 U19174 ( .INP(n11174), .ZN(n11096) );
  NAND2X0 U19175 ( .IN1(n18373), .IN2(n18374), .QN(n11174) );
  NAND2X0 U19176 ( .IN1(g6642), .IN2(g608), .QN(n18374) );
  NOR2X0 U19177 ( .IN1(n18375), .IN2(n18376), .QN(n18373) );
  NOR2X0 U19178 ( .IN1(n9717), .IN2(n4313), .QN(n18376) );
  NOR2X0 U19179 ( .IN1(n9716), .IN2(n4298), .QN(n18375) );
  INVX0 U19180 ( .INP(n18377), .ZN(n18371) );
  NOR2X0 U19181 ( .IN1(n17709), .IN2(n9889), .QN(n18377) );
  NAND2X0 U19182 ( .IN1(n18378), .IN2(n18379), .QN(g20947) );
  NAND2X0 U19183 ( .IN1(n14712), .IN2(g730), .QN(n18379) );
  INVX0 U19184 ( .INP(n14141), .ZN(n14712) );
  NAND2X0 U19185 ( .IN1(n14141), .IN2(n11130), .QN(n18378) );
  NAND2X0 U19186 ( .IN1(n18380), .IN2(n18381), .QN(g20946) );
  NAND2X0 U19187 ( .IN1(n16817), .IN2(n4413), .QN(n18381) );
  NAND2X0 U19188 ( .IN1(n16816), .IN2(g714), .QN(n18380) );
  NAND2X0 U19189 ( .IN1(n18382), .IN2(n18383), .QN(g20945) );
  NAND2X0 U19190 ( .IN1(n16813), .IN2(n4403), .QN(n18383) );
  NAND2X0 U19191 ( .IN1(n16812), .IN2(g712), .QN(n18382) );
  NAND2X0 U19192 ( .IN1(n18384), .IN2(n18385), .QN(g20944) );
  NAND2X0 U19193 ( .IN1(n16707), .IN2(n4414), .QN(n18385) );
  INVX0 U19194 ( .INP(n18386), .ZN(n18384) );
  NOR2X0 U19195 ( .IN1(n16707), .IN2(n10189), .QN(n18386) );
  NAND2X0 U19196 ( .IN1(n18387), .IN2(n18388), .QN(g20941) );
  NAND2X0 U19197 ( .IN1(n16494), .IN2(n4415), .QN(n18388) );
  NAND2X0 U19198 ( .IN1(n16493), .IN2(g2801), .QN(n18387) );
  NAND2X0 U19199 ( .IN1(n18389), .IN2(n18390), .QN(g20940) );
  NAND2X0 U19200 ( .IN1(n16503), .IN2(n4472), .QN(n18390) );
  NAND2X0 U19201 ( .IN1(n16502), .IN2(g2776), .QN(n18389) );
  NAND2X0 U19202 ( .IN1(n18391), .IN2(n18392), .QN(g20939) );
  NAND2X0 U19203 ( .IN1(n16494), .IN2(n4398), .QN(n18392) );
  INVX0 U19204 ( .INP(n16493), .ZN(n16494) );
  NAND2X0 U19205 ( .IN1(n16493), .IN2(g2774), .QN(n18391) );
  NAND2X0 U19206 ( .IN1(n18393), .IN2(n18349), .QN(n16493) );
  NOR2X0 U19207 ( .IN1(n4356), .IN2(g2733), .QN(n18393) );
  NAND2X0 U19208 ( .IN1(n18394), .IN2(n18395), .QN(g20937) );
  NAND2X0 U19209 ( .IN1(n16499), .IN2(n4416), .QN(n18395) );
  NAND2X0 U19210 ( .IN1(n16497), .IN2(g2105), .QN(n18394) );
  NAND2X0 U19211 ( .IN1(n18396), .IN2(n18397), .QN(g20936) );
  NAND2X0 U19212 ( .IN1(n16605), .IN2(n4420), .QN(n18397) );
  NAND2X0 U19213 ( .IN1(n16698), .IN2(g2085), .QN(n18396) );
  NAND2X0 U19214 ( .IN1(n18398), .IN2(n18399), .QN(g20935) );
  NAND2X0 U19215 ( .IN1(n16596), .IN2(n4474), .QN(n18399) );
  NAND2X0 U19216 ( .IN1(n16597), .IN2(g2083), .QN(n18398) );
  NAND2X0 U19217 ( .IN1(n18400), .IN2(n18401), .QN(g20934) );
  NAND2X0 U19218 ( .IN1(n16499), .IN2(n4400), .QN(n18401) );
  INVX0 U19219 ( .INP(n18402), .ZN(n18400) );
  NOR2X0 U19220 ( .IN1(n16499), .IN2(n10172), .QN(n18402) );
  INVX0 U19221 ( .INP(n16497), .ZN(n16499) );
  NAND2X0 U19222 ( .IN1(n18403), .IN2(test_so69), .QN(n16497) );
  NOR2X0 U19223 ( .IN1(n10034), .IN2(n18059), .QN(n18403) );
  NAND2X0 U19224 ( .IN1(n18404), .IN2(n18405), .QN(g20927) );
  NAND2X0 U19225 ( .IN1(n16717), .IN2(n4412), .QN(n18405) );
  NAND2X0 U19226 ( .IN1(n16716), .IN2(g1394), .QN(n18404) );
  NAND2X0 U19227 ( .IN1(n18406), .IN2(n18407), .QN(g20926) );
  NAND2X0 U19228 ( .IN1(n16702), .IN2(n4421), .QN(n18407) );
  NAND2X0 U19229 ( .IN1(n16701), .IN2(g1392), .QN(n18406) );
  NAND2X0 U19230 ( .IN1(n18408), .IN2(n18409), .QN(g20925) );
  NAND2X0 U19231 ( .IN1(n16602), .IN2(n4476), .QN(n18409) );
  INVX0 U19232 ( .INP(n18410), .ZN(n18408) );
  NOR2X0 U19233 ( .IN1(n16602), .IN2(n10181), .QN(n18410) );
  NAND2X0 U19234 ( .IN1(n18411), .IN2(n18412), .QN(g20924) );
  NAND2X0 U19235 ( .IN1(n17709), .IN2(n11130), .QN(n18412) );
  INVX0 U19236 ( .INP(n11183), .ZN(n11130) );
  NAND2X0 U19237 ( .IN1(n18413), .IN2(n18414), .QN(n11183) );
  NAND2X0 U19238 ( .IN1(g6642), .IN2(g617), .QN(n18414) );
  NOR2X0 U19239 ( .IN1(n18415), .IN2(n18416), .QN(n18413) );
  INVX0 U19240 ( .INP(n18417), .ZN(n18416) );
  NAND2X0 U19241 ( .IN1(g550), .IN2(test_so26), .QN(n18417) );
  NOR2X0 U19242 ( .IN1(n9714), .IN2(n17296), .QN(n18415) );
  INVX0 U19243 ( .INP(g6485), .ZN(n17296) );
  INVX0 U19244 ( .INP(n18418), .ZN(n18411) );
  NOR2X0 U19245 ( .IN1(n17709), .IN2(n10297), .QN(n18418) );
  NOR2X0 U19246 ( .IN1(n4309), .IN2(n10075), .QN(n17709) );
  NAND2X0 U19247 ( .IN1(n18419), .IN2(n18420), .QN(g20923) );
  NAND2X0 U19248 ( .IN1(test_so29), .IN2(n16816), .QN(n18420) );
  NAND2X0 U19249 ( .IN1(n16817), .IN2(n4403), .QN(n18419) );
  NAND2X0 U19250 ( .IN1(n18421), .IN2(n18422), .QN(g20922) );
  NAND2X0 U19251 ( .IN1(n16813), .IN2(n4414), .QN(n18422) );
  NAND2X0 U19252 ( .IN1(n16812), .IN2(g709), .QN(n18421) );
  NAND2X0 U19253 ( .IN1(n18423), .IN2(n18424), .QN(g20921) );
  NAND2X0 U19254 ( .IN1(n16707), .IN2(n4422), .QN(n18424) );
  INVX0 U19255 ( .INP(n18425), .ZN(n18423) );
  NOR2X0 U19256 ( .IN1(n16707), .IN2(n10190), .QN(n18425) );
  NAND2X0 U19257 ( .IN1(n18426), .IN2(n18427), .QN(g20919) );
  NAND2X0 U19258 ( .IN1(n16503), .IN2(n4415), .QN(n18427) );
  NAND2X0 U19259 ( .IN1(n16502), .IN2(g2800), .QN(n18426) );
  NAND2X0 U19260 ( .IN1(n18428), .IN2(n18429), .QN(g20918) );
  NAND2X0 U19261 ( .IN1(n16503), .IN2(n4398), .QN(n18429) );
  INVX0 U19262 ( .INP(n16502), .ZN(n16503) );
  NAND2X0 U19263 ( .IN1(n16502), .IN2(g2773), .QN(n18428) );
  NAND2X0 U19264 ( .IN1(n18430), .IN2(n18349), .QN(n16502) );
  NOR2X0 U19265 ( .IN1(n10033), .IN2(n4490), .QN(n18349) );
  NOR2X0 U19266 ( .IN1(n4306), .IN2(g2733), .QN(n18430) );
  NAND2X0 U19267 ( .IN1(n18431), .IN2(n18432), .QN(g20917) );
  NAND2X0 U19268 ( .IN1(test_so72), .IN2(n16597), .QN(n18432) );
  NAND2X0 U19269 ( .IN1(n16596), .IN2(n4416), .QN(n18431) );
  NAND2X0 U19270 ( .IN1(n18433), .IN2(n18434), .QN(g20916) );
  NAND2X0 U19271 ( .IN1(n16605), .IN2(n4474), .QN(n18434) );
  NAND2X0 U19272 ( .IN1(n16698), .IN2(g2082), .QN(n18433) );
  NAND2X0 U19273 ( .IN1(n18435), .IN2(n18436), .QN(g20915) );
  NAND2X0 U19274 ( .IN1(n16596), .IN2(n4400), .QN(n18436) );
  NAND2X0 U19275 ( .IN1(n16597), .IN2(g2080), .QN(n18435) );
  INVX0 U19276 ( .INP(n16596), .ZN(n16597) );
  NOR2X0 U19277 ( .IN1(n18437), .IN2(n4357), .QN(n16596) );
  NAND2X0 U19278 ( .IN1(n18438), .IN2(n18439), .QN(g20913) );
  NAND2X0 U19279 ( .IN1(n16602), .IN2(n4417), .QN(n18439) );
  INVX0 U19280 ( .INP(n18440), .ZN(n18438) );
  NOR2X0 U19281 ( .IN1(n16602), .IN2(n10173), .QN(n18440) );
  NAND2X0 U19282 ( .IN1(n18441), .IN2(n18442), .QN(g20912) );
  NAND2X0 U19283 ( .IN1(n16717), .IN2(n4421), .QN(n18442) );
  NAND2X0 U19284 ( .IN1(n16716), .IN2(g1391), .QN(n18441) );
  NAND2X0 U19285 ( .IN1(n18443), .IN2(n18444), .QN(g20911) );
  NAND2X0 U19286 ( .IN1(n16702), .IN2(n4476), .QN(n18444) );
  NAND2X0 U19287 ( .IN1(n16701), .IN2(g1389), .QN(n18443) );
  NAND2X0 U19288 ( .IN1(n18445), .IN2(n18446), .QN(g20910) );
  NAND2X0 U19289 ( .IN1(n16602), .IN2(n4402), .QN(n18446) );
  INVX0 U19290 ( .INP(n16600), .ZN(n16602) );
  NAND2X0 U19291 ( .IN1(n16600), .IN2(g1384), .QN(n18445) );
  NAND2X0 U19292 ( .IN1(n18447), .IN2(n18069), .QN(n16600) );
  NAND2X0 U19293 ( .IN1(n18448), .IN2(n18449), .QN(g20903) );
  NAND2X0 U19294 ( .IN1(n16817), .IN2(n4414), .QN(n18449) );
  NAND2X0 U19295 ( .IN1(n16816), .IN2(g708), .QN(n18448) );
  NAND2X0 U19296 ( .IN1(n18450), .IN2(n18451), .QN(g20902) );
  NAND2X0 U19297 ( .IN1(n16813), .IN2(n4422), .QN(n18451) );
  NAND2X0 U19298 ( .IN1(n16812), .IN2(g706), .QN(n18450) );
  NAND2X0 U19299 ( .IN1(n18452), .IN2(n18453), .QN(g20901) );
  NAND2X0 U19300 ( .IN1(n16707), .IN2(n4478), .QN(n18453) );
  INVX0 U19301 ( .INP(n18454), .ZN(n18452) );
  NOR2X0 U19302 ( .IN1(n16707), .IN2(n10191), .QN(n18454) );
  NAND2X0 U19303 ( .IN1(n18455), .IN2(n18456), .QN(g20900) );
  NAND2X0 U19304 ( .IN1(n16605), .IN2(n4416), .QN(n18456) );
  NAND2X0 U19305 ( .IN1(n16698), .IN2(g2106), .QN(n18455) );
  NAND2X0 U19306 ( .IN1(n18457), .IN2(n18458), .QN(g20899) );
  NAND2X0 U19307 ( .IN1(n16605), .IN2(n4400), .QN(n18458) );
  NAND2X0 U19308 ( .IN1(n16698), .IN2(g2079), .QN(n18457) );
  INVX0 U19309 ( .INP(n16605), .ZN(n16698) );
  NOR2X0 U19310 ( .IN1(n18437), .IN2(n4307), .QN(n16605) );
  NAND2X0 U19311 ( .IN1(n18459), .IN2(test_so69), .QN(n18437) );
  NOR2X0 U19312 ( .IN1(n10034), .IN2(g2039), .QN(n18459) );
  NAND2X0 U19313 ( .IN1(n18460), .IN2(n18461), .QN(g20898) );
  NAND2X0 U19314 ( .IN1(n16702), .IN2(n4417), .QN(n18461) );
  NAND2X0 U19315 ( .IN1(n16701), .IN2(g1413), .QN(n18460) );
  NAND2X0 U19316 ( .IN1(n18462), .IN2(n18463), .QN(g20897) );
  NAND2X0 U19317 ( .IN1(n16717), .IN2(n4476), .QN(n18463) );
  NAND2X0 U19318 ( .IN1(n16716), .IN2(g1388), .QN(n18462) );
  NAND2X0 U19319 ( .IN1(n18464), .IN2(n18465), .QN(g20896) );
  NAND2X0 U19320 ( .IN1(n16702), .IN2(n4402), .QN(n18465) );
  INVX0 U19321 ( .INP(n16701), .ZN(n16702) );
  NAND2X0 U19322 ( .IN1(n16701), .IN2(g1386), .QN(n18464) );
  NAND2X0 U19323 ( .IN1(n18466), .IN2(n18447), .QN(n16701) );
  NOR2X0 U19324 ( .IN1(n4358), .IN2(g1345), .QN(n18466) );
  NAND2X0 U19325 ( .IN1(n18467), .IN2(n18468), .QN(g20894) );
  NAND2X0 U19326 ( .IN1(n16707), .IN2(n4418), .QN(n18468) );
  NAND2X0 U19327 ( .IN1(n16705), .IN2(g725), .QN(n18467) );
  NAND2X0 U19328 ( .IN1(n18469), .IN2(n18470), .QN(g20893) );
  NAND2X0 U19329 ( .IN1(n16817), .IN2(n4422), .QN(n18470) );
  NAND2X0 U19330 ( .IN1(n16816), .IN2(g705), .QN(n18469) );
  NAND2X0 U19331 ( .IN1(n18471), .IN2(n18472), .QN(g20892) );
  NAND2X0 U19332 ( .IN1(n16813), .IN2(n4478), .QN(n18472) );
  NAND2X0 U19333 ( .IN1(n16812), .IN2(g703), .QN(n18471) );
  NAND2X0 U19334 ( .IN1(n18473), .IN2(n18474), .QN(g20891) );
  NAND2X0 U19335 ( .IN1(n16707), .IN2(n4404), .QN(n18474) );
  INVX0 U19336 ( .INP(n18475), .ZN(n18473) );
  NOR2X0 U19337 ( .IN1(n16707), .IN2(n10192), .QN(n18475) );
  INVX0 U19338 ( .INP(n16705), .ZN(n16707) );
  NAND2X0 U19339 ( .IN1(n18476), .IN2(n17561), .QN(n16705) );
  NOR2X0 U19340 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  NAND2X0 U19341 ( .IN1(n18477), .IN2(n18478), .QN(g20883) );
  NAND2X0 U19342 ( .IN1(n16717), .IN2(n4417), .QN(n18478) );
  NAND2X0 U19343 ( .IN1(n16716), .IN2(g1412), .QN(n18477) );
  NAND2X0 U19344 ( .IN1(n18479), .IN2(n18480), .QN(g20882) );
  NAND2X0 U19345 ( .IN1(test_so49), .IN2(n16716), .QN(n18480) );
  NAND2X0 U19346 ( .IN1(n16717), .IN2(n4402), .QN(n18479) );
  INVX0 U19347 ( .INP(n16716), .ZN(n16717) );
  NAND2X0 U19348 ( .IN1(n18481), .IN2(n18447), .QN(n16716) );
  NOR2X0 U19349 ( .IN1(n10035), .IN2(n4489), .QN(n18447) );
  NOR2X0 U19350 ( .IN1(n4308), .IN2(g1345), .QN(n18481) );
  NAND2X0 U19351 ( .IN1(n18482), .IN2(n18483), .QN(g20881) );
  NAND2X0 U19352 ( .IN1(test_so30), .IN2(n16812), .QN(n18483) );
  NAND2X0 U19353 ( .IN1(n16813), .IN2(n4418), .QN(n18482) );
  NAND2X0 U19354 ( .IN1(n18484), .IN2(n18485), .QN(g20880) );
  NAND2X0 U19355 ( .IN1(n16817), .IN2(n4478), .QN(n18485) );
  NAND2X0 U19356 ( .IN1(n16816), .IN2(g702), .QN(n18484) );
  NAND2X0 U19357 ( .IN1(n18486), .IN2(n18487), .QN(g20879) );
  NAND2X0 U19358 ( .IN1(n16813), .IN2(n4404), .QN(n18487) );
  INVX0 U19359 ( .INP(n16812), .ZN(n16813) );
  NAND2X0 U19360 ( .IN1(n16812), .IN2(g700), .QN(n18486) );
  NAND2X0 U19361 ( .IN1(n18488), .IN2(n18476), .QN(n16812) );
  NOR2X0 U19362 ( .IN1(n4359), .IN2(g659), .QN(n18488) );
  NAND2X0 U19363 ( .IN1(n18489), .IN2(n18490), .QN(g20876) );
  NAND2X0 U19364 ( .IN1(n16817), .IN2(n4418), .QN(n18490) );
  NAND2X0 U19365 ( .IN1(n16816), .IN2(g726), .QN(n18489) );
  NAND2X0 U19366 ( .IN1(n18491), .IN2(n18492), .QN(g20875) );
  NAND2X0 U19367 ( .IN1(n16817), .IN2(n4404), .QN(n18492) );
  INVX0 U19368 ( .INP(n16816), .ZN(n16817) );
  NAND2X0 U19369 ( .IN1(n16816), .IN2(g699), .QN(n18491) );
  NAND2X0 U19370 ( .IN1(n18493), .IN2(n18476), .QN(n16816) );
  NOR2X0 U19371 ( .IN1(n10036), .IN2(n4492), .QN(n18476) );
  NOR2X0 U19372 ( .IN1(n4309), .IN2(g659), .QN(n18493) );
  NAND2X0 U19373 ( .IN1(n18494), .IN2(n18495), .QN(g20874) );
  NAND2X0 U19374 ( .IN1(g2879), .IN2(g8096), .QN(n18495) );
  NAND2X0 U19375 ( .IN1(n18077), .IN2(n4351), .QN(n18494) );
  NAND2X0 U19376 ( .IN1(n18496), .IN2(n18497), .QN(n18077) );
  NAND2X0 U19377 ( .IN1(n18082), .IN2(n10733), .QN(n18497) );
  INVX0 U19378 ( .INP(n18498), .ZN(n18496) );
  NOR2X0 U19379 ( .IN1(n10733), .IN2(n18082), .QN(n18498) );
  NOR2X0 U19380 ( .IN1(g3231), .IN2(n18870), .QN(n18082) );
  NOR2X0 U19381 ( .IN1(n18499), .IN2(n18500), .QN(n10733) );
  INVX0 U19382 ( .INP(n18501), .ZN(n18500) );
  NAND2X0 U19383 ( .IN1(n18502), .IN2(n18503), .QN(n18501) );
  NOR2X0 U19384 ( .IN1(n18503), .IN2(n18502), .QN(n18499) );
  NAND2X0 U19385 ( .IN1(n18504), .IN2(n18505), .QN(n18502) );
  INVX0 U19386 ( .INP(n18506), .ZN(n18505) );
  NOR2X0 U19387 ( .IN1(n18507), .IN2(g2959), .QN(n18506) );
  NAND2X0 U19388 ( .IN1(n18507), .IN2(g2959), .QN(n18504) );
  NAND2X0 U19389 ( .IN1(n18508), .IN2(n18509), .QN(n18507) );
  NAND2X0 U19390 ( .IN1(n10276), .IN2(g2935), .QN(n18509) );
  NAND2X0 U19391 ( .IN1(n10275), .IN2(g2938), .QN(n18508) );
  NOR2X0 U19392 ( .IN1(n18510), .IN2(n18511), .QN(n18503) );
  INVX0 U19393 ( .INP(n18512), .ZN(n18511) );
  NAND2X0 U19394 ( .IN1(n10273), .IN2(n18513), .QN(n18512) );
  NOR2X0 U19395 ( .IN1(n18513), .IN2(n10273), .QN(n18510) );
  NAND2X0 U19396 ( .IN1(n18514), .IN2(n18515), .QN(n18513) );
  NAND2X0 U19397 ( .IN1(n18516), .IN2(n18517), .QN(n18515) );
  NAND2X0 U19398 ( .IN1(n18518), .IN2(n18519), .QN(n18517) );
  NAND2X0 U19399 ( .IN1(n10278), .IN2(g2947), .QN(n18519) );
  NAND2X0 U19400 ( .IN1(n10277), .IN2(g2953), .QN(n18518) );
  NOR2X0 U19401 ( .IN1(n18520), .IN2(n18521), .QN(n18516) );
  NOR2X0 U19402 ( .IN1(n10280), .IN2(g2944), .QN(n18521) );
  NOR2X0 U19403 ( .IN1(n10279), .IN2(g2956), .QN(n18520) );
  NAND2X0 U19404 ( .IN1(n18522), .IN2(n18523), .QN(n18514) );
  NAND2X0 U19405 ( .IN1(n18524), .IN2(n18525), .QN(n18523) );
  NAND2X0 U19406 ( .IN1(n10280), .IN2(g2944), .QN(n18525) );
  NAND2X0 U19407 ( .IN1(n10279), .IN2(g2956), .QN(n18524) );
  NOR2X0 U19408 ( .IN1(n18526), .IN2(n18527), .QN(n18522) );
  NOR2X0 U19409 ( .IN1(n10278), .IN2(g2947), .QN(n18527) );
  NOR2X0 U19410 ( .IN1(n10277), .IN2(g2953), .QN(n18526) );
  NOR2X0 U19411 ( .IN1(n14690), .IN2(n18528), .QN(g20789) );
  NAND2X0 U19412 ( .IN1(n18529), .IN2(n18530), .QN(n18528) );
  NAND2X0 U19413 ( .IN1(n4398), .IN2(n18053), .QN(n18530) );
  INVX0 U19414 ( .INP(n18051), .ZN(n18053) );
  NAND2X0 U19415 ( .IN1(n18051), .IN2(g2714), .QN(n18529) );
  NOR2X0 U19416 ( .IN1(g2733), .IN2(n4292), .QN(n18051) );
  NOR2X0 U19417 ( .IN1(n10072), .IN2(n4356), .QN(n14690) );
  NOR2X0 U19418 ( .IN1(n15735), .IN2(n18531), .QN(g20752) );
  NAND2X0 U19419 ( .IN1(n18532), .IN2(n18533), .QN(n18531) );
  NAND2X0 U19420 ( .IN1(n4400), .IN2(n18059), .QN(n18533) );
  INVX0 U19421 ( .INP(n18057), .ZN(n18059) );
  NAND2X0 U19422 ( .IN1(n18057), .IN2(g2020), .QN(n18532) );
  NOR2X0 U19423 ( .IN1(g2039), .IN2(n4293), .QN(n18057) );
  INVX0 U19424 ( .INP(n14703), .ZN(n15735) );
  NAND2X0 U19425 ( .IN1(g2010), .IN2(g7357), .QN(n14703) );
  NOR2X0 U19426 ( .IN1(n14704), .IN2(n18534), .QN(g20717) );
  NAND2X0 U19427 ( .IN1(n18535), .IN2(n18536), .QN(n18534) );
  NAND2X0 U19428 ( .IN1(n4402), .IN2(n18071), .QN(n18536) );
  INVX0 U19429 ( .INP(n18069), .ZN(n18071) );
  NAND2X0 U19430 ( .IN1(n18069), .IN2(g1326), .QN(n18535) );
  NOR2X0 U19431 ( .IN1(g1345), .IN2(n4294), .QN(n18069) );
  INVX0 U19432 ( .INP(n14834), .ZN(n14704) );
  NAND2X0 U19433 ( .IN1(g1316), .IN2(g7161), .QN(n14834) );
  NOR2X0 U19434 ( .IN1(n14141), .IN2(n18537), .QN(g20682) );
  NAND2X0 U19435 ( .IN1(n18538), .IN2(n18539), .QN(n18537) );
  NAND2X0 U19436 ( .IN1(n4404), .IN2(n17563), .QN(n18539) );
  INVX0 U19437 ( .INP(n17561), .ZN(n17563) );
  NAND2X0 U19438 ( .IN1(n17561), .IN2(g640), .QN(n18538) );
  NOR2X0 U19439 ( .IN1(g659), .IN2(n4295), .QN(n17561) );
  NOR2X0 U19440 ( .IN1(n10075), .IN2(n4359), .QN(n14141) );
  NAND2X0 U19441 ( .IN1(n18540), .IN2(n18541), .QN(g20417) );
  NAND2X0 U19442 ( .IN1(g2879), .IN2(g7334), .QN(n18541) );
  NAND2X0 U19443 ( .IN1(n4351), .IN2(g2963), .QN(n18540) );
  NAND2X0 U19444 ( .IN1(n18542), .IN2(n18543), .QN(g20376) );
  NAND2X0 U19445 ( .IN1(n4351), .IN2(test_so2), .QN(n18543) );
  NAND2X0 U19446 ( .IN1(g2879), .IN2(g6895), .QN(n18542) );
  NAND2X0 U19447 ( .IN1(n18544), .IN2(n18545), .QN(g20375) );
  NAND2X0 U19448 ( .IN1(n4292), .IN2(g2733), .QN(n18545) );
  NAND2X0 U19449 ( .IN1(n18546), .IN2(g2703), .QN(n18544) );
  NAND2X0 U19450 ( .IN1(n18547), .IN2(n18548), .QN(g20353) );
  NAND2X0 U19451 ( .IN1(n4293), .IN2(g2039), .QN(n18548) );
  NAND2X0 U19452 ( .IN1(n18546), .IN2(g2009), .QN(n18547) );
  NAND2X0 U19453 ( .IN1(n18549), .IN2(n18550), .QN(g20343) );
  NAND2X0 U19454 ( .IN1(g2879), .IN2(g6442), .QN(n18550) );
  NAND2X0 U19455 ( .IN1(n4351), .IN2(g2969), .QN(n18549) );
  NAND2X0 U19456 ( .IN1(n18551), .IN2(n18552), .QN(g20333) );
  NAND2X0 U19457 ( .IN1(n4294), .IN2(g1345), .QN(n18552) );
  NAND2X0 U19458 ( .IN1(n18546), .IN2(g1315), .QN(n18551) );
  NAND2X0 U19459 ( .IN1(n18553), .IN2(n18554), .QN(g20314) );
  NAND2X0 U19460 ( .IN1(n4295), .IN2(g659), .QN(n18554) );
  NAND2X0 U19461 ( .IN1(n18546), .IN2(g629), .QN(n18553) );
  INVX0 U19462 ( .INP(n17655), .ZN(n18546) );
  NAND2X0 U19463 ( .IN1(n18555), .IN2(n18556), .QN(n17655) );
  NOR2X0 U19464 ( .IN1(g3002), .IN2(n18557), .QN(n18556) );
  NAND2X0 U19465 ( .IN1(n10305), .IN2(n10327), .QN(n18557) );
  NOR2X0 U19466 ( .IN1(g3013), .IN2(g3024), .QN(n18555) );
  NAND2X0 U19467 ( .IN1(n18558), .IN2(n18559), .QN(g20310) );
  NAND2X0 U19468 ( .IN1(g2879), .IN2(g6225), .QN(n18559) );
  NAND2X0 U19469 ( .IN1(n4351), .IN2(g2972), .QN(n18558) );
  NAND2X0 U19470 ( .IN1(n18560), .IN2(n18561), .QN(g19184) );
  NAND2X0 U19471 ( .IN1(g2879), .IN2(g4590), .QN(n18561) );
  NAND2X0 U19472 ( .IN1(n4351), .IN2(g2975), .QN(n18560) );
  NAND2X0 U19473 ( .IN1(n18562), .IN2(n18563), .QN(g19178) );
  NAND2X0 U19474 ( .IN1(test_so5), .IN2(g2879), .QN(n18563) );
  NAND2X0 U19475 ( .IN1(n4351), .IN2(g2935), .QN(n18562) );
  NAND2X0 U19476 ( .IN1(n18564), .IN2(n18565), .QN(g19173) );
  NAND2X0 U19477 ( .IN1(g2879), .IN2(g4323), .QN(n18565) );
  NAND2X0 U19478 ( .IN1(n4351), .IN2(g2978), .QN(n18564) );
  NAND2X0 U19479 ( .IN1(n18566), .IN2(n18567), .QN(g19172) );
  NAND2X0 U19480 ( .IN1(g2879), .IN2(g4321), .QN(n18567) );
  NAND2X0 U19481 ( .IN1(n4351), .IN2(g2953), .QN(n18566) );
  NAND2X0 U19482 ( .IN1(n18568), .IN2(n18569), .QN(g19167) );
  NAND2X0 U19483 ( .IN1(g2879), .IN2(g4200), .QN(n18569) );
  NAND2X0 U19484 ( .IN1(n4351), .IN2(g2938), .QN(n18568) );
  NAND2X0 U19485 ( .IN1(n18570), .IN2(n18571), .QN(g19163) );
  NAND2X0 U19486 ( .IN1(g2879), .IN2(g4090), .QN(n18571) );
  NAND2X0 U19487 ( .IN1(n4351), .IN2(g2981), .QN(n18570) );
  NAND2X0 U19488 ( .IN1(n18572), .IN2(n18573), .QN(g19162) );
  NAND2X0 U19489 ( .IN1(g2879), .IN2(g4088), .QN(n18573) );
  NAND2X0 U19490 ( .IN1(n4351), .IN2(g2956), .QN(n18572) );
  NAND2X0 U19491 ( .IN1(n18574), .IN2(n18575), .QN(g19157) );
  NAND2X0 U19492 ( .IN1(g2879), .IN2(g3993), .QN(n18575) );
  NAND2X0 U19493 ( .IN1(n4351), .IN2(g2941), .QN(n18574) );
  NAND2X0 U19494 ( .IN1(n18576), .IN2(n18577), .QN(g19154) );
  NAND2X0 U19495 ( .IN1(test_so3), .IN2(g2879), .QN(n18577) );
  NAND2X0 U19496 ( .IN1(n4351), .IN2(g2874), .QN(n18576) );
  NAND2X0 U19497 ( .IN1(n18578), .IN2(n18579), .QN(g19153) );
  NAND2X0 U19498 ( .IN1(g2879), .IN2(g8249), .QN(n18579) );
  NAND2X0 U19499 ( .IN1(n4351), .IN2(g2959), .QN(n18578) );
  NAND2X0 U19500 ( .IN1(n18580), .IN2(n18581), .QN(g19149) );
  NAND2X0 U19501 ( .IN1(g2879), .IN2(g8175), .QN(n18581) );
  NAND2X0 U19502 ( .IN1(n4351), .IN2(g2944), .QN(n18580) );
  NAND2X0 U19503 ( .IN1(n18582), .IN2(n18583), .QN(g19144) );
  NAND2X0 U19504 ( .IN1(g2879), .IN2(g8023), .QN(n18583) );
  NAND2X0 U19505 ( .IN1(n4351), .IN2(g2947), .QN(n18582) );
  NAND2X0 U19506 ( .IN1(n18584), .IN2(n18585), .QN(g18975) );
  NAND2X0 U19507 ( .IN1(n4351), .IN2(g2195), .QN(n18585) );
  NAND2X0 U19508 ( .IN1(g2981), .IN2(g2879), .QN(n18584) );
  NAND2X0 U19509 ( .IN1(n18586), .IN2(n18587), .QN(g18968) );
  NAND2X0 U19510 ( .IN1(n4351), .IN2(g2190), .QN(n18587) );
  NAND2X0 U19511 ( .IN1(g2978), .IN2(g2879), .QN(n18586) );
  NAND2X0 U19512 ( .IN1(n18588), .IN2(n18589), .QN(g18957) );
  NAND2X0 U19513 ( .IN1(n4351), .IN2(g2165), .QN(n18589) );
  NAND2X0 U19514 ( .IN1(g2963), .IN2(g2879), .QN(n18588) );
  NAND2X0 U19515 ( .IN1(n18590), .IN2(n18591), .QN(g18942) );
  NAND2X0 U19516 ( .IN1(n4351), .IN2(g2185), .QN(n18591) );
  NAND2X0 U19517 ( .IN1(g2975), .IN2(g2879), .QN(n18590) );
  NAND2X0 U19518 ( .IN1(n18592), .IN2(n18593), .QN(g18907) );
  NAND2X0 U19519 ( .IN1(n4365), .IN2(g3061), .QN(n18593) );
  NAND2X0 U19520 ( .IN1(g2987), .IN2(g2997), .QN(n18592) );
  NAND2X0 U19521 ( .IN1(n18594), .IN2(n18595), .QN(g18906) );
  NAND2X0 U19522 ( .IN1(n4351), .IN2(g2180), .QN(n18595) );
  NAND2X0 U19523 ( .IN1(g2972), .IN2(g2879), .QN(n18594) );
  NAND2X0 U19524 ( .IN1(n18596), .IN2(n18597), .QN(g18885) );
  NAND2X0 U19525 ( .IN1(n4351), .IN2(g2200), .QN(n18597) );
  NAND2X0 U19526 ( .IN1(g2874), .IN2(g2879), .QN(n18596) );
  NAND2X0 U19527 ( .IN1(n18598), .IN2(n18599), .QN(g18883) );
  NAND2X0 U19528 ( .IN1(n4351), .IN2(g1471), .QN(n18599) );
  NAND2X0 U19529 ( .IN1(g2935), .IN2(g2879), .QN(n18598) );
  NAND2X0 U19530 ( .IN1(n18600), .IN2(n18601), .QN(g18868) );
  NAND2X0 U19531 ( .IN1(n4365), .IN2(g3060), .QN(n18601) );
  NAND2X0 U19532 ( .IN1(g2987), .IN2(g3078), .QN(n18600) );
  NAND2X0 U19533 ( .IN1(n18602), .IN2(n18603), .QN(g18867) );
  NAND2X0 U19534 ( .IN1(n4351), .IN2(g2175), .QN(n18603) );
  NAND2X0 U19535 ( .IN1(g2969), .IN2(g2879), .QN(n18602) );
  NAND2X0 U19536 ( .IN1(n18604), .IN2(n18605), .QN(g18866) );
  NAND2X0 U19537 ( .IN1(n4351), .IN2(g1476), .QN(n18605) );
  NAND2X0 U19538 ( .IN1(g2938), .IN2(g2879), .QN(n18604) );
  NAND2X0 U19539 ( .IN1(n18606), .IN2(n18607), .QN(g18852) );
  NAND2X0 U19540 ( .IN1(n4351), .IN2(g1481), .QN(n18607) );
  NAND2X0 U19541 ( .IN1(g2941), .IN2(g2879), .QN(n18606) );
  NAND2X0 U19542 ( .IN1(n18608), .IN2(n18609), .QN(g18837) );
  NAND2X0 U19543 ( .IN1(n4365), .IN2(g3059), .QN(n18609) );
  NAND2X0 U19544 ( .IN1(g2987), .IN2(g3077), .QN(n18608) );
  NAND2X0 U19545 ( .IN1(n18610), .IN2(n18611), .QN(g18836) );
  NAND2X0 U19546 ( .IN1(n4351), .IN2(g2170), .QN(n18611) );
  NAND2X0 U19547 ( .IN1(test_so2), .IN2(g2879), .QN(n18610) );
  NAND2X0 U19548 ( .IN1(n18612), .IN2(n18613), .QN(g18835) );
  NAND2X0 U19549 ( .IN1(n4351), .IN2(g1486), .QN(n18613) );
  NAND2X0 U19550 ( .IN1(g2944), .IN2(g2879), .QN(n18612) );
  NAND2X0 U19551 ( .IN1(n18614), .IN2(n18615), .QN(g18821) );
  NAND2X0 U19552 ( .IN1(n4351), .IN2(g1491), .QN(n18615) );
  NAND2X0 U19553 ( .IN1(g2947), .IN2(g2879), .QN(n18614) );
  NAND2X0 U19554 ( .IN1(n18616), .IN2(n18617), .QN(g18820) );
  NAND2X0 U19555 ( .IN1(n4299), .IN2(g2584), .QN(n18617) );
  NAND2X0 U19556 ( .IN1(g2624), .IN2(g2631), .QN(n18616) );
  NAND2X0 U19557 ( .IN1(n18618), .IN2(n18619), .QN(g18804) );
  NAND2X0 U19558 ( .IN1(n4365), .IN2(g3058), .QN(n18619) );
  NAND2X0 U19559 ( .IN1(g2987), .IN2(g3076), .QN(n18618) );
  NAND2X0 U19560 ( .IN1(n18620), .IN2(n18621), .QN(g18803) );
  NAND2X0 U19561 ( .IN1(n4351), .IN2(g1496), .QN(n18621) );
  NAND2X0 U19562 ( .IN1(g2953), .IN2(g2879), .QN(n18620) );
  NAND2X0 U19563 ( .IN1(n18622), .IN2(n18623), .QN(g18794) );
  NAND2X0 U19564 ( .IN1(g1937), .IN2(g1930), .QN(n18623) );
  NAND2X0 U19565 ( .IN1(n4366), .IN2(g1890), .QN(n18622) );
  NAND2X0 U19566 ( .IN1(n18624), .IN2(n18625), .QN(g18782) );
  INVX0 U19567 ( .INP(n18626), .ZN(n18625) );
  NOR2X0 U19568 ( .IN1(g3109), .IN2(n4445), .QN(n18626) );
  NAND2X0 U19569 ( .IN1(g559), .IN2(g3109), .QN(n18624) );
  NAND2X0 U19570 ( .IN1(n18627), .IN2(n18628), .QN(g18781) );
  NAND2X0 U19571 ( .IN1(n4351), .IN2(g1501), .QN(n18628) );
  NAND2X0 U19572 ( .IN1(g2956), .IN2(g2879), .QN(n18627) );
  NAND2X0 U19573 ( .IN1(n18629), .IN2(n18630), .QN(g18780) );
  NAND2X0 U19574 ( .IN1(n4299), .IN2(g2631), .QN(n18630) );
  NAND2X0 U19575 ( .IN1(n10264), .IN2(g2624), .QN(n18629) );
  NAND2X0 U19576 ( .IN1(n18631), .IN2(n18632), .QN(g18763) );
  NAND2X0 U19577 ( .IN1(n4300), .IN2(g1196), .QN(n18632) );
  NAND2X0 U19578 ( .IN1(g1236), .IN2(g1243), .QN(n18631) );
  NAND2X0 U19579 ( .IN1(n18633), .IN2(n18634), .QN(g18755) );
  NAND2X0 U19580 ( .IN1(n4365), .IN2(g3057), .QN(n18634) );
  NAND2X0 U19581 ( .IN1(g2987), .IN2(g3075), .QN(n18633) );
  NAND2X0 U19582 ( .IN1(n18635), .IN2(n18636), .QN(g18754) );
  NAND2X0 U19583 ( .IN1(n4351), .IN2(g1506), .QN(n18636) );
  NAND2X0 U19584 ( .IN1(g2959), .IN2(g2879), .QN(n18635) );
  NAND2X0 U19585 ( .IN1(n18637), .IN2(n18638), .QN(g18743) );
  NAND2X0 U19586 ( .IN1(n4366), .IN2(g1937), .QN(n18638) );
  NAND2X0 U19587 ( .IN1(n10265), .IN2(g1930), .QN(n18637) );
  NAND2X0 U19588 ( .IN1(n18639), .IN2(n18640), .QN(g18726) );
  NAND2X0 U19589 ( .IN1(test_so22), .IN2(n4313), .QN(n18640) );
  NAND2X0 U19590 ( .IN1(g550), .IN2(g557), .QN(n18639) );
  NAND2X0 U19591 ( .IN1(n18641), .IN2(n18642), .QN(g18719) );
  NAND2X0 U19592 ( .IN1(n4383), .IN2(g3211), .QN(n18642) );
  NAND2X0 U19593 ( .IN1(g559), .IN2(g8030), .QN(n18641) );
  NAND2X0 U19594 ( .IN1(n18643), .IN2(n18644), .QN(g18707) );
  NAND2X0 U19595 ( .IN1(n4300), .IN2(g1243), .QN(n18644) );
  NAND2X0 U19596 ( .IN1(n10266), .IN2(g1236), .QN(n18643) );
  NAND2X0 U19597 ( .IN1(n18645), .IN2(n18646), .QN(g18678) );
  NAND2X0 U19598 ( .IN1(n4313), .IN2(g557), .QN(n18646) );
  NAND2X0 U19599 ( .IN1(n10267), .IN2(g550), .QN(n18645) );
  NAND2X0 U19600 ( .IN1(n18647), .IN2(n18648), .QN(g18669) );
  NAND2X0 U19601 ( .IN1(n4382), .IN2(test_so6), .QN(n18648) );
  NAND2X0 U19602 ( .IN1(g559), .IN2(g8106), .QN(n18647) );
  NAND2X0 U19603 ( .IN1(n18649), .IN2(n18650), .QN(g17429) );
  NAND2X0 U19604 ( .IN1(g3109), .IN2(g2574), .QN(n18650) );
  INVX0 U19605 ( .INP(n18651), .ZN(n18649) );
  NOR2X0 U19606 ( .IN1(g3109), .IN2(n4341), .QN(n18651) );
  NAND2X0 U19607 ( .IN1(n18652), .IN2(n18653), .QN(g17383) );
  NAND2X0 U19608 ( .IN1(n4494), .IN2(test_so8), .QN(n18653) );
  NAND2X0 U19609 ( .IN1(g3109), .IN2(g1880), .QN(n18652) );
  NAND2X0 U19610 ( .IN1(n18654), .IN2(n18655), .QN(g17341) );
  INVX0 U19611 ( .INP(n18656), .ZN(n18655) );
  NOR2X0 U19612 ( .IN1(g8030), .IN2(n4442), .QN(n18656) );
  NAND2X0 U19613 ( .IN1(g8030), .IN2(g2574), .QN(n18654) );
  NAND2X0 U19614 ( .IN1(n18657), .IN2(n18658), .QN(g17340) );
  NAND2X0 U19615 ( .IN1(g3109), .IN2(g1186), .QN(n18658) );
  INVX0 U19616 ( .INP(n18659), .ZN(n18657) );
  NOR2X0 U19617 ( .IN1(g3109), .IN2(n4441), .QN(n18659) );
  NAND2X0 U19618 ( .IN1(n18660), .IN2(n18661), .QN(g17303) );
  INVX0 U19619 ( .INP(n18662), .ZN(n18661) );
  NOR2X0 U19620 ( .IN1(g8030), .IN2(n4450), .QN(n18662) );
  NAND2X0 U19621 ( .IN1(g8030), .IN2(g1880), .QN(n18660) );
  NAND2X0 U19622 ( .IN1(n18663), .IN2(n18664), .QN(g17302) );
  NAND2X0 U19623 ( .IN1(g3109), .IN2(g499), .QN(n18664) );
  NAND2X0 U19624 ( .IN1(n4494), .IN2(g3161), .QN(n18663) );
  NAND2X0 U19625 ( .IN1(n18665), .IN2(n18666), .QN(g17271) );
  INVX0 U19626 ( .INP(n18667), .ZN(n18666) );
  NOR2X0 U19627 ( .IN1(g8106), .IN2(n4453), .QN(n18667) );
  NAND2X0 U19628 ( .IN1(g8106), .IN2(g2574), .QN(n18665) );
  NAND2X0 U19629 ( .IN1(n18668), .IN2(n18669), .QN(g17270) );
  NAND2X0 U19630 ( .IN1(g8030), .IN2(g1186), .QN(n18669) );
  INVX0 U19631 ( .INP(n18670), .ZN(n18668) );
  NOR2X0 U19632 ( .IN1(g8030), .IN2(n4348), .QN(n18670) );
  NAND2X0 U19633 ( .IN1(n18671), .IN2(n18672), .QN(g17269) );
  NAND2X0 U19634 ( .IN1(n4494), .IN2(g3096), .QN(n18672) );
  NAND2X0 U19635 ( .IN1(g2633), .IN2(g3109), .QN(n18671) );
  NAND2X0 U19636 ( .IN1(n18673), .IN2(n18674), .QN(g17248) );
  NAND2X0 U19637 ( .IN1(g8106), .IN2(g1880), .QN(n18674) );
  INVX0 U19638 ( .INP(n18675), .ZN(n18673) );
  NOR2X0 U19639 ( .IN1(g8106), .IN2(n4338), .QN(n18675) );
  NAND2X0 U19640 ( .IN1(n18676), .IN2(n18677), .QN(g17247) );
  INVX0 U19641 ( .INP(n18678), .ZN(n18677) );
  NOR2X0 U19642 ( .IN1(g8030), .IN2(n4436), .QN(n18678) );
  NAND2X0 U19643 ( .IN1(g8030), .IN2(g499), .QN(n18676) );
  NAND2X0 U19644 ( .IN1(n18679), .IN2(n18680), .QN(g17246) );
  NAND2X0 U19645 ( .IN1(n4494), .IN2(g3093), .QN(n18680) );
  NAND2X0 U19646 ( .IN1(g1939), .IN2(g3109), .QN(n18679) );
  NAND2X0 U19647 ( .IN1(n18681), .IN2(n18682), .QN(g17236) );
  NAND2X0 U19648 ( .IN1(g8106), .IN2(g1186), .QN(n18682) );
  INVX0 U19649 ( .INP(n18683), .ZN(n18681) );
  NOR2X0 U19650 ( .IN1(g8106), .IN2(n4339), .QN(n18683) );
  NAND2X0 U19651 ( .IN1(n18684), .IN2(n18685), .QN(g17235) );
  INVX0 U19652 ( .INP(n18686), .ZN(n18685) );
  NOR2X0 U19653 ( .IN1(g8030), .IN2(n4439), .QN(n18686) );
  NAND2X0 U19654 ( .IN1(g2633), .IN2(g8030), .QN(n18684) );
  NAND2X0 U19655 ( .IN1(n18687), .IN2(n18688), .QN(g17234) );
  INVX0 U19656 ( .INP(n18689), .ZN(n18688) );
  NOR2X0 U19657 ( .IN1(g3109), .IN2(n4344), .QN(n18689) );
  NAND2X0 U19658 ( .IN1(g1245), .IN2(g3109), .QN(n18687) );
  NAND2X0 U19659 ( .IN1(n18690), .IN2(n18691), .QN(g17229) );
  NAND2X0 U19660 ( .IN1(n4382), .IN2(g3155), .QN(n18691) );
  NAND2X0 U19661 ( .IN1(g8106), .IN2(g499), .QN(n18690) );
  NAND2X0 U19662 ( .IN1(n18692), .IN2(n18693), .QN(g17228) );
  NAND2X0 U19663 ( .IN1(n4383), .IN2(g3092), .QN(n18693) );
  NAND2X0 U19664 ( .IN1(g1939), .IN2(g8030), .QN(n18692) );
  NAND2X0 U19665 ( .IN1(n18694), .IN2(n18695), .QN(g17226) );
  NAND2X0 U19666 ( .IN1(n4382), .IN2(g3094), .QN(n18695) );
  NAND2X0 U19667 ( .IN1(g2633), .IN2(g8106), .QN(n18694) );
  NAND2X0 U19668 ( .IN1(n18696), .IN2(n18697), .QN(g17225) );
  INVX0 U19669 ( .INP(n18698), .ZN(n18697) );
  NOR2X0 U19670 ( .IN1(g8030), .IN2(n4337), .QN(n18698) );
  NAND2X0 U19671 ( .IN1(g1245), .IN2(g8030), .QN(n18696) );
  NAND2X0 U19672 ( .IN1(n18699), .IN2(n18700), .QN(g17224) );
  NAND2X0 U19673 ( .IN1(n4382), .IN2(g3091), .QN(n18700) );
  NAND2X0 U19674 ( .IN1(g1939), .IN2(g8106), .QN(n18699) );
  NAND2X0 U19675 ( .IN1(n18701), .IN2(n18702), .QN(g17222) );
  NAND2X0 U19676 ( .IN1(n4382), .IN2(g3085), .QN(n18702) );
  NAND2X0 U19677 ( .IN1(g1245), .IN2(g8106), .QN(n18701) );
  NAND2X0 U19678 ( .IN1(n18703), .IN2(n18704), .QN(g16880) );
  NAND2X0 U19679 ( .IN1(n4365), .IN2(g3056), .QN(n18704) );
  NAND2X0 U19680 ( .IN1(g2987), .IN2(g3074), .QN(n18703) );
  NAND2X0 U19681 ( .IN1(n18705), .IN2(n18706), .QN(g16866) );
  NAND2X0 U19682 ( .IN1(n4365), .IN2(g3051), .QN(n18706) );
  NAND2X0 U19683 ( .IN1(test_so97), .IN2(g2987), .QN(n18705) );
  NAND2X0 U19684 ( .IN1(n18707), .IN2(n18708), .QN(g16861) );
  NAND2X0 U19685 ( .IN1(test_so96), .IN2(n4365), .QN(n18708) );
  NAND2X0 U19686 ( .IN1(g2987), .IN2(g3073), .QN(n18707) );
  NAND2X0 U19687 ( .IN1(n18709), .IN2(n18710), .QN(g16860) );
  NAND2X0 U19688 ( .IN1(n4365), .IN2(g3046), .QN(n18710) );
  NAND2X0 U19689 ( .IN1(g2987), .IN2(g3065), .QN(n18709) );
  NAND2X0 U19690 ( .IN1(n18711), .IN2(n18712), .QN(g16857) );
  NAND2X0 U19691 ( .IN1(n4365), .IN2(g3050), .QN(n18712) );
  NAND2X0 U19692 ( .IN1(g2987), .IN2(g3069), .QN(n18711) );
  NAND2X0 U19693 ( .IN1(n18713), .IN2(n18714), .QN(g16854) );
  NAND2X0 U19694 ( .IN1(n4365), .IN2(g3053), .QN(n18714) );
  NAND2X0 U19695 ( .IN1(g2987), .IN2(g3072), .QN(n18713) );
  NAND2X0 U19696 ( .IN1(n18715), .IN2(n18716), .QN(g16853) );
  NAND2X0 U19697 ( .IN1(n4365), .IN2(g3045), .QN(n18716) );
  NAND2X0 U19698 ( .IN1(g2987), .IN2(g3064), .QN(n18715) );
  NAND2X0 U19699 ( .IN1(n18717), .IN2(n18718), .QN(g16851) );
  NAND2X0 U19700 ( .IN1(n4365), .IN2(g3049), .QN(n18718) );
  NAND2X0 U19701 ( .IN1(g2987), .IN2(g3068), .QN(n18717) );
  NAND2X0 U19702 ( .IN1(n18719), .IN2(n18720), .QN(g16845) );
  NAND2X0 U19703 ( .IN1(n4365), .IN2(g3052), .QN(n18720) );
  NAND2X0 U19704 ( .IN1(g2987), .IN2(g3071), .QN(n18719) );
  NAND2X0 U19705 ( .IN1(n18721), .IN2(n18722), .QN(g16844) );
  NAND2X0 U19706 ( .IN1(n4365), .IN2(g3044), .QN(n18722) );
  NAND2X0 U19707 ( .IN1(g2987), .IN2(g3063), .QN(n18721) );
  NAND2X0 U19708 ( .IN1(n18723), .IN2(n18724), .QN(g16835) );
  NAND2X0 U19709 ( .IN1(n4365), .IN2(g3048), .QN(n18724) );
  NAND2X0 U19710 ( .IN1(g2987), .IN2(g3067), .QN(n18723) );
  NAND2X0 U19711 ( .IN1(n18725), .IN2(n18726), .QN(g16824) );
  NAND2X0 U19712 ( .IN1(n4365), .IN2(g3043), .QN(n18726) );
  NAND2X0 U19713 ( .IN1(g2987), .IN2(g3062), .QN(n18725) );
  NOR2X0 U19714 ( .IN1(g51), .IN2(DFF_1_n1), .QN(g16823) );
  NAND2X0 U19715 ( .IN1(n18727), .IN2(n18728), .QN(g16803) );
  NAND2X0 U19716 ( .IN1(n4365), .IN2(g3047), .QN(n18728) );
  NAND2X0 U19717 ( .IN1(g2987), .IN2(g3066), .QN(n18727) );
  NOR2X0 U19718 ( .IN1(n4423), .IN2(g51), .QN(g16802) );
  NAND2X0 U19719 ( .IN1(n18729), .IN2(n18730), .QN(g16718) );
  NAND2X0 U19720 ( .IN1(g2703), .IN2(g2584), .QN(n18730) );
  INVX0 U19721 ( .INP(n18731), .ZN(n18729) );
  NOR2X0 U19722 ( .IN1(g2703), .IN2(n10072), .QN(n18731) );
  NAND2X0 U19723 ( .IN1(n18732), .IN2(n18733), .QN(g16692) );
  NAND2X0 U19724 ( .IN1(g2009), .IN2(g1890), .QN(n18733) );
  NAND2X0 U19725 ( .IN1(n4293), .IN2(g2010), .QN(n18732) );
  NAND2X0 U19726 ( .IN1(n18734), .IN2(n18735), .QN(g16671) );
  NAND2X0 U19727 ( .IN1(g1315), .IN2(g1196), .QN(n18735) );
  NAND2X0 U19728 ( .IN1(n4294), .IN2(g1316), .QN(n18734) );
  NAND2X0 U19729 ( .IN1(n18736), .IN2(n18737), .QN(g16654) );
  NAND2X0 U19730 ( .IN1(test_so22), .IN2(g629), .QN(n18737) );
  NAND2X0 U19731 ( .IN1(n4295), .IN2(g630), .QN(n18736) );
  NAND2X0 U19732 ( .IN1(n18738), .IN2(g2987), .QN(g16496) );
  NAND2X0 U19733 ( .IN1(DFF_1612_n1), .IN2(g5388), .QN(n18738) );
  NOR2X0 U19734 ( .IN1(n18739), .IN2(n18740), .QN(g13194) );
  NAND2X0 U19735 ( .IN1(n18741), .IN2(n18742), .QN(n18740) );
  NAND2X0 U19736 ( .IN1(n10037), .IN2(g7390), .QN(n18742) );
  INVX0 U19737 ( .INP(n18743), .ZN(n18741) );
  NOR2X0 U19738 ( .IN1(n4314), .IN2(test_so87), .QN(n18743) );
  NOR2X0 U19739 ( .IN1(n4299), .IN2(g2562), .QN(n18739) );
  NOR2X0 U19740 ( .IN1(n18744), .IN2(n18745), .QN(g13182) );
  NAND2X0 U19741 ( .IN1(n18746), .IN2(n18747), .QN(n18745) );
  NAND2X0 U19742 ( .IN1(n10045), .IN2(g7194), .QN(n18747) );
  NAND2X0 U19743 ( .IN1(n10046), .IN2(n14321), .QN(n18746) );
  NOR2X0 U19744 ( .IN1(n4366), .IN2(g1868), .QN(n18744) );
  NOR2X0 U19745 ( .IN1(n18748), .IN2(n18749), .QN(g13175) );
  NAND2X0 U19746 ( .IN1(n18750), .IN2(n18751), .QN(n18749) );
  NAND2X0 U19747 ( .IN1(n10042), .IN2(g7390), .QN(n18751) );
  NAND2X0 U19748 ( .IN1(n10043), .IN2(n13147), .QN(n18750) );
  NOR2X0 U19749 ( .IN1(n4299), .IN2(g2553), .QN(n18748) );
  NOR2X0 U19750 ( .IN1(n18752), .IN2(n18753), .QN(g13171) );
  NAND2X0 U19751 ( .IN1(n18754), .IN2(n18755), .QN(n18753) );
  NAND2X0 U19752 ( .IN1(n10054), .IN2(g6944), .QN(n18755) );
  INVX0 U19753 ( .INP(n18756), .ZN(n18754) );
  NOR2X0 U19754 ( .IN1(n4300), .IN2(test_so44), .QN(n18756) );
  NOR2X0 U19755 ( .IN1(n4371), .IN2(g1175), .QN(n18752) );
  NOR2X0 U19756 ( .IN1(n18757), .IN2(n18758), .QN(g13164) );
  NAND2X0 U19757 ( .IN1(n18759), .IN2(n18760), .QN(n18758) );
  NAND2X0 U19758 ( .IN1(n10051), .IN2(g7194), .QN(n18760) );
  NAND2X0 U19759 ( .IN1(n10052), .IN2(n14321), .QN(n18759) );
  NOR2X0 U19760 ( .IN1(n4366), .IN2(g1859), .QN(n18757) );
  NOR2X0 U19761 ( .IN1(n18761), .IN2(n18762), .QN(g13160) );
  NAND2X0 U19762 ( .IN1(n18763), .IN2(n18764), .QN(n18762) );
  NAND2X0 U19763 ( .IN1(n10062), .IN2(g6642), .QN(n18764) );
  NAND2X0 U19764 ( .IN1(n10063), .IN2(n14574), .QN(n18763) );
  NOR2X0 U19765 ( .IN1(n4313), .IN2(g487), .QN(n18761) );
  NOR2X0 U19766 ( .IN1(n18765), .IN2(n18766), .QN(g13155) );
  NAND2X0 U19767 ( .IN1(n18767), .IN2(n18768), .QN(n18766) );
  NAND2X0 U19768 ( .IN1(n10059), .IN2(g6944), .QN(n18768) );
  NAND2X0 U19769 ( .IN1(n10060), .IN2(n14180), .QN(n18767) );
  NOR2X0 U19770 ( .IN1(n4300), .IN2(g1165), .QN(n18765) );
  NOR2X0 U19771 ( .IN1(n18769), .IN2(n18770), .QN(g13149) );
  NAND2X0 U19772 ( .IN1(n18771), .IN2(n18772), .QN(n18770) );
  NAND2X0 U19773 ( .IN1(n10068), .IN2(g6642), .QN(n18772) );
  NAND2X0 U19774 ( .IN1(n10069), .IN2(n14574), .QN(n18771) );
  NOR2X0 U19775 ( .IN1(n4313), .IN2(g478), .QN(n18769) );
  NOR2X0 U19776 ( .IN1(n18773), .IN2(n18774), .QN(g13143) );
  NAND2X0 U19777 ( .IN1(n18775), .IN2(n18776), .QN(n18774) );
  NAND2X0 U19778 ( .IN1(n10039), .IN2(g7390), .QN(n18776) );
  NAND2X0 U19779 ( .IN1(n10040), .IN2(n13147), .QN(n18775) );
  INVX0 U19780 ( .INP(n4314), .ZN(n13147) );
  NOR2X0 U19781 ( .IN1(n4299), .IN2(g2559), .QN(n18773) );
  NOR2X0 U19782 ( .IN1(n18777), .IN2(n18778), .QN(g13135) );
  NAND2X0 U19783 ( .IN1(n18779), .IN2(n18780), .QN(n18778) );
  NAND2X0 U19784 ( .IN1(n10048), .IN2(g7194), .QN(n18780) );
  NAND2X0 U19785 ( .IN1(n10049), .IN2(n14321), .QN(n18779) );
  INVX0 U19786 ( .INP(n4296), .ZN(n14321) );
  NOR2X0 U19787 ( .IN1(n4366), .IN2(g1865), .QN(n18777) );
  NOR2X0 U19788 ( .IN1(n18781), .IN2(n18782), .QN(g13124) );
  NAND2X0 U19789 ( .IN1(n18783), .IN2(n18784), .QN(n18782) );
  NAND2X0 U19790 ( .IN1(n10056), .IN2(g6944), .QN(n18784) );
  NAND2X0 U19791 ( .IN1(n10057), .IN2(n14180), .QN(n18783) );
  INVX0 U19792 ( .INP(n4371), .ZN(n14180) );
  NOR2X0 U19793 ( .IN1(n4300), .IN2(g1171), .QN(n18781) );
  NOR2X0 U19794 ( .IN1(n18785), .IN2(n18786), .QN(g13111) );
  NAND2X0 U19795 ( .IN1(n18787), .IN2(n18788), .QN(n18786) );
  NAND2X0 U19796 ( .IN1(n10065), .IN2(g6642), .QN(n18788) );
  NAND2X0 U19797 ( .IN1(n10066), .IN2(n14574), .QN(n18787) );
  INVX0 U19798 ( .INP(n4298), .ZN(n14574) );
  NOR2X0 U19799 ( .IN1(n4313), .IN2(g484), .QN(n18785) );
  NAND2X0 U19800 ( .IN1(n18789), .IN2(n18790), .QN(N995) );
  NAND2X0 U19801 ( .IN1(n10293), .IN2(n11071), .QN(n18790) );
  INVX0 U19802 ( .INP(n18791), .ZN(n18789) );
  NOR2X0 U19803 ( .IN1(n11071), .IN2(n10293), .QN(n18791) );
  NOR2X0 U19804 ( .IN1(n18792), .IN2(n18793), .QN(n11071) );
  INVX0 U19805 ( .INP(n18794), .ZN(n18793) );
  NAND2X0 U19806 ( .IN1(n18795), .IN2(n18796), .QN(n18794) );
  NOR2X0 U19807 ( .IN1(n18796), .IN2(n18795), .QN(n18792) );
  NAND2X0 U19808 ( .IN1(n18797), .IN2(n18798), .QN(n18795) );
  NAND2X0 U19809 ( .IN1(n10289), .IN2(n18799), .QN(n18798) );
  INVX0 U19810 ( .INP(n18800), .ZN(n18797) );
  NOR2X0 U19811 ( .IN1(n18799), .IN2(n10289), .QN(n18800) );
  NOR2X0 U19812 ( .IN1(n18801), .IN2(n18802), .QN(n18799) );
  NOR2X0 U19813 ( .IN1(n10330), .IN2(n10290), .QN(n18802) );
  INVX0 U19814 ( .INP(n18803), .ZN(n18801) );
  NAND2X0 U19815 ( .IN1(n10290), .IN2(n10330), .QN(n18803) );
  NOR2X0 U19816 ( .IN1(n18804), .IN2(n18805), .QN(n18796) );
  INVX0 U19817 ( .INP(n18806), .ZN(n18805) );
  NAND2X0 U19818 ( .IN1(n10288), .IN2(n18807), .QN(n18806) );
  NOR2X0 U19819 ( .IN1(n18807), .IN2(n10288), .QN(n18804) );
  NAND2X0 U19820 ( .IN1(n18808), .IN2(n18809), .QN(n18807) );
  NAND2X0 U19821 ( .IN1(n18810), .IN2(n18811), .QN(n18809) );
  NOR2X0 U19822 ( .IN1(n18812), .IN2(n18813), .QN(n18811) );
  NOR2X0 U19823 ( .IN1(n18874), .IN2(g8269), .QN(n18813) );
  NOR2X0 U19824 ( .IN1(n10291), .IN2(g8273), .QN(n18812) );
  NOR2X0 U19825 ( .IN1(n18814), .IN2(n18815), .QN(n18810) );
  NOR2X0 U19826 ( .IN1(n18875), .IN2(g8268), .QN(n18815) );
  NOR2X0 U19827 ( .IN1(n18876), .IN2(g8272), .QN(n18814) );
  NAND2X0 U19828 ( .IN1(n18816), .IN2(n18817), .QN(n18808) );
  NAND2X0 U19829 ( .IN1(n18818), .IN2(n18819), .QN(n18817) );
  NAND2X0 U19830 ( .IN1(n18874), .IN2(g8269), .QN(n18819) );
  NAND2X0 U19831 ( .IN1(n10291), .IN2(g8273), .QN(n18818) );
  NAND2X0 U19832 ( .IN1(n18820), .IN2(n18821), .QN(n18816) );
  NAND2X0 U19833 ( .IN1(n18875), .IN2(g8268), .QN(n18821) );
  NAND2X0 U19834 ( .IN1(n18876), .IN2(g8272), .QN(n18820) );
  NOR2X0 U19835 ( .IN1(n18822), .IN2(n18823), .QN(N690) );
  NOR2X0 U19836 ( .IN1(n10295), .IN2(n11076), .QN(n18823) );
  INVX0 U19837 ( .INP(n18824), .ZN(n18822) );
  NAND2X0 U19838 ( .IN1(n11076), .IN2(n10295), .QN(n18824) );
  NOR2X0 U19839 ( .IN1(n18825), .IN2(n18826), .QN(n11076) );
  INVX0 U19840 ( .INP(n18827), .ZN(n18826) );
  NAND2X0 U19841 ( .IN1(n18828), .IN2(n18829), .QN(n18827) );
  NOR2X0 U19842 ( .IN1(n18829), .IN2(n18828), .QN(n18825) );
  NAND2X0 U19843 ( .IN1(n18830), .IN2(n18831), .QN(n18828) );
  NAND2X0 U19844 ( .IN1(n10269), .IN2(n18832), .QN(n18831) );
  INVX0 U19845 ( .INP(n18833), .ZN(n18830) );
  NOR2X0 U19846 ( .IN1(n18832), .IN2(n10269), .QN(n18833) );
  NOR2X0 U19847 ( .IN1(n18834), .IN2(n18835), .QN(n18832) );
  NOR2X0 U19848 ( .IN1(g8264), .IN2(n10270), .QN(n18835) );
  INVX0 U19849 ( .INP(n18836), .ZN(n18834) );
  NAND2X0 U19850 ( .IN1(n10270), .IN2(g8264), .QN(n18836) );
  NOR2X0 U19851 ( .IN1(n18837), .IN2(n18838), .QN(n18829) );
  INVX0 U19852 ( .INP(n18839), .ZN(n18838) );
  NAND2X0 U19853 ( .IN1(n10268), .IN2(n18840), .QN(n18839) );
  NOR2X0 U19854 ( .IN1(n18840), .IN2(n10268), .QN(n18837) );
  NAND2X0 U19855 ( .IN1(n18841), .IN2(n18842), .QN(n18840) );
  NAND2X0 U19856 ( .IN1(n18843), .IN2(n18844), .QN(n18842) );
  NOR2X0 U19857 ( .IN1(n18845), .IN2(n18846), .QN(n18844) );
  NOR2X0 U19858 ( .IN1(n18877), .IN2(g8263), .QN(n18846) );
  NOR2X0 U19859 ( .IN1(n10272), .IN2(g8266), .QN(n18845) );
  NOR2X0 U19860 ( .IN1(n18847), .IN2(n18848), .QN(n18843) );
  NOR2X0 U19861 ( .IN1(n18878), .IN2(g8262), .QN(n18848) );
  NOR2X0 U19862 ( .IN1(n18879), .IN2(g8265), .QN(n18847) );
  NAND2X0 U19863 ( .IN1(n18849), .IN2(n18850), .QN(n18841) );
  NAND2X0 U19864 ( .IN1(n18851), .IN2(n18852), .QN(n18850) );
  NAND2X0 U19865 ( .IN1(n18877), .IN2(g8263), .QN(n18852) );
  NAND2X0 U19866 ( .IN1(n10272), .IN2(g8266), .QN(n18851) );
  NAND2X0 U19867 ( .IN1(n18853), .IN2(n18854), .QN(n18849) );
  NAND2X0 U19868 ( .IN1(n18878), .IN2(g8262), .QN(n18854) );
  NAND2X0 U19869 ( .IN1(n18879), .IN2(g8265), .QN(n18853) );
  NOR2X0 U3772_U2 ( .IN1(n2230), .IN2(n2217), .QN(U3772_n1) );
  INVX0 U3772_U1 ( .INP(U3772_n1), .ZN(n2231) );
  NOR2X0 U3776_U2 ( .IN1(n2374), .IN2(n2361), .QN(U3776_n1) );
  INVX0 U3776_U1 ( .INP(U3776_n1), .ZN(n2375) );
  NOR2X0 U3777_U2 ( .IN1(g51), .IN2(DFF_2_n1), .QN(U3777_n1) );
  INVX0 U3777_U1 ( .INP(U3777_n1), .ZN(n4264) );
  NOR2X0 U3778_U2 ( .IN1(n2445), .IN2(n2446), .QN(U3778_n1) );
  INVX0 U3778_U1 ( .INP(U3778_n1), .ZN(n2440) );
  NOR2X0 U3779_U2 ( .IN1(n557), .IN2(n2446), .QN(U3779_n1) );
  INVX0 U3779_U1 ( .INP(U3779_n1), .ZN(n2426) );
  NOR2X0 U3780_U2 ( .IN1(n2670), .IN2(n2671), .QN(U3780_n1) );
  INVX0 U3780_U1 ( .INP(U3780_n1), .ZN(n2669) );
  NOR2X0 U3781_U2 ( .IN1(n2685), .IN2(n2686), .QN(U3781_n1) );
  INVX0 U3781_U1 ( .INP(U3781_n1), .ZN(n2684) );
  NOR2X0 U3782_U2 ( .IN1(n2718), .IN2(n2719), .QN(U3782_n1) );
  INVX0 U3782_U1 ( .INP(U3782_n1), .ZN(n2717) );
  NOR2X0 U3783_U2 ( .IN1(n2982), .IN2(g2124), .QN(U3783_n1) );
  INVX0 U3783_U1 ( .INP(U3783_n1), .ZN(n2981) );
  NOR2X0 U3784_U2 ( .IN1(n2985), .IN2(g1430), .QN(U3784_n1) );
  INVX0 U3784_U1 ( .INP(U3784_n1), .ZN(n2984) );
  NOR2X0 U3785_U2 ( .IN1(n2988), .IN2(g744), .QN(U3785_n1) );
  INVX0 U3785_U1 ( .INP(U3785_n1), .ZN(n2987) );
  NOR2X0 U3786_U2 ( .IN1(n2991), .IN2(g56), .QN(U3786_n1) );
  INVX0 U3786_U1 ( .INP(U3786_n1), .ZN(n2990) );
  NOR2X0 U3787_U2 ( .IN1(n3742), .IN2(test_so98), .QN(U3787_n1) );
  INVX0 U3787_U1 ( .INP(U3787_n1), .ZN(n3741) );
  NOR2X0 U3901_U2 ( .IN1(n2302), .IN2(n2289), .QN(U3901_n1) );
  INVX0 U3901_U1 ( .INP(U3901_n1), .ZN(n2303) );
  NOR2X0 U3902_U2 ( .IN1(n602), .IN2(n2289), .QN(U3902_n1) );
  INVX0 U3902_U1 ( .INP(U3902_n1), .ZN(n2275) );
  INVX0 U4467_U2 ( .INP(n1658), .ZN(U4467_n1) );
  NOR2X0 U4467_U1 ( .IN1(n3254), .IN2(U4467_n1), .QN(n3252) );
  INVX0 U4904_U2 ( .INP(n2800), .ZN(U4904_n1) );
  NOR2X0 U4904_U1 ( .IN1(n2617), .IN2(U4904_n1), .QN(n2798) );
  INVX0 U4930_U2 ( .INP(n2616), .ZN(U4930_n1) );
  NOR2X0 U4930_U1 ( .IN1(n2617), .IN2(U4930_n1), .QN(n2594) );
  INVX0 U5128_U2 ( .INP(n3933), .ZN(U5128_n1) );
  NOR2X0 U5128_U1 ( .IN1(n4406), .IN2(U5128_n1), .QN(n3940) );
  INVX0 U5141_U2 ( .INP(n3939), .ZN(U5141_n1) );
  NOR2X0 U5141_U1 ( .IN1(n4405), .IN2(U5141_n1), .QN(n3936) );
  INVX0 U5749_U2 ( .INP(g2133), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3160), .IN2(U5749_n1), .QN(n3159) );
  INVX0 U5750_U2 ( .INP(g1439), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3164), .IN2(U5750_n1), .QN(n3163) );
  INVX0 U5751_U2 ( .INP(g753), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3168), .IN2(U5751_n1), .QN(n3167) );
  INVX0 U5752_U2 ( .INP(g65), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3172), .IN2(U5752_n1), .QN(n3171) );
  INVX0 U5753_U2 ( .INP(g2142), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4522), .IN2(U5753_n1), .QN(n3424) );
  INVX0 U5754_U2 ( .INP(g2151), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4526), .IN2(U5754_n1), .QN(n3683) );
  INVX0 U5755_U2 ( .INP(g2160), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3888), .IN2(U5755_n1), .QN(n3887) );
  INVX0 U5756_U2 ( .INP(g1448), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4523), .IN2(U5756_n1), .QN(n3427) );
  INVX0 U5757_U2 ( .INP(g1457), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(n3686) );
  INVX0 U5758_U2 ( .INP(g1466), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3891), .IN2(U5758_n1), .QN(n3890) );
  INVX0 U5759_U2 ( .INP(g762), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3431), .IN2(U5759_n1), .QN(n3430) );
  INVX0 U5760_U2 ( .INP(g771), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3690), .IN2(U5760_n1), .QN(n3689) );
  INVX0 U5761_U2 ( .INP(g780), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3894), .IN2(U5761_n1), .QN(n3893) );
  INVX0 U5762_U2 ( .INP(g74), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4521), .IN2(U5762_n1), .QN(n3433) );
  INVX0 U5763_U2 ( .INP(g83), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(n3692) );
  INVX0 U5764_U2 ( .INP(g92), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3897), .IN2(U5764_n1), .QN(n3896) );
  INVX0 U5882_U2 ( .INP(n4102), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(g3036), .IN2(U5882_n1), .QN(n4101) );
  INVX0 U5939_U2 ( .INP(g2257), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n1497), .IN2(U5939_n1), .QN(n3038) );
  INVX0 U5940_U2 ( .INP(g1563), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n1146), .IN2(U5940_n1), .QN(n3070) );
  INVX0 U5941_U2 ( .INP(g869), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n795), .IN2(U5941_n1), .QN(n3102) );
  INVX0 U5942_U2 ( .INP(g181), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n372), .IN2(U5942_n1), .QN(n3130) );
  INVX0 U6140_U2 ( .INP(g3002), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4066), .IN2(U6140_n1), .QN(n4065) );
  INVX0 U6460_U2 ( .INP(g3233), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(g3230), .IN2(U6460_n1), .QN(n3700) );
  INVX0 U6470_U2 ( .INP(g2892), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4305), .IN2(U6470_n1), .QN(n4182) );
  INVX0 U6562_U2 ( .INP(n306), .ZN(U6562_n1) );
  NOR2X0 U6562_U1 ( .IN1(g3204), .IN2(U6562_n1), .QN(n3939) );
  INVX0 U6563_U2 ( .INP(n4073), .ZN(U6563_n1) );
  NOR2X0 U6563_U1 ( .IN1(g3204), .IN2(U6563_n1), .QN(n3705) );
  INVX0 U6718_U2 ( .INP(n307), .ZN(U6718_n1) );
  NOR2X0 U6718_U1 ( .IN1(g3197), .IN2(U6718_n1), .QN(n4073) );
  INVX0 U7116_U2 ( .INP(n18), .ZN(U7116_n1) );
  NOR2X0 U7116_U1 ( .IN1(g2903), .IN2(U7116_n1), .QN(n4057) );
  INVX0 U7118_U2 ( .INP(n4123), .ZN(U7118_n1) );
  NOR2X0 U7118_U1 ( .IN1(g2896), .IN2(U7118_n1), .QN(n4122) );
  INVX0 U7293_U2 ( .INP(n4598), .ZN(U7293_n1) );
  NOR2X0 U7293_U1 ( .IN1(g3234), .IN2(U7293_n1), .QN(g20877) );
endmodule

