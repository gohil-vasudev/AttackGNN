module add_mul_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, operation_0_, operation_1_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_
 );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334;

  OR2_X1 U2121 ( .A1(n4241), .A2(n4242), .ZN(n2089) );
  OR2_X1 U2122 ( .A1(n4242), .A2(operation_0_), .ZN(n2090) );
  OR2_X1 U2123 ( .A1(n4241), .A2(operation_1_), .ZN(n2091) );
  OR2_X1 U2124 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2092) );
  INV_X2 U2125 ( .A(n2092), .ZN(n2093) );
  INV_X2 U2126 ( .A(n2091), .ZN(n2094) );
  INV_X2 U2127 ( .A(n2090), .ZN(n2095) );
  INV_X2 U2128 ( .A(n2089), .ZN(n2096) );
  NAND2_X1 U2129 ( .A1(n2097), .A2(n2098), .ZN(Result_9_) );
  NAND2_X1 U2130 ( .A1(n2099), .A2(n2096), .ZN(n2098) );
  XOR2_X1 U2131 ( .A(n2100), .B(n2101), .Z(n2099) );
  AND2_X1 U2132 ( .A1(n2102), .A2(n2103), .ZN(n2101) );
  NAND2_X1 U2133 ( .A1(n2097), .A2(n2104), .ZN(Result_8_) );
  NAND2_X1 U2134 ( .A1(n2105), .A2(n2096), .ZN(n2104) );
  XOR2_X1 U2135 ( .A(n2106), .B(n2107), .Z(n2105) );
  AND2_X1 U2136 ( .A1(n2108), .A2(n2109), .ZN(n2107) );
  NAND2_X1 U2137 ( .A1(n2097), .A2(n2110), .ZN(Result_7_) );
  NAND2_X1 U2138 ( .A1(n2111), .A2(n2096), .ZN(n2110) );
  XOR2_X1 U2139 ( .A(n2112), .B(n2113), .Z(n2111) );
  AND2_X1 U2140 ( .A1(n2114), .A2(n2115), .ZN(n2113) );
  NAND2_X1 U2141 ( .A1(n2097), .A2(n2116), .ZN(Result_6_) );
  NAND2_X1 U2142 ( .A1(n2117), .A2(n2096), .ZN(n2116) );
  XOR2_X1 U2143 ( .A(n2118), .B(n2119), .Z(n2117) );
  AND2_X1 U2144 ( .A1(n2120), .A2(n2121), .ZN(n2119) );
  NAND2_X1 U2145 ( .A1(n2097), .A2(n2122), .ZN(Result_5_) );
  NAND2_X1 U2146 ( .A1(n2123), .A2(n2096), .ZN(n2122) );
  XOR2_X1 U2147 ( .A(n2124), .B(n2125), .Z(n2123) );
  AND2_X1 U2148 ( .A1(n2126), .A2(n2127), .ZN(n2125) );
  NAND2_X1 U2149 ( .A1(n2097), .A2(n2128), .ZN(Result_4_) );
  NAND2_X1 U2150 ( .A1(n2129), .A2(n2096), .ZN(n2128) );
  XOR2_X1 U2151 ( .A(n2130), .B(n2131), .Z(n2129) );
  AND2_X1 U2152 ( .A1(n2132), .A2(n2133), .ZN(n2131) );
  NAND2_X1 U2153 ( .A1(n2097), .A2(n2134), .ZN(Result_3_) );
  NAND2_X1 U2154 ( .A1(n2135), .A2(n2096), .ZN(n2134) );
  XOR2_X1 U2155 ( .A(n2136), .B(n2137), .Z(n2135) );
  AND2_X1 U2156 ( .A1(n2138), .A2(n2139), .ZN(n2137) );
  NAND2_X1 U2157 ( .A1(n2140), .A2(n2141), .ZN(Result_31_) );
  NAND2_X1 U2158 ( .A1(n2142), .A2(n2096), .ZN(n2141) );
  NAND2_X1 U2159 ( .A1(n2143), .A2(n2144), .ZN(n2140) );
  OR3_X1 U2160 ( .A1(n2095), .A2(n2094), .A3(n2093), .ZN(n2144) );
  NAND2_X1 U2161 ( .A1(n2145), .A2(n2146), .ZN(n2143) );
  NAND3_X1 U2162 ( .A1(n2147), .A2(n2148), .A3(n2149), .ZN(Result_30_) );
  NAND3_X1 U2163 ( .A1(a_14_), .A2(n2150), .A3(n2096), .ZN(n2149) );
  NAND2_X1 U2164 ( .A1(b_14_), .A2(n2151), .ZN(n2148) );
  NAND3_X1 U2165 ( .A1(n2152), .A2(n2153), .A3(n2154), .ZN(n2151) );
  NAND2_X1 U2166 ( .A1(n2096), .A2(n2155), .ZN(n2154) );
  NAND2_X1 U2167 ( .A1(n2146), .A2(n2156), .ZN(n2155) );
  NAND2_X1 U2168 ( .A1(n2157), .A2(n2158), .ZN(n2153) );
  NAND2_X1 U2169 ( .A1(a_14_), .A2(n2159), .ZN(n2152) );
  NAND2_X1 U2170 ( .A1(n2160), .A2(n2161), .ZN(n2147) );
  NAND2_X1 U2171 ( .A1(n2162), .A2(n2163), .ZN(n2160) );
  NAND2_X1 U2172 ( .A1(n2159), .A2(n2158), .ZN(n2163) );
  NAND3_X1 U2173 ( .A1(n2164), .A2(n2165), .A3(n2166), .ZN(n2159) );
  NAND2_X1 U2174 ( .A1(n2094), .A2(n2167), .ZN(n2166) );
  NAND2_X1 U2175 ( .A1(n2093), .A2(n2142), .ZN(n2165) );
  INV_X1 U2176 ( .A(n2168), .ZN(n2142) );
  NAND2_X1 U2177 ( .A1(n2095), .A2(n2150), .ZN(n2164) );
  NAND2_X1 U2178 ( .A1(a_14_), .A2(n2169), .ZN(n2162) );
  NAND2_X1 U2179 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
  NAND2_X1 U2180 ( .A1(n2096), .A2(b_15_), .ZN(n2171) );
  INV_X1 U2181 ( .A(n2157), .ZN(n2170) );
  NAND3_X1 U2182 ( .A1(n2172), .A2(n2173), .A3(n2174), .ZN(n2157) );
  NAND2_X1 U2183 ( .A1(n2094), .A2(n2146), .ZN(n2174) );
  NAND2_X1 U2184 ( .A1(n2093), .A2(n2168), .ZN(n2173) );
  NAND2_X1 U2185 ( .A1(n2095), .A2(n2145), .ZN(n2172) );
  NAND2_X1 U2186 ( .A1(n2097), .A2(n2175), .ZN(Result_2_) );
  NAND2_X1 U2187 ( .A1(n2176), .A2(n2096), .ZN(n2175) );
  XOR2_X1 U2188 ( .A(n2177), .B(n2178), .Z(n2176) );
  AND2_X1 U2189 ( .A1(n2179), .A2(n2180), .ZN(n2178) );
  NAND3_X1 U2190 ( .A1(n2181), .A2(n2182), .A3(n2183), .ZN(Result_29_) );
  NAND2_X1 U2191 ( .A1(n2184), .A2(n2096), .ZN(n2183) );
  XOR2_X1 U2192 ( .A(n2185), .B(n2186), .Z(n2184) );
  NOR2_X1 U2193 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
  XOR2_X1 U2194 ( .A(n2189), .B(n2190), .Z(n2185) );
  NAND2_X1 U2195 ( .A1(n2191), .A2(n2192), .ZN(n2182) );
  NAND3_X1 U2196 ( .A1(n2193), .A2(n2194), .A3(n2195), .ZN(n2191) );
  NAND2_X1 U2197 ( .A1(n2094), .A2(n2196), .ZN(n2195) );
  NAND2_X1 U2198 ( .A1(n2093), .A2(n2197), .ZN(n2194) );
  NAND2_X1 U2199 ( .A1(n2095), .A2(n2198), .ZN(n2193) );
  NAND2_X1 U2200 ( .A1(n2199), .A2(n2200), .ZN(n2181) );
  NAND3_X1 U2201 ( .A1(n2201), .A2(n2202), .A3(n2203), .ZN(n2200) );
  NAND2_X1 U2202 ( .A1(n2094), .A2(n2204), .ZN(n2203) );
  NAND2_X1 U2203 ( .A1(n2205), .A2(n2093), .ZN(n2202) );
  INV_X1 U2204 ( .A(n2197), .ZN(n2205) );
  NAND2_X1 U2205 ( .A1(n2095), .A2(n2206), .ZN(n2201) );
  INV_X1 U2206 ( .A(n2192), .ZN(n2199) );
  NAND2_X1 U2207 ( .A1(n2207), .A2(n2208), .ZN(n2192) );
  NAND3_X1 U2208 ( .A1(n2209), .A2(n2210), .A3(n2211), .ZN(Result_28_) );
  NAND2_X1 U2209 ( .A1(n2096), .A2(n2212), .ZN(n2211) );
  XOR2_X1 U2210 ( .A(n2213), .B(n2214), .Z(n2212) );
  XOR2_X1 U2211 ( .A(n2215), .B(n2216), .Z(n2214) );
  NAND2_X1 U2212 ( .A1(n2217), .A2(n2218), .ZN(n2210) );
  NAND3_X1 U2213 ( .A1(n2219), .A2(n2220), .A3(n2221), .ZN(n2217) );
  NAND2_X1 U2214 ( .A1(n2094), .A2(n2222), .ZN(n2221) );
  NAND2_X1 U2215 ( .A1(n2093), .A2(n2223), .ZN(n2220) );
  NAND2_X1 U2216 ( .A1(n2095), .A2(n2224), .ZN(n2219) );
  NAND2_X1 U2217 ( .A1(n2225), .A2(n2226), .ZN(n2209) );
  NAND3_X1 U2218 ( .A1(n2227), .A2(n2228), .A3(n2229), .ZN(n2226) );
  NAND2_X1 U2219 ( .A1(n2094), .A2(n2230), .ZN(n2229) );
  NAND2_X1 U2220 ( .A1(n2231), .A2(n2093), .ZN(n2228) );
  INV_X1 U2221 ( .A(n2223), .ZN(n2231) );
  NAND2_X1 U2222 ( .A1(n2095), .A2(n2232), .ZN(n2227) );
  INV_X1 U2223 ( .A(n2218), .ZN(n2225) );
  NAND2_X1 U2224 ( .A1(n2233), .A2(n2234), .ZN(n2218) );
  NAND3_X1 U2225 ( .A1(n2235), .A2(n2236), .A3(n2237), .ZN(Result_27_) );
  NAND2_X1 U2226 ( .A1(n2096), .A2(n2238), .ZN(n2237) );
  XNOR2_X1 U2227 ( .A(n2239), .B(n2240), .ZN(n2238) );
  NAND2_X1 U2228 ( .A1(n2241), .A2(n2242), .ZN(n2239) );
  NAND2_X1 U2229 ( .A1(n2243), .A2(n2244), .ZN(n2236) );
  NAND3_X1 U2230 ( .A1(n2245), .A2(n2246), .A3(n2247), .ZN(n2243) );
  NAND2_X1 U2231 ( .A1(n2094), .A2(n2248), .ZN(n2247) );
  NAND2_X1 U2232 ( .A1(n2093), .A2(n2249), .ZN(n2246) );
  NAND2_X1 U2233 ( .A1(n2095), .A2(n2250), .ZN(n2245) );
  NAND2_X1 U2234 ( .A1(n2251), .A2(n2252), .ZN(n2235) );
  NAND3_X1 U2235 ( .A1(n2253), .A2(n2254), .A3(n2255), .ZN(n2252) );
  NAND2_X1 U2236 ( .A1(n2094), .A2(n2256), .ZN(n2255) );
  NAND2_X1 U2237 ( .A1(n2257), .A2(n2093), .ZN(n2254) );
  INV_X1 U2238 ( .A(n2249), .ZN(n2257) );
  NAND2_X1 U2239 ( .A1(n2095), .A2(n2258), .ZN(n2253) );
  INV_X1 U2240 ( .A(n2244), .ZN(n2251) );
  NAND2_X1 U2241 ( .A1(n2259), .A2(n2260), .ZN(n2244) );
  NAND3_X1 U2242 ( .A1(n2261), .A2(n2262), .A3(n2263), .ZN(Result_26_) );
  NAND2_X1 U2243 ( .A1(n2096), .A2(n2264), .ZN(n2263) );
  XOR2_X1 U2244 ( .A(n2265), .B(n2266), .Z(n2264) );
  XOR2_X1 U2245 ( .A(n2267), .B(n2268), .Z(n2266) );
  NAND2_X1 U2246 ( .A1(n2269), .A2(n2270), .ZN(n2262) );
  NAND3_X1 U2247 ( .A1(n2271), .A2(n2272), .A3(n2273), .ZN(n2270) );
  NAND2_X1 U2248 ( .A1(n2094), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2249 ( .A1(n2275), .A2(n2093), .ZN(n2272) );
  INV_X1 U2250 ( .A(n2276), .ZN(n2275) );
  NAND2_X1 U2251 ( .A1(n2095), .A2(n2277), .ZN(n2271) );
  NAND2_X1 U2252 ( .A1(n2278), .A2(n2279), .ZN(n2261) );
  NAND3_X1 U2253 ( .A1(n2280), .A2(n2281), .A3(n2282), .ZN(n2279) );
  NAND2_X1 U2254 ( .A1(n2094), .A2(n2283), .ZN(n2282) );
  NAND2_X1 U2255 ( .A1(n2093), .A2(n2276), .ZN(n2281) );
  NAND2_X1 U2256 ( .A1(n2095), .A2(n2284), .ZN(n2280) );
  INV_X1 U2257 ( .A(n2269), .ZN(n2278) );
  XNOR2_X1 U2258 ( .A(n2285), .B(a_10_), .ZN(n2269) );
  NAND3_X1 U2259 ( .A1(n2286), .A2(n2287), .A3(n2288), .ZN(Result_25_) );
  NAND2_X1 U2260 ( .A1(n2289), .A2(n2096), .ZN(n2288) );
  XNOR2_X1 U2261 ( .A(n2290), .B(n2291), .ZN(n2289) );
  NAND2_X1 U2262 ( .A1(n2292), .A2(n2293), .ZN(n2290) );
  NAND2_X1 U2263 ( .A1(n2294), .A2(n2295), .ZN(n2287) );
  NAND3_X1 U2264 ( .A1(n2296), .A2(n2297), .A3(n2298), .ZN(n2295) );
  NAND2_X1 U2265 ( .A1(n2094), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2266 ( .A1(n2300), .A2(n2093), .ZN(n2297) );
  NAND2_X1 U2267 ( .A1(n2095), .A2(n2301), .ZN(n2296) );
  NAND2_X1 U2268 ( .A1(n2302), .A2(n2303), .ZN(n2286) );
  NAND3_X1 U2269 ( .A1(n2304), .A2(n2305), .A3(n2306), .ZN(n2303) );
  NAND2_X1 U2270 ( .A1(n2094), .A2(n2307), .ZN(n2306) );
  NAND2_X1 U2271 ( .A1(n2093), .A2(n2308), .ZN(n2305) );
  NAND2_X1 U2272 ( .A1(n2095), .A2(n2309), .ZN(n2304) );
  INV_X1 U2273 ( .A(n2294), .ZN(n2302) );
  XNOR2_X1 U2274 ( .A(n2310), .B(b_9_), .ZN(n2294) );
  NAND3_X1 U2275 ( .A1(n2311), .A2(n2312), .A3(n2313), .ZN(Result_24_) );
  NAND2_X1 U2276 ( .A1(n2096), .A2(n2314), .ZN(n2313) );
  XNOR2_X1 U2277 ( .A(n2315), .B(n2316), .ZN(n2314) );
  XNOR2_X1 U2278 ( .A(n2317), .B(n2318), .ZN(n2316) );
  NAND2_X1 U2279 ( .A1(n2319), .A2(n2320), .ZN(n2312) );
  NAND3_X1 U2280 ( .A1(n2321), .A2(n2322), .A3(n2323), .ZN(n2320) );
  NAND2_X1 U2281 ( .A1(n2094), .A2(n2324), .ZN(n2323) );
  NAND2_X1 U2282 ( .A1(n2325), .A2(n2093), .ZN(n2322) );
  NAND2_X1 U2283 ( .A1(n2095), .A2(n2326), .ZN(n2321) );
  NAND2_X1 U2284 ( .A1(n2327), .A2(n2328), .ZN(n2311) );
  NAND3_X1 U2285 ( .A1(n2329), .A2(n2330), .A3(n2331), .ZN(n2328) );
  NAND2_X1 U2286 ( .A1(n2094), .A2(n2332), .ZN(n2331) );
  NAND2_X1 U2287 ( .A1(n2093), .A2(n2333), .ZN(n2330) );
  NAND2_X1 U2288 ( .A1(n2095), .A2(n2334), .ZN(n2329) );
  INV_X1 U2289 ( .A(n2319), .ZN(n2327) );
  XNOR2_X1 U2290 ( .A(n2335), .B(a_8_), .ZN(n2319) );
  NAND3_X1 U2291 ( .A1(n2336), .A2(n2337), .A3(n2338), .ZN(Result_23_) );
  NAND2_X1 U2292 ( .A1(n2339), .A2(n2096), .ZN(n2338) );
  XNOR2_X1 U2293 ( .A(n2340), .B(n2341), .ZN(n2339) );
  NAND2_X1 U2294 ( .A1(n2342), .A2(n2343), .ZN(n2340) );
  NAND2_X1 U2295 ( .A1(n2344), .A2(n2345), .ZN(n2337) );
  NAND3_X1 U2296 ( .A1(n2346), .A2(n2347), .A3(n2348), .ZN(n2345) );
  NAND2_X1 U2297 ( .A1(n2094), .A2(n2349), .ZN(n2348) );
  NAND2_X1 U2298 ( .A1(n2350), .A2(n2093), .ZN(n2347) );
  INV_X1 U2299 ( .A(n2351), .ZN(n2350) );
  NAND2_X1 U2300 ( .A1(n2095), .A2(n2352), .ZN(n2346) );
  NAND2_X1 U2301 ( .A1(n2353), .A2(n2354), .ZN(n2336) );
  NAND3_X1 U2302 ( .A1(n2355), .A2(n2356), .A3(n2357), .ZN(n2354) );
  NAND2_X1 U2303 ( .A1(n2094), .A2(n2358), .ZN(n2357) );
  NAND2_X1 U2304 ( .A1(n2093), .A2(n2351), .ZN(n2356) );
  NAND2_X1 U2305 ( .A1(n2095), .A2(n2359), .ZN(n2355) );
  INV_X1 U2306 ( .A(n2344), .ZN(n2353) );
  XNOR2_X1 U2307 ( .A(n2360), .B(b_7_), .ZN(n2344) );
  NAND3_X1 U2308 ( .A1(n2361), .A2(n2362), .A3(n2363), .ZN(Result_22_) );
  NAND2_X1 U2309 ( .A1(n2096), .A2(n2364), .ZN(n2363) );
  XNOR2_X1 U2310 ( .A(n2365), .B(n2366), .ZN(n2364) );
  XNOR2_X1 U2311 ( .A(n2367), .B(n2368), .ZN(n2366) );
  NAND2_X1 U2312 ( .A1(n2369), .A2(n2370), .ZN(n2362) );
  NAND3_X1 U2313 ( .A1(n2371), .A2(n2372), .A3(n2373), .ZN(n2370) );
  NAND2_X1 U2314 ( .A1(n2094), .A2(n2374), .ZN(n2373) );
  NAND2_X1 U2315 ( .A1(n2375), .A2(n2093), .ZN(n2372) );
  INV_X1 U2316 ( .A(n2376), .ZN(n2375) );
  NAND2_X1 U2317 ( .A1(n2095), .A2(n2377), .ZN(n2371) );
  NAND2_X1 U2318 ( .A1(n2378), .A2(n2379), .ZN(n2361) );
  NAND3_X1 U2319 ( .A1(n2380), .A2(n2381), .A3(n2382), .ZN(n2379) );
  NAND2_X1 U2320 ( .A1(n2094), .A2(n2383), .ZN(n2382) );
  NAND2_X1 U2321 ( .A1(n2093), .A2(n2376), .ZN(n2381) );
  NAND2_X1 U2322 ( .A1(n2095), .A2(n2384), .ZN(n2380) );
  INV_X1 U2323 ( .A(n2369), .ZN(n2378) );
  XNOR2_X1 U2324 ( .A(n2385), .B(a_6_), .ZN(n2369) );
  NAND3_X1 U2325 ( .A1(n2386), .A2(n2387), .A3(n2388), .ZN(Result_21_) );
  NAND2_X1 U2326 ( .A1(n2096), .A2(n2389), .ZN(n2388) );
  XNOR2_X1 U2327 ( .A(n2390), .B(n2391), .ZN(n2389) );
  NAND2_X1 U2328 ( .A1(n2392), .A2(n2393), .ZN(n2390) );
  NAND2_X1 U2329 ( .A1(n2394), .A2(n2395), .ZN(n2387) );
  NAND3_X1 U2330 ( .A1(n2396), .A2(n2397), .A3(n2398), .ZN(n2395) );
  NAND2_X1 U2331 ( .A1(n2094), .A2(n2399), .ZN(n2398) );
  NAND2_X1 U2332 ( .A1(n2400), .A2(n2093), .ZN(n2397) );
  INV_X1 U2333 ( .A(n2401), .ZN(n2400) );
  NAND2_X1 U2334 ( .A1(n2095), .A2(n2402), .ZN(n2396) );
  NAND2_X1 U2335 ( .A1(n2403), .A2(n2404), .ZN(n2386) );
  NAND3_X1 U2336 ( .A1(n2405), .A2(n2406), .A3(n2407), .ZN(n2404) );
  NAND2_X1 U2337 ( .A1(n2094), .A2(n2408), .ZN(n2407) );
  NAND2_X1 U2338 ( .A1(n2093), .A2(n2401), .ZN(n2406) );
  NAND2_X1 U2339 ( .A1(n2095), .A2(n2409), .ZN(n2405) );
  INV_X1 U2340 ( .A(n2394), .ZN(n2403) );
  XNOR2_X1 U2341 ( .A(n2410), .B(b_5_), .ZN(n2394) );
  NAND3_X1 U2342 ( .A1(n2411), .A2(n2412), .A3(n2413), .ZN(Result_20_) );
  NAND2_X1 U2343 ( .A1(n2414), .A2(n2096), .ZN(n2413) );
  XNOR2_X1 U2344 ( .A(n2415), .B(n2416), .ZN(n2414) );
  XOR2_X1 U2345 ( .A(n2417), .B(n2418), .Z(n2416) );
  NAND2_X1 U2346 ( .A1(a_4_), .A2(b_15_), .ZN(n2418) );
  NAND2_X1 U2347 ( .A1(n2419), .A2(n2420), .ZN(n2412) );
  NAND3_X1 U2348 ( .A1(n2421), .A2(n2422), .A3(n2423), .ZN(n2420) );
  NAND2_X1 U2349 ( .A1(n2094), .A2(n2424), .ZN(n2423) );
  NAND2_X1 U2350 ( .A1(n2425), .A2(n2093), .ZN(n2422) );
  NAND2_X1 U2351 ( .A1(n2095), .A2(n2426), .ZN(n2421) );
  NAND2_X1 U2352 ( .A1(n2427), .A2(n2428), .ZN(n2411) );
  NAND3_X1 U2353 ( .A1(n2429), .A2(n2430), .A3(n2431), .ZN(n2428) );
  NAND2_X1 U2354 ( .A1(n2094), .A2(n2432), .ZN(n2431) );
  NAND2_X1 U2355 ( .A1(n2093), .A2(n2433), .ZN(n2430) );
  NAND2_X1 U2356 ( .A1(n2095), .A2(n2434), .ZN(n2429) );
  INV_X1 U2357 ( .A(n2419), .ZN(n2427) );
  XNOR2_X1 U2358 ( .A(n2435), .B(b_4_), .ZN(n2419) );
  NAND2_X1 U2359 ( .A1(n2097), .A2(n2436), .ZN(Result_1_) );
  NAND2_X1 U2360 ( .A1(n2437), .A2(n2096), .ZN(n2436) );
  XOR2_X1 U2361 ( .A(n2438), .B(n2439), .Z(n2437) );
  AND2_X1 U2362 ( .A1(n2440), .A2(n2441), .ZN(n2439) );
  NAND3_X1 U2363 ( .A1(n2442), .A2(n2443), .A3(n2444), .ZN(Result_19_) );
  NAND2_X1 U2364 ( .A1(n2445), .A2(n2096), .ZN(n2444) );
  XNOR2_X1 U2365 ( .A(n2446), .B(n2447), .ZN(n2445) );
  XOR2_X1 U2366 ( .A(n2448), .B(n2449), .Z(n2447) );
  NAND2_X1 U2367 ( .A1(a_3_), .A2(b_15_), .ZN(n2449) );
  NAND2_X1 U2368 ( .A1(n2450), .A2(n2451), .ZN(n2443) );
  NAND3_X1 U2369 ( .A1(n2452), .A2(n2453), .A3(n2454), .ZN(n2451) );
  NAND2_X1 U2370 ( .A1(n2094), .A2(n2455), .ZN(n2454) );
  NAND2_X1 U2371 ( .A1(n2456), .A2(n2093), .ZN(n2453) );
  INV_X1 U2372 ( .A(n2457), .ZN(n2456) );
  NAND2_X1 U2373 ( .A1(n2095), .A2(n2458), .ZN(n2452) );
  NAND2_X1 U2374 ( .A1(n2459), .A2(n2460), .ZN(n2442) );
  NAND3_X1 U2375 ( .A1(n2461), .A2(n2462), .A3(n2463), .ZN(n2460) );
  NAND2_X1 U2376 ( .A1(n2094), .A2(n2464), .ZN(n2463) );
  NAND2_X1 U2377 ( .A1(n2093), .A2(n2457), .ZN(n2462) );
  NAND2_X1 U2378 ( .A1(n2095), .A2(n2465), .ZN(n2461) );
  INV_X1 U2379 ( .A(n2450), .ZN(n2459) );
  XNOR2_X1 U2380 ( .A(n2466), .B(b_3_), .ZN(n2450) );
  NAND3_X1 U2381 ( .A1(n2467), .A2(n2468), .A3(n2469), .ZN(Result_18_) );
  NAND2_X1 U2382 ( .A1(n2096), .A2(n2470), .ZN(n2469) );
  XOR2_X1 U2383 ( .A(n2471), .B(n2472), .Z(n2470) );
  XNOR2_X1 U2384 ( .A(n2473), .B(n2474), .ZN(n2472) );
  NAND2_X1 U2385 ( .A1(a_2_), .A2(b_15_), .ZN(n2474) );
  NAND2_X1 U2386 ( .A1(n2475), .A2(n2476), .ZN(n2468) );
  NAND3_X1 U2387 ( .A1(n2477), .A2(n2478), .A3(n2479), .ZN(n2476) );
  NAND2_X1 U2388 ( .A1(n2094), .A2(n2480), .ZN(n2479) );
  NAND2_X1 U2389 ( .A1(n2481), .A2(n2093), .ZN(n2478) );
  INV_X1 U2390 ( .A(n2482), .ZN(n2481) );
  NAND2_X1 U2391 ( .A1(n2095), .A2(n2483), .ZN(n2477) );
  NAND2_X1 U2392 ( .A1(n2484), .A2(n2485), .ZN(n2467) );
  NAND3_X1 U2393 ( .A1(n2486), .A2(n2487), .A3(n2488), .ZN(n2485) );
  NAND2_X1 U2394 ( .A1(n2094), .A2(n2489), .ZN(n2488) );
  NAND2_X1 U2395 ( .A1(n2093), .A2(n2482), .ZN(n2487) );
  NAND2_X1 U2396 ( .A1(n2095), .A2(n2490), .ZN(n2486) );
  INV_X1 U2397 ( .A(n2475), .ZN(n2484) );
  XNOR2_X1 U2398 ( .A(n2491), .B(b_2_), .ZN(n2475) );
  NAND3_X1 U2399 ( .A1(n2492), .A2(n2493), .A3(n2494), .ZN(Result_17_) );
  NAND2_X1 U2400 ( .A1(n2096), .A2(n2495), .ZN(n2494) );
  XOR2_X1 U2401 ( .A(n2496), .B(n2497), .Z(n2495) );
  XNOR2_X1 U2402 ( .A(n2498), .B(n2499), .ZN(n2497) );
  NAND2_X1 U2403 ( .A1(a_1_), .A2(b_15_), .ZN(n2499) );
  NAND2_X1 U2404 ( .A1(n2500), .A2(n2501), .ZN(n2493) );
  NAND3_X1 U2405 ( .A1(n2502), .A2(n2503), .A3(n2504), .ZN(n2501) );
  NAND2_X1 U2406 ( .A1(n2094), .A2(n2505), .ZN(n2504) );
  NAND2_X1 U2407 ( .A1(n2506), .A2(n2093), .ZN(n2503) );
  NAND2_X1 U2408 ( .A1(n2095), .A2(n2507), .ZN(n2502) );
  NAND2_X1 U2409 ( .A1(n2508), .A2(n2509), .ZN(n2492) );
  NAND3_X1 U2410 ( .A1(n2510), .A2(n2511), .A3(n2512), .ZN(n2509) );
  NAND2_X1 U2411 ( .A1(n2094), .A2(n2513), .ZN(n2512) );
  NAND2_X1 U2412 ( .A1(n2093), .A2(n2514), .ZN(n2511) );
  NAND2_X1 U2413 ( .A1(n2095), .A2(n2515), .ZN(n2510) );
  INV_X1 U2414 ( .A(n2500), .ZN(n2508) );
  XNOR2_X1 U2415 ( .A(n2516), .B(b_1_), .ZN(n2500) );
  NAND3_X1 U2416 ( .A1(n2517), .A2(n2518), .A3(n2519), .ZN(Result_16_) );
  NAND2_X1 U2417 ( .A1(n2096), .A2(n2520), .ZN(n2519) );
  XOR2_X1 U2418 ( .A(n2521), .B(n2522), .Z(n2520) );
  XNOR2_X1 U2419 ( .A(n2523), .B(n2524), .ZN(n2522) );
  NAND2_X1 U2420 ( .A1(a_0_), .A2(b_15_), .ZN(n2524) );
  NAND2_X1 U2421 ( .A1(n2525), .A2(n2526), .ZN(n2518) );
  NAND3_X1 U2422 ( .A1(n2527), .A2(n2528), .A3(n2529), .ZN(n2526) );
  NAND2_X1 U2423 ( .A1(n2094), .A2(n2530), .ZN(n2529) );
  NAND2_X1 U2424 ( .A1(n2093), .A2(n2531), .ZN(n2528) );
  NAND2_X1 U2425 ( .A1(n2095), .A2(n2532), .ZN(n2527) );
  NAND2_X1 U2426 ( .A1(n2533), .A2(n2534), .ZN(n2517) );
  NAND3_X1 U2427 ( .A1(n2535), .A2(n2536), .A3(n2537), .ZN(n2534) );
  NAND2_X1 U2428 ( .A1(n2094), .A2(n2538), .ZN(n2537) );
  NAND2_X1 U2429 ( .A1(n2539), .A2(n2093), .ZN(n2536) );
  INV_X1 U2430 ( .A(n2531), .ZN(n2539) );
  NAND2_X1 U2431 ( .A1(n2540), .A2(n2541), .ZN(n2531) );
  NAND2_X1 U2432 ( .A1(n2506), .A2(n2542), .ZN(n2541) );
  INV_X1 U2433 ( .A(n2514), .ZN(n2506) );
  NAND2_X1 U2434 ( .A1(n2543), .A2(n2544), .ZN(n2514) );
  NAND2_X1 U2435 ( .A1(n2545), .A2(n2482), .ZN(n2544) );
  NAND2_X1 U2436 ( .A1(n2546), .A2(n2547), .ZN(n2482) );
  NAND2_X1 U2437 ( .A1(n2548), .A2(n2457), .ZN(n2547) );
  NAND2_X1 U2438 ( .A1(n2549), .A2(n2550), .ZN(n2457) );
  NAND2_X1 U2439 ( .A1(n2551), .A2(n2433), .ZN(n2550) );
  INV_X1 U2440 ( .A(n2425), .ZN(n2433) );
  NOR2_X1 U2441 ( .A1(n2552), .A2(n2553), .ZN(n2425) );
  AND2_X1 U2442 ( .A1(n2554), .A2(n2401), .ZN(n2553) );
  NAND2_X1 U2443 ( .A1(n2555), .A2(n2556), .ZN(n2401) );
  NAND2_X1 U2444 ( .A1(n2557), .A2(n2376), .ZN(n2556) );
  NAND2_X1 U2445 ( .A1(n2558), .A2(n2559), .ZN(n2376) );
  NAND2_X1 U2446 ( .A1(n2560), .A2(n2351), .ZN(n2559) );
  NAND2_X1 U2447 ( .A1(n2561), .A2(n2562), .ZN(n2351) );
  NAND2_X1 U2448 ( .A1(n2563), .A2(n2333), .ZN(n2562) );
  INV_X1 U2449 ( .A(n2325), .ZN(n2333) );
  NOR2_X1 U2450 ( .A1(n2564), .A2(n2565), .ZN(n2325) );
  AND2_X1 U2451 ( .A1(n2566), .A2(n2308), .ZN(n2565) );
  INV_X1 U2452 ( .A(n2300), .ZN(n2308) );
  NOR2_X1 U2453 ( .A1(n2567), .A2(n2568), .ZN(n2300) );
  AND2_X1 U2454 ( .A1(n2569), .A2(n2276), .ZN(n2568) );
  NAND2_X1 U2455 ( .A1(n2259), .A2(n2570), .ZN(n2276) );
  NAND2_X1 U2456 ( .A1(n2260), .A2(n2249), .ZN(n2570) );
  NAND2_X1 U2457 ( .A1(n2233), .A2(n2571), .ZN(n2249) );
  NAND2_X1 U2458 ( .A1(n2234), .A2(n2223), .ZN(n2571) );
  NAND2_X1 U2459 ( .A1(n2207), .A2(n2572), .ZN(n2223) );
  NAND2_X1 U2460 ( .A1(n2208), .A2(n2197), .ZN(n2572) );
  NAND2_X1 U2461 ( .A1(n2573), .A2(n2574), .ZN(n2197) );
  NAND2_X1 U2462 ( .A1(b_14_), .A2(n2575), .ZN(n2574) );
  NAND2_X1 U2463 ( .A1(n2158), .A2(n2168), .ZN(n2575) );
  NAND2_X1 U2464 ( .A1(a_15_), .A2(b_15_), .ZN(n2168) );
  NAND2_X1 U2465 ( .A1(n2576), .A2(b_15_), .ZN(n2573) );
  NAND2_X1 U2466 ( .A1(n2577), .A2(n2188), .ZN(n2208) );
  NAND2_X1 U2467 ( .A1(n2578), .A2(n2579), .ZN(n2234) );
  NAND2_X1 U2468 ( .A1(n2580), .A2(n2581), .ZN(n2260) );
  NAND2_X1 U2469 ( .A1(n2285), .A2(n2582), .ZN(n2569) );
  NAND2_X1 U2470 ( .A1(n2583), .A2(n2310), .ZN(n2566) );
  NAND2_X1 U2471 ( .A1(n2335), .A2(n2584), .ZN(n2563) );
  NAND2_X1 U2472 ( .A1(n2585), .A2(n2360), .ZN(n2560) );
  NAND2_X1 U2473 ( .A1(n2385), .A2(n2586), .ZN(n2557) );
  NAND2_X1 U2474 ( .A1(n2587), .A2(n2410), .ZN(n2554) );
  NAND2_X1 U2475 ( .A1(n2588), .A2(n2435), .ZN(n2551) );
  NAND2_X1 U2476 ( .A1(n2589), .A2(n2466), .ZN(n2548) );
  NAND2_X1 U2477 ( .A1(n2590), .A2(n2491), .ZN(n2545) );
  NAND2_X1 U2478 ( .A1(n2591), .A2(n2516), .ZN(n2540) );
  NAND2_X1 U2479 ( .A1(n2095), .A2(n2592), .ZN(n2535) );
  INV_X1 U2480 ( .A(n2525), .ZN(n2533) );
  XNOR2_X1 U2481 ( .A(n2593), .B(a_0_), .ZN(n2525) );
  NAND2_X1 U2482 ( .A1(n2097), .A2(n2594), .ZN(Result_15_) );
  NAND2_X1 U2483 ( .A1(n2595), .A2(n2096), .ZN(n2594) );
  XOR2_X1 U2484 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND2_X1 U2485 ( .A1(n2097), .A2(n2598), .ZN(Result_14_) );
  NAND3_X1 U2486 ( .A1(n2599), .A2(n2600), .A3(n2096), .ZN(n2598) );
  NAND2_X1 U2487 ( .A1(n2601), .A2(n2602), .ZN(n2599) );
  NAND2_X1 U2488 ( .A1(n2597), .A2(n2596), .ZN(n2602) );
  XNOR2_X1 U2489 ( .A(n2603), .B(n2604), .ZN(n2601) );
  NAND2_X1 U2490 ( .A1(n2097), .A2(n2605), .ZN(Result_13_) );
  NAND2_X1 U2491 ( .A1(n2096), .A2(n2606), .ZN(n2605) );
  XOR2_X1 U2492 ( .A(n2600), .B(n2607), .Z(n2606) );
  NAND2_X1 U2493 ( .A1(n2608), .A2(n2609), .ZN(n2607) );
  NAND2_X1 U2494 ( .A1(n2610), .A2(n2611), .ZN(n2609) );
  NAND2_X1 U2495 ( .A1(n2603), .A2(n2604), .ZN(n2610) );
  NAND2_X1 U2496 ( .A1(n2097), .A2(n2612), .ZN(Result_12_) );
  NAND2_X1 U2497 ( .A1(n2096), .A2(n2613), .ZN(n2612) );
  XOR2_X1 U2498 ( .A(n2614), .B(n2615), .Z(n2613) );
  NAND2_X1 U2499 ( .A1(n2097), .A2(n2616), .ZN(Result_11_) );
  NAND2_X1 U2500 ( .A1(n2096), .A2(n2617), .ZN(n2616) );
  XOR2_X1 U2501 ( .A(n2618), .B(n2619), .Z(n2617) );
  AND2_X1 U2502 ( .A1(n2620), .A2(n2621), .ZN(n2619) );
  NAND2_X1 U2503 ( .A1(n2097), .A2(n2622), .ZN(Result_10_) );
  NAND2_X1 U2504 ( .A1(n2623), .A2(n2096), .ZN(n2622) );
  XOR2_X1 U2505 ( .A(n2624), .B(n2625), .Z(n2623) );
  AND2_X1 U2506 ( .A1(n2626), .A2(n2627), .ZN(n2625) );
  NAND2_X1 U2507 ( .A1(n2097), .A2(n2628), .ZN(Result_0_) );
  NAND2_X1 U2508 ( .A1(n2096), .A2(n2629), .ZN(n2628) );
  NAND3_X1 U2509 ( .A1(n2630), .A2(n2441), .A3(n2631), .ZN(n2629) );
  NAND2_X1 U2510 ( .A1(a_0_), .A2(n2632), .ZN(n2631) );
  NAND4_X1 U2511 ( .A1(n2633), .A2(n2634), .A3(n2635), .A4(n2636), .ZN(n2441)
         );
  NAND2_X1 U2512 ( .A1(n2440), .A2(n2438), .ZN(n2630) );
  NAND2_X1 U2513 ( .A1(n2180), .A2(n2637), .ZN(n2438) );
  NAND2_X1 U2514 ( .A1(n2179), .A2(n2177), .ZN(n2637) );
  NAND2_X1 U2515 ( .A1(n2139), .A2(n2638), .ZN(n2177) );
  NAND2_X1 U2516 ( .A1(n2138), .A2(n2136), .ZN(n2638) );
  NAND2_X1 U2517 ( .A1(n2133), .A2(n2639), .ZN(n2136) );
  NAND2_X1 U2518 ( .A1(n2132), .A2(n2130), .ZN(n2639) );
  NAND2_X1 U2519 ( .A1(n2127), .A2(n2640), .ZN(n2130) );
  NAND2_X1 U2520 ( .A1(n2126), .A2(n2124), .ZN(n2640) );
  NAND2_X1 U2521 ( .A1(n2121), .A2(n2641), .ZN(n2124) );
  NAND2_X1 U2522 ( .A1(n2120), .A2(n2118), .ZN(n2641) );
  NAND2_X1 U2523 ( .A1(n2115), .A2(n2642), .ZN(n2118) );
  NAND2_X1 U2524 ( .A1(n2114), .A2(n2112), .ZN(n2642) );
  NAND2_X1 U2525 ( .A1(n2109), .A2(n2643), .ZN(n2112) );
  NAND2_X1 U2526 ( .A1(n2108), .A2(n2106), .ZN(n2643) );
  NAND2_X1 U2527 ( .A1(n2103), .A2(n2644), .ZN(n2106) );
  NAND2_X1 U2528 ( .A1(n2102), .A2(n2100), .ZN(n2644) );
  NAND2_X1 U2529 ( .A1(n2627), .A2(n2645), .ZN(n2100) );
  NAND2_X1 U2530 ( .A1(n2624), .A2(n2626), .ZN(n2645) );
  NAND2_X1 U2531 ( .A1(n2646), .A2(n2647), .ZN(n2626) );
  XNOR2_X1 U2532 ( .A(n2648), .B(n2649), .ZN(n2646) );
  NAND2_X1 U2533 ( .A1(n2621), .A2(n2650), .ZN(n2624) );
  NAND2_X1 U2534 ( .A1(n2618), .A2(n2620), .ZN(n2650) );
  NAND2_X1 U2535 ( .A1(n2651), .A2(n2652), .ZN(n2620) );
  NAND2_X1 U2536 ( .A1(n2653), .A2(n2647), .ZN(n2652) );
  NAND2_X1 U2537 ( .A1(n2654), .A2(n2655), .ZN(n2651) );
  NOR2_X1 U2538 ( .A1(n2615), .A2(n2614), .ZN(n2618) );
  AND3_X1 U2539 ( .A1(n2656), .A2(n2608), .A3(n2657), .ZN(n2614) );
  OR2_X1 U2540 ( .A1(n2600), .A2(n2611), .ZN(n2657) );
  NAND3_X1 U2541 ( .A1(n2658), .A2(n2596), .A3(n2597), .ZN(n2600) );
  XNOR2_X1 U2542 ( .A(n2659), .B(n2660), .ZN(n2597) );
  XOR2_X1 U2543 ( .A(n2661), .B(n2662), .Z(n2660) );
  NAND2_X1 U2544 ( .A1(b_14_), .A2(a_0_), .ZN(n2662) );
  NAND2_X1 U2545 ( .A1(n2663), .A2(n2664), .ZN(n2596) );
  NAND3_X1 U2546 ( .A1(b_15_), .A2(n2665), .A3(a_0_), .ZN(n2664) );
  NAND2_X1 U2547 ( .A1(n2523), .A2(n2521), .ZN(n2665) );
  OR2_X1 U2548 ( .A1(n2521), .A2(n2523), .ZN(n2663) );
  AND2_X1 U2549 ( .A1(n2666), .A2(n2667), .ZN(n2523) );
  NAND3_X1 U2550 ( .A1(b_15_), .A2(n2668), .A3(a_1_), .ZN(n2667) );
  NAND2_X1 U2551 ( .A1(n2498), .A2(n2496), .ZN(n2668) );
  OR2_X1 U2552 ( .A1(n2496), .A2(n2498), .ZN(n2666) );
  AND2_X1 U2553 ( .A1(n2669), .A2(n2670), .ZN(n2498) );
  NAND3_X1 U2554 ( .A1(b_15_), .A2(n2671), .A3(a_2_), .ZN(n2670) );
  NAND2_X1 U2555 ( .A1(n2473), .A2(n2471), .ZN(n2671) );
  OR2_X1 U2556 ( .A1(n2471), .A2(n2473), .ZN(n2669) );
  AND2_X1 U2557 ( .A1(n2672), .A2(n2673), .ZN(n2473) );
  NAND3_X1 U2558 ( .A1(b_15_), .A2(n2674), .A3(a_3_), .ZN(n2673) );
  OR2_X1 U2559 ( .A1(n2448), .A2(n2446), .ZN(n2674) );
  NAND2_X1 U2560 ( .A1(n2446), .A2(n2448), .ZN(n2672) );
  NAND2_X1 U2561 ( .A1(n2675), .A2(n2676), .ZN(n2448) );
  NAND3_X1 U2562 ( .A1(b_15_), .A2(n2677), .A3(a_4_), .ZN(n2676) );
  OR2_X1 U2563 ( .A1(n2417), .A2(n2415), .ZN(n2677) );
  NAND2_X1 U2564 ( .A1(n2415), .A2(n2417), .ZN(n2675) );
  NAND2_X1 U2565 ( .A1(n2392), .A2(n2678), .ZN(n2417) );
  NAND2_X1 U2566 ( .A1(n2391), .A2(n2393), .ZN(n2678) );
  NAND2_X1 U2567 ( .A1(n2679), .A2(n2680), .ZN(n2393) );
  NAND2_X1 U2568 ( .A1(a_5_), .A2(b_15_), .ZN(n2680) );
  INV_X1 U2569 ( .A(n2681), .ZN(n2679) );
  XNOR2_X1 U2570 ( .A(n2682), .B(n2683), .ZN(n2391) );
  XNOR2_X1 U2571 ( .A(n2684), .B(n2685), .ZN(n2682) );
  NOR2_X1 U2572 ( .A1(n2586), .A2(n2161), .ZN(n2685) );
  NAND2_X1 U2573 ( .A1(a_5_), .A2(n2681), .ZN(n2392) );
  NAND2_X1 U2574 ( .A1(n2686), .A2(n2687), .ZN(n2681) );
  NAND2_X1 U2575 ( .A1(n2365), .A2(n2688), .ZN(n2687) );
  OR2_X1 U2576 ( .A1(n2367), .A2(n2368), .ZN(n2688) );
  XOR2_X1 U2577 ( .A(n2689), .B(n2690), .Z(n2365) );
  XOR2_X1 U2578 ( .A(n2691), .B(n2692), .Z(n2689) );
  NAND2_X1 U2579 ( .A1(n2368), .A2(n2367), .ZN(n2686) );
  NAND2_X1 U2580 ( .A1(n2342), .A2(n2693), .ZN(n2367) );
  NAND2_X1 U2581 ( .A1(n2341), .A2(n2343), .ZN(n2693) );
  NAND2_X1 U2582 ( .A1(n2694), .A2(n2695), .ZN(n2343) );
  NAND2_X1 U2583 ( .A1(a_7_), .A2(b_15_), .ZN(n2695) );
  INV_X1 U2584 ( .A(n2696), .ZN(n2694) );
  XOR2_X1 U2585 ( .A(n2697), .B(n2698), .Z(n2341) );
  XNOR2_X1 U2586 ( .A(n2699), .B(n2700), .ZN(n2697) );
  NAND2_X1 U2587 ( .A1(b_14_), .A2(a_8_), .ZN(n2699) );
  NAND2_X1 U2588 ( .A1(a_7_), .A2(n2696), .ZN(n2342) );
  NAND2_X1 U2589 ( .A1(n2701), .A2(n2702), .ZN(n2696) );
  NAND2_X1 U2590 ( .A1(n2315), .A2(n2703), .ZN(n2702) );
  OR2_X1 U2591 ( .A1(n2317), .A2(n2318), .ZN(n2703) );
  XNOR2_X1 U2592 ( .A(n2704), .B(n2705), .ZN(n2315) );
  XNOR2_X1 U2593 ( .A(n2706), .B(n2707), .ZN(n2705) );
  NAND2_X1 U2594 ( .A1(n2318), .A2(n2317), .ZN(n2701) );
  NAND2_X1 U2595 ( .A1(n2292), .A2(n2708), .ZN(n2317) );
  NAND2_X1 U2596 ( .A1(n2291), .A2(n2293), .ZN(n2708) );
  NAND2_X1 U2597 ( .A1(n2709), .A2(n2710), .ZN(n2293) );
  NAND2_X1 U2598 ( .A1(a_9_), .A2(b_15_), .ZN(n2710) );
  INV_X1 U2599 ( .A(n2711), .ZN(n2709) );
  XNOR2_X1 U2600 ( .A(n2712), .B(n2713), .ZN(n2291) );
  XOR2_X1 U2601 ( .A(n2714), .B(n2715), .Z(n2713) );
  NAND2_X1 U2602 ( .A1(b_14_), .A2(a_10_), .ZN(n2715) );
  NAND2_X1 U2603 ( .A1(a_9_), .A2(n2711), .ZN(n2292) );
  NAND2_X1 U2604 ( .A1(n2716), .A2(n2717), .ZN(n2711) );
  NAND2_X1 U2605 ( .A1(n2265), .A2(n2718), .ZN(n2717) );
  OR2_X1 U2606 ( .A1(n2267), .A2(n2268), .ZN(n2718) );
  XOR2_X1 U2607 ( .A(n2719), .B(n2720), .Z(n2265) );
  XOR2_X1 U2608 ( .A(n2721), .B(n2722), .Z(n2719) );
  NAND2_X1 U2609 ( .A1(n2268), .A2(n2267), .ZN(n2716) );
  NAND2_X1 U2610 ( .A1(n2241), .A2(n2723), .ZN(n2267) );
  NAND2_X1 U2611 ( .A1(n2240), .A2(n2242), .ZN(n2723) );
  NAND2_X1 U2612 ( .A1(n2724), .A2(n2725), .ZN(n2242) );
  NAND2_X1 U2613 ( .A1(a_11_), .A2(b_15_), .ZN(n2725) );
  INV_X1 U2614 ( .A(n2726), .ZN(n2724) );
  XNOR2_X1 U2615 ( .A(n2727), .B(n2728), .ZN(n2240) );
  XOR2_X1 U2616 ( .A(n2729), .B(n2730), .Z(n2727) );
  NAND2_X1 U2617 ( .A1(b_14_), .A2(a_12_), .ZN(n2729) );
  NAND2_X1 U2618 ( .A1(a_11_), .A2(n2726), .ZN(n2241) );
  NAND2_X1 U2619 ( .A1(n2731), .A2(n2732), .ZN(n2726) );
  NAND2_X1 U2620 ( .A1(n2216), .A2(n2733), .ZN(n2732) );
  OR2_X1 U2621 ( .A1(n2215), .A2(n2213), .ZN(n2733) );
  NOR2_X1 U2622 ( .A1(n2579), .A2(n2187), .ZN(n2216) );
  NAND2_X1 U2623 ( .A1(n2213), .A2(n2215), .ZN(n2731) );
  NAND2_X1 U2624 ( .A1(n2734), .A2(n2735), .ZN(n2215) );
  NAND3_X1 U2625 ( .A1(b_15_), .A2(n2736), .A3(a_13_), .ZN(n2735) );
  OR2_X1 U2626 ( .A1(n2189), .A2(n2190), .ZN(n2736) );
  NAND2_X1 U2627 ( .A1(n2190), .A2(n2189), .ZN(n2734) );
  NAND2_X1 U2628 ( .A1(n2737), .A2(n2738), .ZN(n2189) );
  NAND2_X1 U2629 ( .A1(b_13_), .A2(n2739), .ZN(n2738) );
  NAND2_X1 U2630 ( .A1(n2156), .A2(n2740), .ZN(n2739) );
  NAND2_X1 U2631 ( .A1(a_15_), .A2(n2161), .ZN(n2740) );
  NAND2_X1 U2632 ( .A1(b_14_), .A2(n2741), .ZN(n2737) );
  NAND2_X1 U2633 ( .A1(n2742), .A2(n2743), .ZN(n2741) );
  NAND2_X1 U2634 ( .A1(a_14_), .A2(n2577), .ZN(n2743) );
  AND3_X1 U2635 ( .A1(b_14_), .A2(b_15_), .A3(n2576), .ZN(n2190) );
  XOR2_X1 U2636 ( .A(n2744), .B(n2745), .Z(n2213) );
  XOR2_X1 U2637 ( .A(n2746), .B(n2747), .Z(n2744) );
  NOR2_X1 U2638 ( .A1(n2582), .A2(n2187), .ZN(n2268) );
  NOR2_X1 U2639 ( .A1(n2584), .A2(n2187), .ZN(n2318) );
  NOR2_X1 U2640 ( .A1(n2586), .A2(n2187), .ZN(n2368) );
  XNOR2_X1 U2641 ( .A(n2748), .B(n2749), .ZN(n2415) );
  XNOR2_X1 U2642 ( .A(n2750), .B(n2751), .ZN(n2748) );
  XNOR2_X1 U2643 ( .A(n2752), .B(n2753), .ZN(n2446) );
  XNOR2_X1 U2644 ( .A(n2754), .B(n2755), .ZN(n2752) );
  NOR2_X1 U2645 ( .A1(n2435), .A2(n2161), .ZN(n2755) );
  XOR2_X1 U2646 ( .A(n2756), .B(n2757), .Z(n2471) );
  XNOR2_X1 U2647 ( .A(n2758), .B(n2759), .ZN(n2757) );
  XOR2_X1 U2648 ( .A(n2760), .B(n2761), .Z(n2496) );
  XOR2_X1 U2649 ( .A(n2762), .B(n2763), .Z(n2761) );
  NAND2_X1 U2650 ( .A1(b_14_), .A2(a_2_), .ZN(n2763) );
  XNOR2_X1 U2651 ( .A(n2764), .B(n2765), .ZN(n2521) );
  XOR2_X1 U2652 ( .A(n2766), .B(n2767), .Z(n2764) );
  NOR2_X1 U2653 ( .A1(n2516), .A2(n2161), .ZN(n2767) );
  XOR2_X1 U2654 ( .A(n2604), .B(n2603), .Z(n2658) );
  NAND3_X1 U2655 ( .A1(n2603), .A2(n2604), .A3(n2768), .ZN(n2608) );
  INV_X1 U2656 ( .A(n2611), .ZN(n2768) );
  NAND2_X1 U2657 ( .A1(n2656), .A2(n2769), .ZN(n2611) );
  NAND2_X1 U2658 ( .A1(n2770), .A2(n2771), .ZN(n2769) );
  NAND2_X1 U2659 ( .A1(n2772), .A2(n2773), .ZN(n2604) );
  NAND3_X1 U2660 ( .A1(a_0_), .A2(n2774), .A3(b_14_), .ZN(n2773) );
  OR2_X1 U2661 ( .A1(n2661), .A2(n2659), .ZN(n2774) );
  NAND2_X1 U2662 ( .A1(n2659), .A2(n2661), .ZN(n2772) );
  NAND2_X1 U2663 ( .A1(n2775), .A2(n2776), .ZN(n2661) );
  NAND3_X1 U2664 ( .A1(a_1_), .A2(n2777), .A3(b_14_), .ZN(n2776) );
  OR2_X1 U2665 ( .A1(n2766), .A2(n2765), .ZN(n2777) );
  NAND2_X1 U2666 ( .A1(n2765), .A2(n2766), .ZN(n2775) );
  NAND2_X1 U2667 ( .A1(n2778), .A2(n2779), .ZN(n2766) );
  NAND3_X1 U2668 ( .A1(a_2_), .A2(n2780), .A3(b_14_), .ZN(n2779) );
  OR2_X1 U2669 ( .A1(n2762), .A2(n2760), .ZN(n2780) );
  NAND2_X1 U2670 ( .A1(n2760), .A2(n2762), .ZN(n2778) );
  NAND2_X1 U2671 ( .A1(n2781), .A2(n2782), .ZN(n2762) );
  NAND2_X1 U2672 ( .A1(n2759), .A2(n2783), .ZN(n2782) );
  OR2_X1 U2673 ( .A1(n2758), .A2(n2756), .ZN(n2783) );
  NOR2_X1 U2674 ( .A1(n2161), .A2(n2466), .ZN(n2759) );
  NAND2_X1 U2675 ( .A1(n2756), .A2(n2758), .ZN(n2781) );
  NAND2_X1 U2676 ( .A1(n2784), .A2(n2785), .ZN(n2758) );
  NAND3_X1 U2677 ( .A1(a_4_), .A2(n2786), .A3(b_14_), .ZN(n2785) );
  NAND2_X1 U2678 ( .A1(n2754), .A2(n2753), .ZN(n2786) );
  OR2_X1 U2679 ( .A1(n2753), .A2(n2754), .ZN(n2784) );
  AND2_X1 U2680 ( .A1(n2787), .A2(n2788), .ZN(n2754) );
  NAND2_X1 U2681 ( .A1(n2751), .A2(n2789), .ZN(n2788) );
  NAND2_X1 U2682 ( .A1(n2750), .A2(n2749), .ZN(n2789) );
  NOR2_X1 U2683 ( .A1(n2161), .A2(n2410), .ZN(n2751) );
  OR2_X1 U2684 ( .A1(n2749), .A2(n2750), .ZN(n2787) );
  AND2_X1 U2685 ( .A1(n2790), .A2(n2791), .ZN(n2750) );
  NAND3_X1 U2686 ( .A1(a_6_), .A2(n2792), .A3(b_14_), .ZN(n2791) );
  NAND2_X1 U2687 ( .A1(n2684), .A2(n2683), .ZN(n2792) );
  OR2_X1 U2688 ( .A1(n2683), .A2(n2684), .ZN(n2790) );
  AND2_X1 U2689 ( .A1(n2793), .A2(n2794), .ZN(n2684) );
  NAND2_X1 U2690 ( .A1(n2692), .A2(n2795), .ZN(n2794) );
  OR2_X1 U2691 ( .A1(n2691), .A2(n2690), .ZN(n2795) );
  NOR2_X1 U2692 ( .A1(n2161), .A2(n2360), .ZN(n2692) );
  NAND2_X1 U2693 ( .A1(n2690), .A2(n2691), .ZN(n2793) );
  NAND2_X1 U2694 ( .A1(n2796), .A2(n2797), .ZN(n2691) );
  NAND3_X1 U2695 ( .A1(a_8_), .A2(n2798), .A3(b_14_), .ZN(n2797) );
  OR2_X1 U2696 ( .A1(n2700), .A2(n2698), .ZN(n2798) );
  NAND2_X1 U2697 ( .A1(n2698), .A2(n2700), .ZN(n2796) );
  NAND2_X1 U2698 ( .A1(n2799), .A2(n2800), .ZN(n2700) );
  NAND2_X1 U2699 ( .A1(n2707), .A2(n2801), .ZN(n2800) );
  OR2_X1 U2700 ( .A1(n2706), .A2(n2704), .ZN(n2801) );
  NOR2_X1 U2701 ( .A1(n2161), .A2(n2310), .ZN(n2707) );
  NAND2_X1 U2702 ( .A1(n2704), .A2(n2706), .ZN(n2799) );
  NAND2_X1 U2703 ( .A1(n2802), .A2(n2803), .ZN(n2706) );
  NAND3_X1 U2704 ( .A1(a_10_), .A2(n2804), .A3(b_14_), .ZN(n2803) );
  OR2_X1 U2705 ( .A1(n2714), .A2(n2712), .ZN(n2804) );
  NAND2_X1 U2706 ( .A1(n2712), .A2(n2714), .ZN(n2802) );
  NAND2_X1 U2707 ( .A1(n2805), .A2(n2806), .ZN(n2714) );
  NAND2_X1 U2708 ( .A1(n2722), .A2(n2807), .ZN(n2806) );
  OR2_X1 U2709 ( .A1(n2721), .A2(n2720), .ZN(n2807) );
  NOR2_X1 U2710 ( .A1(n2161), .A2(n2581), .ZN(n2722) );
  NAND2_X1 U2711 ( .A1(n2720), .A2(n2721), .ZN(n2805) );
  NAND2_X1 U2712 ( .A1(n2808), .A2(n2809), .ZN(n2721) );
  NAND3_X1 U2713 ( .A1(a_12_), .A2(n2810), .A3(b_14_), .ZN(n2809) );
  NAND2_X1 U2714 ( .A1(n2730), .A2(n2728), .ZN(n2810) );
  OR2_X1 U2715 ( .A1(n2728), .A2(n2730), .ZN(n2808) );
  AND2_X1 U2716 ( .A1(n2811), .A2(n2812), .ZN(n2730) );
  NAND2_X1 U2717 ( .A1(n2745), .A2(n2813), .ZN(n2812) );
  OR2_X1 U2718 ( .A1(n2746), .A2(n2747), .ZN(n2813) );
  NOR2_X1 U2719 ( .A1(n2161), .A2(n2188), .ZN(n2745) );
  NAND2_X1 U2720 ( .A1(n2747), .A2(n2746), .ZN(n2811) );
  NAND2_X1 U2721 ( .A1(n2814), .A2(n2815), .ZN(n2746) );
  NAND2_X1 U2722 ( .A1(b_12_), .A2(n2816), .ZN(n2815) );
  NAND2_X1 U2723 ( .A1(n2156), .A2(n2817), .ZN(n2816) );
  NAND2_X1 U2724 ( .A1(a_15_), .A2(n2577), .ZN(n2817) );
  NAND2_X1 U2725 ( .A1(b_13_), .A2(n2818), .ZN(n2814) );
  NAND2_X1 U2726 ( .A1(n2742), .A2(n2819), .ZN(n2818) );
  NAND2_X1 U2727 ( .A1(a_14_), .A2(n2578), .ZN(n2819) );
  AND3_X1 U2728 ( .A1(b_13_), .A2(b_14_), .A3(n2576), .ZN(n2747) );
  XNOR2_X1 U2729 ( .A(n2820), .B(n2821), .ZN(n2728) );
  XOR2_X1 U2730 ( .A(n2822), .B(n2823), .Z(n2820) );
  XNOR2_X1 U2731 ( .A(n2824), .B(n2825), .ZN(n2720) );
  XOR2_X1 U2732 ( .A(n2826), .B(n2827), .Z(n2824) );
  NAND2_X1 U2733 ( .A1(b_13_), .A2(a_12_), .ZN(n2826) );
  XNOR2_X1 U2734 ( .A(n2828), .B(n2829), .ZN(n2712) );
  NAND2_X1 U2735 ( .A1(n2830), .A2(n2831), .ZN(n2828) );
  XNOR2_X1 U2736 ( .A(n2832), .B(n2833), .ZN(n2704) );
  NAND2_X1 U2737 ( .A1(n2834), .A2(n2835), .ZN(n2832) );
  XNOR2_X1 U2738 ( .A(n2836), .B(n2837), .ZN(n2698) );
  XNOR2_X1 U2739 ( .A(n2838), .B(n2839), .ZN(n2836) );
  XNOR2_X1 U2740 ( .A(n2840), .B(n2841), .ZN(n2690) );
  XOR2_X1 U2741 ( .A(n2842), .B(n2843), .Z(n2841) );
  NAND2_X1 U2742 ( .A1(b_13_), .A2(a_8_), .ZN(n2843) );
  XOR2_X1 U2743 ( .A(n2844), .B(n2845), .Z(n2683) );
  XOR2_X1 U2744 ( .A(n2846), .B(n2847), .Z(n2845) );
  NAND2_X1 U2745 ( .A1(b_13_), .A2(a_7_), .ZN(n2847) );
  XOR2_X1 U2746 ( .A(n2848), .B(n2849), .Z(n2749) );
  NAND2_X1 U2747 ( .A1(n2850), .A2(n2851), .ZN(n2848) );
  XNOR2_X1 U2748 ( .A(n2852), .B(n2853), .ZN(n2753) );
  XOR2_X1 U2749 ( .A(n2854), .B(n2855), .Z(n2852) );
  XNOR2_X1 U2750 ( .A(n2856), .B(n2857), .ZN(n2756) );
  XNOR2_X1 U2751 ( .A(n2858), .B(n2859), .ZN(n2856) );
  NOR2_X1 U2752 ( .A1(n2435), .A2(n2577), .ZN(n2859) );
  XNOR2_X1 U2753 ( .A(n2860), .B(n2861), .ZN(n2760) );
  NAND2_X1 U2754 ( .A1(n2862), .A2(n2863), .ZN(n2860) );
  XNOR2_X1 U2755 ( .A(n2864), .B(n2865), .ZN(n2765) );
  XNOR2_X1 U2756 ( .A(n2866), .B(n2867), .ZN(n2865) );
  XNOR2_X1 U2757 ( .A(n2868), .B(n2869), .ZN(n2659) );
  XOR2_X1 U2758 ( .A(n2870), .B(n2871), .Z(n2869) );
  NAND2_X1 U2759 ( .A1(b_13_), .A2(a_1_), .ZN(n2871) );
  XOR2_X1 U2760 ( .A(n2872), .B(n2873), .Z(n2603) );
  XNOR2_X1 U2761 ( .A(n2874), .B(n2875), .ZN(n2873) );
  OR2_X1 U2762 ( .A1(n2771), .A2(n2770), .ZN(n2656) );
  XOR2_X1 U2763 ( .A(n2876), .B(n2877), .Z(n2770) );
  XOR2_X1 U2764 ( .A(n2878), .B(n2879), .Z(n2876) );
  NAND2_X1 U2765 ( .A1(b_12_), .A2(a_0_), .ZN(n2878) );
  NAND2_X1 U2766 ( .A1(n2880), .A2(n2881), .ZN(n2771) );
  NAND2_X1 U2767 ( .A1(n2874), .A2(n2882), .ZN(n2881) );
  OR2_X1 U2768 ( .A1(n2875), .A2(n2872), .ZN(n2882) );
  AND2_X1 U2769 ( .A1(n2883), .A2(n2884), .ZN(n2874) );
  NAND3_X1 U2770 ( .A1(a_1_), .A2(n2885), .A3(b_13_), .ZN(n2884) );
  OR2_X1 U2771 ( .A1(n2870), .A2(n2868), .ZN(n2885) );
  NAND2_X1 U2772 ( .A1(n2868), .A2(n2870), .ZN(n2883) );
  NAND2_X1 U2773 ( .A1(n2886), .A2(n2887), .ZN(n2870) );
  NAND2_X1 U2774 ( .A1(n2867), .A2(n2888), .ZN(n2887) );
  OR2_X1 U2775 ( .A1(n2866), .A2(n2864), .ZN(n2888) );
  NOR2_X1 U2776 ( .A1(n2577), .A2(n2491), .ZN(n2867) );
  NAND2_X1 U2777 ( .A1(n2864), .A2(n2866), .ZN(n2886) );
  NAND2_X1 U2778 ( .A1(n2862), .A2(n2889), .ZN(n2866) );
  NAND2_X1 U2779 ( .A1(n2861), .A2(n2863), .ZN(n2889) );
  NAND2_X1 U2780 ( .A1(n2890), .A2(n2891), .ZN(n2863) );
  NAND2_X1 U2781 ( .A1(b_13_), .A2(a_3_), .ZN(n2891) );
  INV_X1 U2782 ( .A(n2892), .ZN(n2890) );
  XNOR2_X1 U2783 ( .A(n2893), .B(n2894), .ZN(n2861) );
  XNOR2_X1 U2784 ( .A(n2895), .B(n2896), .ZN(n2893) );
  NOR2_X1 U2785 ( .A1(n2435), .A2(n2578), .ZN(n2896) );
  NAND2_X1 U2786 ( .A1(a_3_), .A2(n2892), .ZN(n2862) );
  NAND2_X1 U2787 ( .A1(n2897), .A2(n2898), .ZN(n2892) );
  NAND3_X1 U2788 ( .A1(a_4_), .A2(n2899), .A3(b_13_), .ZN(n2898) );
  NAND2_X1 U2789 ( .A1(n2858), .A2(n2857), .ZN(n2899) );
  OR2_X1 U2790 ( .A1(n2857), .A2(n2858), .ZN(n2897) );
  AND2_X1 U2791 ( .A1(n2900), .A2(n2901), .ZN(n2858) );
  NAND2_X1 U2792 ( .A1(n2855), .A2(n2902), .ZN(n2901) );
  OR2_X1 U2793 ( .A1(n2854), .A2(n2853), .ZN(n2902) );
  NOR2_X1 U2794 ( .A1(n2577), .A2(n2410), .ZN(n2855) );
  NAND2_X1 U2795 ( .A1(n2853), .A2(n2854), .ZN(n2900) );
  NAND2_X1 U2796 ( .A1(n2850), .A2(n2903), .ZN(n2854) );
  NAND2_X1 U2797 ( .A1(n2849), .A2(n2851), .ZN(n2903) );
  NAND2_X1 U2798 ( .A1(n2904), .A2(n2905), .ZN(n2851) );
  NAND2_X1 U2799 ( .A1(b_13_), .A2(a_6_), .ZN(n2905) );
  INV_X1 U2800 ( .A(n2906), .ZN(n2904) );
  XOR2_X1 U2801 ( .A(n2907), .B(n2908), .Z(n2849) );
  XOR2_X1 U2802 ( .A(n2909), .B(n2910), .Z(n2907) );
  NAND2_X1 U2803 ( .A1(a_6_), .A2(n2906), .ZN(n2850) );
  NAND2_X1 U2804 ( .A1(n2911), .A2(n2912), .ZN(n2906) );
  NAND3_X1 U2805 ( .A1(a_7_), .A2(n2913), .A3(b_13_), .ZN(n2912) );
  OR2_X1 U2806 ( .A1(n2846), .A2(n2844), .ZN(n2913) );
  NAND2_X1 U2807 ( .A1(n2844), .A2(n2846), .ZN(n2911) );
  NAND2_X1 U2808 ( .A1(n2914), .A2(n2915), .ZN(n2846) );
  NAND3_X1 U2809 ( .A1(a_8_), .A2(n2916), .A3(b_13_), .ZN(n2915) );
  OR2_X1 U2810 ( .A1(n2842), .A2(n2840), .ZN(n2916) );
  NAND2_X1 U2811 ( .A1(n2840), .A2(n2842), .ZN(n2914) );
  NAND2_X1 U2812 ( .A1(n2917), .A2(n2918), .ZN(n2842) );
  NAND2_X1 U2813 ( .A1(n2838), .A2(n2919), .ZN(n2918) );
  NAND2_X1 U2814 ( .A1(n2839), .A2(n2837), .ZN(n2919) );
  NOR2_X1 U2815 ( .A1(n2577), .A2(n2310), .ZN(n2838) );
  OR2_X1 U2816 ( .A1(n2837), .A2(n2839), .ZN(n2917) );
  AND2_X1 U2817 ( .A1(n2834), .A2(n2920), .ZN(n2839) );
  NAND2_X1 U2818 ( .A1(n2833), .A2(n2835), .ZN(n2920) );
  NAND2_X1 U2819 ( .A1(n2921), .A2(n2922), .ZN(n2835) );
  NAND2_X1 U2820 ( .A1(b_13_), .A2(a_10_), .ZN(n2922) );
  INV_X1 U2821 ( .A(n2923), .ZN(n2921) );
  XNOR2_X1 U2822 ( .A(n2924), .B(n2925), .ZN(n2833) );
  NAND2_X1 U2823 ( .A1(n2926), .A2(n2927), .ZN(n2924) );
  NAND2_X1 U2824 ( .A1(a_10_), .A2(n2923), .ZN(n2834) );
  NAND2_X1 U2825 ( .A1(n2830), .A2(n2928), .ZN(n2923) );
  NAND2_X1 U2826 ( .A1(n2829), .A2(n2831), .ZN(n2928) );
  NAND2_X1 U2827 ( .A1(n2929), .A2(n2930), .ZN(n2831) );
  NAND2_X1 U2828 ( .A1(b_13_), .A2(a_11_), .ZN(n2930) );
  INV_X1 U2829 ( .A(n2931), .ZN(n2929) );
  XOR2_X1 U2830 ( .A(n2932), .B(n2933), .Z(n2829) );
  XOR2_X1 U2831 ( .A(n2233), .B(n2934), .Z(n2932) );
  NAND2_X1 U2832 ( .A1(a_11_), .A2(n2931), .ZN(n2830) );
  NAND2_X1 U2833 ( .A1(n2935), .A2(n2936), .ZN(n2931) );
  NAND3_X1 U2834 ( .A1(a_12_), .A2(n2937), .A3(b_13_), .ZN(n2936) );
  NAND2_X1 U2835 ( .A1(n2827), .A2(n2825), .ZN(n2937) );
  OR2_X1 U2836 ( .A1(n2825), .A2(n2827), .ZN(n2935) );
  AND2_X1 U2837 ( .A1(n2938), .A2(n2939), .ZN(n2827) );
  NAND2_X1 U2838 ( .A1(n2821), .A2(n2940), .ZN(n2939) );
  OR2_X1 U2839 ( .A1(n2822), .A2(n2823), .ZN(n2940) );
  INV_X1 U2840 ( .A(n2207), .ZN(n2821) );
  NAND2_X1 U2841 ( .A1(b_13_), .A2(a_13_), .ZN(n2207) );
  NAND2_X1 U2842 ( .A1(n2823), .A2(n2822), .ZN(n2938) );
  NAND2_X1 U2843 ( .A1(n2941), .A2(n2942), .ZN(n2822) );
  NAND2_X1 U2844 ( .A1(b_11_), .A2(n2943), .ZN(n2942) );
  NAND2_X1 U2845 ( .A1(n2156), .A2(n2944), .ZN(n2943) );
  NAND2_X1 U2846 ( .A1(a_15_), .A2(n2578), .ZN(n2944) );
  NAND2_X1 U2847 ( .A1(b_12_), .A2(n2945), .ZN(n2941) );
  NAND2_X1 U2848 ( .A1(n2742), .A2(n2946), .ZN(n2945) );
  NAND2_X1 U2849 ( .A1(a_14_), .A2(n2580), .ZN(n2946) );
  AND3_X1 U2850 ( .A1(b_12_), .A2(b_13_), .A3(n2576), .ZN(n2823) );
  XNOR2_X1 U2851 ( .A(n2947), .B(n2948), .ZN(n2825) );
  XOR2_X1 U2852 ( .A(n2949), .B(n2950), .Z(n2947) );
  XNOR2_X1 U2853 ( .A(n2951), .B(n2952), .ZN(n2837) );
  NOR2_X1 U2854 ( .A1(n2953), .A2(n2954), .ZN(n2952) );
  NOR2_X1 U2855 ( .A1(n2955), .A2(n2956), .ZN(n2953) );
  NOR2_X1 U2856 ( .A1(n2582), .A2(n2578), .ZN(n2955) );
  XOR2_X1 U2857 ( .A(n2957), .B(n2958), .Z(n2840) );
  XOR2_X1 U2858 ( .A(n2959), .B(n2960), .Z(n2957) );
  XNOR2_X1 U2859 ( .A(n2961), .B(n2962), .ZN(n2844) );
  XNOR2_X1 U2860 ( .A(n2963), .B(n2964), .ZN(n2961) );
  NOR2_X1 U2861 ( .A1(n2584), .A2(n2578), .ZN(n2964) );
  XNOR2_X1 U2862 ( .A(n2965), .B(n2966), .ZN(n2853) );
  XOR2_X1 U2863 ( .A(n2967), .B(n2968), .Z(n2966) );
  NAND2_X1 U2864 ( .A1(b_12_), .A2(a_6_), .ZN(n2968) );
  XNOR2_X1 U2865 ( .A(n2969), .B(n2970), .ZN(n2857) );
  XOR2_X1 U2866 ( .A(n2971), .B(n2972), .Z(n2969) );
  XNOR2_X1 U2867 ( .A(n2973), .B(n2974), .ZN(n2864) );
  NAND2_X1 U2868 ( .A1(n2975), .A2(n2976), .ZN(n2973) );
  XNOR2_X1 U2869 ( .A(n2977), .B(n2978), .ZN(n2868) );
  XNOR2_X1 U2870 ( .A(n2979), .B(n2980), .ZN(n2978) );
  NAND2_X1 U2871 ( .A1(n2872), .A2(n2875), .ZN(n2880) );
  NAND2_X1 U2872 ( .A1(b_13_), .A2(a_0_), .ZN(n2875) );
  XOR2_X1 U2873 ( .A(n2981), .B(n2982), .Z(n2872) );
  XNOR2_X1 U2874 ( .A(n2983), .B(n2984), .ZN(n2982) );
  XNOR2_X1 U2875 ( .A(n2655), .B(n2654), .ZN(n2615) );
  NAND4_X1 U2876 ( .A1(n2654), .A2(n2653), .A3(n2655), .A4(n2647), .ZN(n2621)
         );
  INV_X1 U2877 ( .A(n2985), .ZN(n2647) );
  NAND2_X1 U2878 ( .A1(n2986), .A2(n2987), .ZN(n2655) );
  NAND3_X1 U2879 ( .A1(a_0_), .A2(n2988), .A3(b_12_), .ZN(n2987) );
  NAND2_X1 U2880 ( .A1(n2879), .A2(n2877), .ZN(n2988) );
  OR2_X1 U2881 ( .A1(n2877), .A2(n2879), .ZN(n2986) );
  AND2_X1 U2882 ( .A1(n2989), .A2(n2990), .ZN(n2879) );
  NAND2_X1 U2883 ( .A1(n2984), .A2(n2991), .ZN(n2990) );
  OR2_X1 U2884 ( .A1(n2983), .A2(n2981), .ZN(n2991) );
  NOR2_X1 U2885 ( .A1(n2578), .A2(n2516), .ZN(n2984) );
  NAND2_X1 U2886 ( .A1(n2981), .A2(n2983), .ZN(n2989) );
  NAND2_X1 U2887 ( .A1(n2992), .A2(n2993), .ZN(n2983) );
  NAND2_X1 U2888 ( .A1(n2980), .A2(n2994), .ZN(n2993) );
  OR2_X1 U2889 ( .A1(n2979), .A2(n2977), .ZN(n2994) );
  NOR2_X1 U2890 ( .A1(n2578), .A2(n2491), .ZN(n2980) );
  NAND2_X1 U2891 ( .A1(n2977), .A2(n2979), .ZN(n2992) );
  NAND2_X1 U2892 ( .A1(n2975), .A2(n2995), .ZN(n2979) );
  NAND2_X1 U2893 ( .A1(n2974), .A2(n2976), .ZN(n2995) );
  NAND2_X1 U2894 ( .A1(n2996), .A2(n2997), .ZN(n2976) );
  NAND2_X1 U2895 ( .A1(b_12_), .A2(a_3_), .ZN(n2997) );
  INV_X1 U2896 ( .A(n2998), .ZN(n2996) );
  XOR2_X1 U2897 ( .A(n2999), .B(n3000), .Z(n2974) );
  XOR2_X1 U2898 ( .A(n3001), .B(n3002), .Z(n2999) );
  NOR2_X1 U2899 ( .A1(n2435), .A2(n2580), .ZN(n3002) );
  NAND2_X1 U2900 ( .A1(a_3_), .A2(n2998), .ZN(n2975) );
  NAND2_X1 U2901 ( .A1(n3003), .A2(n3004), .ZN(n2998) );
  NAND3_X1 U2902 ( .A1(a_4_), .A2(n3005), .A3(b_12_), .ZN(n3004) );
  NAND2_X1 U2903 ( .A1(n2895), .A2(n2894), .ZN(n3005) );
  OR2_X1 U2904 ( .A1(n2894), .A2(n2895), .ZN(n3003) );
  AND2_X1 U2905 ( .A1(n3006), .A2(n3007), .ZN(n2895) );
  NAND2_X1 U2906 ( .A1(n2972), .A2(n3008), .ZN(n3007) );
  OR2_X1 U2907 ( .A1(n2971), .A2(n2970), .ZN(n3008) );
  NOR2_X1 U2908 ( .A1(n2578), .A2(n2410), .ZN(n2972) );
  NAND2_X1 U2909 ( .A1(n2970), .A2(n2971), .ZN(n3006) );
  NAND2_X1 U2910 ( .A1(n3009), .A2(n3010), .ZN(n2971) );
  NAND3_X1 U2911 ( .A1(a_6_), .A2(n3011), .A3(b_12_), .ZN(n3010) );
  OR2_X1 U2912 ( .A1(n2967), .A2(n2965), .ZN(n3011) );
  NAND2_X1 U2913 ( .A1(n2965), .A2(n2967), .ZN(n3009) );
  NAND2_X1 U2914 ( .A1(n3012), .A2(n3013), .ZN(n2967) );
  NAND2_X1 U2915 ( .A1(n2910), .A2(n3014), .ZN(n3013) );
  OR2_X1 U2916 ( .A1(n2909), .A2(n2908), .ZN(n3014) );
  NOR2_X1 U2917 ( .A1(n2578), .A2(n2360), .ZN(n2910) );
  NAND2_X1 U2918 ( .A1(n2908), .A2(n2909), .ZN(n3012) );
  NAND2_X1 U2919 ( .A1(n3015), .A2(n3016), .ZN(n2909) );
  NAND3_X1 U2920 ( .A1(a_8_), .A2(n3017), .A3(b_12_), .ZN(n3016) );
  NAND2_X1 U2921 ( .A1(n2963), .A2(n2962), .ZN(n3017) );
  OR2_X1 U2922 ( .A1(n2962), .A2(n2963), .ZN(n3015) );
  AND2_X1 U2923 ( .A1(n3018), .A2(n3019), .ZN(n2963) );
  NAND2_X1 U2924 ( .A1(n2960), .A2(n3020), .ZN(n3019) );
  OR2_X1 U2925 ( .A1(n2959), .A2(n2958), .ZN(n3020) );
  NOR2_X1 U2926 ( .A1(n2578), .A2(n2310), .ZN(n2960) );
  NAND2_X1 U2927 ( .A1(n2958), .A2(n2959), .ZN(n3018) );
  OR2_X1 U2928 ( .A1(n2954), .A2(n3021), .ZN(n2959) );
  AND2_X1 U2929 ( .A1(n2951), .A2(n3022), .ZN(n3021) );
  NAND2_X1 U2930 ( .A1(n3023), .A2(n3024), .ZN(n3022) );
  NAND2_X1 U2931 ( .A1(b_12_), .A2(a_10_), .ZN(n3024) );
  XOR2_X1 U2932 ( .A(n3025), .B(n3026), .Z(n2951) );
  XOR2_X1 U2933 ( .A(n3027), .B(n3028), .Z(n3025) );
  NOR2_X1 U2934 ( .A1(n2582), .A2(n3023), .ZN(n2954) );
  INV_X1 U2935 ( .A(n2956), .ZN(n3023) );
  NAND2_X1 U2936 ( .A1(n2926), .A2(n3029), .ZN(n2956) );
  NAND2_X1 U2937 ( .A1(n2925), .A2(n2927), .ZN(n3029) );
  NAND2_X1 U2938 ( .A1(n3030), .A2(n3031), .ZN(n2927) );
  NAND2_X1 U2939 ( .A1(b_12_), .A2(a_11_), .ZN(n3031) );
  INV_X1 U2940 ( .A(n3032), .ZN(n3030) );
  XNOR2_X1 U2941 ( .A(n3033), .B(n3034), .ZN(n2925) );
  XOR2_X1 U2942 ( .A(n3035), .B(n3036), .Z(n3033) );
  NAND2_X1 U2943 ( .A1(b_11_), .A2(a_12_), .ZN(n3035) );
  NAND2_X1 U2944 ( .A1(a_11_), .A2(n3032), .ZN(n2926) );
  NAND2_X1 U2945 ( .A1(n3037), .A2(n3038), .ZN(n3032) );
  NAND2_X1 U2946 ( .A1(n2933), .A2(n3039), .ZN(n3038) );
  NAND2_X1 U2947 ( .A1(n2934), .A2(n2233), .ZN(n3039) );
  INV_X1 U2948 ( .A(n3040), .ZN(n2934) );
  XOR2_X1 U2949 ( .A(n3041), .B(n3042), .Z(n2933) );
  XOR2_X1 U2950 ( .A(n3043), .B(n3044), .Z(n3041) );
  NAND2_X1 U2951 ( .A1(n3045), .A2(n3040), .ZN(n3037) );
  NAND2_X1 U2952 ( .A1(n3046), .A2(n3047), .ZN(n3040) );
  NAND2_X1 U2953 ( .A1(n2948), .A2(n3048), .ZN(n3047) );
  OR2_X1 U2954 ( .A1(n2949), .A2(n2950), .ZN(n3048) );
  NOR2_X1 U2955 ( .A1(n2578), .A2(n2188), .ZN(n2948) );
  NAND2_X1 U2956 ( .A1(n2950), .A2(n2949), .ZN(n3046) );
  NAND2_X1 U2957 ( .A1(n3049), .A2(n3050), .ZN(n2949) );
  NAND2_X1 U2958 ( .A1(b_10_), .A2(n3051), .ZN(n3050) );
  NAND2_X1 U2959 ( .A1(n2156), .A2(n3052), .ZN(n3051) );
  NAND2_X1 U2960 ( .A1(a_15_), .A2(n2580), .ZN(n3052) );
  NAND2_X1 U2961 ( .A1(b_11_), .A2(n3053), .ZN(n3049) );
  NAND2_X1 U2962 ( .A1(n2742), .A2(n3054), .ZN(n3053) );
  NAND2_X1 U2963 ( .A1(a_14_), .A2(n2285), .ZN(n3054) );
  AND3_X1 U2964 ( .A1(b_11_), .A2(b_12_), .A3(n2576), .ZN(n2950) );
  INV_X1 U2965 ( .A(n2233), .ZN(n3045) );
  NAND2_X1 U2966 ( .A1(b_12_), .A2(a_12_), .ZN(n2233) );
  XNOR2_X1 U2967 ( .A(n3055), .B(n3056), .ZN(n2958) );
  XOR2_X1 U2968 ( .A(n3057), .B(n3058), .Z(n3056) );
  NAND2_X1 U2969 ( .A1(b_11_), .A2(a_10_), .ZN(n3058) );
  XOR2_X1 U2970 ( .A(n3059), .B(n3060), .Z(n2962) );
  XNOR2_X1 U2971 ( .A(n3061), .B(n3062), .ZN(n3060) );
  XNOR2_X1 U2972 ( .A(n3063), .B(n3064), .ZN(n2908) );
  XNOR2_X1 U2973 ( .A(n3065), .B(n3066), .ZN(n3063) );
  NOR2_X1 U2974 ( .A1(n2584), .A2(n2580), .ZN(n3066) );
  XNOR2_X1 U2975 ( .A(n3067), .B(n3068), .ZN(n2965) );
  XNOR2_X1 U2976 ( .A(n3069), .B(n3070), .ZN(n3068) );
  XNOR2_X1 U2977 ( .A(n3071), .B(n3072), .ZN(n2970) );
  XOR2_X1 U2978 ( .A(n3073), .B(n3074), .Z(n3072) );
  NAND2_X1 U2979 ( .A1(b_11_), .A2(a_6_), .ZN(n3074) );
  XOR2_X1 U2980 ( .A(n3075), .B(n3076), .Z(n2894) );
  XNOR2_X1 U2981 ( .A(n3077), .B(n3078), .ZN(n3076) );
  XNOR2_X1 U2982 ( .A(n3079), .B(n3080), .ZN(n2977) );
  NAND2_X1 U2983 ( .A1(n3081), .A2(n3082), .ZN(n3079) );
  XNOR2_X1 U2984 ( .A(n3083), .B(n3084), .ZN(n2981) );
  NAND2_X1 U2985 ( .A1(n3085), .A2(n3086), .ZN(n3083) );
  XNOR2_X1 U2986 ( .A(n3087), .B(n3088), .ZN(n2877) );
  XOR2_X1 U2987 ( .A(n3089), .B(n3090), .Z(n3087) );
  NOR2_X1 U2988 ( .A1(n2516), .A2(n2580), .ZN(n3090) );
  NAND2_X1 U2989 ( .A1(n3091), .A2(n3092), .ZN(n2653) );
  XOR2_X1 U2990 ( .A(n3093), .B(n3094), .Z(n2654) );
  XNOR2_X1 U2991 ( .A(n3095), .B(n3096), .ZN(n3094) );
  NAND2_X1 U2992 ( .A1(n2985), .A2(n3097), .ZN(n2627) );
  XOR2_X1 U2993 ( .A(n2648), .B(n2649), .Z(n3097) );
  NOR2_X1 U2994 ( .A1(n3092), .A2(n3091), .ZN(n2985) );
  XNOR2_X1 U2995 ( .A(n3098), .B(n3099), .ZN(n3091) );
  XOR2_X1 U2996 ( .A(n3100), .B(n3101), .Z(n3098) );
  NOR2_X1 U2997 ( .A1(n3102), .A2(n2285), .ZN(n3101) );
  NAND2_X1 U2998 ( .A1(n3103), .A2(n3104), .ZN(n3092) );
  NAND2_X1 U2999 ( .A1(n3093), .A2(n3105), .ZN(n3104) );
  NAND2_X1 U3000 ( .A1(n3096), .A2(n3095), .ZN(n3105) );
  XOR2_X1 U3001 ( .A(n3106), .B(n3107), .Z(n3093) );
  XNOR2_X1 U3002 ( .A(n3108), .B(n3109), .ZN(n3107) );
  OR2_X1 U3003 ( .A1(n3095), .A2(n3096), .ZN(n3103) );
  NOR2_X1 U3004 ( .A1(n2580), .A2(n3102), .ZN(n3096) );
  NAND2_X1 U3005 ( .A1(n3110), .A2(n3111), .ZN(n3095) );
  NAND3_X1 U3006 ( .A1(a_1_), .A2(n3112), .A3(b_11_), .ZN(n3111) );
  OR2_X1 U3007 ( .A1(n3089), .A2(n3088), .ZN(n3112) );
  NAND2_X1 U3008 ( .A1(n3088), .A2(n3089), .ZN(n3110) );
  NAND2_X1 U3009 ( .A1(n3085), .A2(n3113), .ZN(n3089) );
  NAND2_X1 U3010 ( .A1(n3084), .A2(n3086), .ZN(n3113) );
  NAND2_X1 U3011 ( .A1(n3114), .A2(n3115), .ZN(n3086) );
  NAND2_X1 U3012 ( .A1(b_11_), .A2(a_2_), .ZN(n3115) );
  INV_X1 U3013 ( .A(n3116), .ZN(n3114) );
  XOR2_X1 U3014 ( .A(n3117), .B(n3118), .Z(n3084) );
  XOR2_X1 U3015 ( .A(n3119), .B(n3120), .Z(n3117) );
  NAND2_X1 U3016 ( .A1(a_2_), .A2(n3116), .ZN(n3085) );
  NAND2_X1 U3017 ( .A1(n3081), .A2(n3121), .ZN(n3116) );
  NAND2_X1 U3018 ( .A1(n3080), .A2(n3082), .ZN(n3121) );
  NAND2_X1 U3019 ( .A1(n3122), .A2(n3123), .ZN(n3082) );
  NAND2_X1 U3020 ( .A1(b_11_), .A2(a_3_), .ZN(n3123) );
  INV_X1 U3021 ( .A(n3124), .ZN(n3122) );
  XOR2_X1 U3022 ( .A(n3125), .B(n3126), .Z(n3080) );
  XOR2_X1 U3023 ( .A(n3127), .B(n3128), .Z(n3125) );
  NAND2_X1 U3024 ( .A1(a_3_), .A2(n3124), .ZN(n3081) );
  NAND2_X1 U3025 ( .A1(n3129), .A2(n3130), .ZN(n3124) );
  NAND3_X1 U3026 ( .A1(a_4_), .A2(n3131), .A3(b_11_), .ZN(n3130) );
  OR2_X1 U3027 ( .A1(n3001), .A2(n3000), .ZN(n3131) );
  NAND2_X1 U3028 ( .A1(n3000), .A2(n3001), .ZN(n3129) );
  NAND2_X1 U3029 ( .A1(n3132), .A2(n3133), .ZN(n3001) );
  NAND2_X1 U3030 ( .A1(n3078), .A2(n3134), .ZN(n3133) );
  OR2_X1 U3031 ( .A1(n3077), .A2(n3075), .ZN(n3134) );
  NOR2_X1 U3032 ( .A1(n2580), .A2(n2410), .ZN(n3078) );
  NAND2_X1 U3033 ( .A1(n3075), .A2(n3077), .ZN(n3132) );
  NAND2_X1 U3034 ( .A1(n3135), .A2(n3136), .ZN(n3077) );
  NAND3_X1 U3035 ( .A1(a_6_), .A2(n3137), .A3(b_11_), .ZN(n3136) );
  OR2_X1 U3036 ( .A1(n3073), .A2(n3071), .ZN(n3137) );
  NAND2_X1 U3037 ( .A1(n3071), .A2(n3073), .ZN(n3135) );
  NAND2_X1 U3038 ( .A1(n3138), .A2(n3139), .ZN(n3073) );
  NAND2_X1 U3039 ( .A1(n3070), .A2(n3140), .ZN(n3139) );
  OR2_X1 U3040 ( .A1(n3069), .A2(n3067), .ZN(n3140) );
  NOR2_X1 U3041 ( .A1(n2580), .A2(n2360), .ZN(n3070) );
  NAND2_X1 U3042 ( .A1(n3067), .A2(n3069), .ZN(n3138) );
  NAND2_X1 U3043 ( .A1(n3141), .A2(n3142), .ZN(n3069) );
  NAND3_X1 U3044 ( .A1(a_8_), .A2(n3143), .A3(b_11_), .ZN(n3142) );
  NAND2_X1 U3045 ( .A1(n3065), .A2(n3064), .ZN(n3143) );
  OR2_X1 U3046 ( .A1(n3064), .A2(n3065), .ZN(n3141) );
  AND2_X1 U3047 ( .A1(n3144), .A2(n3145), .ZN(n3065) );
  NAND2_X1 U3048 ( .A1(n3062), .A2(n3146), .ZN(n3145) );
  OR2_X1 U3049 ( .A1(n3061), .A2(n3059), .ZN(n3146) );
  NOR2_X1 U3050 ( .A1(n2580), .A2(n2310), .ZN(n3062) );
  NAND2_X1 U3051 ( .A1(n3059), .A2(n3061), .ZN(n3144) );
  NAND2_X1 U3052 ( .A1(n3147), .A2(n3148), .ZN(n3061) );
  NAND3_X1 U3053 ( .A1(a_10_), .A2(n3149), .A3(b_11_), .ZN(n3148) );
  OR2_X1 U3054 ( .A1(n3057), .A2(n3055), .ZN(n3149) );
  NAND2_X1 U3055 ( .A1(n3055), .A2(n3057), .ZN(n3147) );
  NAND2_X1 U3056 ( .A1(n3150), .A2(n3151), .ZN(n3057) );
  NAND2_X1 U3057 ( .A1(n3028), .A2(n3152), .ZN(n3151) );
  OR2_X1 U3058 ( .A1(n3027), .A2(n3026), .ZN(n3152) );
  INV_X1 U3059 ( .A(n2259), .ZN(n3028) );
  NAND2_X1 U3060 ( .A1(b_11_), .A2(a_11_), .ZN(n2259) );
  NAND2_X1 U3061 ( .A1(n3026), .A2(n3027), .ZN(n3150) );
  NAND2_X1 U3062 ( .A1(n3153), .A2(n3154), .ZN(n3027) );
  NAND3_X1 U3063 ( .A1(a_12_), .A2(n3155), .A3(b_11_), .ZN(n3154) );
  NAND2_X1 U3064 ( .A1(n3036), .A2(n3034), .ZN(n3155) );
  OR2_X1 U3065 ( .A1(n3034), .A2(n3036), .ZN(n3153) );
  AND2_X1 U3066 ( .A1(n3156), .A2(n3157), .ZN(n3036) );
  NAND2_X1 U3067 ( .A1(n3042), .A2(n3158), .ZN(n3157) );
  OR2_X1 U3068 ( .A1(n3043), .A2(n3044), .ZN(n3158) );
  NOR2_X1 U3069 ( .A1(n2580), .A2(n2188), .ZN(n3042) );
  NAND2_X1 U3070 ( .A1(n3044), .A2(n3043), .ZN(n3156) );
  NAND2_X1 U3071 ( .A1(n3159), .A2(n3160), .ZN(n3043) );
  NAND2_X1 U3072 ( .A1(b_10_), .A2(n3161), .ZN(n3160) );
  NAND2_X1 U3073 ( .A1(n2742), .A2(n3162), .ZN(n3161) );
  NAND2_X1 U3074 ( .A1(a_14_), .A2(n2583), .ZN(n3162) );
  NAND2_X1 U3075 ( .A1(b_9_), .A2(n3163), .ZN(n3159) );
  NAND2_X1 U3076 ( .A1(n2156), .A2(n3164), .ZN(n3163) );
  NAND2_X1 U3077 ( .A1(a_15_), .A2(n2285), .ZN(n3164) );
  AND3_X1 U3078 ( .A1(b_10_), .A2(b_11_), .A3(n2576), .ZN(n3044) );
  XNOR2_X1 U3079 ( .A(n3165), .B(n3166), .ZN(n3034) );
  XOR2_X1 U3080 ( .A(n3167), .B(n3168), .Z(n3165) );
  XNOR2_X1 U3081 ( .A(n3169), .B(n3170), .ZN(n3026) );
  XOR2_X1 U3082 ( .A(n3171), .B(n3172), .Z(n3169) );
  NAND2_X1 U3083 ( .A1(b_10_), .A2(a_12_), .ZN(n3171) );
  XOR2_X1 U3084 ( .A(n3173), .B(n3174), .Z(n3055) );
  XOR2_X1 U3085 ( .A(n3175), .B(n3176), .Z(n3173) );
  XNOR2_X1 U3086 ( .A(n3177), .B(n3178), .ZN(n3059) );
  XNOR2_X1 U3087 ( .A(n3179), .B(n2567), .ZN(n3178) );
  XNOR2_X1 U3088 ( .A(n3180), .B(n3181), .ZN(n3064) );
  XOR2_X1 U3089 ( .A(n3182), .B(n3183), .Z(n3180) );
  XNOR2_X1 U3090 ( .A(n3184), .B(n3185), .ZN(n3067) );
  XNOR2_X1 U3091 ( .A(n3186), .B(n3187), .ZN(n3184) );
  NOR2_X1 U3092 ( .A1(n2584), .A2(n2285), .ZN(n3187) );
  XOR2_X1 U3093 ( .A(n3188), .B(n3189), .Z(n3071) );
  XOR2_X1 U3094 ( .A(n3190), .B(n3191), .Z(n3188) );
  XNOR2_X1 U3095 ( .A(n3192), .B(n3193), .ZN(n3075) );
  XOR2_X1 U3096 ( .A(n3194), .B(n3195), .Z(n3193) );
  NAND2_X1 U3097 ( .A1(b_10_), .A2(a_6_), .ZN(n3195) );
  XNOR2_X1 U3098 ( .A(n3196), .B(n3197), .ZN(n3000) );
  XOR2_X1 U3099 ( .A(n3198), .B(n3199), .Z(n3197) );
  NAND2_X1 U3100 ( .A1(b_10_), .A2(a_5_), .ZN(n3199) );
  XOR2_X1 U3101 ( .A(n3200), .B(n3201), .Z(n3088) );
  XOR2_X1 U3102 ( .A(n3202), .B(n3203), .Z(n3200) );
  NAND2_X1 U3103 ( .A1(n3204), .A2(n3205), .ZN(n2102) );
  NAND2_X1 U3104 ( .A1(n2649), .A2(n2648), .ZN(n3205) );
  XNOR2_X1 U3105 ( .A(n3206), .B(n3207), .ZN(n3204) );
  NAND3_X1 U3106 ( .A1(n2649), .A2(n2648), .A3(n3208), .ZN(n2103) );
  XOR2_X1 U3107 ( .A(n3206), .B(n3207), .Z(n3208) );
  NAND2_X1 U3108 ( .A1(n3209), .A2(n3210), .ZN(n2648) );
  NAND3_X1 U3109 ( .A1(a_0_), .A2(n3211), .A3(b_10_), .ZN(n3210) );
  OR2_X1 U3110 ( .A1(n3099), .A2(n3100), .ZN(n3211) );
  NAND2_X1 U3111 ( .A1(n3099), .A2(n3100), .ZN(n3209) );
  NAND2_X1 U3112 ( .A1(n3212), .A2(n3213), .ZN(n3100) );
  NAND2_X1 U3113 ( .A1(n3109), .A2(n3214), .ZN(n3213) );
  OR2_X1 U3114 ( .A1(n3106), .A2(n3108), .ZN(n3214) );
  NOR2_X1 U3115 ( .A1(n2285), .A2(n2516), .ZN(n3109) );
  NAND2_X1 U3116 ( .A1(n3106), .A2(n3108), .ZN(n3212) );
  NAND2_X1 U3117 ( .A1(n3215), .A2(n3216), .ZN(n3108) );
  NAND2_X1 U3118 ( .A1(n3203), .A2(n3217), .ZN(n3216) );
  OR2_X1 U3119 ( .A1(n3202), .A2(n3201), .ZN(n3217) );
  NOR2_X1 U3120 ( .A1(n2285), .A2(n2491), .ZN(n3203) );
  NAND2_X1 U3121 ( .A1(n3201), .A2(n3202), .ZN(n3215) );
  NAND2_X1 U3122 ( .A1(n3218), .A2(n3219), .ZN(n3202) );
  NAND2_X1 U3123 ( .A1(n3120), .A2(n3220), .ZN(n3219) );
  OR2_X1 U3124 ( .A1(n3118), .A2(n3119), .ZN(n3220) );
  NOR2_X1 U3125 ( .A1(n2285), .A2(n2466), .ZN(n3120) );
  NAND2_X1 U3126 ( .A1(n3118), .A2(n3119), .ZN(n3218) );
  NAND2_X1 U3127 ( .A1(n3221), .A2(n3222), .ZN(n3119) );
  NAND2_X1 U3128 ( .A1(n3128), .A2(n3223), .ZN(n3222) );
  OR2_X1 U3129 ( .A1(n3126), .A2(n3127), .ZN(n3223) );
  NOR2_X1 U3130 ( .A1(n2285), .A2(n2435), .ZN(n3128) );
  NAND2_X1 U3131 ( .A1(n3126), .A2(n3127), .ZN(n3221) );
  NAND2_X1 U3132 ( .A1(n3224), .A2(n3225), .ZN(n3127) );
  NAND3_X1 U3133 ( .A1(a_5_), .A2(n3226), .A3(b_10_), .ZN(n3225) );
  OR2_X1 U3134 ( .A1(n3198), .A2(n3196), .ZN(n3226) );
  NAND2_X1 U3135 ( .A1(n3196), .A2(n3198), .ZN(n3224) );
  NAND2_X1 U3136 ( .A1(n3227), .A2(n3228), .ZN(n3198) );
  NAND3_X1 U3137 ( .A1(a_6_), .A2(n3229), .A3(b_10_), .ZN(n3228) );
  OR2_X1 U3138 ( .A1(n3194), .A2(n3192), .ZN(n3229) );
  NAND2_X1 U3139 ( .A1(n3192), .A2(n3194), .ZN(n3227) );
  NAND2_X1 U3140 ( .A1(n3230), .A2(n3231), .ZN(n3194) );
  NAND2_X1 U3141 ( .A1(n3191), .A2(n3232), .ZN(n3231) );
  OR2_X1 U3142 ( .A1(n3189), .A2(n3190), .ZN(n3232) );
  NOR2_X1 U3143 ( .A1(n2285), .A2(n2360), .ZN(n3191) );
  NAND2_X1 U3144 ( .A1(n3189), .A2(n3190), .ZN(n3230) );
  NAND2_X1 U3145 ( .A1(n3233), .A2(n3234), .ZN(n3190) );
  NAND3_X1 U3146 ( .A1(a_8_), .A2(n3235), .A3(b_10_), .ZN(n3234) );
  NAND2_X1 U3147 ( .A1(n3186), .A2(n3185), .ZN(n3235) );
  OR2_X1 U3148 ( .A1(n3185), .A2(n3186), .ZN(n3233) );
  AND2_X1 U3149 ( .A1(n3236), .A2(n3237), .ZN(n3186) );
  NAND2_X1 U3150 ( .A1(n3183), .A2(n3238), .ZN(n3237) );
  OR2_X1 U3151 ( .A1(n3181), .A2(n3182), .ZN(n3238) );
  NOR2_X1 U3152 ( .A1(n2285), .A2(n2310), .ZN(n3183) );
  NAND2_X1 U3153 ( .A1(n3181), .A2(n3182), .ZN(n3236) );
  NAND2_X1 U3154 ( .A1(n3239), .A2(n3240), .ZN(n3182) );
  NAND2_X1 U3155 ( .A1(n3177), .A2(n3241), .ZN(n3240) );
  OR2_X1 U3156 ( .A1(n3179), .A2(n2567), .ZN(n3241) );
  XOR2_X1 U3157 ( .A(n3242), .B(n3243), .Z(n3177) );
  XOR2_X1 U3158 ( .A(n3244), .B(n3245), .Z(n3242) );
  NAND2_X1 U3159 ( .A1(n2567), .A2(n3179), .ZN(n3239) );
  NAND2_X1 U3160 ( .A1(n3246), .A2(n3247), .ZN(n3179) );
  NAND2_X1 U3161 ( .A1(n3176), .A2(n3248), .ZN(n3247) );
  OR2_X1 U3162 ( .A1(n3174), .A2(n3175), .ZN(n3248) );
  NOR2_X1 U3163 ( .A1(n2285), .A2(n2581), .ZN(n3176) );
  NAND2_X1 U3164 ( .A1(n3174), .A2(n3175), .ZN(n3246) );
  NAND2_X1 U3165 ( .A1(n3249), .A2(n3250), .ZN(n3175) );
  NAND3_X1 U3166 ( .A1(a_12_), .A2(n3251), .A3(b_10_), .ZN(n3250) );
  NAND2_X1 U3167 ( .A1(n3172), .A2(n3170), .ZN(n3251) );
  OR2_X1 U3168 ( .A1(n3170), .A2(n3172), .ZN(n3249) );
  AND2_X1 U3169 ( .A1(n3252), .A2(n3253), .ZN(n3172) );
  NAND2_X1 U3170 ( .A1(n3166), .A2(n3254), .ZN(n3253) );
  OR2_X1 U3171 ( .A1(n3167), .A2(n3168), .ZN(n3254) );
  NOR2_X1 U3172 ( .A1(n2285), .A2(n2188), .ZN(n3166) );
  NAND2_X1 U3173 ( .A1(n3168), .A2(n3167), .ZN(n3252) );
  NAND2_X1 U3174 ( .A1(n3255), .A2(n3256), .ZN(n3167) );
  NAND2_X1 U3175 ( .A1(b_8_), .A2(n3257), .ZN(n3256) );
  NAND2_X1 U3176 ( .A1(n2156), .A2(n3258), .ZN(n3257) );
  NAND2_X1 U3177 ( .A1(a_15_), .A2(n2583), .ZN(n3258) );
  NAND2_X1 U3178 ( .A1(b_9_), .A2(n3259), .ZN(n3255) );
  NAND2_X1 U3179 ( .A1(n2742), .A2(n3260), .ZN(n3259) );
  NAND2_X1 U3180 ( .A1(a_14_), .A2(n2335), .ZN(n3260) );
  AND3_X1 U3181 ( .A1(b_9_), .A2(b_10_), .A3(n2576), .ZN(n3168) );
  XNOR2_X1 U3182 ( .A(n3261), .B(n3262), .ZN(n3170) );
  XOR2_X1 U3183 ( .A(n3263), .B(n3264), .Z(n3261) );
  XNOR2_X1 U3184 ( .A(n3265), .B(n3266), .ZN(n3174) );
  XOR2_X1 U3185 ( .A(n3267), .B(n3268), .Z(n3265) );
  NAND2_X1 U3186 ( .A1(b_9_), .A2(a_12_), .ZN(n3267) );
  NOR2_X1 U3187 ( .A1(n2285), .A2(n2582), .ZN(n2567) );
  XNOR2_X1 U3188 ( .A(n3269), .B(n3270), .ZN(n3181) );
  XOR2_X1 U3189 ( .A(n3271), .B(n3272), .Z(n3270) );
  NAND2_X1 U3190 ( .A1(b_9_), .A2(a_10_), .ZN(n3272) );
  XOR2_X1 U3191 ( .A(n3273), .B(n3274), .Z(n3185) );
  XNOR2_X1 U3192 ( .A(n3275), .B(n2564), .ZN(n3274) );
  XNOR2_X1 U3193 ( .A(n3276), .B(n3277), .ZN(n3189) );
  XNOR2_X1 U3194 ( .A(n3278), .B(n3279), .ZN(n3276) );
  NOR2_X1 U3195 ( .A1(n2584), .A2(n2583), .ZN(n3279) );
  XOR2_X1 U3196 ( .A(n3280), .B(n3281), .Z(n3192) );
  XOR2_X1 U3197 ( .A(n3282), .B(n3283), .Z(n3280) );
  XNOR2_X1 U3198 ( .A(n3284), .B(n3285), .ZN(n3196) );
  XNOR2_X1 U3199 ( .A(n3286), .B(n3287), .ZN(n3285) );
  XNOR2_X1 U3200 ( .A(n3288), .B(n3289), .ZN(n3126) );
  XOR2_X1 U3201 ( .A(n3290), .B(n3291), .Z(n3288) );
  NAND2_X1 U3202 ( .A1(b_9_), .A2(a_5_), .ZN(n3290) );
  XOR2_X1 U3203 ( .A(n3292), .B(n3293), .Z(n3118) );
  XNOR2_X1 U3204 ( .A(n3294), .B(n3295), .ZN(n3293) );
  NAND2_X1 U3205 ( .A1(b_9_), .A2(a_4_), .ZN(n3295) );
  XOR2_X1 U3206 ( .A(n3296), .B(n3297), .Z(n3201) );
  XOR2_X1 U3207 ( .A(n3298), .B(n3299), .Z(n3296) );
  NOR2_X1 U3208 ( .A1(n2466), .A2(n2583), .ZN(n3299) );
  XOR2_X1 U3209 ( .A(n3300), .B(n3301), .Z(n3106) );
  XOR2_X1 U3210 ( .A(n3302), .B(n3303), .Z(n3300) );
  NOR2_X1 U3211 ( .A1(n2491), .A2(n2583), .ZN(n3303) );
  XOR2_X1 U3212 ( .A(n3304), .B(n3305), .Z(n3099) );
  XNOR2_X1 U3213 ( .A(n3306), .B(n3307), .ZN(n3305) );
  NAND2_X1 U3214 ( .A1(b_9_), .A2(a_1_), .ZN(n3307) );
  XNOR2_X1 U3215 ( .A(n3308), .B(n3309), .ZN(n2649) );
  XOR2_X1 U3216 ( .A(n3310), .B(n3311), .Z(n3309) );
  NAND2_X1 U3217 ( .A1(b_9_), .A2(a_0_), .ZN(n3311) );
  NAND2_X1 U3218 ( .A1(n3312), .A2(n3313), .ZN(n2108) );
  NAND2_X1 U3219 ( .A1(n3207), .A2(n3206), .ZN(n3313) );
  XNOR2_X1 U3220 ( .A(n3314), .B(n3315), .ZN(n3312) );
  NAND3_X1 U3221 ( .A1(n3207), .A2(n3206), .A3(n3316), .ZN(n2109) );
  XOR2_X1 U3222 ( .A(n3315), .B(n3314), .Z(n3316) );
  NAND2_X1 U3223 ( .A1(n3317), .A2(n3318), .ZN(n3206) );
  NAND3_X1 U3224 ( .A1(a_0_), .A2(n3319), .A3(b_9_), .ZN(n3318) );
  OR2_X1 U3225 ( .A1(n3308), .A2(n3310), .ZN(n3319) );
  NAND2_X1 U3226 ( .A1(n3308), .A2(n3310), .ZN(n3317) );
  NAND2_X1 U3227 ( .A1(n3320), .A2(n3321), .ZN(n3310) );
  NAND3_X1 U3228 ( .A1(a_1_), .A2(n3322), .A3(b_9_), .ZN(n3321) );
  NAND2_X1 U3229 ( .A1(n3306), .A2(n3304), .ZN(n3322) );
  OR2_X1 U3230 ( .A1(n3304), .A2(n3306), .ZN(n3320) );
  AND2_X1 U3231 ( .A1(n3323), .A2(n3324), .ZN(n3306) );
  NAND3_X1 U3232 ( .A1(a_2_), .A2(n3325), .A3(b_9_), .ZN(n3324) );
  OR2_X1 U3233 ( .A1(n3302), .A2(n3301), .ZN(n3325) );
  NAND2_X1 U3234 ( .A1(n3301), .A2(n3302), .ZN(n3323) );
  NAND2_X1 U3235 ( .A1(n3326), .A2(n3327), .ZN(n3302) );
  NAND3_X1 U3236 ( .A1(a_3_), .A2(n3328), .A3(b_9_), .ZN(n3327) );
  OR2_X1 U3237 ( .A1(n3297), .A2(n3298), .ZN(n3328) );
  NAND2_X1 U3238 ( .A1(n3297), .A2(n3298), .ZN(n3326) );
  NAND2_X1 U3239 ( .A1(n3329), .A2(n3330), .ZN(n3298) );
  NAND3_X1 U3240 ( .A1(a_4_), .A2(n3331), .A3(b_9_), .ZN(n3330) );
  NAND2_X1 U3241 ( .A1(n3294), .A2(n3292), .ZN(n3331) );
  OR2_X1 U3242 ( .A1(n3292), .A2(n3294), .ZN(n3329) );
  AND2_X1 U3243 ( .A1(n3332), .A2(n3333), .ZN(n3294) );
  NAND3_X1 U3244 ( .A1(a_5_), .A2(n3334), .A3(b_9_), .ZN(n3333) );
  NAND2_X1 U3245 ( .A1(n3291), .A2(n3289), .ZN(n3334) );
  OR2_X1 U3246 ( .A1(n3289), .A2(n3291), .ZN(n3332) );
  AND2_X1 U3247 ( .A1(n3335), .A2(n3336), .ZN(n3291) );
  NAND2_X1 U3248 ( .A1(n3287), .A2(n3337), .ZN(n3336) );
  OR2_X1 U3249 ( .A1(n3284), .A2(n3286), .ZN(n3337) );
  NOR2_X1 U3250 ( .A1(n2583), .A2(n2586), .ZN(n3287) );
  NAND2_X1 U3251 ( .A1(n3284), .A2(n3286), .ZN(n3335) );
  NAND2_X1 U3252 ( .A1(n3338), .A2(n3339), .ZN(n3286) );
  NAND2_X1 U3253 ( .A1(n3283), .A2(n3340), .ZN(n3339) );
  OR2_X1 U3254 ( .A1(n3281), .A2(n3282), .ZN(n3340) );
  NOR2_X1 U3255 ( .A1(n2583), .A2(n2360), .ZN(n3283) );
  NAND2_X1 U3256 ( .A1(n3281), .A2(n3282), .ZN(n3338) );
  NAND2_X1 U3257 ( .A1(n3341), .A2(n3342), .ZN(n3282) );
  NAND3_X1 U3258 ( .A1(a_8_), .A2(n3343), .A3(b_9_), .ZN(n3342) );
  NAND2_X1 U3259 ( .A1(n3278), .A2(n3277), .ZN(n3343) );
  OR2_X1 U3260 ( .A1(n3277), .A2(n3278), .ZN(n3341) );
  AND2_X1 U3261 ( .A1(n3344), .A2(n3345), .ZN(n3278) );
  NAND2_X1 U3262 ( .A1(n2564), .A2(n3346), .ZN(n3345) );
  OR2_X1 U3263 ( .A1(n3273), .A2(n3275), .ZN(n3346) );
  NOR2_X1 U3264 ( .A1(n2583), .A2(n2310), .ZN(n2564) );
  NAND2_X1 U3265 ( .A1(n3273), .A2(n3275), .ZN(n3344) );
  NAND2_X1 U3266 ( .A1(n3347), .A2(n3348), .ZN(n3275) );
  NAND3_X1 U3267 ( .A1(a_10_), .A2(n3349), .A3(b_9_), .ZN(n3348) );
  OR2_X1 U3268 ( .A1(n3271), .A2(n3269), .ZN(n3349) );
  NAND2_X1 U3269 ( .A1(n3269), .A2(n3271), .ZN(n3347) );
  NAND2_X1 U3270 ( .A1(n3350), .A2(n3351), .ZN(n3271) );
  NAND2_X1 U3271 ( .A1(n3245), .A2(n3352), .ZN(n3351) );
  OR2_X1 U3272 ( .A1(n3243), .A2(n3244), .ZN(n3352) );
  NOR2_X1 U3273 ( .A1(n2583), .A2(n2581), .ZN(n3245) );
  NAND2_X1 U3274 ( .A1(n3243), .A2(n3244), .ZN(n3350) );
  NAND2_X1 U3275 ( .A1(n3353), .A2(n3354), .ZN(n3244) );
  NAND3_X1 U3276 ( .A1(a_12_), .A2(n3355), .A3(b_9_), .ZN(n3354) );
  NAND2_X1 U3277 ( .A1(n3268), .A2(n3266), .ZN(n3355) );
  OR2_X1 U3278 ( .A1(n3266), .A2(n3268), .ZN(n3353) );
  AND2_X1 U3279 ( .A1(n3356), .A2(n3357), .ZN(n3268) );
  NAND2_X1 U3280 ( .A1(n3262), .A2(n3358), .ZN(n3357) );
  OR2_X1 U3281 ( .A1(n3263), .A2(n3264), .ZN(n3358) );
  NOR2_X1 U3282 ( .A1(n2583), .A2(n2188), .ZN(n3262) );
  NAND2_X1 U3283 ( .A1(n3264), .A2(n3263), .ZN(n3356) );
  NAND2_X1 U3284 ( .A1(n3359), .A2(n3360), .ZN(n3263) );
  NAND2_X1 U3285 ( .A1(b_7_), .A2(n3361), .ZN(n3360) );
  NAND2_X1 U3286 ( .A1(n2156), .A2(n3362), .ZN(n3361) );
  NAND2_X1 U3287 ( .A1(a_15_), .A2(n2335), .ZN(n3362) );
  NAND2_X1 U3288 ( .A1(b_8_), .A2(n3363), .ZN(n3359) );
  NAND2_X1 U3289 ( .A1(n2742), .A2(n3364), .ZN(n3363) );
  NAND2_X1 U3290 ( .A1(a_14_), .A2(n2585), .ZN(n3364) );
  AND3_X1 U3291 ( .A1(b_8_), .A2(b_9_), .A3(n2576), .ZN(n3264) );
  XNOR2_X1 U3292 ( .A(n3365), .B(n3366), .ZN(n3266) );
  XOR2_X1 U3293 ( .A(n3367), .B(n3368), .Z(n3365) );
  XNOR2_X1 U3294 ( .A(n3369), .B(n3370), .ZN(n3243) );
  XOR2_X1 U3295 ( .A(n3371), .B(n3372), .Z(n3369) );
  NAND2_X1 U3296 ( .A1(b_8_), .A2(a_12_), .ZN(n3371) );
  XOR2_X1 U3297 ( .A(n3373), .B(n3374), .Z(n3269) );
  XOR2_X1 U3298 ( .A(n3375), .B(n3376), .Z(n3373) );
  XNOR2_X1 U3299 ( .A(n3377), .B(n3378), .ZN(n3273) );
  XOR2_X1 U3300 ( .A(n3379), .B(n3380), .Z(n3378) );
  NAND2_X1 U3301 ( .A1(b_8_), .A2(a_10_), .ZN(n3380) );
  XOR2_X1 U3302 ( .A(n3381), .B(n3382), .Z(n3277) );
  XNOR2_X1 U3303 ( .A(n3383), .B(n3384), .ZN(n3382) );
  XOR2_X1 U3304 ( .A(n3385), .B(n3386), .Z(n3281) );
  XOR2_X1 U3305 ( .A(n3387), .B(n3388), .Z(n3385) );
  XNOR2_X1 U3306 ( .A(n3389), .B(n3390), .ZN(n3284) );
  NAND2_X1 U3307 ( .A1(n3391), .A2(n3392), .ZN(n3389) );
  XOR2_X1 U3308 ( .A(n3393), .B(n3394), .Z(n3289) );
  XNOR2_X1 U3309 ( .A(n3395), .B(n3396), .ZN(n3394) );
  XOR2_X1 U3310 ( .A(n3397), .B(n3398), .Z(n3292) );
  XNOR2_X1 U3311 ( .A(n3399), .B(n3400), .ZN(n3398) );
  XOR2_X1 U3312 ( .A(n3401), .B(n3402), .Z(n3297) );
  XOR2_X1 U3313 ( .A(n3403), .B(n3404), .Z(n3401) );
  XNOR2_X1 U3314 ( .A(n3405), .B(n3406), .ZN(n3301) );
  XOR2_X1 U3315 ( .A(n3407), .B(n3408), .Z(n3406) );
  NAND2_X1 U3316 ( .A1(b_8_), .A2(a_3_), .ZN(n3408) );
  XNOR2_X1 U3317 ( .A(n3409), .B(n3410), .ZN(n3304) );
  XOR2_X1 U3318 ( .A(n3411), .B(n3412), .Z(n3409) );
  XNOR2_X1 U3319 ( .A(n3413), .B(n3414), .ZN(n3308) );
  NAND2_X1 U3320 ( .A1(n3415), .A2(n3416), .ZN(n3413) );
  XNOR2_X1 U3321 ( .A(n3417), .B(n3418), .ZN(n3207) );
  NAND2_X1 U3322 ( .A1(n3419), .A2(n3420), .ZN(n3417) );
  NAND2_X1 U3323 ( .A1(n3421), .A2(n3422), .ZN(n2114) );
  NAND2_X1 U3324 ( .A1(n3314), .A2(n3315), .ZN(n3422) );
  XOR2_X1 U3325 ( .A(n3423), .B(n3424), .Z(n3421) );
  INV_X1 U3326 ( .A(n3425), .ZN(n3424) );
  NAND3_X1 U3327 ( .A1(n3426), .A2(n3315), .A3(n3314), .ZN(n2115) );
  XOR2_X1 U3328 ( .A(n3427), .B(n3428), .Z(n3314) );
  XOR2_X1 U3329 ( .A(n3429), .B(n3430), .Z(n3427) );
  NOR2_X1 U3330 ( .A1(n3102), .A2(n2585), .ZN(n3430) );
  NAND2_X1 U3331 ( .A1(n3419), .A2(n3431), .ZN(n3315) );
  NAND2_X1 U3332 ( .A1(n3418), .A2(n3420), .ZN(n3431) );
  NAND2_X1 U3333 ( .A1(n3432), .A2(n3433), .ZN(n3420) );
  NAND2_X1 U3334 ( .A1(b_8_), .A2(a_0_), .ZN(n3433) );
  INV_X1 U3335 ( .A(n3434), .ZN(n3432) );
  XNOR2_X1 U3336 ( .A(n3435), .B(n3436), .ZN(n3418) );
  XOR2_X1 U3337 ( .A(n3437), .B(n3438), .Z(n3435) );
  NAND2_X1 U3338 ( .A1(b_7_), .A2(a_1_), .ZN(n3437) );
  NAND2_X1 U3339 ( .A1(a_0_), .A2(n3434), .ZN(n3419) );
  NAND2_X1 U3340 ( .A1(n3415), .A2(n3439), .ZN(n3434) );
  NAND2_X1 U3341 ( .A1(n3414), .A2(n3416), .ZN(n3439) );
  NAND2_X1 U3342 ( .A1(n3440), .A2(n3441), .ZN(n3416) );
  NAND2_X1 U3343 ( .A1(b_8_), .A2(a_1_), .ZN(n3441) );
  INV_X1 U3344 ( .A(n3442), .ZN(n3440) );
  XNOR2_X1 U3345 ( .A(n3443), .B(n3444), .ZN(n3414) );
  XNOR2_X1 U3346 ( .A(n3445), .B(n3446), .ZN(n3443) );
  NAND2_X1 U3347 ( .A1(a_1_), .A2(n3442), .ZN(n3415) );
  NAND2_X1 U3348 ( .A1(n3447), .A2(n3448), .ZN(n3442) );
  NAND2_X1 U3349 ( .A1(n3412), .A2(n3449), .ZN(n3448) );
  OR2_X1 U3350 ( .A1(n3410), .A2(n3411), .ZN(n3449) );
  NOR2_X1 U3351 ( .A1(n2335), .A2(n2491), .ZN(n3412) );
  NAND2_X1 U3352 ( .A1(n3410), .A2(n3411), .ZN(n3447) );
  NAND2_X1 U3353 ( .A1(n3450), .A2(n3451), .ZN(n3411) );
  NAND3_X1 U3354 ( .A1(a_3_), .A2(n3452), .A3(b_8_), .ZN(n3451) );
  OR2_X1 U3355 ( .A1(n3405), .A2(n3407), .ZN(n3452) );
  NAND2_X1 U3356 ( .A1(n3405), .A2(n3407), .ZN(n3450) );
  NAND2_X1 U3357 ( .A1(n3453), .A2(n3454), .ZN(n3407) );
  NAND2_X1 U3358 ( .A1(n3403), .A2(n3455), .ZN(n3454) );
  OR2_X1 U3359 ( .A1(n3404), .A2(n3402), .ZN(n3455) );
  NOR2_X1 U3360 ( .A1(n2335), .A2(n2435), .ZN(n3403) );
  NAND2_X1 U3361 ( .A1(n3402), .A2(n3404), .ZN(n3453) );
  NAND2_X1 U3362 ( .A1(n3456), .A2(n3457), .ZN(n3404) );
  NAND2_X1 U3363 ( .A1(n3400), .A2(n3458), .ZN(n3457) );
  OR2_X1 U3364 ( .A1(n3397), .A2(n3399), .ZN(n3458) );
  NOR2_X1 U3365 ( .A1(n2335), .A2(n2410), .ZN(n3400) );
  NAND2_X1 U3366 ( .A1(n3397), .A2(n3399), .ZN(n3456) );
  NAND2_X1 U3367 ( .A1(n3459), .A2(n3460), .ZN(n3399) );
  NAND2_X1 U3368 ( .A1(n3396), .A2(n3461), .ZN(n3460) );
  OR2_X1 U3369 ( .A1(n3393), .A2(n3395), .ZN(n3461) );
  NOR2_X1 U3370 ( .A1(n2335), .A2(n2586), .ZN(n3396) );
  NAND2_X1 U3371 ( .A1(n3393), .A2(n3395), .ZN(n3459) );
  NAND2_X1 U3372 ( .A1(n3391), .A2(n3462), .ZN(n3395) );
  NAND2_X1 U3373 ( .A1(n3390), .A2(n3392), .ZN(n3462) );
  NAND2_X1 U3374 ( .A1(n3463), .A2(n3464), .ZN(n3392) );
  NAND2_X1 U3375 ( .A1(b_8_), .A2(a_7_), .ZN(n3464) );
  INV_X1 U3376 ( .A(n3465), .ZN(n3463) );
  XNOR2_X1 U3377 ( .A(n3466), .B(n3467), .ZN(n3390) );
  XNOR2_X1 U3378 ( .A(n3468), .B(n3469), .ZN(n3466) );
  NOR2_X1 U3379 ( .A1(n2584), .A2(n2585), .ZN(n3469) );
  NAND2_X1 U3380 ( .A1(a_7_), .A2(n3465), .ZN(n3391) );
  NAND2_X1 U3381 ( .A1(n3470), .A2(n3471), .ZN(n3465) );
  NAND2_X1 U3382 ( .A1(n3386), .A2(n3472), .ZN(n3471) );
  OR2_X1 U3383 ( .A1(n3387), .A2(n3388), .ZN(n3472) );
  XNOR2_X1 U3384 ( .A(n3473), .B(n3474), .ZN(n3386) );
  XNOR2_X1 U3385 ( .A(n3475), .B(n3476), .ZN(n3474) );
  NAND2_X1 U3386 ( .A1(n3388), .A2(n3387), .ZN(n3470) );
  NAND2_X1 U3387 ( .A1(n3477), .A2(n3478), .ZN(n3387) );
  NAND2_X1 U3388 ( .A1(n3384), .A2(n3479), .ZN(n3478) );
  OR2_X1 U3389 ( .A1(n3381), .A2(n3383), .ZN(n3479) );
  NOR2_X1 U3390 ( .A1(n2335), .A2(n2310), .ZN(n3384) );
  NAND2_X1 U3391 ( .A1(n3381), .A2(n3383), .ZN(n3477) );
  NAND2_X1 U3392 ( .A1(n3480), .A2(n3481), .ZN(n3383) );
  NAND3_X1 U3393 ( .A1(a_10_), .A2(n3482), .A3(b_8_), .ZN(n3481) );
  OR2_X1 U3394 ( .A1(n3379), .A2(n3377), .ZN(n3482) );
  NAND2_X1 U3395 ( .A1(n3377), .A2(n3379), .ZN(n3480) );
  NAND2_X1 U3396 ( .A1(n3483), .A2(n3484), .ZN(n3379) );
  NAND2_X1 U3397 ( .A1(n3376), .A2(n3485), .ZN(n3484) );
  OR2_X1 U3398 ( .A1(n3374), .A2(n3375), .ZN(n3485) );
  NOR2_X1 U3399 ( .A1(n2335), .A2(n2581), .ZN(n3376) );
  NAND2_X1 U3400 ( .A1(n3374), .A2(n3375), .ZN(n3483) );
  NAND2_X1 U3401 ( .A1(n3486), .A2(n3487), .ZN(n3375) );
  NAND3_X1 U3402 ( .A1(a_12_), .A2(n3488), .A3(b_8_), .ZN(n3487) );
  NAND2_X1 U3403 ( .A1(n3372), .A2(n3370), .ZN(n3488) );
  OR2_X1 U3404 ( .A1(n3370), .A2(n3372), .ZN(n3486) );
  AND2_X1 U3405 ( .A1(n3489), .A2(n3490), .ZN(n3372) );
  NAND2_X1 U3406 ( .A1(n3366), .A2(n3491), .ZN(n3490) );
  OR2_X1 U3407 ( .A1(n3367), .A2(n3368), .ZN(n3491) );
  NOR2_X1 U3408 ( .A1(n2335), .A2(n2188), .ZN(n3366) );
  NAND2_X1 U3409 ( .A1(n3368), .A2(n3367), .ZN(n3489) );
  NAND2_X1 U3410 ( .A1(n3492), .A2(n3493), .ZN(n3367) );
  NAND2_X1 U3411 ( .A1(b_6_), .A2(n3494), .ZN(n3493) );
  NAND2_X1 U3412 ( .A1(n2156), .A2(n3495), .ZN(n3494) );
  NAND2_X1 U3413 ( .A1(a_15_), .A2(n2585), .ZN(n3495) );
  NAND2_X1 U3414 ( .A1(b_7_), .A2(n3496), .ZN(n3492) );
  NAND2_X1 U3415 ( .A1(n2742), .A2(n3497), .ZN(n3496) );
  NAND2_X1 U3416 ( .A1(a_14_), .A2(n2385), .ZN(n3497) );
  AND3_X1 U3417 ( .A1(b_7_), .A2(b_8_), .A3(n2576), .ZN(n3368) );
  XNOR2_X1 U3418 ( .A(n3498), .B(n3499), .ZN(n3370) );
  XOR2_X1 U3419 ( .A(n3500), .B(n3501), .Z(n3498) );
  XNOR2_X1 U3420 ( .A(n3502), .B(n3503), .ZN(n3374) );
  XOR2_X1 U3421 ( .A(n3504), .B(n3505), .Z(n3502) );
  NAND2_X1 U3422 ( .A1(b_7_), .A2(a_12_), .ZN(n3504) );
  XOR2_X1 U3423 ( .A(n3506), .B(n3507), .Z(n3377) );
  XOR2_X1 U3424 ( .A(n3508), .B(n3509), .Z(n3506) );
  XNOR2_X1 U3425 ( .A(n3510), .B(n3511), .ZN(n3381) );
  XOR2_X1 U3426 ( .A(n3512), .B(n3513), .Z(n3511) );
  NAND2_X1 U3427 ( .A1(b_7_), .A2(a_10_), .ZN(n3513) );
  INV_X1 U3428 ( .A(n2561), .ZN(n3388) );
  NAND2_X1 U3429 ( .A1(b_8_), .A2(a_8_), .ZN(n2561) );
  XOR2_X1 U3430 ( .A(n3514), .B(n3515), .Z(n3393) );
  XOR2_X1 U3431 ( .A(n3516), .B(n3517), .Z(n3514) );
  XNOR2_X1 U3432 ( .A(n3518), .B(n3519), .ZN(n3397) );
  NAND2_X1 U3433 ( .A1(n3520), .A2(n3521), .ZN(n3518) );
  XOR2_X1 U3434 ( .A(n3522), .B(n3523), .Z(n3402) );
  XOR2_X1 U3435 ( .A(n3524), .B(n3525), .Z(n3522) );
  NOR2_X1 U3436 ( .A1(n2410), .A2(n2585), .ZN(n3525) );
  XOR2_X1 U3437 ( .A(n3526), .B(n3527), .Z(n3405) );
  XNOR2_X1 U3438 ( .A(n3528), .B(n3529), .ZN(n3527) );
  NAND2_X1 U3439 ( .A1(b_7_), .A2(a_4_), .ZN(n3529) );
  XOR2_X1 U3440 ( .A(n3530), .B(n3531), .Z(n3410) );
  XOR2_X1 U3441 ( .A(n3532), .B(n3533), .Z(n3530) );
  NOR2_X1 U3442 ( .A1(n2466), .A2(n2585), .ZN(n3533) );
  XOR2_X1 U3443 ( .A(n3423), .B(n3425), .Z(n3426) );
  NAND2_X1 U3444 ( .A1(n3534), .A2(n3535), .ZN(n2120) );
  NAND2_X1 U3445 ( .A1(n3425), .A2(n3423), .ZN(n3535) );
  XNOR2_X1 U3446 ( .A(n3536), .B(n3537), .ZN(n3534) );
  NAND3_X1 U3447 ( .A1(n3425), .A2(n3423), .A3(n3538), .ZN(n2121) );
  XOR2_X1 U3448 ( .A(n3536), .B(n3537), .Z(n3538) );
  NAND2_X1 U3449 ( .A1(n3539), .A2(n3540), .ZN(n3423) );
  NAND3_X1 U3450 ( .A1(a_0_), .A2(n3541), .A3(b_7_), .ZN(n3540) );
  OR2_X1 U3451 ( .A1(n3428), .A2(n3429), .ZN(n3541) );
  NAND2_X1 U3452 ( .A1(n3428), .A2(n3429), .ZN(n3539) );
  NAND2_X1 U3453 ( .A1(n3542), .A2(n3543), .ZN(n3429) );
  NAND3_X1 U3454 ( .A1(a_1_), .A2(n3544), .A3(b_7_), .ZN(n3543) );
  NAND2_X1 U3455 ( .A1(n3438), .A2(n3436), .ZN(n3544) );
  OR2_X1 U3456 ( .A1(n3436), .A2(n3438), .ZN(n3542) );
  AND2_X1 U3457 ( .A1(n3545), .A2(n3546), .ZN(n3438) );
  NAND2_X1 U3458 ( .A1(n3446), .A2(n3547), .ZN(n3546) );
  NAND2_X1 U3459 ( .A1(n3445), .A2(n3444), .ZN(n3547) );
  NOR2_X1 U3460 ( .A1(n2585), .A2(n2491), .ZN(n3446) );
  OR2_X1 U3461 ( .A1(n3444), .A2(n3445), .ZN(n3545) );
  AND2_X1 U3462 ( .A1(n3548), .A2(n3549), .ZN(n3445) );
  NAND3_X1 U3463 ( .A1(a_3_), .A2(n3550), .A3(b_7_), .ZN(n3549) );
  OR2_X1 U3464 ( .A1(n3532), .A2(n3531), .ZN(n3550) );
  NAND2_X1 U3465 ( .A1(n3531), .A2(n3532), .ZN(n3548) );
  NAND2_X1 U3466 ( .A1(n3551), .A2(n3552), .ZN(n3532) );
  NAND3_X1 U3467 ( .A1(a_4_), .A2(n3553), .A3(b_7_), .ZN(n3552) );
  NAND2_X1 U3468 ( .A1(n3528), .A2(n3526), .ZN(n3553) );
  OR2_X1 U3469 ( .A1(n3526), .A2(n3528), .ZN(n3551) );
  AND2_X1 U3470 ( .A1(n3554), .A2(n3555), .ZN(n3528) );
  NAND3_X1 U3471 ( .A1(a_5_), .A2(n3556), .A3(b_7_), .ZN(n3555) );
  OR2_X1 U3472 ( .A1(n3523), .A2(n3524), .ZN(n3556) );
  NAND2_X1 U3473 ( .A1(n3523), .A2(n3524), .ZN(n3554) );
  NAND2_X1 U3474 ( .A1(n3520), .A2(n3557), .ZN(n3524) );
  NAND2_X1 U3475 ( .A1(n3519), .A2(n3521), .ZN(n3557) );
  NAND2_X1 U3476 ( .A1(n3558), .A2(n3559), .ZN(n3521) );
  NAND2_X1 U3477 ( .A1(b_7_), .A2(a_6_), .ZN(n3559) );
  INV_X1 U3478 ( .A(n3560), .ZN(n3558) );
  XNOR2_X1 U3479 ( .A(n3561), .B(n3562), .ZN(n3519) );
  XNOR2_X1 U3480 ( .A(n3563), .B(n3564), .ZN(n3561) );
  NAND2_X1 U3481 ( .A1(a_6_), .A2(n3560), .ZN(n3520) );
  NAND2_X1 U3482 ( .A1(n3565), .A2(n3566), .ZN(n3560) );
  NAND2_X1 U3483 ( .A1(n3515), .A2(n3567), .ZN(n3566) );
  OR2_X1 U3484 ( .A1(n3516), .A2(n3517), .ZN(n3567) );
  XNOR2_X1 U3485 ( .A(n3568), .B(n3569), .ZN(n3515) );
  XNOR2_X1 U3486 ( .A(n3570), .B(n3571), .ZN(n3568) );
  NAND2_X1 U3487 ( .A1(n3517), .A2(n3516), .ZN(n3565) );
  NAND2_X1 U3488 ( .A1(n3572), .A2(n3573), .ZN(n3516) );
  NAND3_X1 U3489 ( .A1(a_8_), .A2(n3574), .A3(b_7_), .ZN(n3573) );
  NAND2_X1 U3490 ( .A1(n3468), .A2(n3467), .ZN(n3574) );
  OR2_X1 U3491 ( .A1(n3467), .A2(n3468), .ZN(n3572) );
  AND2_X1 U3492 ( .A1(n3575), .A2(n3576), .ZN(n3468) );
  NAND2_X1 U3493 ( .A1(n3476), .A2(n3577), .ZN(n3576) );
  OR2_X1 U3494 ( .A1(n3473), .A2(n3475), .ZN(n3577) );
  NOR2_X1 U3495 ( .A1(n2585), .A2(n2310), .ZN(n3476) );
  NAND2_X1 U3496 ( .A1(n3473), .A2(n3475), .ZN(n3575) );
  NAND2_X1 U3497 ( .A1(n3578), .A2(n3579), .ZN(n3475) );
  NAND3_X1 U3498 ( .A1(a_10_), .A2(n3580), .A3(b_7_), .ZN(n3579) );
  OR2_X1 U3499 ( .A1(n3512), .A2(n3510), .ZN(n3580) );
  NAND2_X1 U3500 ( .A1(n3510), .A2(n3512), .ZN(n3578) );
  NAND2_X1 U3501 ( .A1(n3581), .A2(n3582), .ZN(n3512) );
  NAND2_X1 U3502 ( .A1(n3509), .A2(n3583), .ZN(n3582) );
  OR2_X1 U3503 ( .A1(n3507), .A2(n3508), .ZN(n3583) );
  NOR2_X1 U3504 ( .A1(n2585), .A2(n2581), .ZN(n3509) );
  NAND2_X1 U3505 ( .A1(n3507), .A2(n3508), .ZN(n3581) );
  NAND2_X1 U3506 ( .A1(n3584), .A2(n3585), .ZN(n3508) );
  NAND3_X1 U3507 ( .A1(a_12_), .A2(n3586), .A3(b_7_), .ZN(n3585) );
  NAND2_X1 U3508 ( .A1(n3505), .A2(n3503), .ZN(n3586) );
  OR2_X1 U3509 ( .A1(n3503), .A2(n3505), .ZN(n3584) );
  AND2_X1 U3510 ( .A1(n3587), .A2(n3588), .ZN(n3505) );
  NAND2_X1 U3511 ( .A1(n3499), .A2(n3589), .ZN(n3588) );
  OR2_X1 U3512 ( .A1(n3500), .A2(n3501), .ZN(n3589) );
  NOR2_X1 U3513 ( .A1(n2585), .A2(n2188), .ZN(n3499) );
  NAND2_X1 U3514 ( .A1(n3501), .A2(n3500), .ZN(n3587) );
  NAND2_X1 U3515 ( .A1(n3590), .A2(n3591), .ZN(n3500) );
  NAND2_X1 U3516 ( .A1(b_5_), .A2(n3592), .ZN(n3591) );
  NAND2_X1 U3517 ( .A1(n2156), .A2(n3593), .ZN(n3592) );
  NAND2_X1 U3518 ( .A1(a_15_), .A2(n2385), .ZN(n3593) );
  NAND2_X1 U3519 ( .A1(b_6_), .A2(n3594), .ZN(n3590) );
  NAND2_X1 U3520 ( .A1(n2742), .A2(n3595), .ZN(n3594) );
  NAND2_X1 U3521 ( .A1(a_14_), .A2(n2587), .ZN(n3595) );
  AND3_X1 U3522 ( .A1(b_6_), .A2(b_7_), .A3(n2576), .ZN(n3501) );
  XNOR2_X1 U3523 ( .A(n3596), .B(n3597), .ZN(n3503) );
  XOR2_X1 U3524 ( .A(n3598), .B(n3599), .Z(n3596) );
  XNOR2_X1 U3525 ( .A(n3600), .B(n3601), .ZN(n3507) );
  XOR2_X1 U3526 ( .A(n3602), .B(n3603), .Z(n3600) );
  NAND2_X1 U3527 ( .A1(b_6_), .A2(a_12_), .ZN(n3602) );
  XOR2_X1 U3528 ( .A(n3604), .B(n3605), .Z(n3510) );
  XOR2_X1 U3529 ( .A(n3606), .B(n3607), .Z(n3604) );
  XNOR2_X1 U3530 ( .A(n3608), .B(n3609), .ZN(n3473) );
  XOR2_X1 U3531 ( .A(n3610), .B(n3611), .Z(n3609) );
  NAND2_X1 U3532 ( .A1(b_6_), .A2(a_10_), .ZN(n3611) );
  XOR2_X1 U3533 ( .A(n3612), .B(n3613), .Z(n3467) );
  NAND2_X1 U3534 ( .A1(n3614), .A2(n3615), .ZN(n3612) );
  INV_X1 U3535 ( .A(n2558), .ZN(n3517) );
  NAND2_X1 U3536 ( .A1(b_7_), .A2(a_7_), .ZN(n2558) );
  XOR2_X1 U3537 ( .A(n3616), .B(n3617), .Z(n3523) );
  XOR2_X1 U3538 ( .A(n3618), .B(n3619), .Z(n3616) );
  XOR2_X1 U3539 ( .A(n3620), .B(n3621), .Z(n3526) );
  NAND2_X1 U3540 ( .A1(n3622), .A2(n3623), .ZN(n3620) );
  XNOR2_X1 U3541 ( .A(n3624), .B(n3625), .ZN(n3531) );
  XNOR2_X1 U3542 ( .A(n3626), .B(n3627), .ZN(n3625) );
  XOR2_X1 U3543 ( .A(n3628), .B(n3629), .Z(n3444) );
  NAND2_X1 U3544 ( .A1(n3630), .A2(n3631), .ZN(n3628) );
  XNOR2_X1 U3545 ( .A(n3632), .B(n3633), .ZN(n3436) );
  XNOR2_X1 U3546 ( .A(n3634), .B(n3635), .ZN(n3632) );
  NAND2_X1 U3547 ( .A1(b_6_), .A2(a_2_), .ZN(n3634) );
  XOR2_X1 U3548 ( .A(n3636), .B(n3637), .Z(n3428) );
  XOR2_X1 U3549 ( .A(n3638), .B(n3639), .Z(n3636) );
  XNOR2_X1 U3550 ( .A(n3640), .B(n3641), .ZN(n3425) );
  XOR2_X1 U3551 ( .A(n3642), .B(n3643), .Z(n3641) );
  NAND2_X1 U3552 ( .A1(b_6_), .A2(a_0_), .ZN(n3643) );
  NAND2_X1 U3553 ( .A1(n3644), .A2(n3645), .ZN(n2126) );
  NAND2_X1 U3554 ( .A1(n3537), .A2(n3536), .ZN(n3645) );
  XNOR2_X1 U3555 ( .A(n3646), .B(n3647), .ZN(n3644) );
  NAND3_X1 U3556 ( .A1(n3537), .A2(n3536), .A3(n3648), .ZN(n2127) );
  XOR2_X1 U3557 ( .A(n3646), .B(n3647), .Z(n3648) );
  NAND2_X1 U3558 ( .A1(n3649), .A2(n3650), .ZN(n3536) );
  NAND3_X1 U3559 ( .A1(a_0_), .A2(n3651), .A3(b_6_), .ZN(n3650) );
  OR2_X1 U3560 ( .A1(n3640), .A2(n3642), .ZN(n3651) );
  NAND2_X1 U3561 ( .A1(n3640), .A2(n3642), .ZN(n3649) );
  NAND2_X1 U3562 ( .A1(n3652), .A2(n3653), .ZN(n3642) );
  NAND2_X1 U3563 ( .A1(n3639), .A2(n3654), .ZN(n3653) );
  OR2_X1 U3564 ( .A1(n3638), .A2(n3637), .ZN(n3654) );
  NOR2_X1 U3565 ( .A1(n2385), .A2(n2516), .ZN(n3639) );
  NAND2_X1 U3566 ( .A1(n3637), .A2(n3638), .ZN(n3652) );
  NAND2_X1 U3567 ( .A1(n3655), .A2(n3656), .ZN(n3638) );
  NAND3_X1 U3568 ( .A1(a_2_), .A2(n3657), .A3(b_6_), .ZN(n3656) );
  OR2_X1 U3569 ( .A1(n3633), .A2(n3635), .ZN(n3657) );
  NAND2_X1 U3570 ( .A1(n3633), .A2(n3635), .ZN(n3655) );
  NAND2_X1 U3571 ( .A1(n3630), .A2(n3658), .ZN(n3635) );
  NAND2_X1 U3572 ( .A1(n3629), .A2(n3631), .ZN(n3658) );
  NAND2_X1 U3573 ( .A1(n3659), .A2(n3660), .ZN(n3631) );
  NAND2_X1 U3574 ( .A1(b_6_), .A2(a_3_), .ZN(n3660) );
  INV_X1 U3575 ( .A(n3661), .ZN(n3659) );
  XNOR2_X1 U3576 ( .A(n3662), .B(n3663), .ZN(n3629) );
  XNOR2_X1 U3577 ( .A(n3664), .B(n3665), .ZN(n3662) );
  NOR2_X1 U3578 ( .A1(n2435), .A2(n2587), .ZN(n3665) );
  NAND2_X1 U3579 ( .A1(a_3_), .A2(n3661), .ZN(n3630) );
  NAND2_X1 U3580 ( .A1(n3666), .A2(n3667), .ZN(n3661) );
  NAND2_X1 U3581 ( .A1(n3627), .A2(n3668), .ZN(n3667) );
  OR2_X1 U3582 ( .A1(n3624), .A2(n3626), .ZN(n3668) );
  NOR2_X1 U3583 ( .A1(n2385), .A2(n2435), .ZN(n3627) );
  NAND2_X1 U3584 ( .A1(n3624), .A2(n3626), .ZN(n3666) );
  NAND2_X1 U3585 ( .A1(n3622), .A2(n3669), .ZN(n3626) );
  NAND2_X1 U3586 ( .A1(n3621), .A2(n3623), .ZN(n3669) );
  NAND2_X1 U3587 ( .A1(n3670), .A2(n3671), .ZN(n3623) );
  NAND2_X1 U3588 ( .A1(b_6_), .A2(a_5_), .ZN(n3671) );
  INV_X1 U3589 ( .A(n3672), .ZN(n3670) );
  XNOR2_X1 U3590 ( .A(n3673), .B(n3674), .ZN(n3621) );
  XOR2_X1 U3591 ( .A(n3675), .B(n3676), .Z(n3674) );
  NAND2_X1 U3592 ( .A1(b_5_), .A2(a_6_), .ZN(n3676) );
  NAND2_X1 U3593 ( .A1(a_5_), .A2(n3672), .ZN(n3622) );
  NAND2_X1 U3594 ( .A1(n3677), .A2(n3678), .ZN(n3672) );
  NAND2_X1 U3595 ( .A1(n3617), .A2(n3679), .ZN(n3678) );
  OR2_X1 U3596 ( .A1(n3618), .A2(n3619), .ZN(n3679) );
  XNOR2_X1 U3597 ( .A(n3680), .B(n3681), .ZN(n3617) );
  XNOR2_X1 U3598 ( .A(n3682), .B(n3683), .ZN(n3680) );
  NOR2_X1 U3599 ( .A1(n2360), .A2(n2587), .ZN(n3683) );
  NAND2_X1 U3600 ( .A1(n3619), .A2(n3618), .ZN(n3677) );
  NAND2_X1 U3601 ( .A1(n3684), .A2(n3685), .ZN(n3618) );
  NAND2_X1 U3602 ( .A1(n3563), .A2(n3686), .ZN(n3685) );
  NAND2_X1 U3603 ( .A1(n3564), .A2(n3562), .ZN(n3686) );
  NOR2_X1 U3604 ( .A1(n2385), .A2(n2360), .ZN(n3563) );
  OR2_X1 U3605 ( .A1(n3562), .A2(n3564), .ZN(n3684) );
  AND2_X1 U3606 ( .A1(n3687), .A2(n3688), .ZN(n3564) );
  NAND2_X1 U3607 ( .A1(n3570), .A2(n3689), .ZN(n3688) );
  NAND2_X1 U3608 ( .A1(n3569), .A2(n3571), .ZN(n3689) );
  NOR2_X1 U3609 ( .A1(n2385), .A2(n2584), .ZN(n3570) );
  OR2_X1 U3610 ( .A1(n3569), .A2(n3571), .ZN(n3687) );
  AND2_X1 U3611 ( .A1(n3614), .A2(n3690), .ZN(n3571) );
  NAND2_X1 U3612 ( .A1(n3613), .A2(n3615), .ZN(n3690) );
  NAND2_X1 U3613 ( .A1(n3691), .A2(n3692), .ZN(n3615) );
  NAND2_X1 U3614 ( .A1(b_6_), .A2(a_9_), .ZN(n3692) );
  INV_X1 U3615 ( .A(n3693), .ZN(n3691) );
  XNOR2_X1 U3616 ( .A(n3694), .B(n3695), .ZN(n3613) );
  XOR2_X1 U3617 ( .A(n3696), .B(n3697), .Z(n3695) );
  NAND2_X1 U3618 ( .A1(b_5_), .A2(a_10_), .ZN(n3697) );
  NAND2_X1 U3619 ( .A1(a_9_), .A2(n3693), .ZN(n3614) );
  NAND2_X1 U3620 ( .A1(n3698), .A2(n3699), .ZN(n3693) );
  NAND3_X1 U3621 ( .A1(a_10_), .A2(n3700), .A3(b_6_), .ZN(n3699) );
  OR2_X1 U3622 ( .A1(n3610), .A2(n3608), .ZN(n3700) );
  NAND2_X1 U3623 ( .A1(n3608), .A2(n3610), .ZN(n3698) );
  NAND2_X1 U3624 ( .A1(n3701), .A2(n3702), .ZN(n3610) );
  NAND2_X1 U3625 ( .A1(n3607), .A2(n3703), .ZN(n3702) );
  OR2_X1 U3626 ( .A1(n3605), .A2(n3606), .ZN(n3703) );
  NOR2_X1 U3627 ( .A1(n2385), .A2(n2581), .ZN(n3607) );
  NAND2_X1 U3628 ( .A1(n3605), .A2(n3606), .ZN(n3701) );
  NAND2_X1 U3629 ( .A1(n3704), .A2(n3705), .ZN(n3606) );
  NAND3_X1 U3630 ( .A1(a_12_), .A2(n3706), .A3(b_6_), .ZN(n3705) );
  NAND2_X1 U3631 ( .A1(n3603), .A2(n3601), .ZN(n3706) );
  OR2_X1 U3632 ( .A1(n3601), .A2(n3603), .ZN(n3704) );
  AND2_X1 U3633 ( .A1(n3707), .A2(n3708), .ZN(n3603) );
  NAND2_X1 U3634 ( .A1(n3597), .A2(n3709), .ZN(n3708) );
  OR2_X1 U3635 ( .A1(n3598), .A2(n3599), .ZN(n3709) );
  NOR2_X1 U3636 ( .A1(n2385), .A2(n2188), .ZN(n3597) );
  NAND2_X1 U3637 ( .A1(n3599), .A2(n3598), .ZN(n3707) );
  NAND2_X1 U3638 ( .A1(n3710), .A2(n3711), .ZN(n3598) );
  NAND2_X1 U3639 ( .A1(b_4_), .A2(n3712), .ZN(n3711) );
  NAND2_X1 U3640 ( .A1(n2156), .A2(n3713), .ZN(n3712) );
  NAND2_X1 U3641 ( .A1(a_15_), .A2(n2587), .ZN(n3713) );
  NAND2_X1 U3642 ( .A1(b_5_), .A2(n3714), .ZN(n3710) );
  NAND2_X1 U3643 ( .A1(n2742), .A2(n3715), .ZN(n3714) );
  NAND2_X1 U3644 ( .A1(a_14_), .A2(n2588), .ZN(n3715) );
  AND3_X1 U3645 ( .A1(b_5_), .A2(b_6_), .A3(n2576), .ZN(n3599) );
  XNOR2_X1 U3646 ( .A(n3716), .B(n3717), .ZN(n3601) );
  XOR2_X1 U3647 ( .A(n3718), .B(n3719), .Z(n3716) );
  XNOR2_X1 U3648 ( .A(n3720), .B(n3721), .ZN(n3605) );
  XOR2_X1 U3649 ( .A(n3722), .B(n3723), .Z(n3720) );
  NAND2_X1 U3650 ( .A1(b_5_), .A2(a_12_), .ZN(n3722) );
  XOR2_X1 U3651 ( .A(n3724), .B(n3725), .Z(n3608) );
  XOR2_X1 U3652 ( .A(n3726), .B(n3727), .Z(n3724) );
  XOR2_X1 U3653 ( .A(n3728), .B(n3729), .Z(n3569) );
  NAND2_X1 U3654 ( .A1(n3730), .A2(n3731), .ZN(n3728) );
  XNOR2_X1 U3655 ( .A(n3732), .B(n3733), .ZN(n3562) );
  XNOR2_X1 U3656 ( .A(n3734), .B(n3735), .ZN(n3732) );
  NAND2_X1 U3657 ( .A1(b_5_), .A2(a_8_), .ZN(n3734) );
  INV_X1 U3658 ( .A(n2555), .ZN(n3619) );
  NAND2_X1 U3659 ( .A1(b_6_), .A2(a_6_), .ZN(n2555) );
  XNOR2_X1 U3660 ( .A(n3736), .B(n3737), .ZN(n3624) );
  XNOR2_X1 U3661 ( .A(n2552), .B(n3738), .ZN(n3737) );
  XOR2_X1 U3662 ( .A(n3739), .B(n3740), .Z(n3633) );
  XOR2_X1 U3663 ( .A(n3741), .B(n3742), .Z(n3739) );
  NOR2_X1 U3664 ( .A1(n2466), .A2(n2587), .ZN(n3742) );
  XNOR2_X1 U3665 ( .A(n3743), .B(n3744), .ZN(n3637) );
  XOR2_X1 U3666 ( .A(n3745), .B(n3746), .Z(n3744) );
  NAND2_X1 U3667 ( .A1(b_5_), .A2(a_2_), .ZN(n3746) );
  XOR2_X1 U3668 ( .A(n3747), .B(n3748), .Z(n3640) );
  XOR2_X1 U3669 ( .A(n3749), .B(n3750), .Z(n3747) );
  NOR2_X1 U3670 ( .A1(n2516), .A2(n2587), .ZN(n3750) );
  XNOR2_X1 U3671 ( .A(n3751), .B(n3752), .ZN(n3537) );
  NAND2_X1 U3672 ( .A1(n3753), .A2(n3754), .ZN(n3751) );
  NAND2_X1 U3673 ( .A1(n3755), .A2(n3756), .ZN(n2132) );
  NAND2_X1 U3674 ( .A1(n3647), .A2(n3646), .ZN(n3756) );
  XOR2_X1 U3675 ( .A(n3757), .B(n3758), .Z(n3755) );
  INV_X1 U3676 ( .A(n3759), .ZN(n3758) );
  NAND3_X1 U3677 ( .A1(n3647), .A2(n3646), .A3(n3760), .ZN(n2133) );
  XOR2_X1 U3678 ( .A(n3757), .B(n3759), .Z(n3760) );
  NAND2_X1 U3679 ( .A1(n3753), .A2(n3761), .ZN(n3646) );
  NAND2_X1 U3680 ( .A1(n3752), .A2(n3754), .ZN(n3761) );
  NAND2_X1 U3681 ( .A1(n3762), .A2(n3763), .ZN(n3754) );
  NAND2_X1 U3682 ( .A1(b_5_), .A2(a_0_), .ZN(n3763) );
  INV_X1 U3683 ( .A(n3764), .ZN(n3762) );
  XNOR2_X1 U3684 ( .A(n3765), .B(n3766), .ZN(n3752) );
  XNOR2_X1 U3685 ( .A(n3767), .B(n3768), .ZN(n3765) );
  NAND2_X1 U3686 ( .A1(a_0_), .A2(n3764), .ZN(n3753) );
  NAND2_X1 U3687 ( .A1(n3769), .A2(n3770), .ZN(n3764) );
  NAND3_X1 U3688 ( .A1(a_1_), .A2(n3771), .A3(b_5_), .ZN(n3770) );
  OR2_X1 U3689 ( .A1(n3749), .A2(n3748), .ZN(n3771) );
  NAND2_X1 U3690 ( .A1(n3748), .A2(n3749), .ZN(n3769) );
  NAND2_X1 U3691 ( .A1(n3772), .A2(n3773), .ZN(n3749) );
  NAND3_X1 U3692 ( .A1(a_2_), .A2(n3774), .A3(b_5_), .ZN(n3773) );
  OR2_X1 U3693 ( .A1(n3743), .A2(n3745), .ZN(n3774) );
  NAND2_X1 U3694 ( .A1(n3743), .A2(n3745), .ZN(n3772) );
  NAND2_X1 U3695 ( .A1(n3775), .A2(n3776), .ZN(n3745) );
  NAND3_X1 U3696 ( .A1(a_3_), .A2(n3777), .A3(b_5_), .ZN(n3776) );
  OR2_X1 U3697 ( .A1(n3741), .A2(n3740), .ZN(n3777) );
  NAND2_X1 U3698 ( .A1(n3740), .A2(n3741), .ZN(n3775) );
  NAND2_X1 U3699 ( .A1(n3778), .A2(n3779), .ZN(n3741) );
  NAND3_X1 U3700 ( .A1(a_4_), .A2(n3780), .A3(b_5_), .ZN(n3779) );
  NAND2_X1 U3701 ( .A1(n3663), .A2(n3664), .ZN(n3780) );
  OR2_X1 U3702 ( .A1(n3663), .A2(n3664), .ZN(n3778) );
  AND2_X1 U3703 ( .A1(n3781), .A2(n3782), .ZN(n3664) );
  NAND2_X1 U3704 ( .A1(n3736), .A2(n3783), .ZN(n3782) );
  OR2_X1 U3705 ( .A1(n3738), .A2(n2552), .ZN(n3783) );
  XOR2_X1 U3706 ( .A(n3784), .B(n3785), .Z(n3736) );
  XNOR2_X1 U3707 ( .A(n3786), .B(n3787), .ZN(n3784) );
  NAND2_X1 U3708 ( .A1(b_4_), .A2(a_6_), .ZN(n3786) );
  NAND2_X1 U3709 ( .A1(n2552), .A2(n3738), .ZN(n3781) );
  NAND2_X1 U3710 ( .A1(n3788), .A2(n3789), .ZN(n3738) );
  NAND3_X1 U3711 ( .A1(a_6_), .A2(n3790), .A3(b_5_), .ZN(n3789) );
  OR2_X1 U3712 ( .A1(n3673), .A2(n3675), .ZN(n3790) );
  NAND2_X1 U3713 ( .A1(n3673), .A2(n3675), .ZN(n3788) );
  NAND2_X1 U3714 ( .A1(n3791), .A2(n3792), .ZN(n3675) );
  NAND3_X1 U3715 ( .A1(a_7_), .A2(n3793), .A3(b_5_), .ZN(n3792) );
  NAND2_X1 U3716 ( .A1(n3681), .A2(n3682), .ZN(n3793) );
  OR2_X1 U3717 ( .A1(n3681), .A2(n3682), .ZN(n3791) );
  AND2_X1 U3718 ( .A1(n3794), .A2(n3795), .ZN(n3682) );
  NAND3_X1 U3719 ( .A1(a_8_), .A2(n3796), .A3(b_5_), .ZN(n3795) );
  OR2_X1 U3720 ( .A1(n3733), .A2(n3735), .ZN(n3796) );
  NAND2_X1 U3721 ( .A1(n3733), .A2(n3735), .ZN(n3794) );
  NAND2_X1 U3722 ( .A1(n3730), .A2(n3797), .ZN(n3735) );
  NAND2_X1 U3723 ( .A1(n3729), .A2(n3731), .ZN(n3797) );
  NAND2_X1 U3724 ( .A1(n3798), .A2(n3799), .ZN(n3731) );
  NAND2_X1 U3725 ( .A1(b_5_), .A2(a_9_), .ZN(n3799) );
  INV_X1 U3726 ( .A(n3800), .ZN(n3798) );
  XNOR2_X1 U3727 ( .A(n3801), .B(n3802), .ZN(n3729) );
  XOR2_X1 U3728 ( .A(n3803), .B(n3804), .Z(n3802) );
  NAND2_X1 U3729 ( .A1(b_4_), .A2(a_10_), .ZN(n3804) );
  NAND2_X1 U3730 ( .A1(a_9_), .A2(n3800), .ZN(n3730) );
  NAND2_X1 U3731 ( .A1(n3805), .A2(n3806), .ZN(n3800) );
  NAND3_X1 U3732 ( .A1(a_10_), .A2(n3807), .A3(b_5_), .ZN(n3806) );
  OR2_X1 U3733 ( .A1(n3694), .A2(n3696), .ZN(n3807) );
  NAND2_X1 U3734 ( .A1(n3694), .A2(n3696), .ZN(n3805) );
  NAND2_X1 U3735 ( .A1(n3808), .A2(n3809), .ZN(n3696) );
  NAND2_X1 U3736 ( .A1(n3727), .A2(n3810), .ZN(n3809) );
  OR2_X1 U3737 ( .A1(n3725), .A2(n3726), .ZN(n3810) );
  NOR2_X1 U3738 ( .A1(n2587), .A2(n2581), .ZN(n3727) );
  NAND2_X1 U3739 ( .A1(n3725), .A2(n3726), .ZN(n3808) );
  NAND2_X1 U3740 ( .A1(n3811), .A2(n3812), .ZN(n3726) );
  NAND3_X1 U3741 ( .A1(a_12_), .A2(n3813), .A3(b_5_), .ZN(n3812) );
  NAND2_X1 U3742 ( .A1(n3723), .A2(n3721), .ZN(n3813) );
  OR2_X1 U3743 ( .A1(n3721), .A2(n3723), .ZN(n3811) );
  AND2_X1 U3744 ( .A1(n3814), .A2(n3815), .ZN(n3723) );
  NAND2_X1 U3745 ( .A1(n3717), .A2(n3816), .ZN(n3815) );
  OR2_X1 U3746 ( .A1(n3718), .A2(n3719), .ZN(n3816) );
  NOR2_X1 U3747 ( .A1(n2587), .A2(n2188), .ZN(n3717) );
  NAND2_X1 U3748 ( .A1(n3719), .A2(n3718), .ZN(n3814) );
  NAND2_X1 U3749 ( .A1(n3817), .A2(n3818), .ZN(n3718) );
  NAND2_X1 U3750 ( .A1(b_3_), .A2(n3819), .ZN(n3818) );
  NAND2_X1 U3751 ( .A1(n2156), .A2(n3820), .ZN(n3819) );
  NAND2_X1 U3752 ( .A1(a_15_), .A2(n2588), .ZN(n3820) );
  NAND2_X1 U3753 ( .A1(b_4_), .A2(n3821), .ZN(n3817) );
  NAND2_X1 U3754 ( .A1(n2742), .A2(n3822), .ZN(n3821) );
  NAND2_X1 U3755 ( .A1(a_14_), .A2(n2589), .ZN(n3822) );
  AND3_X1 U3756 ( .A1(b_4_), .A2(b_5_), .A3(n2576), .ZN(n3719) );
  XNOR2_X1 U3757 ( .A(n3823), .B(n3824), .ZN(n3721) );
  XOR2_X1 U3758 ( .A(n3825), .B(n3826), .Z(n3823) );
  XOR2_X1 U3759 ( .A(n3827), .B(n3828), .Z(n3725) );
  XNOR2_X1 U3760 ( .A(n3829), .B(n3830), .ZN(n3827) );
  NAND2_X1 U3761 ( .A1(b_4_), .A2(a_12_), .ZN(n3829) );
  XNOR2_X1 U3762 ( .A(n3831), .B(n3832), .ZN(n3694) );
  NAND2_X1 U3763 ( .A1(n3833), .A2(n3834), .ZN(n3831) );
  XNOR2_X1 U3764 ( .A(n3835), .B(n3836), .ZN(n3733) );
  NAND2_X1 U3765 ( .A1(n3837), .A2(n3838), .ZN(n3835) );
  XNOR2_X1 U3766 ( .A(n3839), .B(n3840), .ZN(n3681) );
  XNOR2_X1 U3767 ( .A(n3841), .B(n3842), .ZN(n3839) );
  NAND2_X1 U3768 ( .A1(b_4_), .A2(a_8_), .ZN(n3841) );
  XOR2_X1 U3769 ( .A(n3843), .B(n3844), .Z(n3673) );
  XOR2_X1 U3770 ( .A(n3845), .B(n3846), .Z(n3843) );
  NOR2_X1 U3771 ( .A1(n2360), .A2(n2588), .ZN(n3846) );
  NOR2_X1 U3772 ( .A1(n2587), .A2(n2410), .ZN(n2552) );
  XNOR2_X1 U3773 ( .A(n3847), .B(n3848), .ZN(n3663) );
  XOR2_X1 U3774 ( .A(n3849), .B(n3850), .Z(n3847) );
  NOR2_X1 U3775 ( .A1(n2410), .A2(n2588), .ZN(n3850) );
  XOR2_X1 U3776 ( .A(n3851), .B(n3852), .Z(n3740) );
  XOR2_X1 U3777 ( .A(n3853), .B(n3854), .Z(n3851) );
  XOR2_X1 U3778 ( .A(n3855), .B(n3856), .Z(n3743) );
  XOR2_X1 U3779 ( .A(n3857), .B(n3858), .Z(n3855) );
  NOR2_X1 U3780 ( .A1(n2466), .A2(n2588), .ZN(n3858) );
  XOR2_X1 U3781 ( .A(n3859), .B(n3860), .Z(n3748) );
  XOR2_X1 U3782 ( .A(n3861), .B(n3862), .Z(n3859) );
  NOR2_X1 U3783 ( .A1(n2491), .A2(n2588), .ZN(n3862) );
  XOR2_X1 U3784 ( .A(n3863), .B(n3864), .Z(n3647) );
  XOR2_X1 U3785 ( .A(n3865), .B(n3866), .Z(n3863) );
  NOR2_X1 U3786 ( .A1(n3102), .A2(n2588), .ZN(n3866) );
  NAND2_X1 U3787 ( .A1(n3867), .A2(n3868), .ZN(n2138) );
  NAND2_X1 U3788 ( .A1(n3759), .A2(n3757), .ZN(n3868) );
  XOR2_X1 U3789 ( .A(n3869), .B(n3870), .Z(n3867) );
  INV_X1 U3790 ( .A(n3871), .ZN(n3870) );
  NAND3_X1 U3791 ( .A1(n3872), .A2(n3757), .A3(n3759), .ZN(n2139) );
  XOR2_X1 U3792 ( .A(n3873), .B(n3874), .Z(n3759) );
  XOR2_X1 U3793 ( .A(n3875), .B(n3876), .Z(n3873) );
  NOR2_X1 U3794 ( .A1(n3102), .A2(n2589), .ZN(n3876) );
  NAND2_X1 U3795 ( .A1(n3877), .A2(n3878), .ZN(n3757) );
  NAND3_X1 U3796 ( .A1(a_0_), .A2(n3879), .A3(b_4_), .ZN(n3878) );
  OR2_X1 U3797 ( .A1(n3865), .A2(n3864), .ZN(n3879) );
  NAND2_X1 U3798 ( .A1(n3864), .A2(n3865), .ZN(n3877) );
  NAND2_X1 U3799 ( .A1(n3880), .A2(n3881), .ZN(n3865) );
  NAND2_X1 U3800 ( .A1(n3768), .A2(n3882), .ZN(n3881) );
  NAND2_X1 U3801 ( .A1(n3767), .A2(n3766), .ZN(n3882) );
  NOR2_X1 U3802 ( .A1(n2588), .A2(n2516), .ZN(n3768) );
  OR2_X1 U3803 ( .A1(n3766), .A2(n3767), .ZN(n3880) );
  AND2_X1 U3804 ( .A1(n3883), .A2(n3884), .ZN(n3767) );
  NAND3_X1 U3805 ( .A1(a_2_), .A2(n3885), .A3(b_4_), .ZN(n3884) );
  OR2_X1 U3806 ( .A1(n3860), .A2(n3861), .ZN(n3885) );
  NAND2_X1 U3807 ( .A1(n3860), .A2(n3861), .ZN(n3883) );
  NAND2_X1 U3808 ( .A1(n3886), .A2(n3887), .ZN(n3861) );
  NAND3_X1 U3809 ( .A1(a_3_), .A2(n3888), .A3(b_4_), .ZN(n3887) );
  OR2_X1 U3810 ( .A1(n3857), .A2(n3856), .ZN(n3888) );
  NAND2_X1 U3811 ( .A1(n3856), .A2(n3857), .ZN(n3886) );
  NAND2_X1 U3812 ( .A1(n3889), .A2(n3890), .ZN(n3857) );
  NAND2_X1 U3813 ( .A1(n3852), .A2(n3891), .ZN(n3890) );
  OR2_X1 U3814 ( .A1(n3853), .A2(n3854), .ZN(n3891) );
  XNOR2_X1 U3815 ( .A(n3892), .B(n3893), .ZN(n3852) );
  XNOR2_X1 U3816 ( .A(n3894), .B(n3895), .ZN(n3892) );
  NOR2_X1 U3817 ( .A1(n2410), .A2(n2589), .ZN(n3895) );
  NAND2_X1 U3818 ( .A1(n3854), .A2(n3853), .ZN(n3889) );
  NAND2_X1 U3819 ( .A1(n3896), .A2(n3897), .ZN(n3853) );
  NAND3_X1 U3820 ( .A1(a_5_), .A2(n3898), .A3(b_4_), .ZN(n3897) );
  OR2_X1 U3821 ( .A1(n3849), .A2(n3848), .ZN(n3898) );
  NAND2_X1 U3822 ( .A1(n3848), .A2(n3849), .ZN(n3896) );
  NAND2_X1 U3823 ( .A1(n3899), .A2(n3900), .ZN(n3849) );
  NAND3_X1 U3824 ( .A1(a_6_), .A2(n3901), .A3(b_4_), .ZN(n3900) );
  OR2_X1 U3825 ( .A1(n3785), .A2(n3787), .ZN(n3901) );
  NAND2_X1 U3826 ( .A1(n3785), .A2(n3787), .ZN(n3899) );
  NAND2_X1 U3827 ( .A1(n3902), .A2(n3903), .ZN(n3787) );
  NAND3_X1 U3828 ( .A1(a_7_), .A2(n3904), .A3(b_4_), .ZN(n3903) );
  OR2_X1 U3829 ( .A1(n3845), .A2(n3844), .ZN(n3904) );
  NAND2_X1 U3830 ( .A1(n3844), .A2(n3845), .ZN(n3902) );
  NAND2_X1 U3831 ( .A1(n3905), .A2(n3906), .ZN(n3845) );
  NAND3_X1 U3832 ( .A1(a_8_), .A2(n3907), .A3(b_4_), .ZN(n3906) );
  OR2_X1 U3833 ( .A1(n3842), .A2(n3840), .ZN(n3907) );
  NAND2_X1 U3834 ( .A1(n3840), .A2(n3842), .ZN(n3905) );
  NAND2_X1 U3835 ( .A1(n3837), .A2(n3908), .ZN(n3842) );
  NAND2_X1 U3836 ( .A1(n3836), .A2(n3838), .ZN(n3908) );
  NAND2_X1 U3837 ( .A1(n3909), .A2(n3910), .ZN(n3838) );
  NAND2_X1 U3838 ( .A1(b_4_), .A2(a_9_), .ZN(n3910) );
  INV_X1 U3839 ( .A(n3911), .ZN(n3909) );
  XNOR2_X1 U3840 ( .A(n3912), .B(n3913), .ZN(n3836) );
  NAND2_X1 U3841 ( .A1(n3914), .A2(n3915), .ZN(n3912) );
  NAND2_X1 U3842 ( .A1(a_9_), .A2(n3911), .ZN(n3837) );
  NAND2_X1 U3843 ( .A1(n3916), .A2(n3917), .ZN(n3911) );
  NAND3_X1 U3844 ( .A1(a_10_), .A2(n3918), .A3(b_4_), .ZN(n3917) );
  OR2_X1 U3845 ( .A1(n3803), .A2(n3801), .ZN(n3918) );
  NAND2_X1 U3846 ( .A1(n3801), .A2(n3803), .ZN(n3916) );
  NAND2_X1 U3847 ( .A1(n3833), .A2(n3919), .ZN(n3803) );
  NAND2_X1 U3848 ( .A1(n3832), .A2(n3834), .ZN(n3919) );
  NAND2_X1 U3849 ( .A1(n3920), .A2(n3921), .ZN(n3834) );
  NAND2_X1 U3850 ( .A1(b_4_), .A2(a_11_), .ZN(n3921) );
  INV_X1 U3851 ( .A(n3922), .ZN(n3920) );
  XNOR2_X1 U3852 ( .A(n3923), .B(n3924), .ZN(n3832) );
  XOR2_X1 U3853 ( .A(n3925), .B(n3926), .Z(n3923) );
  NAND2_X1 U3854 ( .A1(b_3_), .A2(a_12_), .ZN(n3925) );
  NAND2_X1 U3855 ( .A1(a_11_), .A2(n3922), .ZN(n3833) );
  NAND2_X1 U3856 ( .A1(n3927), .A2(n3928), .ZN(n3922) );
  NAND3_X1 U3857 ( .A1(a_12_), .A2(n3929), .A3(b_4_), .ZN(n3928) );
  OR2_X1 U3858 ( .A1(n3830), .A2(n3828), .ZN(n3929) );
  NAND2_X1 U3859 ( .A1(n3828), .A2(n3830), .ZN(n3927) );
  NAND2_X1 U3860 ( .A1(n3930), .A2(n3931), .ZN(n3830) );
  NAND2_X1 U3861 ( .A1(n3824), .A2(n3932), .ZN(n3931) );
  OR2_X1 U3862 ( .A1(n3825), .A2(n3826), .ZN(n3932) );
  NOR2_X1 U3863 ( .A1(n2588), .A2(n2188), .ZN(n3824) );
  NAND2_X1 U3864 ( .A1(n3826), .A2(n3825), .ZN(n3930) );
  NAND2_X1 U3865 ( .A1(n3933), .A2(n3934), .ZN(n3825) );
  NAND2_X1 U3866 ( .A1(b_2_), .A2(n3935), .ZN(n3934) );
  NAND2_X1 U3867 ( .A1(n2156), .A2(n3936), .ZN(n3935) );
  NAND2_X1 U3868 ( .A1(a_15_), .A2(n2589), .ZN(n3936) );
  NAND2_X1 U3869 ( .A1(b_3_), .A2(n3937), .ZN(n3933) );
  NAND2_X1 U3870 ( .A1(n2742), .A2(n3938), .ZN(n3937) );
  NAND2_X1 U3871 ( .A1(a_14_), .A2(n2590), .ZN(n3938) );
  AND3_X1 U3872 ( .A1(b_3_), .A2(b_4_), .A3(n2576), .ZN(n3826) );
  XOR2_X1 U3873 ( .A(n3939), .B(n3940), .Z(n3828) );
  XOR2_X1 U3874 ( .A(n3941), .B(n3942), .Z(n3939) );
  XNOR2_X1 U3875 ( .A(n3943), .B(n3944), .ZN(n3801) );
  NAND2_X1 U3876 ( .A1(n3945), .A2(n3946), .ZN(n3943) );
  XNOR2_X1 U3877 ( .A(n3947), .B(n3948), .ZN(n3840) );
  NAND2_X1 U3878 ( .A1(n3949), .A2(n3950), .ZN(n3947) );
  XOR2_X1 U3879 ( .A(n3951), .B(n3952), .Z(n3844) );
  XOR2_X1 U3880 ( .A(n3953), .B(n3954), .Z(n3951) );
  NOR2_X1 U3881 ( .A1(n2584), .A2(n2589), .ZN(n3954) );
  XOR2_X1 U3882 ( .A(n3955), .B(n3956), .Z(n3785) );
  XOR2_X1 U3883 ( .A(n3957), .B(n3958), .Z(n3955) );
  NOR2_X1 U3884 ( .A1(n2360), .A2(n2589), .ZN(n3958) );
  XOR2_X1 U3885 ( .A(n3959), .B(n3960), .Z(n3848) );
  XOR2_X1 U3886 ( .A(n3961), .B(n3962), .Z(n3959) );
  NOR2_X1 U3887 ( .A1(n2586), .A2(n2589), .ZN(n3962) );
  INV_X1 U3888 ( .A(n2549), .ZN(n3854) );
  NAND2_X1 U3889 ( .A1(b_4_), .A2(a_4_), .ZN(n2549) );
  XOR2_X1 U3890 ( .A(n3963), .B(n3964), .Z(n3856) );
  XOR2_X1 U3891 ( .A(n3965), .B(n3966), .Z(n3963) );
  NOR2_X1 U3892 ( .A1(n2435), .A2(n2589), .ZN(n3966) );
  XOR2_X1 U3893 ( .A(n3967), .B(n3968), .Z(n3860) );
  XOR2_X1 U3894 ( .A(n3969), .B(n3970), .Z(n3967) );
  XNOR2_X1 U3895 ( .A(n3971), .B(n3972), .ZN(n3766) );
  XOR2_X1 U3896 ( .A(n3973), .B(n3974), .Z(n3971) );
  NOR2_X1 U3897 ( .A1(n2491), .A2(n2589), .ZN(n3974) );
  XOR2_X1 U3898 ( .A(n3975), .B(n3976), .Z(n3864) );
  XOR2_X1 U3899 ( .A(n3977), .B(n3978), .Z(n3975) );
  NOR2_X1 U3900 ( .A1(n2516), .A2(n2589), .ZN(n3978) );
  XOR2_X1 U3901 ( .A(n3869), .B(n3871), .Z(n3872) );
  NAND2_X1 U3902 ( .A1(n3979), .A2(n3980), .ZN(n2179) );
  NAND2_X1 U3903 ( .A1(n3871), .A2(n3869), .ZN(n3980) );
  XOR2_X1 U3904 ( .A(n2636), .B(n3981), .Z(n3979) );
  INV_X1 U3905 ( .A(n2635), .ZN(n3981) );
  NAND3_X1 U3906 ( .A1(n3982), .A2(n3869), .A3(n3871), .ZN(n2180) );
  XNOR2_X1 U3907 ( .A(n3983), .B(n3984), .ZN(n3871) );
  NAND2_X1 U3908 ( .A1(n3985), .A2(n3986), .ZN(n3983) );
  NAND2_X1 U3909 ( .A1(n3987), .A2(n3988), .ZN(n3869) );
  NAND3_X1 U3910 ( .A1(a_0_), .A2(n3989), .A3(b_3_), .ZN(n3988) );
  OR2_X1 U3911 ( .A1(n3874), .A2(n3875), .ZN(n3989) );
  NAND2_X1 U3912 ( .A1(n3874), .A2(n3875), .ZN(n3987) );
  NAND2_X1 U3913 ( .A1(n3990), .A2(n3991), .ZN(n3875) );
  NAND3_X1 U3914 ( .A1(a_1_), .A2(n3992), .A3(b_3_), .ZN(n3991) );
  OR2_X1 U3915 ( .A1(n3976), .A2(n3977), .ZN(n3992) );
  NAND2_X1 U3916 ( .A1(n3976), .A2(n3977), .ZN(n3990) );
  NAND2_X1 U3917 ( .A1(n3993), .A2(n3994), .ZN(n3977) );
  NAND3_X1 U3918 ( .A1(a_2_), .A2(n3995), .A3(b_3_), .ZN(n3994) );
  OR2_X1 U3919 ( .A1(n3972), .A2(n3973), .ZN(n3995) );
  NAND2_X1 U3920 ( .A1(n3972), .A2(n3973), .ZN(n3993) );
  NAND2_X1 U3921 ( .A1(n3996), .A2(n3997), .ZN(n3973) );
  NAND2_X1 U3922 ( .A1(n3968), .A2(n3998), .ZN(n3997) );
  OR2_X1 U3923 ( .A1(n3969), .A2(n3970), .ZN(n3998) );
  XNOR2_X1 U3924 ( .A(n3999), .B(n4000), .ZN(n3968) );
  NAND2_X1 U3925 ( .A1(n4001), .A2(n4002), .ZN(n3999) );
  NAND2_X1 U3926 ( .A1(n3970), .A2(n3969), .ZN(n3996) );
  NAND2_X1 U3927 ( .A1(n4003), .A2(n4004), .ZN(n3969) );
  NAND3_X1 U3928 ( .A1(a_4_), .A2(n4005), .A3(b_3_), .ZN(n4004) );
  OR2_X1 U3929 ( .A1(n3964), .A2(n3965), .ZN(n4005) );
  NAND2_X1 U3930 ( .A1(n3964), .A2(n3965), .ZN(n4003) );
  NAND2_X1 U3931 ( .A1(n4006), .A2(n4007), .ZN(n3965) );
  NAND3_X1 U3932 ( .A1(a_5_), .A2(n4008), .A3(b_3_), .ZN(n4007) );
  NAND2_X1 U3933 ( .A1(n3894), .A2(n3893), .ZN(n4008) );
  OR2_X1 U3934 ( .A1(n3893), .A2(n3894), .ZN(n4006) );
  AND2_X1 U3935 ( .A1(n4009), .A2(n4010), .ZN(n3894) );
  NAND3_X1 U3936 ( .A1(a_6_), .A2(n4011), .A3(b_3_), .ZN(n4010) );
  OR2_X1 U3937 ( .A1(n3960), .A2(n3961), .ZN(n4011) );
  NAND2_X1 U3938 ( .A1(n3960), .A2(n3961), .ZN(n4009) );
  NAND2_X1 U3939 ( .A1(n4012), .A2(n4013), .ZN(n3961) );
  NAND3_X1 U3940 ( .A1(a_7_), .A2(n4014), .A3(b_3_), .ZN(n4013) );
  OR2_X1 U3941 ( .A1(n3957), .A2(n3956), .ZN(n4014) );
  NAND2_X1 U3942 ( .A1(n3956), .A2(n3957), .ZN(n4012) );
  NAND2_X1 U3943 ( .A1(n4015), .A2(n4016), .ZN(n3957) );
  NAND3_X1 U3944 ( .A1(a_8_), .A2(n4017), .A3(b_3_), .ZN(n4016) );
  OR2_X1 U3945 ( .A1(n3952), .A2(n3953), .ZN(n4017) );
  NAND2_X1 U3946 ( .A1(n3952), .A2(n3953), .ZN(n4015) );
  NAND2_X1 U3947 ( .A1(n3949), .A2(n4018), .ZN(n3953) );
  NAND2_X1 U3948 ( .A1(n3948), .A2(n3950), .ZN(n4018) );
  NAND2_X1 U3949 ( .A1(n4019), .A2(n4020), .ZN(n3950) );
  NAND2_X1 U3950 ( .A1(b_3_), .A2(a_9_), .ZN(n4020) );
  INV_X1 U3951 ( .A(n4021), .ZN(n4019) );
  XNOR2_X1 U3952 ( .A(n4022), .B(n4023), .ZN(n3948) );
  NAND2_X1 U3953 ( .A1(n4024), .A2(n4025), .ZN(n4022) );
  NAND2_X1 U3954 ( .A1(a_9_), .A2(n4021), .ZN(n3949) );
  NAND2_X1 U3955 ( .A1(n3914), .A2(n4026), .ZN(n4021) );
  NAND2_X1 U3956 ( .A1(n3913), .A2(n3915), .ZN(n4026) );
  NAND2_X1 U3957 ( .A1(n4027), .A2(n4028), .ZN(n3915) );
  NAND2_X1 U3958 ( .A1(b_3_), .A2(a_10_), .ZN(n4028) );
  INV_X1 U3959 ( .A(n4029), .ZN(n4027) );
  XNOR2_X1 U3960 ( .A(n4030), .B(n4031), .ZN(n3913) );
  XNOR2_X1 U3961 ( .A(n4032), .B(n4033), .ZN(n4031) );
  NAND2_X1 U3962 ( .A1(a_10_), .A2(n4029), .ZN(n3914) );
  NAND2_X1 U3963 ( .A1(n3945), .A2(n4034), .ZN(n4029) );
  NAND2_X1 U3964 ( .A1(n3944), .A2(n3946), .ZN(n4034) );
  NAND2_X1 U3965 ( .A1(n4035), .A2(n4036), .ZN(n3946) );
  NAND2_X1 U3966 ( .A1(b_3_), .A2(a_11_), .ZN(n4036) );
  INV_X1 U3967 ( .A(n4037), .ZN(n4035) );
  XNOR2_X1 U3968 ( .A(n4038), .B(n4039), .ZN(n3944) );
  XNOR2_X1 U3969 ( .A(n4040), .B(n4041), .ZN(n4039) );
  NOR2_X1 U3970 ( .A1(n2579), .A2(n2590), .ZN(n4041) );
  NAND2_X1 U3971 ( .A1(a_11_), .A2(n4037), .ZN(n3945) );
  NAND2_X1 U3972 ( .A1(n4042), .A2(n4043), .ZN(n4037) );
  NAND3_X1 U3973 ( .A1(a_12_), .A2(n4044), .A3(b_3_), .ZN(n4043) );
  NAND2_X1 U3974 ( .A1(n3926), .A2(n3924), .ZN(n4044) );
  OR2_X1 U3975 ( .A1(n3924), .A2(n3926), .ZN(n4042) );
  AND2_X1 U3976 ( .A1(n4045), .A2(n4046), .ZN(n3926) );
  NAND2_X1 U3977 ( .A1(n3940), .A2(n4047), .ZN(n4046) );
  OR2_X1 U3978 ( .A1(n3941), .A2(n3942), .ZN(n4047) );
  NOR2_X1 U3979 ( .A1(n2589), .A2(n2188), .ZN(n3940) );
  NAND2_X1 U3980 ( .A1(n3942), .A2(n3941), .ZN(n4045) );
  NAND2_X1 U3981 ( .A1(n4048), .A2(n4049), .ZN(n3941) );
  NAND2_X1 U3982 ( .A1(b_1_), .A2(n4050), .ZN(n4049) );
  NAND2_X1 U3983 ( .A1(n2156), .A2(n4051), .ZN(n4050) );
  NAND2_X1 U3984 ( .A1(a_15_), .A2(n2590), .ZN(n4051) );
  NAND2_X1 U3985 ( .A1(b_2_), .A2(n4052), .ZN(n4048) );
  NAND2_X1 U3986 ( .A1(n2742), .A2(n4053), .ZN(n4052) );
  NAND2_X1 U3987 ( .A1(a_14_), .A2(n2591), .ZN(n4053) );
  AND3_X1 U3988 ( .A1(b_2_), .A2(b_3_), .A3(n2576), .ZN(n3942) );
  XNOR2_X1 U3989 ( .A(n4054), .B(n4055), .ZN(n3924) );
  NOR2_X1 U3990 ( .A1(n2188), .A2(n2590), .ZN(n4055) );
  XOR2_X1 U3991 ( .A(n4056), .B(n4057), .Z(n4054) );
  XOR2_X1 U3992 ( .A(n4058), .B(n4059), .Z(n3952) );
  XOR2_X1 U3993 ( .A(n4060), .B(n4061), .Z(n4058) );
  XNOR2_X1 U3994 ( .A(n4062), .B(n4063), .ZN(n3956) );
  NAND2_X1 U3995 ( .A1(n4064), .A2(n4065), .ZN(n4062) );
  XOR2_X1 U3996 ( .A(n4066), .B(n4067), .Z(n3960) );
  XOR2_X1 U3997 ( .A(n4068), .B(n4069), .Z(n4066) );
  XOR2_X1 U3998 ( .A(n4070), .B(n4071), .Z(n3893) );
  NAND2_X1 U3999 ( .A1(n4072), .A2(n4073), .ZN(n4070) );
  XOR2_X1 U4000 ( .A(n4074), .B(n4075), .Z(n3964) );
  XOR2_X1 U4001 ( .A(n4076), .B(n4077), .Z(n4074) );
  INV_X1 U4002 ( .A(n2546), .ZN(n3970) );
  NAND2_X1 U4003 ( .A1(b_3_), .A2(a_3_), .ZN(n2546) );
  XOR2_X1 U4004 ( .A(n4078), .B(n4079), .Z(n3972) );
  XOR2_X1 U4005 ( .A(n4080), .B(n4081), .Z(n4078) );
  XOR2_X1 U4006 ( .A(n4082), .B(n4083), .Z(n3976) );
  XOR2_X1 U4007 ( .A(n2543), .B(n4084), .Z(n4082) );
  XOR2_X1 U4008 ( .A(n4085), .B(n4086), .Z(n3874) );
  XOR2_X1 U4009 ( .A(n4087), .B(n4088), .Z(n4085) );
  NOR2_X1 U4010 ( .A1(n2516), .A2(n2590), .ZN(n4088) );
  XOR2_X1 U4011 ( .A(n2636), .B(n2635), .Z(n3982) );
  NAND2_X1 U4012 ( .A1(n4089), .A2(n4090), .ZN(n2440) );
  NAND2_X1 U4013 ( .A1(n2635), .A2(n2636), .ZN(n4090) );
  NAND2_X1 U4014 ( .A1(n3985), .A2(n4091), .ZN(n2636) );
  NAND2_X1 U4015 ( .A1(n3984), .A2(n3986), .ZN(n4091) );
  NAND2_X1 U4016 ( .A1(n4092), .A2(n4093), .ZN(n3986) );
  NAND2_X1 U4017 ( .A1(b_2_), .A2(a_0_), .ZN(n4093) );
  INV_X1 U4018 ( .A(n4094), .ZN(n4092) );
  XOR2_X1 U4019 ( .A(n4095), .B(n4096), .Z(n3984) );
  NOR2_X1 U4020 ( .A1(n2491), .A2(n2593), .ZN(n4096) );
  XOR2_X1 U4021 ( .A(n2542), .B(n4097), .Z(n4095) );
  NAND2_X1 U4022 ( .A1(a_0_), .A2(n4094), .ZN(n3985) );
  NAND2_X1 U4023 ( .A1(n4098), .A2(n4099), .ZN(n4094) );
  NAND3_X1 U4024 ( .A1(a_1_), .A2(n4100), .A3(b_2_), .ZN(n4099) );
  OR2_X1 U4025 ( .A1(n4087), .A2(n4086), .ZN(n4100) );
  NAND2_X1 U4026 ( .A1(n4086), .A2(n4087), .ZN(n4098) );
  NAND2_X1 U4027 ( .A1(n4101), .A2(n4102), .ZN(n4087) );
  NAND2_X1 U4028 ( .A1(n4083), .A2(n4103), .ZN(n4102) );
  NAND2_X1 U4029 ( .A1(n4084), .A2(n2543), .ZN(n4103) );
  XOR2_X1 U4030 ( .A(n4104), .B(n4105), .Z(n4083) );
  NOR2_X1 U4031 ( .A1(n2466), .A2(n2591), .ZN(n4105) );
  XOR2_X1 U4032 ( .A(n4106), .B(n4107), .Z(n4104) );
  OR2_X1 U4033 ( .A1(n2543), .A2(n4084), .ZN(n4101) );
  AND2_X1 U4034 ( .A1(n4108), .A2(n4109), .ZN(n4084) );
  NAND2_X1 U4035 ( .A1(n4081), .A2(n4110), .ZN(n4109) );
  OR2_X1 U4036 ( .A1(n4080), .A2(n4079), .ZN(n4110) );
  NOR2_X1 U4037 ( .A1(n2590), .A2(n2466), .ZN(n4081) );
  NAND2_X1 U4038 ( .A1(n4079), .A2(n4080), .ZN(n4108) );
  NAND2_X1 U4039 ( .A1(n4001), .A2(n4111), .ZN(n4080) );
  NAND2_X1 U4040 ( .A1(n4000), .A2(n4002), .ZN(n4111) );
  NAND2_X1 U4041 ( .A1(n4112), .A2(n4113), .ZN(n4002) );
  NAND2_X1 U4042 ( .A1(b_2_), .A2(a_4_), .ZN(n4113) );
  INV_X1 U4043 ( .A(n4114), .ZN(n4112) );
  XOR2_X1 U4044 ( .A(n4115), .B(n4116), .Z(n4000) );
  NOR2_X1 U4045 ( .A1(n2410), .A2(n2591), .ZN(n4116) );
  XOR2_X1 U4046 ( .A(n4117), .B(n4118), .Z(n4115) );
  NAND2_X1 U4047 ( .A1(a_4_), .A2(n4114), .ZN(n4001) );
  NAND2_X1 U4048 ( .A1(n4119), .A2(n4120), .ZN(n4114) );
  NAND2_X1 U4049 ( .A1(n4077), .A2(n4121), .ZN(n4120) );
  OR2_X1 U4050 ( .A1(n4076), .A2(n4075), .ZN(n4121) );
  NOR2_X1 U4051 ( .A1(n2590), .A2(n2410), .ZN(n4077) );
  NAND2_X1 U4052 ( .A1(n4075), .A2(n4076), .ZN(n4119) );
  NAND2_X1 U4053 ( .A1(n4072), .A2(n4122), .ZN(n4076) );
  NAND2_X1 U4054 ( .A1(n4071), .A2(n4073), .ZN(n4122) );
  NAND2_X1 U4055 ( .A1(n4123), .A2(n4124), .ZN(n4073) );
  NAND2_X1 U4056 ( .A1(b_2_), .A2(a_6_), .ZN(n4124) );
  INV_X1 U4057 ( .A(n4125), .ZN(n4123) );
  XOR2_X1 U4058 ( .A(n4126), .B(n4127), .Z(n4071) );
  NOR2_X1 U4059 ( .A1(n2360), .A2(n2591), .ZN(n4127) );
  XOR2_X1 U4060 ( .A(n4128), .B(n4129), .Z(n4126) );
  NAND2_X1 U4061 ( .A1(a_6_), .A2(n4125), .ZN(n4072) );
  NAND2_X1 U4062 ( .A1(n4130), .A2(n4131), .ZN(n4125) );
  NAND2_X1 U4063 ( .A1(n4069), .A2(n4132), .ZN(n4131) );
  OR2_X1 U4064 ( .A1(n4068), .A2(n4067), .ZN(n4132) );
  NOR2_X1 U4065 ( .A1(n2590), .A2(n2360), .ZN(n4069) );
  NAND2_X1 U4066 ( .A1(n4067), .A2(n4068), .ZN(n4130) );
  NAND2_X1 U4067 ( .A1(n4064), .A2(n4133), .ZN(n4068) );
  NAND2_X1 U4068 ( .A1(n4063), .A2(n4065), .ZN(n4133) );
  NAND2_X1 U4069 ( .A1(n4134), .A2(n4135), .ZN(n4065) );
  NAND2_X1 U4070 ( .A1(b_2_), .A2(a_8_), .ZN(n4135) );
  INV_X1 U4071 ( .A(n4136), .ZN(n4134) );
  XOR2_X1 U4072 ( .A(n4137), .B(n4138), .Z(n4063) );
  NOR2_X1 U4073 ( .A1(n2310), .A2(n2591), .ZN(n4138) );
  XOR2_X1 U4074 ( .A(n4139), .B(n4140), .Z(n4137) );
  NAND2_X1 U4075 ( .A1(a_8_), .A2(n4136), .ZN(n4064) );
  NAND2_X1 U4076 ( .A1(n4141), .A2(n4142), .ZN(n4136) );
  NAND2_X1 U4077 ( .A1(n4061), .A2(n4143), .ZN(n4142) );
  OR2_X1 U4078 ( .A1(n4060), .A2(n4059), .ZN(n4143) );
  NOR2_X1 U4079 ( .A1(n2590), .A2(n2310), .ZN(n4061) );
  NAND2_X1 U4080 ( .A1(n4059), .A2(n4060), .ZN(n4141) );
  NAND2_X1 U4081 ( .A1(n4024), .A2(n4144), .ZN(n4060) );
  NAND2_X1 U4082 ( .A1(n4023), .A2(n4025), .ZN(n4144) );
  NAND2_X1 U4083 ( .A1(n4145), .A2(n4146), .ZN(n4025) );
  NAND2_X1 U4084 ( .A1(b_2_), .A2(a_10_), .ZN(n4146) );
  INV_X1 U4085 ( .A(n4147), .ZN(n4145) );
  XOR2_X1 U4086 ( .A(n4148), .B(n4149), .Z(n4023) );
  NOR2_X1 U4087 ( .A1(n2581), .A2(n2591), .ZN(n4149) );
  XOR2_X1 U4088 ( .A(n4150), .B(n4151), .Z(n4148) );
  NAND2_X1 U4089 ( .A1(a_10_), .A2(n4147), .ZN(n4024) );
  NAND2_X1 U4090 ( .A1(n4152), .A2(n4153), .ZN(n4147) );
  NAND2_X1 U4091 ( .A1(n4033), .A2(n4154), .ZN(n4153) );
  OR2_X1 U4092 ( .A1(n4032), .A2(n4030), .ZN(n4154) );
  NOR2_X1 U4093 ( .A1(n2590), .A2(n2581), .ZN(n4033) );
  NAND2_X1 U4094 ( .A1(n4030), .A2(n4032), .ZN(n4152) );
  NAND2_X1 U4095 ( .A1(n4155), .A2(n4156), .ZN(n4032) );
  NAND3_X1 U4096 ( .A1(a_12_), .A2(n4157), .A3(b_2_), .ZN(n4156) );
  OR2_X1 U4097 ( .A1(n4038), .A2(n4040), .ZN(n4157) );
  NAND2_X1 U4098 ( .A1(n4038), .A2(n4040), .ZN(n4155) );
  NAND2_X1 U4099 ( .A1(n4158), .A2(n4159), .ZN(n4040) );
  NAND3_X1 U4100 ( .A1(a_13_), .A2(n4160), .A3(b_2_), .ZN(n4159) );
  OR2_X1 U4101 ( .A1(n4056), .A2(n4057), .ZN(n4160) );
  NAND2_X1 U4102 ( .A1(n4057), .A2(n4056), .ZN(n4158) );
  NAND2_X1 U4103 ( .A1(n4161), .A2(n4162), .ZN(n4056) );
  NAND2_X1 U4104 ( .A1(b_0_), .A2(n4163), .ZN(n4162) );
  NAND2_X1 U4105 ( .A1(n2156), .A2(n4164), .ZN(n4163) );
  NAND2_X1 U4106 ( .A1(a_15_), .A2(n2591), .ZN(n4164) );
  NAND2_X1 U4107 ( .A1(a_15_), .A2(n2158), .ZN(n2156) );
  NAND2_X1 U4108 ( .A1(b_1_), .A2(n4165), .ZN(n4161) );
  NAND2_X1 U4109 ( .A1(n2742), .A2(n4166), .ZN(n4165) );
  NAND2_X1 U4110 ( .A1(a_14_), .A2(n2593), .ZN(n4166) );
  NAND2_X1 U4111 ( .A1(a_14_), .A2(n4167), .ZN(n2742) );
  AND3_X1 U4112 ( .A1(b_1_), .A2(b_2_), .A3(n2576), .ZN(n4057) );
  XNOR2_X1 U4113 ( .A(n4168), .B(n4169), .ZN(n4038) );
  XNOR2_X1 U4114 ( .A(n4170), .B(n4171), .ZN(n4169) );
  NAND2_X1 U4115 ( .A1(b_0_), .A2(a_14_), .ZN(n4168) );
  XNOR2_X1 U4116 ( .A(n4172), .B(n4173), .ZN(n4030) );
  NAND2_X1 U4117 ( .A1(n4174), .A2(n4175), .ZN(n4172) );
  NAND2_X1 U4118 ( .A1(n4176), .A2(n4177), .ZN(n4175) );
  NAND2_X1 U4119 ( .A1(b_1_), .A2(a_12_), .ZN(n4176) );
  XOR2_X1 U4120 ( .A(n4178), .B(n4179), .Z(n4059) );
  XNOR2_X1 U4121 ( .A(n4180), .B(n4181), .ZN(n4179) );
  NAND2_X1 U4122 ( .A1(b_1_), .A2(a_10_), .ZN(n4178) );
  XOR2_X1 U4123 ( .A(n4182), .B(n4183), .Z(n4067) );
  XNOR2_X1 U4124 ( .A(n4184), .B(n4185), .ZN(n4183) );
  NAND2_X1 U4125 ( .A1(b_1_), .A2(a_8_), .ZN(n4182) );
  XOR2_X1 U4126 ( .A(n4186), .B(n4187), .Z(n4075) );
  XNOR2_X1 U4127 ( .A(n4188), .B(n4189), .ZN(n4187) );
  NAND2_X1 U4128 ( .A1(b_1_), .A2(a_6_), .ZN(n4186) );
  XOR2_X1 U4129 ( .A(n4190), .B(n4191), .Z(n4079) );
  XNOR2_X1 U4130 ( .A(n4192), .B(n4193), .ZN(n4191) );
  NAND2_X1 U4131 ( .A1(b_1_), .A2(a_4_), .ZN(n4190) );
  NAND2_X1 U4132 ( .A1(b_2_), .A2(a_2_), .ZN(n2543) );
  XOR2_X1 U4133 ( .A(n4194), .B(n4195), .Z(n4086) );
  XNOR2_X1 U4134 ( .A(n4196), .B(n4197), .ZN(n4195) );
  NAND2_X1 U4135 ( .A1(b_1_), .A2(a_2_), .ZN(n4194) );
  XOR2_X1 U4136 ( .A(n4198), .B(n4199), .Z(n2635) );
  XNOR2_X1 U4137 ( .A(n4200), .B(n4201), .ZN(n4199) );
  NAND2_X1 U4138 ( .A1(b_0_), .A2(a_1_), .ZN(n4198) );
  XOR2_X1 U4139 ( .A(n2634), .B(n2633), .Z(n4089) );
  NOR2_X1 U4140 ( .A1(n2593), .A2(n3102), .ZN(n2633) );
  INV_X1 U4141 ( .A(n2632), .ZN(n2634) );
  NAND2_X1 U4142 ( .A1(n4202), .A2(n4203), .ZN(n2632) );
  NAND3_X1 U4143 ( .A1(a_1_), .A2(n4204), .A3(b_0_), .ZN(n4203) );
  OR2_X1 U4144 ( .A1(n4201), .A2(n4200), .ZN(n4204) );
  NAND2_X1 U4145 ( .A1(n4200), .A2(n4201), .ZN(n4202) );
  NAND2_X1 U4146 ( .A1(n4205), .A2(n4206), .ZN(n4201) );
  NAND3_X1 U4147 ( .A1(a_2_), .A2(n4207), .A3(b_0_), .ZN(n4206) );
  NAND2_X1 U4148 ( .A1(n4097), .A2(n2542), .ZN(n4207) );
  OR2_X1 U4149 ( .A1(n2542), .A2(n4097), .ZN(n4205) );
  AND2_X1 U4150 ( .A1(n4208), .A2(n4209), .ZN(n4097) );
  NAND3_X1 U4151 ( .A1(a_2_), .A2(n4210), .A3(b_1_), .ZN(n4209) );
  OR2_X1 U4152 ( .A1(n4197), .A2(n4196), .ZN(n4210) );
  NAND2_X1 U4153 ( .A1(n4196), .A2(n4197), .ZN(n4208) );
  NAND2_X1 U4154 ( .A1(n4211), .A2(n4212), .ZN(n4197) );
  NAND3_X1 U4155 ( .A1(a_3_), .A2(n4213), .A3(b_1_), .ZN(n4212) );
  OR2_X1 U4156 ( .A1(n4107), .A2(n4106), .ZN(n4213) );
  NAND2_X1 U4157 ( .A1(n4106), .A2(n4107), .ZN(n4211) );
  NAND2_X1 U4158 ( .A1(n4214), .A2(n4215), .ZN(n4107) );
  NAND3_X1 U4159 ( .A1(a_4_), .A2(n4216), .A3(b_1_), .ZN(n4215) );
  OR2_X1 U4160 ( .A1(n4193), .A2(n4192), .ZN(n4216) );
  NAND2_X1 U4161 ( .A1(n4192), .A2(n4193), .ZN(n4214) );
  NAND2_X1 U4162 ( .A1(n4217), .A2(n4218), .ZN(n4193) );
  NAND3_X1 U4163 ( .A1(a_5_), .A2(n4219), .A3(b_1_), .ZN(n4218) );
  OR2_X1 U4164 ( .A1(n4118), .A2(n4117), .ZN(n4219) );
  NAND2_X1 U4165 ( .A1(n4117), .A2(n4118), .ZN(n4217) );
  NAND2_X1 U4166 ( .A1(n4220), .A2(n4221), .ZN(n4118) );
  NAND3_X1 U4167 ( .A1(a_6_), .A2(n4222), .A3(b_1_), .ZN(n4221) );
  OR2_X1 U4168 ( .A1(n4189), .A2(n4188), .ZN(n4222) );
  NAND2_X1 U4169 ( .A1(n4188), .A2(n4189), .ZN(n4220) );
  NAND2_X1 U4170 ( .A1(n4223), .A2(n4224), .ZN(n4189) );
  NAND3_X1 U4171 ( .A1(a_7_), .A2(n4225), .A3(b_1_), .ZN(n4224) );
  OR2_X1 U4172 ( .A1(n4129), .A2(n4128), .ZN(n4225) );
  NAND2_X1 U4173 ( .A1(n4128), .A2(n4129), .ZN(n4223) );
  NAND2_X1 U4174 ( .A1(n4226), .A2(n4227), .ZN(n4129) );
  NAND3_X1 U4175 ( .A1(a_8_), .A2(n4228), .A3(b_1_), .ZN(n4227) );
  OR2_X1 U4176 ( .A1(n4185), .A2(n4184), .ZN(n4228) );
  NAND2_X1 U4177 ( .A1(n4184), .A2(n4185), .ZN(n4226) );
  NAND2_X1 U4178 ( .A1(n4229), .A2(n4230), .ZN(n4185) );
  NAND3_X1 U4179 ( .A1(a_9_), .A2(n4231), .A3(b_1_), .ZN(n4230) );
  OR2_X1 U4180 ( .A1(n4140), .A2(n4139), .ZN(n4231) );
  NAND2_X1 U4181 ( .A1(n4139), .A2(n4140), .ZN(n4229) );
  NAND2_X1 U4182 ( .A1(n4232), .A2(n4233), .ZN(n4140) );
  NAND3_X1 U4183 ( .A1(a_10_), .A2(n4234), .A3(b_1_), .ZN(n4233) );
  OR2_X1 U4184 ( .A1(n4181), .A2(n4180), .ZN(n4234) );
  NAND2_X1 U4185 ( .A1(n4180), .A2(n4181), .ZN(n4232) );
  NAND2_X1 U4186 ( .A1(n4235), .A2(n4236), .ZN(n4181) );
  NAND3_X1 U4187 ( .A1(a_11_), .A2(n4237), .A3(b_1_), .ZN(n4236) );
  OR2_X1 U4188 ( .A1(n4151), .A2(n4150), .ZN(n4237) );
  NAND2_X1 U4189 ( .A1(n4150), .A2(n4151), .ZN(n4235) );
  NAND2_X1 U4190 ( .A1(n4174), .A2(n4238), .ZN(n4151) );
  NAND2_X1 U4191 ( .A1(n4239), .A2(n4173), .ZN(n4238) );
  NAND2_X1 U4192 ( .A1(n4171), .A2(n4240), .ZN(n4173) );
  NAND3_X1 U4193 ( .A1(b_0_), .A2(a_14_), .A3(n4170), .ZN(n4240) );
  NOR2_X1 U4194 ( .A1(n2591), .A2(n2188), .ZN(n4170) );
  NAND3_X1 U4195 ( .A1(b_0_), .A2(b_1_), .A3(n2576), .ZN(n4171) );
  NOR2_X1 U4196 ( .A1(n4167), .A2(n2158), .ZN(n2576) );
  NAND2_X1 U4197 ( .A1(n4177), .A2(n2579), .ZN(n4239) );
  OR3_X1 U4198 ( .A1(n2591), .A2(n2579), .A3(n4177), .ZN(n4174) );
  NAND2_X1 U4199 ( .A1(b_0_), .A2(a_13_), .ZN(n4177) );
  NOR2_X1 U4200 ( .A1(n2593), .A2(n2579), .ZN(n4150) );
  NOR2_X1 U4201 ( .A1(n2593), .A2(n2581), .ZN(n4180) );
  NOR2_X1 U4202 ( .A1(n2593), .A2(n2582), .ZN(n4139) );
  NOR2_X1 U4203 ( .A1(n2593), .A2(n2310), .ZN(n4184) );
  NOR2_X1 U4204 ( .A1(n2593), .A2(n2584), .ZN(n4128) );
  NOR2_X1 U4205 ( .A1(n2593), .A2(n2360), .ZN(n4188) );
  NOR2_X1 U4206 ( .A1(n2593), .A2(n2586), .ZN(n4117) );
  NOR2_X1 U4207 ( .A1(n2593), .A2(n2410), .ZN(n4192) );
  NOR2_X1 U4208 ( .A1(n2593), .A2(n2435), .ZN(n4106) );
  NOR2_X1 U4209 ( .A1(n2593), .A2(n2466), .ZN(n4196) );
  NAND2_X1 U4210 ( .A1(b_1_), .A2(a_1_), .ZN(n2542) );
  NOR2_X1 U4211 ( .A1(n2591), .A2(n3102), .ZN(n4200) );
  AND2_X1 U4212 ( .A1(n4243), .A2(n4244), .ZN(n2097) );
  NAND3_X1 U4213 ( .A1(n4245), .A2(n4246), .A3(n2095), .ZN(n4244) );
  INV_X1 U4214 ( .A(operation_1_), .ZN(n4242) );
  NAND2_X1 U4215 ( .A1(n4247), .A2(n2593), .ZN(n4246) );
  INV_X1 U4216 ( .A(b_0_), .ZN(n2593) );
  NAND2_X1 U4217 ( .A1(n2592), .A2(n3102), .ZN(n4247) );
  INV_X1 U4218 ( .A(n2532), .ZN(n2592) );
  NAND2_X1 U4219 ( .A1(a_0_), .A2(n2532), .ZN(n4245) );
  NAND2_X1 U4220 ( .A1(n4248), .A2(n4249), .ZN(n2532) );
  NAND2_X1 U4221 ( .A1(n4250), .A2(n2591), .ZN(n4249) );
  INV_X1 U4222 ( .A(b_1_), .ZN(n2591) );
  NAND2_X1 U4223 ( .A1(n2515), .A2(n2516), .ZN(n4250) );
  INV_X1 U4224 ( .A(n2507), .ZN(n2515) );
  NAND2_X1 U4225 ( .A1(a_1_), .A2(n2507), .ZN(n4248) );
  NAND2_X1 U4226 ( .A1(n4251), .A2(n4252), .ZN(n2507) );
  NAND2_X1 U4227 ( .A1(n4253), .A2(n2590), .ZN(n4252) );
  INV_X1 U4228 ( .A(b_2_), .ZN(n2590) );
  NAND2_X1 U4229 ( .A1(n2490), .A2(n2491), .ZN(n4253) );
  INV_X1 U4230 ( .A(n2483), .ZN(n2490) );
  NAND2_X1 U4231 ( .A1(a_2_), .A2(n2483), .ZN(n4251) );
  NAND2_X1 U4232 ( .A1(n4254), .A2(n4255), .ZN(n2483) );
  NAND2_X1 U4233 ( .A1(n4256), .A2(n2589), .ZN(n4255) );
  INV_X1 U4234 ( .A(b_3_), .ZN(n2589) );
  NAND2_X1 U4235 ( .A1(n2465), .A2(n2466), .ZN(n4256) );
  INV_X1 U4236 ( .A(n2458), .ZN(n2465) );
  NAND2_X1 U4237 ( .A1(a_3_), .A2(n2458), .ZN(n4254) );
  NAND2_X1 U4238 ( .A1(n4257), .A2(n4258), .ZN(n2458) );
  NAND2_X1 U4239 ( .A1(n4259), .A2(n2588), .ZN(n4258) );
  INV_X1 U4240 ( .A(b_4_), .ZN(n2588) );
  NAND2_X1 U4241 ( .A1(n2434), .A2(n2435), .ZN(n4259) );
  INV_X1 U4242 ( .A(n2426), .ZN(n2434) );
  NAND2_X1 U4243 ( .A1(a_4_), .A2(n2426), .ZN(n4257) );
  NAND2_X1 U4244 ( .A1(n4260), .A2(n4261), .ZN(n2426) );
  NAND2_X1 U4245 ( .A1(n4262), .A2(n2587), .ZN(n4261) );
  INV_X1 U4246 ( .A(b_5_), .ZN(n2587) );
  NAND2_X1 U4247 ( .A1(n2409), .A2(n2410), .ZN(n4262) );
  INV_X1 U4248 ( .A(n2402), .ZN(n2409) );
  NAND2_X1 U4249 ( .A1(a_5_), .A2(n2402), .ZN(n4260) );
  NAND2_X1 U4250 ( .A1(n4263), .A2(n4264), .ZN(n2402) );
  NAND2_X1 U4251 ( .A1(n4265), .A2(n2385), .ZN(n4264) );
  INV_X1 U4252 ( .A(b_6_), .ZN(n2385) );
  NAND2_X1 U4253 ( .A1(n2384), .A2(n2586), .ZN(n4265) );
  INV_X1 U4254 ( .A(n2377), .ZN(n2384) );
  NAND2_X1 U4255 ( .A1(a_6_), .A2(n2377), .ZN(n4263) );
  NAND2_X1 U4256 ( .A1(n4266), .A2(n4267), .ZN(n2377) );
  NAND2_X1 U4257 ( .A1(n4268), .A2(n2585), .ZN(n4267) );
  INV_X1 U4258 ( .A(b_7_), .ZN(n2585) );
  NAND2_X1 U4259 ( .A1(n2359), .A2(n2360), .ZN(n4268) );
  INV_X1 U4260 ( .A(n2352), .ZN(n2359) );
  NAND2_X1 U4261 ( .A1(a_7_), .A2(n2352), .ZN(n4266) );
  NAND2_X1 U4262 ( .A1(n4269), .A2(n4270), .ZN(n2352) );
  NAND2_X1 U4263 ( .A1(n4271), .A2(n2335), .ZN(n4270) );
  INV_X1 U4264 ( .A(b_8_), .ZN(n2335) );
  NAND2_X1 U4265 ( .A1(n2334), .A2(n2584), .ZN(n4271) );
  INV_X1 U4266 ( .A(n2326), .ZN(n2334) );
  NAND2_X1 U4267 ( .A1(a_8_), .A2(n2326), .ZN(n4269) );
  NAND2_X1 U4268 ( .A1(n4272), .A2(n4273), .ZN(n2326) );
  NAND2_X1 U4269 ( .A1(n4274), .A2(n2583), .ZN(n4273) );
  INV_X1 U4270 ( .A(b_9_), .ZN(n2583) );
  NAND2_X1 U4271 ( .A1(n2309), .A2(n2310), .ZN(n4274) );
  INV_X1 U4272 ( .A(n2301), .ZN(n2309) );
  NAND2_X1 U4273 ( .A1(a_9_), .A2(n2301), .ZN(n4272) );
  NAND2_X1 U4274 ( .A1(n4275), .A2(n4276), .ZN(n2301) );
  NAND2_X1 U4275 ( .A1(n4277), .A2(n2285), .ZN(n4276) );
  INV_X1 U4276 ( .A(b_10_), .ZN(n2285) );
  NAND2_X1 U4277 ( .A1(n2284), .A2(n2582), .ZN(n4277) );
  INV_X1 U4278 ( .A(n2277), .ZN(n2284) );
  NAND2_X1 U4279 ( .A1(a_10_), .A2(n2277), .ZN(n4275) );
  NAND2_X1 U4280 ( .A1(n4278), .A2(n4279), .ZN(n2277) );
  NAND2_X1 U4281 ( .A1(n4280), .A2(n2580), .ZN(n4279) );
  INV_X1 U4282 ( .A(b_11_), .ZN(n2580) );
  NAND2_X1 U4283 ( .A1(n2250), .A2(n2581), .ZN(n4280) );
  INV_X1 U4284 ( .A(n2258), .ZN(n2250) );
  NAND2_X1 U4285 ( .A1(a_11_), .A2(n2258), .ZN(n4278) );
  NAND2_X1 U4286 ( .A1(n4281), .A2(n4282), .ZN(n2258) );
  NAND2_X1 U4287 ( .A1(n4283), .A2(n2578), .ZN(n4282) );
  INV_X1 U4288 ( .A(b_12_), .ZN(n2578) );
  NAND2_X1 U4289 ( .A1(n2224), .A2(n2579), .ZN(n4283) );
  INV_X1 U4290 ( .A(n2232), .ZN(n2224) );
  NAND2_X1 U4291 ( .A1(a_12_), .A2(n2232), .ZN(n4281) );
  NAND2_X1 U4292 ( .A1(n4284), .A2(n4285), .ZN(n2232) );
  NAND2_X1 U4293 ( .A1(n4286), .A2(n2577), .ZN(n4285) );
  INV_X1 U4294 ( .A(b_13_), .ZN(n2577) );
  NAND2_X1 U4295 ( .A1(n2198), .A2(n2188), .ZN(n4286) );
  INV_X1 U4296 ( .A(n2206), .ZN(n2198) );
  NAND2_X1 U4297 ( .A1(a_13_), .A2(n2206), .ZN(n4284) );
  NAND2_X1 U4298 ( .A1(n4287), .A2(n4288), .ZN(n2206) );
  NAND2_X1 U4299 ( .A1(n4289), .A2(n2161), .ZN(n4288) );
  INV_X1 U4300 ( .A(b_14_), .ZN(n2161) );
  NAND2_X1 U4301 ( .A1(n2150), .A2(n2158), .ZN(n4289) );
  INV_X1 U4302 ( .A(n2145), .ZN(n2150) );
  NAND2_X1 U4303 ( .A1(a_14_), .A2(n2145), .ZN(n4287) );
  NAND2_X1 U4304 ( .A1(b_15_), .A2(n4167), .ZN(n2145) );
  INV_X1 U4305 ( .A(a_15_), .ZN(n4167) );
  NAND3_X1 U4306 ( .A1(n4290), .A2(n4291), .A3(n2094), .ZN(n4243) );
  INV_X1 U4307 ( .A(operation_0_), .ZN(n4241) );
  NAND2_X1 U4308 ( .A1(b_0_), .A2(n4292), .ZN(n4291) );
  NAND2_X1 U4309 ( .A1(n2538), .A2(a_0_), .ZN(n4292) );
  INV_X1 U4310 ( .A(n2530), .ZN(n2538) );
  NAND2_X1 U4311 ( .A1(n2530), .A2(n3102), .ZN(n4290) );
  INV_X1 U4312 ( .A(a_0_), .ZN(n3102) );
  NAND2_X1 U4313 ( .A1(n4293), .A2(n4294), .ZN(n2530) );
  NAND2_X1 U4314 ( .A1(b_1_), .A2(n4295), .ZN(n4294) );
  NAND2_X1 U4315 ( .A1(n2513), .A2(a_1_), .ZN(n4295) );
  INV_X1 U4316 ( .A(n2505), .ZN(n2513) );
  NAND2_X1 U4317 ( .A1(n2505), .A2(n2516), .ZN(n4293) );
  INV_X1 U4318 ( .A(a_1_), .ZN(n2516) );
  NAND2_X1 U4319 ( .A1(n4296), .A2(n4297), .ZN(n2505) );
  NAND2_X1 U4320 ( .A1(b_2_), .A2(n4298), .ZN(n4297) );
  NAND2_X1 U4321 ( .A1(n2489), .A2(a_2_), .ZN(n4298) );
  INV_X1 U4322 ( .A(n2480), .ZN(n2489) );
  NAND2_X1 U4323 ( .A1(n2480), .A2(n2491), .ZN(n4296) );
  INV_X1 U4324 ( .A(a_2_), .ZN(n2491) );
  NAND2_X1 U4325 ( .A1(n4299), .A2(n4300), .ZN(n2480) );
  NAND2_X1 U4326 ( .A1(b_3_), .A2(n4301), .ZN(n4300) );
  NAND2_X1 U4327 ( .A1(n2464), .A2(a_3_), .ZN(n4301) );
  INV_X1 U4328 ( .A(n2455), .ZN(n2464) );
  NAND2_X1 U4329 ( .A1(n2455), .A2(n2466), .ZN(n4299) );
  INV_X1 U4330 ( .A(a_3_), .ZN(n2466) );
  NAND2_X1 U4331 ( .A1(n4302), .A2(n4303), .ZN(n2455) );
  NAND2_X1 U4332 ( .A1(b_4_), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U4333 ( .A1(n2432), .A2(a_4_), .ZN(n4304) );
  INV_X1 U4334 ( .A(n2424), .ZN(n2432) );
  NAND2_X1 U4335 ( .A1(n2424), .A2(n2435), .ZN(n4302) );
  INV_X1 U4336 ( .A(a_4_), .ZN(n2435) );
  NAND2_X1 U4337 ( .A1(n4305), .A2(n4306), .ZN(n2424) );
  NAND2_X1 U4338 ( .A1(b_5_), .A2(n4307), .ZN(n4306) );
  NAND2_X1 U4339 ( .A1(n2408), .A2(a_5_), .ZN(n4307) );
  INV_X1 U4340 ( .A(n2399), .ZN(n2408) );
  NAND2_X1 U4341 ( .A1(n2399), .A2(n2410), .ZN(n4305) );
  INV_X1 U4342 ( .A(a_5_), .ZN(n2410) );
  NAND2_X1 U4343 ( .A1(n4308), .A2(n4309), .ZN(n2399) );
  NAND2_X1 U4344 ( .A1(b_6_), .A2(n4310), .ZN(n4309) );
  NAND2_X1 U4345 ( .A1(n2383), .A2(a_6_), .ZN(n4310) );
  INV_X1 U4346 ( .A(n2374), .ZN(n2383) );
  NAND2_X1 U4347 ( .A1(n2374), .A2(n2586), .ZN(n4308) );
  INV_X1 U4348 ( .A(a_6_), .ZN(n2586) );
  NAND2_X1 U4349 ( .A1(n4311), .A2(n4312), .ZN(n2374) );
  NAND2_X1 U4350 ( .A1(b_7_), .A2(n4313), .ZN(n4312) );
  NAND2_X1 U4351 ( .A1(n2358), .A2(a_7_), .ZN(n4313) );
  INV_X1 U4352 ( .A(n2349), .ZN(n2358) );
  NAND2_X1 U4353 ( .A1(n2349), .A2(n2360), .ZN(n4311) );
  INV_X1 U4354 ( .A(a_7_), .ZN(n2360) );
  NAND2_X1 U4355 ( .A1(n4314), .A2(n4315), .ZN(n2349) );
  NAND2_X1 U4356 ( .A1(b_8_), .A2(n4316), .ZN(n4315) );
  NAND2_X1 U4357 ( .A1(n2332), .A2(a_8_), .ZN(n4316) );
  INV_X1 U4358 ( .A(n2324), .ZN(n2332) );
  NAND2_X1 U4359 ( .A1(n2324), .A2(n2584), .ZN(n4314) );
  INV_X1 U4360 ( .A(a_8_), .ZN(n2584) );
  NAND2_X1 U4361 ( .A1(n4317), .A2(n4318), .ZN(n2324) );
  NAND2_X1 U4362 ( .A1(b_9_), .A2(n4319), .ZN(n4318) );
  NAND2_X1 U4363 ( .A1(n2307), .A2(a_9_), .ZN(n4319) );
  INV_X1 U4364 ( .A(n2299), .ZN(n2307) );
  NAND2_X1 U4365 ( .A1(n2299), .A2(n2310), .ZN(n4317) );
  INV_X1 U4366 ( .A(a_9_), .ZN(n2310) );
  NAND2_X1 U4367 ( .A1(n4320), .A2(n4321), .ZN(n2299) );
  NAND2_X1 U4368 ( .A1(b_10_), .A2(n4322), .ZN(n4321) );
  NAND2_X1 U4369 ( .A1(n2283), .A2(a_10_), .ZN(n4322) );
  INV_X1 U4370 ( .A(n2274), .ZN(n2283) );
  NAND2_X1 U4371 ( .A1(n2274), .A2(n2582), .ZN(n4320) );
  INV_X1 U4372 ( .A(a_10_), .ZN(n2582) );
  NAND2_X1 U4373 ( .A1(n4323), .A2(n4324), .ZN(n2274) );
  NAND2_X1 U4374 ( .A1(b_11_), .A2(n4325), .ZN(n4324) );
  NAND2_X1 U4375 ( .A1(n2248), .A2(a_11_), .ZN(n4325) );
  INV_X1 U4376 ( .A(n2256), .ZN(n2248) );
  NAND2_X1 U4377 ( .A1(n2256), .A2(n2581), .ZN(n4323) );
  INV_X1 U4378 ( .A(a_11_), .ZN(n2581) );
  NAND2_X1 U4379 ( .A1(n4326), .A2(n4327), .ZN(n2256) );
  NAND2_X1 U4380 ( .A1(b_12_), .A2(n4328), .ZN(n4327) );
  NAND2_X1 U4381 ( .A1(n2222), .A2(a_12_), .ZN(n4328) );
  INV_X1 U4382 ( .A(n2230), .ZN(n2222) );
  NAND2_X1 U4383 ( .A1(n2230), .A2(n2579), .ZN(n4326) );
  INV_X1 U4384 ( .A(a_12_), .ZN(n2579) );
  NAND2_X1 U4385 ( .A1(n4329), .A2(n4330), .ZN(n2230) );
  NAND2_X1 U4386 ( .A1(b_13_), .A2(n4331), .ZN(n4330) );
  NAND2_X1 U4387 ( .A1(n2196), .A2(a_13_), .ZN(n4331) );
  INV_X1 U4388 ( .A(n2204), .ZN(n2196) );
  NAND2_X1 U4389 ( .A1(n2204), .A2(n2188), .ZN(n4329) );
  INV_X1 U4390 ( .A(a_13_), .ZN(n2188) );
  NAND2_X1 U4391 ( .A1(n4332), .A2(n4333), .ZN(n2204) );
  NAND2_X1 U4392 ( .A1(b_14_), .A2(n4334), .ZN(n4333) );
  NAND2_X1 U4393 ( .A1(n2167), .A2(a_14_), .ZN(n4334) );
  INV_X1 U4394 ( .A(n2146), .ZN(n2167) );
  NAND2_X1 U4395 ( .A1(n2146), .A2(n2158), .ZN(n4332) );
  INV_X1 U4396 ( .A(a_14_), .ZN(n2158) );
  NAND2_X1 U4397 ( .A1(a_15_), .A2(n2187), .ZN(n2146) );
  INV_X1 U4398 ( .A(b_15_), .ZN(n2187) );
endmodule

