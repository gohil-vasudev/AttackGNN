module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245;

  NOR2_X2 U2143 ( .A1(n4142), .A2(n2415), .ZN(n2416) );
  INV_X2 U2144 ( .A(operation), .ZN(n2112) );
  NOR2_X1 U2145 ( .A1(n2111), .A2(n2112), .ZN(Result_9_) );
  XNOR2_X1 U2146 ( .A(n2113), .B(n2114), .ZN(n2111) );
  NAND2_X1 U2147 ( .A1(n2115), .A2(n2116), .ZN(n2114) );
  NAND2_X1 U2148 ( .A1(n2117), .A2(n2118), .ZN(n2113) );
  NAND2_X1 U2149 ( .A1(n2119), .A2(n2120), .ZN(n2117) );
  NAND2_X1 U2150 ( .A1(n2121), .A2(n2122), .ZN(n2120) );
  NOR2_X1 U2151 ( .A1(n2123), .A2(n2112), .ZN(Result_8_) );
  XNOR2_X1 U2152 ( .A(n2124), .B(n2125), .ZN(n2123) );
  NOR2_X1 U2153 ( .A1(n2126), .A2(n2112), .ZN(Result_7_) );
  XOR2_X1 U2154 ( .A(n2127), .B(n2128), .Z(n2126) );
  NOR2_X1 U2155 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
  NOR2_X1 U2156 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
  NOR2_X1 U2157 ( .A1(n2133), .A2(n2134), .ZN(n2131) );
  NAND2_X1 U2158 ( .A1(n2125), .A2(n2124), .ZN(n2127) );
  NOR2_X1 U2159 ( .A1(n2135), .A2(n2112), .ZN(Result_6_) );
  XNOR2_X1 U2160 ( .A(n2136), .B(n2137), .ZN(n2135) );
  NOR2_X1 U2161 ( .A1(n2138), .A2(n2112), .ZN(Result_5_) );
  XOR2_X1 U2162 ( .A(n2139), .B(n2140), .Z(n2138) );
  NOR2_X1 U2163 ( .A1(n2141), .A2(n2142), .ZN(n2140) );
  NOR2_X1 U2164 ( .A1(n2143), .A2(n2144), .ZN(n2142) );
  NOR2_X1 U2165 ( .A1(n2145), .A2(n2146), .ZN(n2143) );
  NAND2_X1 U2166 ( .A1(n2137), .A2(n2136), .ZN(n2139) );
  NOR2_X1 U2167 ( .A1(n2147), .A2(n2112), .ZN(Result_4_) );
  XNOR2_X1 U2168 ( .A(n2148), .B(n2149), .ZN(n2147) );
  NOR2_X1 U2169 ( .A1(n2150), .A2(n2112), .ZN(Result_3_) );
  XOR2_X1 U2170 ( .A(n2151), .B(n2152), .Z(n2150) );
  NOR2_X1 U2171 ( .A1(n2153), .A2(n2154), .ZN(n2152) );
  NOR2_X1 U2172 ( .A1(n2155), .A2(n2156), .ZN(n2154) );
  NOR2_X1 U2173 ( .A1(n2157), .A2(n2158), .ZN(n2155) );
  NAND2_X1 U2174 ( .A1(n2149), .A2(n2148), .ZN(n2151) );
  NAND2_X1 U2175 ( .A1(n2159), .A2(n2160), .ZN(Result_31_) );
  NAND2_X1 U2176 ( .A1(n2161), .A2(n2112), .ZN(n2160) );
  XNOR2_X1 U2177 ( .A(n2162), .B(a_15_), .ZN(n2161) );
  NAND2_X1 U2178 ( .A1(n2163), .A2(operation), .ZN(n2159) );
  NAND2_X1 U2179 ( .A1(n2164), .A2(n2165), .ZN(Result_30_) );
  NAND2_X1 U2180 ( .A1(operation), .A2(n2166), .ZN(n2165) );
  NAND2_X1 U2181 ( .A1(n2167), .A2(n2168), .ZN(n2166) );
  NAND2_X1 U2182 ( .A1(b_14_), .A2(n2169), .ZN(n2168) );
  NAND2_X1 U2183 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
  NAND2_X1 U2184 ( .A1(a_15_), .A2(n2162), .ZN(n2171) );
  NAND2_X1 U2185 ( .A1(b_15_), .A2(n2172), .ZN(n2167) );
  NAND2_X1 U2186 ( .A1(n2173), .A2(n2174), .ZN(n2172) );
  NAND2_X1 U2187 ( .A1(a_14_), .A2(n2175), .ZN(n2174) );
  NAND2_X1 U2188 ( .A1(n2176), .A2(n2112), .ZN(n2164) );
  XOR2_X1 U2189 ( .A(n2163), .B(n2177), .Z(n2176) );
  XNOR2_X1 U2190 ( .A(n2175), .B(a_14_), .ZN(n2177) );
  INV_X1 U2191 ( .A(n2178), .ZN(n2163) );
  NOR2_X1 U2192 ( .A1(n2112), .A2(n2179), .ZN(Result_2_) );
  XNOR2_X1 U2193 ( .A(n2180), .B(n2181), .ZN(n2179) );
  NAND2_X1 U2194 ( .A1(n2182), .A2(n2183), .ZN(Result_29_) );
  NAND2_X1 U2195 ( .A1(n2184), .A2(n2112), .ZN(n2183) );
  NAND3_X1 U2196 ( .A1(n2185), .A2(n2186), .A3(n2187), .ZN(n2184) );
  NAND2_X1 U2197 ( .A1(n2188), .A2(n2189), .ZN(n2187) );
  NAND3_X1 U2198 ( .A1(n2190), .A2(n2191), .A3(b_13_), .ZN(n2186) );
  NAND2_X1 U2199 ( .A1(n2192), .A2(n2193), .ZN(n2185) );
  XNOR2_X1 U2200 ( .A(a_13_), .B(n2190), .ZN(n2192) );
  INV_X1 U2201 ( .A(n2189), .ZN(n2190) );
  NAND2_X1 U2202 ( .A1(n2194), .A2(operation), .ZN(n2182) );
  XNOR2_X1 U2203 ( .A(n2195), .B(n2196), .ZN(n2194) );
  XOR2_X1 U2204 ( .A(n2197), .B(n2198), .Z(n2196) );
  NAND2_X1 U2205 ( .A1(n2199), .A2(n2200), .ZN(Result_28_) );
  NAND2_X1 U2206 ( .A1(n2201), .A2(n2112), .ZN(n2200) );
  XNOR2_X1 U2207 ( .A(n2202), .B(n2203), .ZN(n2201) );
  NAND2_X1 U2208 ( .A1(n2204), .A2(n2205), .ZN(n2203) );
  NAND2_X1 U2209 ( .A1(n2206), .A2(operation), .ZN(n2199) );
  XOR2_X1 U2210 ( .A(n2207), .B(n2208), .Z(n2206) );
  XOR2_X1 U2211 ( .A(n2209), .B(n2210), .Z(n2207) );
  NOR2_X1 U2212 ( .A1(n2211), .A2(n2162), .ZN(n2210) );
  NAND2_X1 U2213 ( .A1(n2212), .A2(n2213), .ZN(Result_27_) );
  NAND2_X1 U2214 ( .A1(n2214), .A2(n2112), .ZN(n2213) );
  NAND3_X1 U2215 ( .A1(n2215), .A2(n2216), .A3(n2217), .ZN(n2214) );
  INV_X1 U2216 ( .A(n2218), .ZN(n2217) );
  NOR2_X1 U2217 ( .A1(n2219), .A2(n2220), .ZN(n2218) );
  NAND3_X1 U2218 ( .A1(n2220), .A2(n2221), .A3(b_11_), .ZN(n2216) );
  NAND2_X1 U2219 ( .A1(n2222), .A2(n2223), .ZN(n2215) );
  XNOR2_X1 U2220 ( .A(n2220), .B(a_11_), .ZN(n2222) );
  INV_X1 U2221 ( .A(n2224), .ZN(n2220) );
  NAND2_X1 U2222 ( .A1(n2225), .A2(operation), .ZN(n2212) );
  XNOR2_X1 U2223 ( .A(n2226), .B(n2227), .ZN(n2225) );
  XNOR2_X1 U2224 ( .A(n2228), .B(n2229), .ZN(n2226) );
  NAND2_X1 U2225 ( .A1(n2230), .A2(n2231), .ZN(Result_26_) );
  NAND2_X1 U2226 ( .A1(n2232), .A2(n2112), .ZN(n2231) );
  XNOR2_X1 U2227 ( .A(n2233), .B(n2234), .ZN(n2232) );
  NAND2_X1 U2228 ( .A1(n2235), .A2(n2236), .ZN(n2234) );
  NAND2_X1 U2229 ( .A1(n2237), .A2(operation), .ZN(n2230) );
  XNOR2_X1 U2230 ( .A(n2238), .B(n2239), .ZN(n2237) );
  XOR2_X1 U2231 ( .A(n2240), .B(n2241), .Z(n2239) );
  NAND2_X1 U2232 ( .A1(n2242), .A2(n2243), .ZN(Result_25_) );
  NAND2_X1 U2233 ( .A1(n2244), .A2(n2112), .ZN(n2243) );
  NAND3_X1 U2234 ( .A1(n2245), .A2(n2246), .A3(n2247), .ZN(n2244) );
  NAND2_X1 U2235 ( .A1(n2248), .A2(n2249), .ZN(n2247) );
  NAND3_X1 U2236 ( .A1(n2250), .A2(n2251), .A3(b_9_), .ZN(n2246) );
  INV_X1 U2237 ( .A(n2249), .ZN(n2250) );
  NAND2_X1 U2238 ( .A1(n2252), .A2(n2253), .ZN(n2245) );
  XNOR2_X1 U2239 ( .A(n2249), .B(n2251), .ZN(n2252) );
  NAND2_X1 U2240 ( .A1(n2254), .A2(operation), .ZN(n2242) );
  XNOR2_X1 U2241 ( .A(n2255), .B(n2256), .ZN(n2254) );
  XNOR2_X1 U2242 ( .A(n2257), .B(n2258), .ZN(n2255) );
  NAND2_X1 U2243 ( .A1(n2259), .A2(n2260), .ZN(Result_24_) );
  NAND2_X1 U2244 ( .A1(n2261), .A2(n2112), .ZN(n2260) );
  XNOR2_X1 U2245 ( .A(n2262), .B(n2263), .ZN(n2261) );
  NOR2_X1 U2246 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  NAND2_X1 U2247 ( .A1(n2266), .A2(operation), .ZN(n2259) );
  XOR2_X1 U2248 ( .A(n2267), .B(n2268), .Z(n2266) );
  XNOR2_X1 U2249 ( .A(n2269), .B(n2270), .ZN(n2267) );
  NAND2_X1 U2250 ( .A1(n2271), .A2(n2272), .ZN(Result_23_) );
  NAND2_X1 U2251 ( .A1(n2273), .A2(n2112), .ZN(n2272) );
  NAND3_X1 U2252 ( .A1(n2274), .A2(n2275), .A3(n2276), .ZN(n2273) );
  NAND2_X1 U2253 ( .A1(n2277), .A2(n2278), .ZN(n2276) );
  NAND3_X1 U2254 ( .A1(n2279), .A2(n2280), .A3(b_7_), .ZN(n2275) );
  NAND2_X1 U2255 ( .A1(n2281), .A2(n2282), .ZN(n2274) );
  XNOR2_X1 U2256 ( .A(n2279), .B(a_7_), .ZN(n2281) );
  NAND2_X1 U2257 ( .A1(n2283), .A2(operation), .ZN(n2271) );
  XNOR2_X1 U2258 ( .A(n2284), .B(n2285), .ZN(n2283) );
  NAND2_X1 U2259 ( .A1(n2286), .A2(n2287), .ZN(n2284) );
  NAND2_X1 U2260 ( .A1(n2288), .A2(n2289), .ZN(Result_22_) );
  NAND2_X1 U2261 ( .A1(n2290), .A2(n2112), .ZN(n2289) );
  XNOR2_X1 U2262 ( .A(n2291), .B(n2292), .ZN(n2290) );
  NAND2_X1 U2263 ( .A1(n2293), .A2(n2294), .ZN(n2292) );
  NAND2_X1 U2264 ( .A1(n2295), .A2(operation), .ZN(n2288) );
  XNOR2_X1 U2265 ( .A(n2296), .B(n2297), .ZN(n2295) );
  XOR2_X1 U2266 ( .A(n2298), .B(n2299), .Z(n2297) );
  NAND2_X1 U2267 ( .A1(n2300), .A2(n2301), .ZN(Result_21_) );
  NAND2_X1 U2268 ( .A1(n2302), .A2(n2112), .ZN(n2301) );
  NAND3_X1 U2269 ( .A1(n2303), .A2(n2304), .A3(n2305), .ZN(n2302) );
  INV_X1 U2270 ( .A(n2306), .ZN(n2305) );
  NOR2_X1 U2271 ( .A1(n2307), .A2(n2308), .ZN(n2306) );
  NAND3_X1 U2272 ( .A1(n2308), .A2(n2309), .A3(b_5_), .ZN(n2304) );
  NAND2_X1 U2273 ( .A1(n2310), .A2(n2311), .ZN(n2303) );
  XNOR2_X1 U2274 ( .A(n2308), .B(a_5_), .ZN(n2310) );
  INV_X1 U2275 ( .A(n2312), .ZN(n2308) );
  NAND2_X1 U2276 ( .A1(n2313), .A2(operation), .ZN(n2300) );
  XNOR2_X1 U2277 ( .A(n2314), .B(n2315), .ZN(n2313) );
  NAND2_X1 U2278 ( .A1(n2316), .A2(n2317), .ZN(n2314) );
  NAND2_X1 U2279 ( .A1(n2318), .A2(n2319), .ZN(Result_20_) );
  NAND2_X1 U2280 ( .A1(n2320), .A2(n2112), .ZN(n2319) );
  XNOR2_X1 U2281 ( .A(n2321), .B(n2322), .ZN(n2320) );
  NAND2_X1 U2282 ( .A1(n2323), .A2(n2324), .ZN(n2322) );
  NAND2_X1 U2283 ( .A1(n2325), .A2(operation), .ZN(n2318) );
  XOR2_X1 U2284 ( .A(n2326), .B(n2327), .Z(n2325) );
  XOR2_X1 U2285 ( .A(n2328), .B(n2329), .Z(n2327) );
  NOR2_X1 U2286 ( .A1(n2330), .A2(n2112), .ZN(Result_1_) );
  XOR2_X1 U2287 ( .A(n2331), .B(n2332), .Z(n2330) );
  NOR2_X1 U2288 ( .A1(n2333), .A2(n2334), .ZN(n2332) );
  NAND2_X1 U2289 ( .A1(n2335), .A2(n2336), .ZN(Result_19_) );
  NAND2_X1 U2290 ( .A1(n2337), .A2(n2112), .ZN(n2336) );
  NAND3_X1 U2291 ( .A1(n2338), .A2(n2339), .A3(n2340), .ZN(n2337) );
  NAND2_X1 U2292 ( .A1(n2341), .A2(n2342), .ZN(n2340) );
  NAND3_X1 U2293 ( .A1(n2343), .A2(n2344), .A3(b_3_), .ZN(n2339) );
  INV_X1 U2294 ( .A(n2342), .ZN(n2343) );
  NAND2_X1 U2295 ( .A1(n2345), .A2(n2346), .ZN(n2338) );
  XNOR2_X1 U2296 ( .A(n2342), .B(n2344), .ZN(n2345) );
  NAND2_X1 U2297 ( .A1(n2347), .A2(operation), .ZN(n2335) );
  XOR2_X1 U2298 ( .A(n2348), .B(n2349), .Z(n2347) );
  XOR2_X1 U2299 ( .A(n2350), .B(n2351), .Z(n2348) );
  NAND2_X1 U2300 ( .A1(n2352), .A2(n2353), .ZN(Result_18_) );
  NAND2_X1 U2301 ( .A1(n2354), .A2(n2112), .ZN(n2353) );
  XNOR2_X1 U2302 ( .A(n2355), .B(n2356), .ZN(n2354) );
  NAND2_X1 U2303 ( .A1(n2357), .A2(n2358), .ZN(n2356) );
  NAND2_X1 U2304 ( .A1(n2359), .A2(operation), .ZN(n2352) );
  XNOR2_X1 U2305 ( .A(n2360), .B(n2361), .ZN(n2359) );
  XOR2_X1 U2306 ( .A(n2362), .B(n2363), .Z(n2361) );
  NAND2_X1 U2307 ( .A1(b_15_), .A2(a_2_), .ZN(n2363) );
  NAND2_X1 U2308 ( .A1(n2364), .A2(n2365), .ZN(Result_17_) );
  NAND2_X1 U2309 ( .A1(n2366), .A2(n2112), .ZN(n2365) );
  NAND2_X1 U2310 ( .A1(n2367), .A2(n2368), .ZN(n2366) );
  NAND2_X1 U2311 ( .A1(n2369), .A2(n2370), .ZN(n2368) );
  NAND2_X1 U2312 ( .A1(n2371), .A2(n2372), .ZN(n2369) );
  NAND2_X1 U2313 ( .A1(n2373), .A2(n2374), .ZN(n2367) );
  XNOR2_X1 U2314 ( .A(n2375), .B(a_1_), .ZN(n2373) );
  NAND2_X1 U2315 ( .A1(n2376), .A2(operation), .ZN(n2364) );
  XOR2_X1 U2316 ( .A(n2377), .B(n2378), .Z(n2376) );
  XNOR2_X1 U2317 ( .A(n2379), .B(n2380), .ZN(n2378) );
  NAND2_X1 U2318 ( .A1(b_15_), .A2(a_1_), .ZN(n2380) );
  NAND2_X1 U2319 ( .A1(n2381), .A2(n2382), .ZN(Result_16_) );
  NAND2_X1 U2320 ( .A1(n2383), .A2(n2112), .ZN(n2382) );
  XNOR2_X1 U2321 ( .A(n2384), .B(n2385), .ZN(n2383) );
  NOR2_X1 U2322 ( .A1(n2386), .A2(n2387), .ZN(n2385) );
  NOR2_X1 U2323 ( .A1(b_0_), .A2(a_0_), .ZN(n2386) );
  NAND2_X1 U2324 ( .A1(n2372), .A2(n2388), .ZN(n2384) );
  NAND2_X1 U2325 ( .A1(n2371), .A2(n2374), .ZN(n2388) );
  INV_X1 U2326 ( .A(n2370), .ZN(n2374) );
  NAND2_X1 U2327 ( .A1(n2358), .A2(n2389), .ZN(n2370) );
  NAND2_X1 U2328 ( .A1(n2357), .A2(n2355), .ZN(n2389) );
  NAND2_X1 U2329 ( .A1(n2390), .A2(n2391), .ZN(n2355) );
  NAND2_X1 U2330 ( .A1(n2392), .A2(n2342), .ZN(n2391) );
  NAND2_X1 U2331 ( .A1(n2324), .A2(n2393), .ZN(n2342) );
  NAND2_X1 U2332 ( .A1(n2323), .A2(n2321), .ZN(n2393) );
  NAND2_X1 U2333 ( .A1(n2307), .A2(n2394), .ZN(n2321) );
  NAND2_X1 U2334 ( .A1(n2395), .A2(n2312), .ZN(n2394) );
  NAND2_X1 U2335 ( .A1(n2294), .A2(n2396), .ZN(n2312) );
  NAND2_X1 U2336 ( .A1(n2293), .A2(n2291), .ZN(n2396) );
  NAND2_X1 U2337 ( .A1(n2397), .A2(n2398), .ZN(n2291) );
  NAND2_X1 U2338 ( .A1(n2399), .A2(n2278), .ZN(n2398) );
  INV_X1 U2339 ( .A(n2279), .ZN(n2278) );
  NOR2_X1 U2340 ( .A1(n2265), .A2(n2400), .ZN(n2279) );
  NOR2_X1 U2341 ( .A1(n2264), .A2(n2262), .ZN(n2400) );
  INV_X1 U2342 ( .A(n2401), .ZN(n2262) );
  NAND2_X1 U2343 ( .A1(n2402), .A2(n2403), .ZN(n2401) );
  NAND2_X1 U2344 ( .A1(n2404), .A2(n2249), .ZN(n2403) );
  NAND2_X1 U2345 ( .A1(n2236), .A2(n2405), .ZN(n2249) );
  NAND2_X1 U2346 ( .A1(n2235), .A2(n2233), .ZN(n2405) );
  NAND2_X1 U2347 ( .A1(n2219), .A2(n2406), .ZN(n2233) );
  NAND2_X1 U2348 ( .A1(n2407), .A2(n2224), .ZN(n2406) );
  NAND2_X1 U2349 ( .A1(n2205), .A2(n2408), .ZN(n2224) );
  NAND2_X1 U2350 ( .A1(n2204), .A2(n2202), .ZN(n2408) );
  NAND2_X1 U2351 ( .A1(n2409), .A2(n2410), .ZN(n2202) );
  NAND2_X1 U2352 ( .A1(n2411), .A2(n2189), .ZN(n2410) );
  NAND2_X1 U2353 ( .A1(n2412), .A2(n2413), .ZN(n2189) );
  NAND2_X1 U2354 ( .A1(b_14_), .A2(n2414), .ZN(n2413) );
  NAND2_X1 U2355 ( .A1(n2415), .A2(n2178), .ZN(n2414) );
  NAND2_X1 U2356 ( .A1(b_15_), .A2(a_15_), .ZN(n2178) );
  NAND2_X1 U2357 ( .A1(b_15_), .A2(n2416), .ZN(n2412) );
  NAND2_X1 U2358 ( .A1(n2193), .A2(n2191), .ZN(n2411) );
  NAND2_X1 U2359 ( .A1(n2417), .A2(n2211), .ZN(n2204) );
  NAND2_X1 U2360 ( .A1(n2223), .A2(n2221), .ZN(n2407) );
  NAND2_X1 U2361 ( .A1(n2418), .A2(n2419), .ZN(n2235) );
  INV_X1 U2362 ( .A(n2420), .ZN(n2236) );
  NAND2_X1 U2363 ( .A1(n2253), .A2(n2251), .ZN(n2404) );
  NOR2_X1 U2364 ( .A1(b_8_), .A2(a_8_), .ZN(n2264) );
  NAND2_X1 U2365 ( .A1(n2282), .A2(n2280), .ZN(n2399) );
  NAND2_X1 U2366 ( .A1(n2421), .A2(n2422), .ZN(n2293) );
  NAND2_X1 U2367 ( .A1(n2311), .A2(n2309), .ZN(n2395) );
  NAND2_X1 U2368 ( .A1(n2423), .A2(n2424), .ZN(n2323) );
  NAND2_X1 U2369 ( .A1(n2346), .A2(n2344), .ZN(n2392) );
  NAND2_X1 U2370 ( .A1(n2425), .A2(n2426), .ZN(n2357) );
  NAND2_X1 U2371 ( .A1(n2375), .A2(n2427), .ZN(n2372) );
  NAND2_X1 U2372 ( .A1(n2428), .A2(operation), .ZN(n2381) );
  XNOR2_X1 U2373 ( .A(n2429), .B(n2430), .ZN(n2428) );
  XNOR2_X1 U2374 ( .A(n2431), .B(n2432), .ZN(n2429) );
  NOR2_X1 U2375 ( .A1(n2433), .A2(n2162), .ZN(n2432) );
  NOR2_X1 U2376 ( .A1(n2434), .A2(n2112), .ZN(Result_15_) );
  XNOR2_X1 U2377 ( .A(n2435), .B(n2436), .ZN(n2434) );
  NOR3_X1 U2378 ( .A1(n2112), .A2(n2437), .A3(n2438), .ZN(Result_14_) );
  NOR2_X1 U2379 ( .A1(n2439), .A2(n2440), .ZN(n2438) );
  XOR2_X1 U2380 ( .A(n2441), .B(n2442), .Z(n2440) );
  NOR2_X1 U2381 ( .A1(n2435), .A2(n2436), .ZN(n2439) );
  NOR2_X1 U2382 ( .A1(n2443), .A2(n2112), .ZN(Result_13_) );
  XNOR2_X1 U2383 ( .A(n2437), .B(n2444), .ZN(n2443) );
  NOR2_X1 U2384 ( .A1(n2445), .A2(n2446), .ZN(n2444) );
  NOR2_X1 U2385 ( .A1(n2447), .A2(n2448), .ZN(n2446) );
  NOR2_X1 U2386 ( .A1(n2112), .A2(n2449), .ZN(Result_12_) );
  XNOR2_X1 U2387 ( .A(n2450), .B(n2451), .ZN(n2449) );
  NOR2_X1 U2388 ( .A1(n2452), .A2(n2112), .ZN(Result_11_) );
  XNOR2_X1 U2389 ( .A(n2453), .B(n2454), .ZN(n2452) );
  NAND2_X1 U2390 ( .A1(n2450), .A2(n2451), .ZN(n2454) );
  NAND2_X1 U2391 ( .A1(n2455), .A2(n2456), .ZN(n2453) );
  NAND2_X1 U2392 ( .A1(n2457), .A2(n2458), .ZN(n2455) );
  NAND2_X1 U2393 ( .A1(n2459), .A2(n2460), .ZN(n2458) );
  NOR2_X1 U2394 ( .A1(n2461), .A2(n2112), .ZN(Result_10_) );
  XNOR2_X1 U2395 ( .A(n2116), .B(n2115), .ZN(n2461) );
  NOR2_X1 U2396 ( .A1(n2462), .A2(n2112), .ZN(Result_0_) );
  NOR3_X1 U2397 ( .A1(n2463), .A2(n2333), .A3(n2464), .ZN(n2462) );
  NOR2_X1 U2398 ( .A1(n2334), .A2(n2331), .ZN(n2464) );
  NAND2_X1 U2399 ( .A1(n2181), .A2(n2180), .ZN(n2331) );
  NAND3_X1 U2400 ( .A1(n2465), .A2(n2466), .A3(n2467), .ZN(n2180) );
  NAND3_X1 U2401 ( .A1(n2149), .A2(n2148), .A3(n2156), .ZN(n2467) );
  INV_X1 U2402 ( .A(n2468), .ZN(n2156) );
  NAND3_X1 U2403 ( .A1(n2469), .A2(n2470), .A3(n2471), .ZN(n2148) );
  NAND3_X1 U2404 ( .A1(n2137), .A2(n2136), .A3(n2144), .ZN(n2471) );
  INV_X1 U2405 ( .A(n2472), .ZN(n2144) );
  NAND3_X1 U2406 ( .A1(n2473), .A2(n2474), .A3(n2475), .ZN(n2136) );
  NAND3_X1 U2407 ( .A1(n2125), .A2(n2124), .A3(n2132), .ZN(n2475) );
  INV_X1 U2408 ( .A(n2476), .ZN(n2132) );
  NAND3_X1 U2409 ( .A1(n2477), .A2(n2118), .A3(n2478), .ZN(n2124) );
  NAND3_X1 U2410 ( .A1(n2479), .A2(n2115), .A3(n2116), .ZN(n2478) );
  XOR2_X1 U2411 ( .A(n2121), .B(n2122), .Z(n2116) );
  NAND3_X1 U2412 ( .A1(n2480), .A2(n2456), .A3(n2481), .ZN(n2115) );
  NAND2_X1 U2413 ( .A1(n2482), .A2(n2483), .ZN(n2481) );
  NAND3_X1 U2414 ( .A1(n2459), .A2(n2460), .A3(n2484), .ZN(n2456) );
  NAND3_X1 U2415 ( .A1(n2451), .A2(n2450), .A3(n2484), .ZN(n2480) );
  INV_X1 U2416 ( .A(n2457), .ZN(n2484) );
  XNOR2_X1 U2417 ( .A(n2483), .B(n2482), .ZN(n2457) );
  XNOR2_X1 U2418 ( .A(n2485), .B(n2486), .ZN(n2482) );
  XNOR2_X1 U2419 ( .A(n2487), .B(n2488), .ZN(n2485) );
  NAND2_X1 U2420 ( .A1(n2489), .A2(n2490), .ZN(n2483) );
  NAND2_X1 U2421 ( .A1(n2491), .A2(n2492), .ZN(n2490) );
  NAND2_X1 U2422 ( .A1(n2493), .A2(n2494), .ZN(n2492) );
  INV_X1 U2423 ( .A(n2495), .ZN(n2489) );
  NOR2_X1 U2424 ( .A1(n2494), .A2(n2493), .ZN(n2495) );
  NAND3_X1 U2425 ( .A1(n2496), .A2(n2497), .A3(n2498), .ZN(n2450) );
  NAND2_X1 U2426 ( .A1(n2437), .A2(n2448), .ZN(n2498) );
  INV_X1 U2427 ( .A(n2499), .ZN(n2448) );
  NOR4_X1 U2428 ( .A1(n2436), .A2(n2500), .A3(n2435), .A4(n2447), .ZN(n2437)
         );
  INV_X1 U2429 ( .A(n2501), .ZN(n2447) );
  NOR2_X1 U2430 ( .A1(n2502), .A2(n2503), .ZN(n2435) );
  NOR3_X1 U2431 ( .A1(n2433), .A2(n2504), .A3(n2162), .ZN(n2503) );
  INV_X1 U2432 ( .A(n2505), .ZN(n2504) );
  NAND2_X1 U2433 ( .A1(n2431), .A2(n2430), .ZN(n2505) );
  NOR2_X1 U2434 ( .A1(n2430), .A2(n2431), .ZN(n2502) );
  NOR2_X1 U2435 ( .A1(n2506), .A2(n2507), .ZN(n2431) );
  INV_X1 U2436 ( .A(n2508), .ZN(n2507) );
  NAND3_X1 U2437 ( .A1(a_1_), .A2(n2509), .A3(b_15_), .ZN(n2508) );
  NAND2_X1 U2438 ( .A1(n2379), .A2(n2377), .ZN(n2509) );
  NOR2_X1 U2439 ( .A1(n2377), .A2(n2379), .ZN(n2506) );
  NOR2_X1 U2440 ( .A1(n2510), .A2(n2511), .ZN(n2379) );
  NOR3_X1 U2441 ( .A1(n2426), .A2(n2512), .A3(n2162), .ZN(n2511) );
  NOR2_X1 U2442 ( .A1(n2362), .A2(n2360), .ZN(n2512) );
  INV_X1 U2443 ( .A(n2513), .ZN(n2510) );
  NAND2_X1 U2444 ( .A1(n2360), .A2(n2362), .ZN(n2513) );
  NAND2_X1 U2445 ( .A1(n2514), .A2(n2515), .ZN(n2362) );
  NAND2_X1 U2446 ( .A1(n2351), .A2(n2516), .ZN(n2515) );
  INV_X1 U2447 ( .A(n2517), .ZN(n2516) );
  NOR2_X1 U2448 ( .A1(n2350), .A2(n2349), .ZN(n2517) );
  NOR2_X1 U2449 ( .A1(n2162), .A2(n2344), .ZN(n2351) );
  NAND2_X1 U2450 ( .A1(n2349), .A2(n2350), .ZN(n2514) );
  NAND2_X1 U2451 ( .A1(n2518), .A2(n2519), .ZN(n2350) );
  NAND2_X1 U2452 ( .A1(n2329), .A2(n2520), .ZN(n2519) );
  INV_X1 U2453 ( .A(n2521), .ZN(n2520) );
  NOR2_X1 U2454 ( .A1(n2328), .A2(n2326), .ZN(n2521) );
  NOR2_X1 U2455 ( .A1(n2162), .A2(n2424), .ZN(n2329) );
  NAND2_X1 U2456 ( .A1(n2326), .A2(n2328), .ZN(n2518) );
  NAND2_X1 U2457 ( .A1(n2316), .A2(n2522), .ZN(n2328) );
  NAND2_X1 U2458 ( .A1(n2315), .A2(n2317), .ZN(n2522) );
  NAND2_X1 U2459 ( .A1(n2523), .A2(n2524), .ZN(n2317) );
  NAND2_X1 U2460 ( .A1(b_15_), .A2(a_5_), .ZN(n2523) );
  XNOR2_X1 U2461 ( .A(n2525), .B(n2526), .ZN(n2315) );
  XNOR2_X1 U2462 ( .A(n2527), .B(n2528), .ZN(n2525) );
  NOR2_X1 U2463 ( .A1(n2422), .A2(n2175), .ZN(n2528) );
  NAND2_X1 U2464 ( .A1(n2529), .A2(a_5_), .ZN(n2316) );
  INV_X1 U2465 ( .A(n2524), .ZN(n2529) );
  NAND2_X1 U2466 ( .A1(n2530), .A2(n2531), .ZN(n2524) );
  NAND2_X1 U2467 ( .A1(n2532), .A2(n2298), .ZN(n2531) );
  NAND2_X1 U2468 ( .A1(b_15_), .A2(a_6_), .ZN(n2298) );
  NAND2_X1 U2469 ( .A1(n2296), .A2(n2299), .ZN(n2532) );
  INV_X1 U2470 ( .A(n2533), .ZN(n2530) );
  NOR2_X1 U2471 ( .A1(n2299), .A2(n2296), .ZN(n2533) );
  XOR2_X1 U2472 ( .A(n2534), .B(n2535), .Z(n2296) );
  XNOR2_X1 U2473 ( .A(n2536), .B(n2537), .ZN(n2535) );
  NAND2_X1 U2474 ( .A1(b_14_), .A2(a_7_), .ZN(n2537) );
  NAND2_X1 U2475 ( .A1(n2286), .A2(n2538), .ZN(n2299) );
  NAND2_X1 U2476 ( .A1(n2285), .A2(n2287), .ZN(n2538) );
  NAND2_X1 U2477 ( .A1(n2539), .A2(n2540), .ZN(n2287) );
  NAND2_X1 U2478 ( .A1(b_15_), .A2(a_7_), .ZN(n2539) );
  XNOR2_X1 U2479 ( .A(n2541), .B(n2542), .ZN(n2285) );
  XOR2_X1 U2480 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND2_X1 U2481 ( .A1(b_14_), .A2(a_8_), .ZN(n2544) );
  NAND2_X1 U2482 ( .A1(n2545), .A2(a_7_), .ZN(n2286) );
  INV_X1 U2483 ( .A(n2540), .ZN(n2545) );
  NAND2_X1 U2484 ( .A1(n2546), .A2(n2547), .ZN(n2540) );
  NAND2_X1 U2485 ( .A1(n2548), .A2(n2270), .ZN(n2547) );
  NAND2_X1 U2486 ( .A1(b_15_), .A2(a_8_), .ZN(n2270) );
  NAND2_X1 U2487 ( .A1(n2268), .A2(n2269), .ZN(n2548) );
  INV_X1 U2488 ( .A(n2549), .ZN(n2546) );
  NOR2_X1 U2489 ( .A1(n2269), .A2(n2268), .ZN(n2549) );
  XNOR2_X1 U2490 ( .A(n2550), .B(n2551), .ZN(n2268) );
  NAND2_X1 U2491 ( .A1(n2552), .A2(n2553), .ZN(n2550) );
  NAND2_X1 U2492 ( .A1(n2554), .A2(n2555), .ZN(n2269) );
  NAND2_X1 U2493 ( .A1(n2258), .A2(n2556), .ZN(n2555) );
  NAND2_X1 U2494 ( .A1(n2257), .A2(n2256), .ZN(n2556) );
  NOR2_X1 U2495 ( .A1(n2162), .A2(n2251), .ZN(n2258) );
  INV_X1 U2496 ( .A(n2557), .ZN(n2554) );
  NOR2_X1 U2497 ( .A1(n2256), .A2(n2257), .ZN(n2557) );
  NOR2_X1 U2498 ( .A1(n2558), .A2(n2559), .ZN(n2257) );
  NOR2_X1 U2499 ( .A1(n2240), .A2(n2560), .ZN(n2559) );
  NOR2_X1 U2500 ( .A1(n2241), .A2(n2238), .ZN(n2560) );
  NAND2_X1 U2501 ( .A1(b_15_), .A2(a_10_), .ZN(n2240) );
  INV_X1 U2502 ( .A(n2561), .ZN(n2558) );
  NAND2_X1 U2503 ( .A1(n2238), .A2(n2241), .ZN(n2561) );
  NAND2_X1 U2504 ( .A1(n2562), .A2(n2563), .ZN(n2241) );
  NAND2_X1 U2505 ( .A1(n2229), .A2(n2564), .ZN(n2563) );
  NAND2_X1 U2506 ( .A1(n2228), .A2(n2227), .ZN(n2564) );
  NOR2_X1 U2507 ( .A1(n2162), .A2(n2221), .ZN(n2229) );
  INV_X1 U2508 ( .A(n2565), .ZN(n2562) );
  NOR2_X1 U2509 ( .A1(n2227), .A2(n2228), .ZN(n2565) );
  NOR2_X1 U2510 ( .A1(n2566), .A2(n2567), .ZN(n2228) );
  NOR3_X1 U2511 ( .A1(n2211), .A2(n2568), .A3(n2162), .ZN(n2567) );
  INV_X1 U2512 ( .A(b_15_), .ZN(n2162) );
  INV_X1 U2513 ( .A(n2569), .ZN(n2568) );
  NAND2_X1 U2514 ( .A1(n2208), .A2(n2209), .ZN(n2569) );
  NOR2_X1 U2515 ( .A1(n2209), .A2(n2208), .ZN(n2566) );
  XNOR2_X1 U2516 ( .A(n2570), .B(n2571), .ZN(n2208) );
  XNOR2_X1 U2517 ( .A(n2572), .B(n2573), .ZN(n2570) );
  NAND2_X1 U2518 ( .A1(n2574), .A2(n2575), .ZN(n2209) );
  NAND2_X1 U2519 ( .A1(n2576), .A2(n2197), .ZN(n2575) );
  NAND2_X1 U2520 ( .A1(b_15_), .A2(a_13_), .ZN(n2197) );
  NAND2_X1 U2521 ( .A1(n2195), .A2(n2198), .ZN(n2576) );
  INV_X1 U2522 ( .A(n2577), .ZN(n2574) );
  NOR2_X1 U2523 ( .A1(n2198), .A2(n2195), .ZN(n2577) );
  INV_X1 U2524 ( .A(n2578), .ZN(n2195) );
  NAND3_X1 U2525 ( .A1(b_14_), .A2(n2416), .A3(b_15_), .ZN(n2578) );
  NAND2_X1 U2526 ( .A1(n2579), .A2(n2580), .ZN(n2198) );
  NAND2_X1 U2527 ( .A1(b_13_), .A2(n2581), .ZN(n2580) );
  NAND2_X1 U2528 ( .A1(n2170), .A2(n2582), .ZN(n2581) );
  NAND2_X1 U2529 ( .A1(a_15_), .A2(n2175), .ZN(n2582) );
  NAND2_X1 U2530 ( .A1(b_14_), .A2(n2583), .ZN(n2579) );
  NAND2_X1 U2531 ( .A1(n2173), .A2(n2584), .ZN(n2583) );
  NAND2_X1 U2532 ( .A1(a_14_), .A2(n2193), .ZN(n2584) );
  XOR2_X1 U2533 ( .A(n2585), .B(n2586), .Z(n2227) );
  XNOR2_X1 U2534 ( .A(n2587), .B(n2588), .ZN(n2585) );
  XNOR2_X1 U2535 ( .A(n2589), .B(n2590), .ZN(n2238) );
  XOR2_X1 U2536 ( .A(n2591), .B(n2592), .Z(n2589) );
  NAND2_X1 U2537 ( .A1(b_14_), .A2(a_11_), .ZN(n2591) );
  XNOR2_X1 U2538 ( .A(n2593), .B(n2594), .ZN(n2256) );
  XNOR2_X1 U2539 ( .A(n2595), .B(n2596), .ZN(n2594) );
  XNOR2_X1 U2540 ( .A(n2597), .B(n2598), .ZN(n2326) );
  NAND2_X1 U2541 ( .A1(n2599), .A2(n2600), .ZN(n2597) );
  XOR2_X1 U2542 ( .A(n2601), .B(n2602), .Z(n2349) );
  XOR2_X1 U2543 ( .A(n2603), .B(n2604), .Z(n2601) );
  NOR2_X1 U2544 ( .A1(n2424), .A2(n2175), .ZN(n2604) );
  XNOR2_X1 U2545 ( .A(n2605), .B(n2606), .ZN(n2360) );
  XNOR2_X1 U2546 ( .A(n2607), .B(n2608), .ZN(n2605) );
  NOR2_X1 U2547 ( .A1(n2344), .A2(n2175), .ZN(n2608) );
  XNOR2_X1 U2548 ( .A(n2609), .B(n2610), .ZN(n2377) );
  XNOR2_X1 U2549 ( .A(n2611), .B(n2612), .ZN(n2610) );
  NAND2_X1 U2550 ( .A1(b_14_), .A2(a_2_), .ZN(n2612) );
  XOR2_X1 U2551 ( .A(n2613), .B(n2614), .Z(n2430) );
  NAND2_X1 U2552 ( .A1(n2615), .A2(n2616), .ZN(n2613) );
  NOR2_X1 U2553 ( .A1(n2441), .A2(n2442), .ZN(n2500) );
  XNOR2_X1 U2554 ( .A(n2617), .B(n2618), .ZN(n2436) );
  XNOR2_X1 U2555 ( .A(n2619), .B(n2620), .ZN(n2617) );
  NAND2_X1 U2556 ( .A1(b_14_), .A2(a_0_), .ZN(n2619) );
  INV_X1 U2557 ( .A(n2445), .ZN(n2497) );
  NOR2_X1 U2558 ( .A1(n2499), .A2(n2501), .ZN(n2445) );
  NAND2_X1 U2559 ( .A1(n2442), .A2(n2441), .ZN(n2501) );
  NAND2_X1 U2560 ( .A1(n2621), .A2(n2622), .ZN(n2441) );
  INV_X1 U2561 ( .A(n2623), .ZN(n2622) );
  NOR3_X1 U2562 ( .A1(n2433), .A2(n2624), .A3(n2175), .ZN(n2623) );
  NOR2_X1 U2563 ( .A1(n2620), .A2(n2618), .ZN(n2624) );
  NAND2_X1 U2564 ( .A1(n2618), .A2(n2620), .ZN(n2621) );
  NAND2_X1 U2565 ( .A1(n2615), .A2(n2625), .ZN(n2620) );
  NAND2_X1 U2566 ( .A1(n2614), .A2(n2616), .ZN(n2625) );
  NAND2_X1 U2567 ( .A1(n2626), .A2(n2627), .ZN(n2616) );
  NAND2_X1 U2568 ( .A1(b_14_), .A2(a_1_), .ZN(n2627) );
  INV_X1 U2569 ( .A(n2628), .ZN(n2626) );
  XOR2_X1 U2570 ( .A(n2629), .B(n2630), .Z(n2614) );
  XNOR2_X1 U2571 ( .A(n2631), .B(n2632), .ZN(n2630) );
  NAND2_X1 U2572 ( .A1(b_13_), .A2(a_2_), .ZN(n2632) );
  NAND2_X1 U2573 ( .A1(a_1_), .A2(n2628), .ZN(n2615) );
  NAND2_X1 U2574 ( .A1(n2633), .A2(n2634), .ZN(n2628) );
  NAND3_X1 U2575 ( .A1(a_2_), .A2(n2635), .A3(b_14_), .ZN(n2634) );
  NAND2_X1 U2576 ( .A1(n2611), .A2(n2609), .ZN(n2635) );
  INV_X1 U2577 ( .A(n2636), .ZN(n2633) );
  NOR2_X1 U2578 ( .A1(n2609), .A2(n2611), .ZN(n2636) );
  NOR2_X1 U2579 ( .A1(n2637), .A2(n2638), .ZN(n2611) );
  INV_X1 U2580 ( .A(n2639), .ZN(n2638) );
  NAND3_X1 U2581 ( .A1(a_3_), .A2(n2640), .A3(b_14_), .ZN(n2639) );
  NAND2_X1 U2582 ( .A1(n2607), .A2(n2606), .ZN(n2640) );
  NOR2_X1 U2583 ( .A1(n2606), .A2(n2607), .ZN(n2637) );
  NOR2_X1 U2584 ( .A1(n2641), .A2(n2642), .ZN(n2607) );
  NOR3_X1 U2585 ( .A1(n2424), .A2(n2643), .A3(n2175), .ZN(n2642) );
  NOR2_X1 U2586 ( .A1(n2603), .A2(n2602), .ZN(n2643) );
  INV_X1 U2587 ( .A(n2644), .ZN(n2641) );
  NAND2_X1 U2588 ( .A1(n2602), .A2(n2603), .ZN(n2644) );
  NAND2_X1 U2589 ( .A1(n2599), .A2(n2645), .ZN(n2603) );
  NAND2_X1 U2590 ( .A1(n2598), .A2(n2600), .ZN(n2645) );
  NAND2_X1 U2591 ( .A1(n2646), .A2(n2647), .ZN(n2600) );
  NAND2_X1 U2592 ( .A1(b_14_), .A2(a_5_), .ZN(n2647) );
  INV_X1 U2593 ( .A(n2648), .ZN(n2646) );
  XNOR2_X1 U2594 ( .A(n2649), .B(n2650), .ZN(n2598) );
  XOR2_X1 U2595 ( .A(n2651), .B(n2652), .Z(n2650) );
  NAND2_X1 U2596 ( .A1(b_13_), .A2(a_6_), .ZN(n2652) );
  NAND2_X1 U2597 ( .A1(a_5_), .A2(n2648), .ZN(n2599) );
  NAND2_X1 U2598 ( .A1(n2653), .A2(n2654), .ZN(n2648) );
  NAND3_X1 U2599 ( .A1(a_6_), .A2(n2655), .A3(b_14_), .ZN(n2654) );
  NAND2_X1 U2600 ( .A1(n2527), .A2(n2526), .ZN(n2655) );
  INV_X1 U2601 ( .A(n2656), .ZN(n2653) );
  NOR2_X1 U2602 ( .A1(n2526), .A2(n2527), .ZN(n2656) );
  NOR2_X1 U2603 ( .A1(n2657), .A2(n2658), .ZN(n2527) );
  NOR3_X1 U2604 ( .A1(n2280), .A2(n2659), .A3(n2175), .ZN(n2658) );
  INV_X1 U2605 ( .A(n2660), .ZN(n2659) );
  NAND2_X1 U2606 ( .A1(n2536), .A2(n2534), .ZN(n2660) );
  NOR2_X1 U2607 ( .A1(n2534), .A2(n2536), .ZN(n2657) );
  NOR2_X1 U2608 ( .A1(n2661), .A2(n2662), .ZN(n2536) );
  NOR3_X1 U2609 ( .A1(n2663), .A2(n2664), .A3(n2175), .ZN(n2662) );
  NOR2_X1 U2610 ( .A1(n2543), .A2(n2541), .ZN(n2664) );
  INV_X1 U2611 ( .A(n2665), .ZN(n2661) );
  NAND2_X1 U2612 ( .A1(n2541), .A2(n2543), .ZN(n2665) );
  NAND2_X1 U2613 ( .A1(n2552), .A2(n2666), .ZN(n2543) );
  NAND2_X1 U2614 ( .A1(n2551), .A2(n2553), .ZN(n2666) );
  NAND2_X1 U2615 ( .A1(n2667), .A2(n2668), .ZN(n2553) );
  NAND2_X1 U2616 ( .A1(b_14_), .A2(a_9_), .ZN(n2667) );
  XNOR2_X1 U2617 ( .A(n2669), .B(n2670), .ZN(n2551) );
  NAND2_X1 U2618 ( .A1(n2671), .A2(n2672), .ZN(n2669) );
  INV_X1 U2619 ( .A(n2673), .ZN(n2552) );
  NOR2_X1 U2620 ( .A1(n2668), .A2(n2251), .ZN(n2673) );
  NAND2_X1 U2621 ( .A1(n2674), .A2(n2675), .ZN(n2668) );
  NAND2_X1 U2622 ( .A1(n2593), .A2(n2676), .ZN(n2675) );
  INV_X1 U2623 ( .A(n2677), .ZN(n2676) );
  NOR2_X1 U2624 ( .A1(n2596), .A2(n2595), .ZN(n2677) );
  XOR2_X1 U2625 ( .A(n2678), .B(n2679), .Z(n2593) );
  XNOR2_X1 U2626 ( .A(n2680), .B(n2681), .ZN(n2678) );
  NOR2_X1 U2627 ( .A1(n2221), .A2(n2193), .ZN(n2681) );
  NAND2_X1 U2628 ( .A1(n2595), .A2(n2596), .ZN(n2674) );
  NAND2_X1 U2629 ( .A1(b_14_), .A2(a_10_), .ZN(n2596) );
  NOR2_X1 U2630 ( .A1(n2682), .A2(n2683), .ZN(n2595) );
  INV_X1 U2631 ( .A(n2684), .ZN(n2683) );
  NAND3_X1 U2632 ( .A1(a_11_), .A2(n2685), .A3(b_14_), .ZN(n2684) );
  NAND2_X1 U2633 ( .A1(n2592), .A2(n2590), .ZN(n2685) );
  NOR2_X1 U2634 ( .A1(n2590), .A2(n2592), .ZN(n2682) );
  NOR2_X1 U2635 ( .A1(n2686), .A2(n2687), .ZN(n2592) );
  INV_X1 U2636 ( .A(n2688), .ZN(n2687) );
  NAND2_X1 U2637 ( .A1(n2587), .A2(n2689), .ZN(n2688) );
  NAND2_X1 U2638 ( .A1(n2588), .A2(n2586), .ZN(n2689) );
  NOR2_X1 U2639 ( .A1(n2175), .A2(n2211), .ZN(n2587) );
  NOR2_X1 U2640 ( .A1(n2586), .A2(n2588), .ZN(n2686) );
  NOR2_X1 U2641 ( .A1(n2690), .A2(n2691), .ZN(n2588) );
  INV_X1 U2642 ( .A(n2692), .ZN(n2691) );
  NAND2_X1 U2643 ( .A1(n2571), .A2(n2693), .ZN(n2692) );
  NAND2_X1 U2644 ( .A1(n2694), .A2(n2573), .ZN(n2693) );
  NOR2_X1 U2645 ( .A1(n2175), .A2(n2191), .ZN(n2571) );
  INV_X1 U2646 ( .A(b_14_), .ZN(n2175) );
  NOR2_X1 U2647 ( .A1(n2573), .A2(n2694), .ZN(n2690) );
  INV_X1 U2648 ( .A(n2572), .ZN(n2694) );
  NAND2_X1 U2649 ( .A1(n2695), .A2(n2696), .ZN(n2572) );
  NAND2_X1 U2650 ( .A1(b_12_), .A2(n2697), .ZN(n2696) );
  NAND2_X1 U2651 ( .A1(n2170), .A2(n2698), .ZN(n2697) );
  NAND2_X1 U2652 ( .A1(a_15_), .A2(n2193), .ZN(n2698) );
  NAND2_X1 U2653 ( .A1(b_13_), .A2(n2699), .ZN(n2695) );
  NAND2_X1 U2654 ( .A1(n2173), .A2(n2700), .ZN(n2699) );
  NAND2_X1 U2655 ( .A1(a_14_), .A2(n2417), .ZN(n2700) );
  NAND3_X1 U2656 ( .A1(b_13_), .A2(n2416), .A3(b_14_), .ZN(n2573) );
  XOR2_X1 U2657 ( .A(n2701), .B(n2409), .Z(n2586) );
  XOR2_X1 U2658 ( .A(n2702), .B(n2703), .Z(n2701) );
  XNOR2_X1 U2659 ( .A(n2704), .B(n2705), .ZN(n2590) );
  XOR2_X1 U2660 ( .A(n2706), .B(n2707), .Z(n2704) );
  XNOR2_X1 U2661 ( .A(n2708), .B(n2709), .ZN(n2541) );
  NAND2_X1 U2662 ( .A1(n2710), .A2(n2711), .ZN(n2708) );
  XOR2_X1 U2663 ( .A(n2712), .B(n2713), .Z(n2534) );
  XOR2_X1 U2664 ( .A(n2714), .B(n2715), .Z(n2713) );
  NAND2_X1 U2665 ( .A1(b_13_), .A2(a_8_), .ZN(n2715) );
  XNOR2_X1 U2666 ( .A(n2716), .B(n2717), .ZN(n2526) );
  XNOR2_X1 U2667 ( .A(n2718), .B(n2719), .ZN(n2717) );
  NAND2_X1 U2668 ( .A1(b_13_), .A2(a_7_), .ZN(n2719) );
  XNOR2_X1 U2669 ( .A(n2720), .B(n2721), .ZN(n2602) );
  NAND2_X1 U2670 ( .A1(n2722), .A2(n2723), .ZN(n2720) );
  XNOR2_X1 U2671 ( .A(n2724), .B(n2725), .ZN(n2606) );
  XOR2_X1 U2672 ( .A(n2726), .B(n2727), .Z(n2724) );
  NOR2_X1 U2673 ( .A1(n2424), .A2(n2193), .ZN(n2727) );
  XOR2_X1 U2674 ( .A(n2728), .B(n2729), .Z(n2609) );
  XNOR2_X1 U2675 ( .A(n2730), .B(n2731), .ZN(n2728) );
  NOR2_X1 U2676 ( .A1(n2344), .A2(n2193), .ZN(n2731) );
  XNOR2_X1 U2677 ( .A(n2732), .B(n2733), .ZN(n2618) );
  NAND2_X1 U2678 ( .A1(n2734), .A2(n2735), .ZN(n2732) );
  XNOR2_X1 U2679 ( .A(n2736), .B(n2737), .ZN(n2442) );
  NAND2_X1 U2680 ( .A1(n2738), .A2(n2739), .ZN(n2736) );
  NAND2_X1 U2681 ( .A1(n2740), .A2(n2496), .ZN(n2499) );
  NAND2_X1 U2682 ( .A1(n2741), .A2(n2742), .ZN(n2740) );
  XNOR2_X1 U2683 ( .A(n2743), .B(n2744), .ZN(n2742) );
  INV_X1 U2684 ( .A(n2745), .ZN(n2741) );
  NAND2_X1 U2685 ( .A1(n2746), .A2(n2745), .ZN(n2496) );
  NAND2_X1 U2686 ( .A1(n2738), .A2(n2747), .ZN(n2745) );
  NAND2_X1 U2687 ( .A1(n2737), .A2(n2739), .ZN(n2747) );
  NAND2_X1 U2688 ( .A1(n2748), .A2(n2749), .ZN(n2739) );
  NAND2_X1 U2689 ( .A1(b_13_), .A2(a_0_), .ZN(n2749) );
  INV_X1 U2690 ( .A(n2750), .ZN(n2748) );
  XNOR2_X1 U2691 ( .A(n2751), .B(n2752), .ZN(n2737) );
  XOR2_X1 U2692 ( .A(n2753), .B(n2754), .Z(n2752) );
  NAND2_X1 U2693 ( .A1(a_0_), .A2(n2750), .ZN(n2738) );
  NAND2_X1 U2694 ( .A1(n2734), .A2(n2755), .ZN(n2750) );
  NAND2_X1 U2695 ( .A1(n2733), .A2(n2735), .ZN(n2755) );
  NAND2_X1 U2696 ( .A1(n2756), .A2(n2757), .ZN(n2735) );
  NAND2_X1 U2697 ( .A1(b_13_), .A2(a_1_), .ZN(n2757) );
  XOR2_X1 U2698 ( .A(n2758), .B(n2759), .Z(n2733) );
  XNOR2_X1 U2699 ( .A(n2760), .B(n2761), .ZN(n2759) );
  NAND2_X1 U2700 ( .A1(b_12_), .A2(a_2_), .ZN(n2761) );
  NAND2_X1 U2701 ( .A1(a_1_), .A2(n2762), .ZN(n2734) );
  INV_X1 U2702 ( .A(n2756), .ZN(n2762) );
  NOR2_X1 U2703 ( .A1(n2763), .A2(n2764), .ZN(n2756) );
  NOR3_X1 U2704 ( .A1(n2426), .A2(n2765), .A3(n2193), .ZN(n2764) );
  INV_X1 U2705 ( .A(n2766), .ZN(n2765) );
  NAND2_X1 U2706 ( .A1(n2631), .A2(n2629), .ZN(n2766) );
  NOR2_X1 U2707 ( .A1(n2629), .A2(n2631), .ZN(n2763) );
  NOR2_X1 U2708 ( .A1(n2767), .A2(n2768), .ZN(n2631) );
  INV_X1 U2709 ( .A(n2769), .ZN(n2768) );
  NAND3_X1 U2710 ( .A1(a_3_), .A2(n2770), .A3(b_13_), .ZN(n2769) );
  NAND2_X1 U2711 ( .A1(n2730), .A2(n2729), .ZN(n2770) );
  NOR2_X1 U2712 ( .A1(n2729), .A2(n2730), .ZN(n2767) );
  NOR2_X1 U2713 ( .A1(n2771), .A2(n2772), .ZN(n2730) );
  NOR3_X1 U2714 ( .A1(n2424), .A2(n2773), .A3(n2193), .ZN(n2772) );
  NOR2_X1 U2715 ( .A1(n2726), .A2(n2725), .ZN(n2773) );
  INV_X1 U2716 ( .A(n2774), .ZN(n2771) );
  NAND2_X1 U2717 ( .A1(n2725), .A2(n2726), .ZN(n2774) );
  NAND2_X1 U2718 ( .A1(n2722), .A2(n2775), .ZN(n2726) );
  NAND2_X1 U2719 ( .A1(n2721), .A2(n2723), .ZN(n2775) );
  NAND2_X1 U2720 ( .A1(n2776), .A2(n2777), .ZN(n2723) );
  NAND2_X1 U2721 ( .A1(b_13_), .A2(a_5_), .ZN(n2777) );
  XNOR2_X1 U2722 ( .A(n2778), .B(n2779), .ZN(n2721) );
  XOR2_X1 U2723 ( .A(n2780), .B(n2781), .Z(n2779) );
  NAND2_X1 U2724 ( .A1(b_12_), .A2(a_6_), .ZN(n2781) );
  INV_X1 U2725 ( .A(n2782), .ZN(n2722) );
  NOR2_X1 U2726 ( .A1(n2309), .A2(n2776), .ZN(n2782) );
  NOR2_X1 U2727 ( .A1(n2783), .A2(n2784), .ZN(n2776) );
  NOR3_X1 U2728 ( .A1(n2422), .A2(n2785), .A3(n2193), .ZN(n2784) );
  NOR2_X1 U2729 ( .A1(n2651), .A2(n2649), .ZN(n2785) );
  INV_X1 U2730 ( .A(n2786), .ZN(n2783) );
  NAND2_X1 U2731 ( .A1(n2649), .A2(n2651), .ZN(n2786) );
  NAND2_X1 U2732 ( .A1(n2787), .A2(n2788), .ZN(n2651) );
  NAND3_X1 U2733 ( .A1(a_7_), .A2(n2789), .A3(b_13_), .ZN(n2788) );
  NAND2_X1 U2734 ( .A1(n2718), .A2(n2716), .ZN(n2789) );
  INV_X1 U2735 ( .A(n2790), .ZN(n2787) );
  NOR2_X1 U2736 ( .A1(n2716), .A2(n2718), .ZN(n2790) );
  NOR2_X1 U2737 ( .A1(n2791), .A2(n2792), .ZN(n2718) );
  NOR3_X1 U2738 ( .A1(n2663), .A2(n2793), .A3(n2193), .ZN(n2792) );
  NOR2_X1 U2739 ( .A1(n2714), .A2(n2712), .ZN(n2793) );
  INV_X1 U2740 ( .A(n2794), .ZN(n2791) );
  NAND2_X1 U2741 ( .A1(n2712), .A2(n2714), .ZN(n2794) );
  NAND2_X1 U2742 ( .A1(n2710), .A2(n2795), .ZN(n2714) );
  NAND2_X1 U2743 ( .A1(n2709), .A2(n2711), .ZN(n2795) );
  NAND2_X1 U2744 ( .A1(n2796), .A2(n2797), .ZN(n2711) );
  NAND2_X1 U2745 ( .A1(b_13_), .A2(a_9_), .ZN(n2797) );
  INV_X1 U2746 ( .A(n2798), .ZN(n2796) );
  XNOR2_X1 U2747 ( .A(n2799), .B(n2800), .ZN(n2709) );
  NAND2_X1 U2748 ( .A1(n2801), .A2(n2802), .ZN(n2799) );
  NAND2_X1 U2749 ( .A1(a_9_), .A2(n2798), .ZN(n2710) );
  NAND2_X1 U2750 ( .A1(n2671), .A2(n2803), .ZN(n2798) );
  NAND2_X1 U2751 ( .A1(n2670), .A2(n2672), .ZN(n2803) );
  NAND2_X1 U2752 ( .A1(n2804), .A2(n2805), .ZN(n2672) );
  NAND2_X1 U2753 ( .A1(b_13_), .A2(a_10_), .ZN(n2805) );
  INV_X1 U2754 ( .A(n2806), .ZN(n2804) );
  XNOR2_X1 U2755 ( .A(n2807), .B(n2808), .ZN(n2670) );
  XOR2_X1 U2756 ( .A(n2809), .B(n2810), .Z(n2808) );
  NAND2_X1 U2757 ( .A1(b_12_), .A2(a_11_), .ZN(n2810) );
  NAND2_X1 U2758 ( .A1(a_10_), .A2(n2806), .ZN(n2671) );
  NAND2_X1 U2759 ( .A1(n2811), .A2(n2812), .ZN(n2806) );
  NAND3_X1 U2760 ( .A1(a_11_), .A2(n2813), .A3(b_13_), .ZN(n2812) );
  NAND2_X1 U2761 ( .A1(n2680), .A2(n2679), .ZN(n2813) );
  INV_X1 U2762 ( .A(n2814), .ZN(n2811) );
  NOR2_X1 U2763 ( .A1(n2679), .A2(n2680), .ZN(n2814) );
  NOR2_X1 U2764 ( .A1(n2815), .A2(n2816), .ZN(n2680) );
  INV_X1 U2765 ( .A(n2817), .ZN(n2816) );
  NAND2_X1 U2766 ( .A1(n2707), .A2(n2818), .ZN(n2817) );
  NAND2_X1 U2767 ( .A1(n2705), .A2(n2706), .ZN(n2818) );
  NOR2_X1 U2768 ( .A1(n2193), .A2(n2211), .ZN(n2707) );
  NOR2_X1 U2769 ( .A1(n2706), .A2(n2705), .ZN(n2815) );
  XNOR2_X1 U2770 ( .A(n2819), .B(n2820), .ZN(n2705) );
  XNOR2_X1 U2771 ( .A(n2821), .B(n2822), .ZN(n2819) );
  NAND2_X1 U2772 ( .A1(n2823), .A2(n2824), .ZN(n2706) );
  NAND2_X1 U2773 ( .A1(n2825), .A2(n2703), .ZN(n2824) );
  NAND3_X1 U2774 ( .A1(b_12_), .A2(n2416), .A3(b_13_), .ZN(n2703) );
  NAND2_X1 U2775 ( .A1(n2188), .A2(n2826), .ZN(n2825) );
  NAND2_X1 U2776 ( .A1(n2702), .A2(n2409), .ZN(n2823) );
  INV_X1 U2777 ( .A(n2188), .ZN(n2409) );
  NOR2_X1 U2778 ( .A1(n2193), .A2(n2191), .ZN(n2188) );
  INV_X1 U2779 ( .A(b_13_), .ZN(n2193) );
  INV_X1 U2780 ( .A(n2826), .ZN(n2702) );
  NAND2_X1 U2781 ( .A1(n2827), .A2(n2828), .ZN(n2826) );
  NAND2_X1 U2782 ( .A1(b_11_), .A2(n2829), .ZN(n2828) );
  NAND2_X1 U2783 ( .A1(n2170), .A2(n2830), .ZN(n2829) );
  NAND2_X1 U2784 ( .A1(a_15_), .A2(n2417), .ZN(n2830) );
  NAND2_X1 U2785 ( .A1(b_12_), .A2(n2831), .ZN(n2827) );
  NAND2_X1 U2786 ( .A1(n2173), .A2(n2832), .ZN(n2831) );
  NAND2_X1 U2787 ( .A1(a_14_), .A2(n2223), .ZN(n2832) );
  XOR2_X1 U2788 ( .A(n2833), .B(n2834), .Z(n2679) );
  XOR2_X1 U2789 ( .A(n2205), .B(n2835), .Z(n2833) );
  XNOR2_X1 U2790 ( .A(n2836), .B(n2837), .ZN(n2712) );
  NAND2_X1 U2791 ( .A1(n2838), .A2(n2839), .ZN(n2836) );
  XOR2_X1 U2792 ( .A(n2840), .B(n2841), .Z(n2716) );
  XOR2_X1 U2793 ( .A(n2842), .B(n2843), .Z(n2841) );
  NAND2_X1 U2794 ( .A1(b_12_), .A2(a_8_), .ZN(n2843) );
  XNOR2_X1 U2795 ( .A(n2844), .B(n2845), .ZN(n2649) );
  XOR2_X1 U2796 ( .A(n2846), .B(n2847), .Z(n2845) );
  NAND2_X1 U2797 ( .A1(b_12_), .A2(a_7_), .ZN(n2847) );
  XNOR2_X1 U2798 ( .A(n2848), .B(n2849), .ZN(n2725) );
  NAND2_X1 U2799 ( .A1(n2850), .A2(n2851), .ZN(n2848) );
  XNOR2_X1 U2800 ( .A(n2852), .B(n2853), .ZN(n2729) );
  XNOR2_X1 U2801 ( .A(n2854), .B(n2855), .ZN(n2852) );
  NAND2_X1 U2802 ( .A1(b_12_), .A2(a_4_), .ZN(n2854) );
  XNOR2_X1 U2803 ( .A(n2856), .B(n2857), .ZN(n2629) );
  XOR2_X1 U2804 ( .A(n2858), .B(n2859), .Z(n2856) );
  NOR2_X1 U2805 ( .A1(n2344), .A2(n2417), .ZN(n2859) );
  XOR2_X1 U2806 ( .A(n2744), .B(n2743), .Z(n2746) );
  XOR2_X1 U2807 ( .A(n2860), .B(n2861), .Z(n2744) );
  XOR2_X1 U2808 ( .A(n2460), .B(n2459), .Z(n2451) );
  XNOR2_X1 U2809 ( .A(n2493), .B(n2862), .ZN(n2459) );
  XNOR2_X1 U2810 ( .A(n2494), .B(n2491), .ZN(n2862) );
  NOR2_X1 U2811 ( .A1(n2223), .A2(n2433), .ZN(n2491) );
  NAND2_X1 U2812 ( .A1(n2863), .A2(n2864), .ZN(n2494) );
  NAND2_X1 U2813 ( .A1(n2865), .A2(n2866), .ZN(n2864) );
  INV_X1 U2814 ( .A(n2867), .ZN(n2866) );
  NOR2_X1 U2815 ( .A1(n2868), .A2(n2869), .ZN(n2867) );
  NAND2_X1 U2816 ( .A1(n2869), .A2(n2868), .ZN(n2863) );
  XOR2_X1 U2817 ( .A(n2870), .B(n2871), .Z(n2493) );
  NAND2_X1 U2818 ( .A1(n2872), .A2(n2873), .ZN(n2870) );
  NAND2_X1 U2819 ( .A1(n2874), .A2(n2875), .ZN(n2460) );
  NAND2_X1 U2820 ( .A1(n2861), .A2(n2876), .ZN(n2875) );
  NAND2_X1 U2821 ( .A1(n2860), .A2(n2743), .ZN(n2876) );
  NOR2_X1 U2822 ( .A1(n2417), .A2(n2433), .ZN(n2861) );
  INV_X1 U2823 ( .A(n2877), .ZN(n2874) );
  NOR2_X1 U2824 ( .A1(n2743), .A2(n2860), .ZN(n2877) );
  NOR2_X1 U2825 ( .A1(n2878), .A2(n2879), .ZN(n2860) );
  NOR2_X1 U2826 ( .A1(n2754), .A2(n2880), .ZN(n2879) );
  NOR2_X1 U2827 ( .A1(n2753), .A2(n2751), .ZN(n2880) );
  NAND2_X1 U2828 ( .A1(b_12_), .A2(a_1_), .ZN(n2754) );
  INV_X1 U2829 ( .A(n2881), .ZN(n2878) );
  NAND2_X1 U2830 ( .A1(n2751), .A2(n2753), .ZN(n2881) );
  NAND2_X1 U2831 ( .A1(n2882), .A2(n2883), .ZN(n2753) );
  NAND3_X1 U2832 ( .A1(a_2_), .A2(n2884), .A3(b_12_), .ZN(n2883) );
  NAND2_X1 U2833 ( .A1(n2760), .A2(n2758), .ZN(n2884) );
  INV_X1 U2834 ( .A(n2885), .ZN(n2882) );
  NOR2_X1 U2835 ( .A1(n2758), .A2(n2760), .ZN(n2885) );
  NOR2_X1 U2836 ( .A1(n2886), .A2(n2887), .ZN(n2760) );
  NOR3_X1 U2837 ( .A1(n2344), .A2(n2888), .A3(n2417), .ZN(n2887) );
  NOR2_X1 U2838 ( .A1(n2858), .A2(n2857), .ZN(n2888) );
  INV_X1 U2839 ( .A(n2889), .ZN(n2886) );
  NAND2_X1 U2840 ( .A1(n2857), .A2(n2858), .ZN(n2889) );
  NAND2_X1 U2841 ( .A1(n2890), .A2(n2891), .ZN(n2858) );
  NAND3_X1 U2842 ( .A1(a_4_), .A2(n2892), .A3(b_12_), .ZN(n2891) );
  INV_X1 U2843 ( .A(n2893), .ZN(n2892) );
  NOR2_X1 U2844 ( .A1(n2855), .A2(n2853), .ZN(n2893) );
  NAND2_X1 U2845 ( .A1(n2853), .A2(n2855), .ZN(n2890) );
  NAND2_X1 U2846 ( .A1(n2850), .A2(n2894), .ZN(n2855) );
  NAND2_X1 U2847 ( .A1(n2849), .A2(n2851), .ZN(n2894) );
  NAND2_X1 U2848 ( .A1(n2895), .A2(n2896), .ZN(n2851) );
  NAND2_X1 U2849 ( .A1(b_12_), .A2(a_5_), .ZN(n2896) );
  XNOR2_X1 U2850 ( .A(n2897), .B(n2898), .ZN(n2849) );
  XNOR2_X1 U2851 ( .A(n2899), .B(n2900), .ZN(n2897) );
  NOR2_X1 U2852 ( .A1(n2422), .A2(n2223), .ZN(n2900) );
  INV_X1 U2853 ( .A(n2901), .ZN(n2850) );
  NOR2_X1 U2854 ( .A1(n2309), .A2(n2895), .ZN(n2901) );
  NOR2_X1 U2855 ( .A1(n2902), .A2(n2903), .ZN(n2895) );
  NOR3_X1 U2856 ( .A1(n2422), .A2(n2904), .A3(n2417), .ZN(n2903) );
  NOR2_X1 U2857 ( .A1(n2780), .A2(n2778), .ZN(n2904) );
  INV_X1 U2858 ( .A(n2905), .ZN(n2902) );
  NAND2_X1 U2859 ( .A1(n2778), .A2(n2780), .ZN(n2905) );
  NAND2_X1 U2860 ( .A1(n2906), .A2(n2907), .ZN(n2780) );
  NAND3_X1 U2861 ( .A1(a_7_), .A2(n2908), .A3(b_12_), .ZN(n2907) );
  INV_X1 U2862 ( .A(n2909), .ZN(n2908) );
  NOR2_X1 U2863 ( .A1(n2846), .A2(n2844), .ZN(n2909) );
  NAND2_X1 U2864 ( .A1(n2844), .A2(n2846), .ZN(n2906) );
  NAND2_X1 U2865 ( .A1(n2910), .A2(n2911), .ZN(n2846) );
  NAND3_X1 U2866 ( .A1(a_8_), .A2(n2912), .A3(b_12_), .ZN(n2911) );
  INV_X1 U2867 ( .A(n2913), .ZN(n2912) );
  NOR2_X1 U2868 ( .A1(n2842), .A2(n2840), .ZN(n2913) );
  NAND2_X1 U2869 ( .A1(n2840), .A2(n2842), .ZN(n2910) );
  NAND2_X1 U2870 ( .A1(n2838), .A2(n2914), .ZN(n2842) );
  NAND2_X1 U2871 ( .A1(n2837), .A2(n2839), .ZN(n2914) );
  NAND2_X1 U2872 ( .A1(n2915), .A2(n2916), .ZN(n2839) );
  NAND2_X1 U2873 ( .A1(b_12_), .A2(a_9_), .ZN(n2916) );
  INV_X1 U2874 ( .A(n2917), .ZN(n2915) );
  XNOR2_X1 U2875 ( .A(n2918), .B(n2919), .ZN(n2837) );
  NAND2_X1 U2876 ( .A1(n2920), .A2(n2921), .ZN(n2918) );
  NAND2_X1 U2877 ( .A1(a_9_), .A2(n2917), .ZN(n2838) );
  NAND2_X1 U2878 ( .A1(n2801), .A2(n2922), .ZN(n2917) );
  NAND2_X1 U2879 ( .A1(n2800), .A2(n2802), .ZN(n2922) );
  NAND2_X1 U2880 ( .A1(n2923), .A2(n2924), .ZN(n2802) );
  NAND2_X1 U2881 ( .A1(b_12_), .A2(a_10_), .ZN(n2924) );
  INV_X1 U2882 ( .A(n2925), .ZN(n2923) );
  XOR2_X1 U2883 ( .A(n2926), .B(n2927), .Z(n2800) );
  XOR2_X1 U2884 ( .A(n2219), .B(n2928), .Z(n2926) );
  NAND2_X1 U2885 ( .A1(a_10_), .A2(n2925), .ZN(n2801) );
  NAND2_X1 U2886 ( .A1(n2929), .A2(n2930), .ZN(n2925) );
  NAND3_X1 U2887 ( .A1(a_11_), .A2(n2931), .A3(b_12_), .ZN(n2930) );
  NAND2_X1 U2888 ( .A1(n2807), .A2(n2809), .ZN(n2931) );
  INV_X1 U2889 ( .A(n2932), .ZN(n2929) );
  NOR2_X1 U2890 ( .A1(n2809), .A2(n2807), .ZN(n2932) );
  XOR2_X1 U2891 ( .A(n2933), .B(n2934), .Z(n2807) );
  XNOR2_X1 U2892 ( .A(n2935), .B(n2936), .ZN(n2933) );
  NAND2_X1 U2893 ( .A1(n2937), .A2(n2938), .ZN(n2809) );
  NAND2_X1 U2894 ( .A1(n2834), .A2(n2939), .ZN(n2938) );
  INV_X1 U2895 ( .A(n2940), .ZN(n2939) );
  NOR2_X1 U2896 ( .A1(n2205), .A2(n2835), .ZN(n2940) );
  XNOR2_X1 U2897 ( .A(n2941), .B(n2942), .ZN(n2834) );
  XNOR2_X1 U2898 ( .A(n2943), .B(n2944), .ZN(n2941) );
  NAND2_X1 U2899 ( .A1(n2835), .A2(n2205), .ZN(n2937) );
  NAND2_X1 U2900 ( .A1(b_12_), .A2(a_12_), .ZN(n2205) );
  NOR2_X1 U2901 ( .A1(n2945), .A2(n2946), .ZN(n2835) );
  INV_X1 U2902 ( .A(n2947), .ZN(n2946) );
  NAND2_X1 U2903 ( .A1(n2820), .A2(n2948), .ZN(n2947) );
  NAND2_X1 U2904 ( .A1(n2949), .A2(n2822), .ZN(n2948) );
  NOR2_X1 U2905 ( .A1(n2417), .A2(n2191), .ZN(n2820) );
  INV_X1 U2906 ( .A(b_12_), .ZN(n2417) );
  NOR2_X1 U2907 ( .A1(n2822), .A2(n2949), .ZN(n2945) );
  INV_X1 U2908 ( .A(n2821), .ZN(n2949) );
  NAND2_X1 U2909 ( .A1(n2950), .A2(n2951), .ZN(n2821) );
  NAND2_X1 U2910 ( .A1(b_10_), .A2(n2952), .ZN(n2951) );
  NAND2_X1 U2911 ( .A1(n2170), .A2(n2953), .ZN(n2952) );
  NAND2_X1 U2912 ( .A1(a_15_), .A2(n2223), .ZN(n2953) );
  NAND2_X1 U2913 ( .A1(b_11_), .A2(n2954), .ZN(n2950) );
  NAND2_X1 U2914 ( .A1(n2173), .A2(n2955), .ZN(n2954) );
  NAND2_X1 U2915 ( .A1(a_14_), .A2(n2418), .ZN(n2955) );
  NAND3_X1 U2916 ( .A1(b_12_), .A2(n2416), .A3(b_11_), .ZN(n2822) );
  XOR2_X1 U2917 ( .A(n2956), .B(n2957), .Z(n2840) );
  XNOR2_X1 U2918 ( .A(n2958), .B(n2959), .ZN(n2957) );
  XNOR2_X1 U2919 ( .A(n2960), .B(n2961), .ZN(n2844) );
  XNOR2_X1 U2920 ( .A(n2962), .B(n2963), .ZN(n2961) );
  XNOR2_X1 U2921 ( .A(n2964), .B(n2965), .ZN(n2778) );
  XNOR2_X1 U2922 ( .A(n2966), .B(n2967), .ZN(n2964) );
  NOR2_X1 U2923 ( .A1(n2280), .A2(n2223), .ZN(n2967) );
  XNOR2_X1 U2924 ( .A(n2968), .B(n2969), .ZN(n2853) );
  NAND2_X1 U2925 ( .A1(n2970), .A2(n2971), .ZN(n2968) );
  XOR2_X1 U2926 ( .A(n2972), .B(n2973), .Z(n2857) );
  XOR2_X1 U2927 ( .A(n2974), .B(n2975), .Z(n2972) );
  XNOR2_X1 U2928 ( .A(n2976), .B(n2977), .ZN(n2758) );
  XOR2_X1 U2929 ( .A(n2978), .B(n2979), .Z(n2976) );
  XNOR2_X1 U2930 ( .A(n2980), .B(n2981), .ZN(n2751) );
  XOR2_X1 U2931 ( .A(n2982), .B(n2983), .Z(n2981) );
  NAND2_X1 U2932 ( .A1(b_11_), .A2(a_2_), .ZN(n2983) );
  XNOR2_X1 U2933 ( .A(n2865), .B(n2984), .ZN(n2743) );
  XNOR2_X1 U2934 ( .A(n2869), .B(n2868), .ZN(n2984) );
  NAND2_X1 U2935 ( .A1(b_11_), .A2(a_1_), .ZN(n2868) );
  NOR2_X1 U2936 ( .A1(n2985), .A2(n2986), .ZN(n2869) );
  NOR3_X1 U2937 ( .A1(n2426), .A2(n2987), .A3(n2223), .ZN(n2986) );
  NOR2_X1 U2938 ( .A1(n2980), .A2(n2982), .ZN(n2987) );
  INV_X1 U2939 ( .A(n2988), .ZN(n2985) );
  NAND2_X1 U2940 ( .A1(n2980), .A2(n2982), .ZN(n2988) );
  NAND2_X1 U2941 ( .A1(n2989), .A2(n2990), .ZN(n2982) );
  NAND2_X1 U2942 ( .A1(n2979), .A2(n2991), .ZN(n2990) );
  INV_X1 U2943 ( .A(n2992), .ZN(n2991) );
  NOR2_X1 U2944 ( .A1(n2977), .A2(n2978), .ZN(n2992) );
  NOR2_X1 U2945 ( .A1(n2223), .A2(n2344), .ZN(n2979) );
  NAND2_X1 U2946 ( .A1(n2977), .A2(n2978), .ZN(n2989) );
  NAND2_X1 U2947 ( .A1(n2993), .A2(n2994), .ZN(n2978) );
  NAND2_X1 U2948 ( .A1(n2974), .A2(n2995), .ZN(n2994) );
  INV_X1 U2949 ( .A(n2996), .ZN(n2995) );
  NOR2_X1 U2950 ( .A1(n2975), .A2(n2973), .ZN(n2996) );
  NOR2_X1 U2951 ( .A1(n2223), .A2(n2424), .ZN(n2974) );
  NAND2_X1 U2952 ( .A1(n2973), .A2(n2975), .ZN(n2993) );
  NAND2_X1 U2953 ( .A1(n2970), .A2(n2997), .ZN(n2975) );
  NAND2_X1 U2954 ( .A1(n2969), .A2(n2971), .ZN(n2997) );
  NAND2_X1 U2955 ( .A1(n2998), .A2(n2999), .ZN(n2971) );
  NAND2_X1 U2956 ( .A1(b_11_), .A2(a_5_), .ZN(n2999) );
  XNOR2_X1 U2957 ( .A(n3000), .B(n3001), .ZN(n2969) );
  XOR2_X1 U2958 ( .A(n3002), .B(n3003), .Z(n3001) );
  NAND2_X1 U2959 ( .A1(b_10_), .A2(a_6_), .ZN(n3003) );
  INV_X1 U2960 ( .A(n3004), .ZN(n2970) );
  NOR2_X1 U2961 ( .A1(n2309), .A2(n2998), .ZN(n3004) );
  NOR2_X1 U2962 ( .A1(n3005), .A2(n3006), .ZN(n2998) );
  NOR3_X1 U2963 ( .A1(n2422), .A2(n3007), .A3(n2223), .ZN(n3006) );
  INV_X1 U2964 ( .A(n3008), .ZN(n3007) );
  NAND2_X1 U2965 ( .A1(n2898), .A2(n2899), .ZN(n3008) );
  NOR2_X1 U2966 ( .A1(n2898), .A2(n2899), .ZN(n3005) );
  NOR2_X1 U2967 ( .A1(n3009), .A2(n3010), .ZN(n2899) );
  INV_X1 U2968 ( .A(n3011), .ZN(n3010) );
  NAND3_X1 U2969 ( .A1(a_7_), .A2(n3012), .A3(b_11_), .ZN(n3011) );
  NAND2_X1 U2970 ( .A1(n2966), .A2(n2965), .ZN(n3012) );
  NOR2_X1 U2971 ( .A1(n2965), .A2(n2966), .ZN(n3009) );
  NOR2_X1 U2972 ( .A1(n3013), .A2(n3014), .ZN(n2966) );
  INV_X1 U2973 ( .A(n3015), .ZN(n3014) );
  NAND2_X1 U2974 ( .A1(n2963), .A2(n3016), .ZN(n3015) );
  NAND2_X1 U2975 ( .A1(n2960), .A2(n2962), .ZN(n3016) );
  NOR2_X1 U2976 ( .A1(n2223), .A2(n2663), .ZN(n2963) );
  NOR2_X1 U2977 ( .A1(n2960), .A2(n2962), .ZN(n3013) );
  NAND2_X1 U2978 ( .A1(n3017), .A2(n3018), .ZN(n2962) );
  NAND2_X1 U2979 ( .A1(n2956), .A2(n3019), .ZN(n3018) );
  NAND2_X1 U2980 ( .A1(n2959), .A2(n2958), .ZN(n3019) );
  XNOR2_X1 U2981 ( .A(n3020), .B(n3021), .ZN(n2956) );
  XNOR2_X1 U2982 ( .A(n2420), .B(n3022), .ZN(n3021) );
  INV_X1 U2983 ( .A(n3023), .ZN(n3017) );
  NOR2_X1 U2984 ( .A1(n2958), .A2(n2959), .ZN(n3023) );
  NOR2_X1 U2985 ( .A1(n2223), .A2(n2251), .ZN(n2959) );
  NAND2_X1 U2986 ( .A1(n2920), .A2(n3024), .ZN(n2958) );
  NAND2_X1 U2987 ( .A1(n2919), .A2(n2921), .ZN(n3024) );
  NAND2_X1 U2988 ( .A1(n3025), .A2(n3026), .ZN(n2921) );
  NAND2_X1 U2989 ( .A1(b_11_), .A2(a_10_), .ZN(n3025) );
  XNOR2_X1 U2990 ( .A(n3027), .B(n3028), .ZN(n2919) );
  XOR2_X1 U2991 ( .A(n3029), .B(n3030), .Z(n3027) );
  NAND2_X1 U2992 ( .A1(b_10_), .A2(a_11_), .ZN(n3029) );
  INV_X1 U2993 ( .A(n3031), .ZN(n2920) );
  NOR2_X1 U2994 ( .A1(n3026), .A2(n2419), .ZN(n3031) );
  NAND2_X1 U2995 ( .A1(n3032), .A2(n3033), .ZN(n3026) );
  INV_X1 U2996 ( .A(n3034), .ZN(n3033) );
  NOR2_X1 U2997 ( .A1(n2927), .A2(n3035), .ZN(n3034) );
  NOR2_X1 U2998 ( .A1(n2219), .A2(n2928), .ZN(n3035) );
  XNOR2_X1 U2999 ( .A(n3036), .B(n3037), .ZN(n2927) );
  XNOR2_X1 U3000 ( .A(n3038), .B(n3039), .ZN(n3036) );
  NAND2_X1 U3001 ( .A1(n2928), .A2(n2219), .ZN(n3032) );
  NAND2_X1 U3002 ( .A1(b_11_), .A2(a_11_), .ZN(n2219) );
  NOR2_X1 U3003 ( .A1(n3040), .A2(n3041), .ZN(n2928) );
  INV_X1 U3004 ( .A(n3042), .ZN(n3041) );
  NAND2_X1 U3005 ( .A1(n2935), .A2(n3043), .ZN(n3042) );
  NAND2_X1 U3006 ( .A1(n2936), .A2(n2934), .ZN(n3043) );
  NOR2_X1 U3007 ( .A1(n2223), .A2(n2211), .ZN(n2935) );
  NOR2_X1 U3008 ( .A1(n2934), .A2(n2936), .ZN(n3040) );
  NOR2_X1 U3009 ( .A1(n3044), .A2(n3045), .ZN(n2936) );
  INV_X1 U3010 ( .A(n3046), .ZN(n3045) );
  NAND2_X1 U3011 ( .A1(n2942), .A2(n3047), .ZN(n3046) );
  NAND2_X1 U3012 ( .A1(n3048), .A2(n2944), .ZN(n3047) );
  NOR2_X1 U3013 ( .A1(n2223), .A2(n2191), .ZN(n2942) );
  INV_X1 U3014 ( .A(b_11_), .ZN(n2223) );
  NOR2_X1 U3015 ( .A1(n2944), .A2(n3048), .ZN(n3044) );
  INV_X1 U3016 ( .A(n2943), .ZN(n3048) );
  NAND2_X1 U3017 ( .A1(n3049), .A2(n3050), .ZN(n2943) );
  NAND2_X1 U3018 ( .A1(b_10_), .A2(n3051), .ZN(n3050) );
  NAND2_X1 U3019 ( .A1(n2173), .A2(n3052), .ZN(n3051) );
  NAND2_X1 U3020 ( .A1(a_14_), .A2(n2253), .ZN(n3052) );
  NAND2_X1 U3021 ( .A1(b_9_), .A2(n3053), .ZN(n3049) );
  NAND2_X1 U3022 ( .A1(n2170), .A2(n3054), .ZN(n3053) );
  NAND2_X1 U3023 ( .A1(a_15_), .A2(n2418), .ZN(n3054) );
  NAND3_X1 U3024 ( .A1(b_10_), .A2(n2416), .A3(b_11_), .ZN(n2944) );
  XNOR2_X1 U3025 ( .A(n3055), .B(n3056), .ZN(n2934) );
  XNOR2_X1 U3026 ( .A(n3057), .B(n3058), .ZN(n3055) );
  XOR2_X1 U3027 ( .A(n3059), .B(n3060), .Z(n2960) );
  NAND2_X1 U3028 ( .A1(n3061), .A2(n3062), .ZN(n3059) );
  XOR2_X1 U3029 ( .A(n3063), .B(n3064), .Z(n2965) );
  XOR2_X1 U3030 ( .A(n3065), .B(n3066), .Z(n3064) );
  NAND2_X1 U3031 ( .A1(b_10_), .A2(a_8_), .ZN(n3066) );
  XOR2_X1 U3032 ( .A(n3067), .B(n3068), .Z(n2898) );
  XOR2_X1 U3033 ( .A(n3069), .B(n3070), .Z(n3068) );
  NAND2_X1 U3034 ( .A1(b_10_), .A2(a_7_), .ZN(n3070) );
  XNOR2_X1 U3035 ( .A(n3071), .B(n3072), .ZN(n2973) );
  NAND2_X1 U3036 ( .A1(n3073), .A2(n3074), .ZN(n3071) );
  XOR2_X1 U3037 ( .A(n3075), .B(n3076), .Z(n2977) );
  XOR2_X1 U3038 ( .A(n3077), .B(n3078), .Z(n3075) );
  NOR2_X1 U3039 ( .A1(n2424), .A2(n2418), .ZN(n3078) );
  XNOR2_X1 U3040 ( .A(n3079), .B(n3080), .ZN(n2980) );
  XNOR2_X1 U3041 ( .A(n3081), .B(n3082), .ZN(n3079) );
  XOR2_X1 U3042 ( .A(n3083), .B(n3084), .Z(n2865) );
  XOR2_X1 U3043 ( .A(n3085), .B(n3086), .Z(n3083) );
  NAND2_X1 U3044 ( .A1(b_10_), .A2(a_2_), .ZN(n3085) );
  NAND3_X1 U3045 ( .A1(n2122), .A2(n2121), .A3(n2479), .ZN(n2118) );
  INV_X1 U3046 ( .A(n2119), .ZN(n2479) );
  NAND2_X1 U3047 ( .A1(n3087), .A2(n2477), .ZN(n2119) );
  NAND2_X1 U3048 ( .A1(n3088), .A2(n3089), .ZN(n3087) );
  XNOR2_X1 U3049 ( .A(n3090), .B(n3091), .ZN(n3089) );
  INV_X1 U3050 ( .A(n3092), .ZN(n2121) );
  NAND2_X1 U3051 ( .A1(n3093), .A2(n3094), .ZN(n3092) );
  NAND2_X1 U3052 ( .A1(n2486), .A2(n3095), .ZN(n3094) );
  NAND2_X1 U3053 ( .A1(n2487), .A2(n3096), .ZN(n3095) );
  XNOR2_X1 U3054 ( .A(n3097), .B(n3098), .ZN(n2486) );
  XOR2_X1 U3055 ( .A(n3099), .B(n3100), .Z(n3097) );
  NOR2_X1 U3056 ( .A1(n2253), .A2(n2427), .ZN(n3100) );
  NAND2_X1 U3057 ( .A1(n2488), .A2(n3101), .ZN(n3093) );
  INV_X1 U3058 ( .A(n2487), .ZN(n3101) );
  NOR2_X1 U3059 ( .A1(n2418), .A2(n2433), .ZN(n2487) );
  INV_X1 U3060 ( .A(n3096), .ZN(n2488) );
  NAND2_X1 U3061 ( .A1(n2872), .A2(n3102), .ZN(n3096) );
  NAND2_X1 U3062 ( .A1(n2871), .A2(n2873), .ZN(n3102) );
  NAND2_X1 U3063 ( .A1(n3103), .A2(n3104), .ZN(n2873) );
  NAND2_X1 U3064 ( .A1(b_10_), .A2(a_1_), .ZN(n3104) );
  INV_X1 U3065 ( .A(n3105), .ZN(n3103) );
  XOR2_X1 U3066 ( .A(n3106), .B(n3107), .Z(n2871) );
  XNOR2_X1 U3067 ( .A(n3108), .B(n3109), .ZN(n3107) );
  NAND2_X1 U3068 ( .A1(a_2_), .A2(b_9_), .ZN(n3109) );
  NAND2_X1 U3069 ( .A1(a_1_), .A2(n3105), .ZN(n2872) );
  NAND2_X1 U3070 ( .A1(n3110), .A2(n3111), .ZN(n3105) );
  NAND3_X1 U3071 ( .A1(a_2_), .A2(n3112), .A3(b_10_), .ZN(n3111) );
  NAND2_X1 U3072 ( .A1(n3086), .A2(n3084), .ZN(n3112) );
  INV_X1 U3073 ( .A(n3113), .ZN(n3110) );
  NOR2_X1 U3074 ( .A1(n3084), .A2(n3086), .ZN(n3113) );
  NOR2_X1 U3075 ( .A1(n3114), .A2(n3115), .ZN(n3086) );
  INV_X1 U3076 ( .A(n3116), .ZN(n3115) );
  NAND2_X1 U3077 ( .A1(n3082), .A2(n3117), .ZN(n3116) );
  NAND2_X1 U3078 ( .A1(n3081), .A2(n3080), .ZN(n3117) );
  NOR2_X1 U3079 ( .A1(n2418), .A2(n2344), .ZN(n3082) );
  NOR2_X1 U3080 ( .A1(n3080), .A2(n3081), .ZN(n3114) );
  NOR2_X1 U3081 ( .A1(n3118), .A2(n3119), .ZN(n3081) );
  NOR3_X1 U3082 ( .A1(n2424), .A2(n3120), .A3(n2418), .ZN(n3119) );
  NOR2_X1 U3083 ( .A1(n3077), .A2(n3076), .ZN(n3120) );
  INV_X1 U3084 ( .A(n3121), .ZN(n3118) );
  NAND2_X1 U3085 ( .A1(n3076), .A2(n3077), .ZN(n3121) );
  NAND2_X1 U3086 ( .A1(n3073), .A2(n3122), .ZN(n3077) );
  NAND2_X1 U3087 ( .A1(n3072), .A2(n3074), .ZN(n3122) );
  NAND2_X1 U3088 ( .A1(n3123), .A2(n3124), .ZN(n3074) );
  NAND2_X1 U3089 ( .A1(b_10_), .A2(a_5_), .ZN(n3124) );
  XNOR2_X1 U3090 ( .A(n3125), .B(n3126), .ZN(n3072) );
  XNOR2_X1 U3091 ( .A(n3127), .B(n3128), .ZN(n3125) );
  INV_X1 U3092 ( .A(n3129), .ZN(n3073) );
  NOR2_X1 U3093 ( .A1(n2309), .A2(n3123), .ZN(n3129) );
  NOR2_X1 U3094 ( .A1(n3130), .A2(n3131), .ZN(n3123) );
  NOR3_X1 U3095 ( .A1(n2422), .A2(n3132), .A3(n2418), .ZN(n3131) );
  NOR2_X1 U3096 ( .A1(n3002), .A2(n3000), .ZN(n3132) );
  INV_X1 U3097 ( .A(n3133), .ZN(n3130) );
  NAND2_X1 U3098 ( .A1(n3000), .A2(n3002), .ZN(n3133) );
  NAND2_X1 U3099 ( .A1(n3134), .A2(n3135), .ZN(n3002) );
  INV_X1 U3100 ( .A(n3136), .ZN(n3135) );
  NOR3_X1 U3101 ( .A1(n2280), .A2(n3137), .A3(n2418), .ZN(n3136) );
  NOR2_X1 U3102 ( .A1(n3069), .A2(n3067), .ZN(n3137) );
  NAND2_X1 U3103 ( .A1(n3067), .A2(n3069), .ZN(n3134) );
  NAND2_X1 U3104 ( .A1(n3138), .A2(n3139), .ZN(n3069) );
  NAND3_X1 U3105 ( .A1(a_8_), .A2(n3140), .A3(b_10_), .ZN(n3139) );
  INV_X1 U3106 ( .A(n3141), .ZN(n3140) );
  NOR2_X1 U3107 ( .A1(n3065), .A2(n3063), .ZN(n3141) );
  NAND2_X1 U3108 ( .A1(n3063), .A2(n3065), .ZN(n3138) );
  NAND2_X1 U3109 ( .A1(n3061), .A2(n3142), .ZN(n3065) );
  NAND2_X1 U3110 ( .A1(n3060), .A2(n3062), .ZN(n3142) );
  NAND2_X1 U3111 ( .A1(n3143), .A2(n3144), .ZN(n3062) );
  NAND2_X1 U3112 ( .A1(b_10_), .A2(a_9_), .ZN(n3143) );
  XNOR2_X1 U3113 ( .A(n3145), .B(n3146), .ZN(n3060) );
  NAND2_X1 U3114 ( .A1(n3147), .A2(n3148), .ZN(n3145) );
  INV_X1 U3115 ( .A(n3149), .ZN(n3061) );
  NOR2_X1 U3116 ( .A1(n3144), .A2(n2251), .ZN(n3149) );
  NAND2_X1 U3117 ( .A1(n3150), .A2(n3151), .ZN(n3144) );
  NAND2_X1 U3118 ( .A1(n3020), .A2(n3152), .ZN(n3151) );
  NAND2_X1 U3119 ( .A1(n2420), .A2(n3022), .ZN(n3152) );
  XOR2_X1 U3120 ( .A(n3153), .B(n3154), .Z(n3020) );
  XOR2_X1 U3121 ( .A(n3155), .B(n3156), .Z(n3153) );
  NAND2_X1 U3122 ( .A1(a_11_), .A2(b_9_), .ZN(n3155) );
  INV_X1 U3123 ( .A(n3157), .ZN(n3150) );
  NOR2_X1 U3124 ( .A1(n3022), .A2(n2420), .ZN(n3157) );
  NOR2_X1 U3125 ( .A1(n2418), .A2(n2419), .ZN(n2420) );
  NAND2_X1 U3126 ( .A1(n3158), .A2(n3159), .ZN(n3022) );
  NAND3_X1 U3127 ( .A1(a_11_), .A2(n3160), .A3(b_10_), .ZN(n3159) );
  NAND2_X1 U3128 ( .A1(n3030), .A2(n3028), .ZN(n3160) );
  INV_X1 U3129 ( .A(n3161), .ZN(n3158) );
  NOR2_X1 U3130 ( .A1(n3028), .A2(n3030), .ZN(n3161) );
  NOR2_X1 U3131 ( .A1(n3162), .A2(n3163), .ZN(n3030) );
  INV_X1 U3132 ( .A(n3164), .ZN(n3163) );
  NAND2_X1 U3133 ( .A1(n3038), .A2(n3165), .ZN(n3164) );
  NAND2_X1 U3134 ( .A1(n3039), .A2(n3037), .ZN(n3165) );
  NOR2_X1 U3135 ( .A1(n2418), .A2(n2211), .ZN(n3038) );
  NOR2_X1 U3136 ( .A1(n3037), .A2(n3039), .ZN(n3162) );
  NOR2_X1 U3137 ( .A1(n3166), .A2(n3167), .ZN(n3039) );
  INV_X1 U3138 ( .A(n3168), .ZN(n3167) );
  NAND2_X1 U3139 ( .A1(n3056), .A2(n3169), .ZN(n3168) );
  NAND2_X1 U3140 ( .A1(n3170), .A2(n3058), .ZN(n3169) );
  NOR2_X1 U3141 ( .A1(n2418), .A2(n2191), .ZN(n3056) );
  INV_X1 U3142 ( .A(b_10_), .ZN(n2418) );
  NOR2_X1 U3143 ( .A1(n3058), .A2(n3170), .ZN(n3166) );
  INV_X1 U3144 ( .A(n3057), .ZN(n3170) );
  NAND2_X1 U3145 ( .A1(n3171), .A2(n3172), .ZN(n3057) );
  NAND2_X1 U3146 ( .A1(b_8_), .A2(n3173), .ZN(n3172) );
  NAND2_X1 U3147 ( .A1(n2170), .A2(n3174), .ZN(n3173) );
  NAND2_X1 U3148 ( .A1(a_15_), .A2(n2253), .ZN(n3174) );
  NAND2_X1 U3149 ( .A1(b_9_), .A2(n3175), .ZN(n3171) );
  NAND2_X1 U3150 ( .A1(n2173), .A2(n3176), .ZN(n3175) );
  NAND2_X1 U3151 ( .A1(a_14_), .A2(n3177), .ZN(n3176) );
  NAND3_X1 U3152 ( .A1(n2416), .A2(b_9_), .A3(b_10_), .ZN(n3058) );
  XNOR2_X1 U3153 ( .A(n3178), .B(n3179), .ZN(n3037) );
  XNOR2_X1 U3154 ( .A(n3180), .B(n3181), .ZN(n3178) );
  XOR2_X1 U3155 ( .A(n3182), .B(n3183), .Z(n3028) );
  XNOR2_X1 U3156 ( .A(n3184), .B(n3185), .ZN(n3182) );
  XNOR2_X1 U3157 ( .A(n3186), .B(n3187), .ZN(n3063) );
  XNOR2_X1 U3158 ( .A(n2248), .B(n3188), .ZN(n3186) );
  XNOR2_X1 U3159 ( .A(n3189), .B(n3190), .ZN(n3067) );
  XNOR2_X1 U3160 ( .A(n3191), .B(n3192), .ZN(n3190) );
  XNOR2_X1 U3161 ( .A(n3193), .B(n3194), .ZN(n3000) );
  XNOR2_X1 U3162 ( .A(n3195), .B(n3196), .ZN(n3193) );
  NOR2_X1 U3163 ( .A1(n2253), .A2(n2280), .ZN(n3196) );
  XNOR2_X1 U3164 ( .A(n3197), .B(n3198), .ZN(n3076) );
  XOR2_X1 U3165 ( .A(n3199), .B(n3200), .Z(n3198) );
  XOR2_X1 U3166 ( .A(n3201), .B(n3202), .Z(n3080) );
  NAND2_X1 U3167 ( .A1(n3203), .A2(n3204), .ZN(n3201) );
  XNOR2_X1 U3168 ( .A(n3205), .B(n3206), .ZN(n3084) );
  XOR2_X1 U3169 ( .A(n3207), .B(n3208), .Z(n3205) );
  NOR2_X1 U3170 ( .A1(n2253), .A2(n2344), .ZN(n3208) );
  XNOR2_X1 U3171 ( .A(n3209), .B(n3210), .ZN(n2122) );
  XOR2_X1 U3172 ( .A(n3211), .B(n3212), .Z(n3210) );
  NAND2_X1 U3173 ( .A1(a_0_), .A2(b_9_), .ZN(n3212) );
  NAND2_X1 U3174 ( .A1(n3213), .A2(n3214), .ZN(n2477) );
  INV_X1 U3175 ( .A(n3088), .ZN(n3214) );
  NOR2_X1 U3176 ( .A1(n3215), .A2(n3216), .ZN(n3088) );
  NOR3_X1 U3177 ( .A1(n2253), .A2(n3217), .A3(n2433), .ZN(n3216) );
  NOR2_X1 U3178 ( .A1(n3211), .A2(n3209), .ZN(n3217) );
  INV_X1 U3179 ( .A(n3218), .ZN(n3215) );
  NAND2_X1 U3180 ( .A1(n3209), .A2(n3211), .ZN(n3218) );
  NAND2_X1 U3181 ( .A1(n3219), .A2(n3220), .ZN(n3211) );
  NAND3_X1 U3182 ( .A1(b_9_), .A2(n3221), .A3(a_1_), .ZN(n3220) );
  INV_X1 U3183 ( .A(n3222), .ZN(n3221) );
  NOR2_X1 U3184 ( .A1(n3099), .A2(n3098), .ZN(n3222) );
  NAND2_X1 U3185 ( .A1(n3098), .A2(n3099), .ZN(n3219) );
  NAND2_X1 U3186 ( .A1(n3223), .A2(n3224), .ZN(n3099) );
  NAND3_X1 U3187 ( .A1(b_9_), .A2(n3225), .A3(a_2_), .ZN(n3224) );
  NAND2_X1 U3188 ( .A1(n3108), .A2(n3106), .ZN(n3225) );
  INV_X1 U3189 ( .A(n3226), .ZN(n3223) );
  NOR2_X1 U3190 ( .A1(n3106), .A2(n3108), .ZN(n3226) );
  NOR2_X1 U3191 ( .A1(n3227), .A2(n3228), .ZN(n3108) );
  NOR3_X1 U3192 ( .A1(n2253), .A2(n3229), .A3(n2344), .ZN(n3228) );
  NOR2_X1 U3193 ( .A1(n3207), .A2(n3206), .ZN(n3229) );
  INV_X1 U3194 ( .A(n3230), .ZN(n3227) );
  NAND2_X1 U3195 ( .A1(n3206), .A2(n3207), .ZN(n3230) );
  NAND2_X1 U3196 ( .A1(n3203), .A2(n3231), .ZN(n3207) );
  NAND2_X1 U3197 ( .A1(n3202), .A2(n3204), .ZN(n3231) );
  NAND2_X1 U3198 ( .A1(n3232), .A2(n3233), .ZN(n3204) );
  NAND2_X1 U3199 ( .A1(a_4_), .A2(b_9_), .ZN(n3233) );
  INV_X1 U3200 ( .A(n3234), .ZN(n3232) );
  XOR2_X1 U3201 ( .A(n3235), .B(n3236), .Z(n3202) );
  XOR2_X1 U3202 ( .A(n3237), .B(n3238), .Z(n3236) );
  NAND2_X1 U3203 ( .A1(a_4_), .A2(n3234), .ZN(n3203) );
  NAND2_X1 U3204 ( .A1(n3239), .A2(n3240), .ZN(n3234) );
  INV_X1 U3205 ( .A(n3241), .ZN(n3240) );
  NOR2_X1 U3206 ( .A1(n3200), .A2(n3242), .ZN(n3241) );
  NOR2_X1 U3207 ( .A1(n3199), .A2(n3197), .ZN(n3242) );
  NAND2_X1 U3208 ( .A1(b_9_), .A2(a_5_), .ZN(n3200) );
  NAND2_X1 U3209 ( .A1(n3197), .A2(n3199), .ZN(n3239) );
  NAND2_X1 U3210 ( .A1(n3243), .A2(n3244), .ZN(n3199) );
  NAND2_X1 U3211 ( .A1(n3128), .A2(n3245), .ZN(n3244) );
  NAND2_X1 U3212 ( .A1(n3127), .A2(n3126), .ZN(n3245) );
  NOR2_X1 U3213 ( .A1(n2422), .A2(n2253), .ZN(n3128) );
  INV_X1 U3214 ( .A(n3246), .ZN(n3243) );
  NOR2_X1 U3215 ( .A1(n3126), .A2(n3127), .ZN(n3246) );
  NOR2_X1 U3216 ( .A1(n3247), .A2(n3248), .ZN(n3127) );
  NOR3_X1 U3217 ( .A1(n2253), .A2(n3249), .A3(n2280), .ZN(n3248) );
  NOR2_X1 U3218 ( .A1(n3250), .A2(n3251), .ZN(n3249) );
  INV_X1 U3219 ( .A(n3194), .ZN(n3251) );
  INV_X1 U3220 ( .A(n3195), .ZN(n3250) );
  NOR2_X1 U3221 ( .A1(n3194), .A2(n3195), .ZN(n3247) );
  NOR2_X1 U3222 ( .A1(n3252), .A2(n3253), .ZN(n3195) );
  INV_X1 U3223 ( .A(n3254), .ZN(n3253) );
  NAND2_X1 U3224 ( .A1(n3192), .A2(n3255), .ZN(n3254) );
  NAND2_X1 U3225 ( .A1(n3189), .A2(n3191), .ZN(n3255) );
  NOR2_X1 U3226 ( .A1(n2663), .A2(n2253), .ZN(n3192) );
  NOR2_X1 U3227 ( .A1(n3191), .A2(n3189), .ZN(n3252) );
  XOR2_X1 U3228 ( .A(n3256), .B(n3257), .Z(n3189) );
  NAND2_X1 U3229 ( .A1(n3258), .A2(n3259), .ZN(n3256) );
  NAND2_X1 U3230 ( .A1(n3260), .A2(n3261), .ZN(n3191) );
  NAND2_X1 U3231 ( .A1(n3187), .A2(n3262), .ZN(n3261) );
  NAND2_X1 U3232 ( .A1(n2248), .A2(n3263), .ZN(n3262) );
  XOR2_X1 U3233 ( .A(n3264), .B(n3265), .Z(n3187) );
  NAND2_X1 U3234 ( .A1(n3266), .A2(n3267), .ZN(n3264) );
  NAND2_X1 U3235 ( .A1(n3188), .A2(n2402), .ZN(n3260) );
  INV_X1 U3236 ( .A(n2248), .ZN(n2402) );
  NOR2_X1 U3237 ( .A1(n2251), .A2(n2253), .ZN(n2248) );
  INV_X1 U3238 ( .A(n3263), .ZN(n3188) );
  NAND2_X1 U3239 ( .A1(n3147), .A2(n3268), .ZN(n3263) );
  NAND2_X1 U3240 ( .A1(n3146), .A2(n3148), .ZN(n3268) );
  NAND2_X1 U3241 ( .A1(n3269), .A2(n3270), .ZN(n3148) );
  NAND2_X1 U3242 ( .A1(a_10_), .A2(b_9_), .ZN(n3270) );
  INV_X1 U3243 ( .A(n3271), .ZN(n3269) );
  XNOR2_X1 U3244 ( .A(n3272), .B(n3273), .ZN(n3146) );
  XOR2_X1 U3245 ( .A(n3274), .B(n3275), .Z(n3272) );
  NAND2_X1 U3246 ( .A1(a_11_), .A2(b_8_), .ZN(n3274) );
  NAND2_X1 U3247 ( .A1(a_10_), .A2(n3271), .ZN(n3147) );
  NAND2_X1 U3248 ( .A1(n3276), .A2(n3277), .ZN(n3271) );
  NAND3_X1 U3249 ( .A1(b_9_), .A2(n3278), .A3(a_11_), .ZN(n3277) );
  NAND2_X1 U3250 ( .A1(n3156), .A2(n3154), .ZN(n3278) );
  INV_X1 U3251 ( .A(n3279), .ZN(n3276) );
  NOR2_X1 U3252 ( .A1(n3154), .A2(n3156), .ZN(n3279) );
  NOR2_X1 U3253 ( .A1(n3280), .A2(n3281), .ZN(n3156) );
  INV_X1 U3254 ( .A(n3282), .ZN(n3281) );
  NAND2_X1 U3255 ( .A1(n3184), .A2(n3283), .ZN(n3282) );
  NAND2_X1 U3256 ( .A1(n3185), .A2(n3183), .ZN(n3283) );
  NOR2_X1 U3257 ( .A1(n2211), .A2(n2253), .ZN(n3184) );
  NOR2_X1 U3258 ( .A1(n3183), .A2(n3185), .ZN(n3280) );
  NOR2_X1 U3259 ( .A1(n3284), .A2(n3285), .ZN(n3185) );
  INV_X1 U3260 ( .A(n3286), .ZN(n3285) );
  NAND2_X1 U3261 ( .A1(n3179), .A2(n3287), .ZN(n3286) );
  NAND2_X1 U3262 ( .A1(n3288), .A2(n3181), .ZN(n3287) );
  NOR2_X1 U3263 ( .A1(n2191), .A2(n2253), .ZN(n3179) );
  INV_X1 U3264 ( .A(b_9_), .ZN(n2253) );
  NOR2_X1 U3265 ( .A1(n3181), .A2(n3288), .ZN(n3284) );
  INV_X1 U3266 ( .A(n3180), .ZN(n3288) );
  NAND2_X1 U3267 ( .A1(n3289), .A2(n3290), .ZN(n3180) );
  NAND2_X1 U3268 ( .A1(b_7_), .A2(n3291), .ZN(n3290) );
  NAND2_X1 U3269 ( .A1(n2170), .A2(n3292), .ZN(n3291) );
  NAND2_X1 U3270 ( .A1(a_15_), .A2(n3177), .ZN(n3292) );
  NAND2_X1 U3271 ( .A1(b_8_), .A2(n3293), .ZN(n3289) );
  NAND2_X1 U3272 ( .A1(n2173), .A2(n3294), .ZN(n3293) );
  NAND2_X1 U3273 ( .A1(a_14_), .A2(n2282), .ZN(n3294) );
  NAND3_X1 U3274 ( .A1(n2416), .A2(b_9_), .A3(b_8_), .ZN(n3181) );
  XNOR2_X1 U3275 ( .A(n3295), .B(n3296), .ZN(n3183) );
  XNOR2_X1 U3276 ( .A(n3297), .B(n3298), .ZN(n3295) );
  XOR2_X1 U3277 ( .A(n3299), .B(n3300), .Z(n3154) );
  XNOR2_X1 U3278 ( .A(n3301), .B(n3302), .ZN(n3299) );
  XNOR2_X1 U3279 ( .A(n3303), .B(n3304), .ZN(n3194) );
  XNOR2_X1 U3280 ( .A(n2265), .B(n3305), .ZN(n3304) );
  XNOR2_X1 U3281 ( .A(n3306), .B(n3307), .ZN(n3126) );
  XNOR2_X1 U3282 ( .A(n3308), .B(n3309), .ZN(n3307) );
  NAND2_X1 U3283 ( .A1(a_7_), .A2(b_8_), .ZN(n3309) );
  XOR2_X1 U3284 ( .A(n3310), .B(n3311), .Z(n3197) );
  XOR2_X1 U3285 ( .A(n3312), .B(n3313), .Z(n3310) );
  NOR2_X1 U3286 ( .A1(n2422), .A2(n3177), .ZN(n3313) );
  XOR2_X1 U3287 ( .A(n3314), .B(n3315), .Z(n3206) );
  XNOR2_X1 U3288 ( .A(n3316), .B(n3317), .ZN(n3314) );
  NAND2_X1 U3289 ( .A1(a_4_), .A2(b_8_), .ZN(n3316) );
  XOR2_X1 U3290 ( .A(n3318), .B(n3319), .Z(n3106) );
  NAND2_X1 U3291 ( .A1(n3320), .A2(n3321), .ZN(n3318) );
  XNOR2_X1 U3292 ( .A(n3322), .B(n3323), .ZN(n3098) );
  NAND2_X1 U3293 ( .A1(n3324), .A2(n3325), .ZN(n3322) );
  XOR2_X1 U3294 ( .A(n3326), .B(n3327), .Z(n3209) );
  XOR2_X1 U3295 ( .A(n3328), .B(n3329), .Z(n3326) );
  XNOR2_X1 U3296 ( .A(n3091), .B(n3330), .ZN(n3213) );
  XNOR2_X1 U3297 ( .A(n3331), .B(n3332), .ZN(n3091) );
  XNOR2_X1 U3298 ( .A(n3333), .B(n2134), .ZN(n2125) );
  INV_X1 U3299 ( .A(n2129), .ZN(n2474) );
  NOR3_X1 U3300 ( .A1(n2134), .A2(n2133), .A3(n2476), .ZN(n2129) );
  NAND2_X1 U3301 ( .A1(n3334), .A2(n2473), .ZN(n2476) );
  NAND2_X1 U3302 ( .A1(n3335), .A2(n3336), .ZN(n3334) );
  INV_X1 U3303 ( .A(n3337), .ZN(n3336) );
  XOR2_X1 U3304 ( .A(n3338), .B(n3339), .Z(n3335) );
  INV_X1 U3305 ( .A(n3333), .ZN(n2133) );
  NAND2_X1 U3306 ( .A1(n3340), .A2(n3341), .ZN(n3333) );
  NAND2_X1 U3307 ( .A1(n3332), .A2(n3342), .ZN(n3341) );
  NAND2_X1 U3308 ( .A1(n3090), .A2(n3343), .ZN(n3342) );
  INV_X1 U3309 ( .A(n3331), .ZN(n3343) );
  INV_X1 U3310 ( .A(n3330), .ZN(n3090) );
  NOR2_X1 U3311 ( .A1(n2433), .A2(n3177), .ZN(n3332) );
  NAND2_X1 U3312 ( .A1(n3330), .A2(n3331), .ZN(n3340) );
  NAND2_X1 U3313 ( .A1(n3344), .A2(n3345), .ZN(n3331) );
  NAND2_X1 U3314 ( .A1(n3329), .A2(n3346), .ZN(n3345) );
  INV_X1 U3315 ( .A(n3347), .ZN(n3346) );
  NOR2_X1 U3316 ( .A1(n3328), .A2(n3327), .ZN(n3347) );
  NOR2_X1 U3317 ( .A1(n2427), .A2(n3177), .ZN(n3329) );
  NAND2_X1 U3318 ( .A1(n3327), .A2(n3328), .ZN(n3344) );
  NAND2_X1 U3319 ( .A1(n3324), .A2(n3348), .ZN(n3328) );
  NAND2_X1 U3320 ( .A1(n3323), .A2(n3325), .ZN(n3348) );
  NAND2_X1 U3321 ( .A1(n3349), .A2(n3350), .ZN(n3325) );
  NAND2_X1 U3322 ( .A1(a_2_), .A2(b_8_), .ZN(n3350) );
  INV_X1 U3323 ( .A(n3351), .ZN(n3349) );
  XNOR2_X1 U3324 ( .A(n3352), .B(n3353), .ZN(n3323) );
  XNOR2_X1 U3325 ( .A(n3354), .B(n3355), .ZN(n3352) );
  NOR2_X1 U3326 ( .A1(n2282), .A2(n2344), .ZN(n3355) );
  NAND2_X1 U3327 ( .A1(a_2_), .A2(n3351), .ZN(n3324) );
  NAND2_X1 U3328 ( .A1(n3320), .A2(n3356), .ZN(n3351) );
  NAND2_X1 U3329 ( .A1(n3319), .A2(n3321), .ZN(n3356) );
  NAND2_X1 U3330 ( .A1(n3357), .A2(n3358), .ZN(n3321) );
  NAND2_X1 U3331 ( .A1(a_3_), .A2(b_8_), .ZN(n3358) );
  XOR2_X1 U3332 ( .A(n3359), .B(n3360), .Z(n3319) );
  XNOR2_X1 U3333 ( .A(n3361), .B(n3362), .ZN(n3360) );
  NAND2_X1 U3334 ( .A1(a_4_), .A2(b_7_), .ZN(n3362) );
  INV_X1 U3335 ( .A(n3363), .ZN(n3320) );
  NOR2_X1 U3336 ( .A1(n2344), .A2(n3357), .ZN(n3363) );
  NOR2_X1 U3337 ( .A1(n3364), .A2(n3365), .ZN(n3357) );
  NOR3_X1 U3338 ( .A1(n3177), .A2(n3366), .A3(n2424), .ZN(n3365) );
  NOR2_X1 U3339 ( .A1(n3315), .A2(n3317), .ZN(n3366) );
  INV_X1 U3340 ( .A(n3367), .ZN(n3364) );
  NAND2_X1 U3341 ( .A1(n3315), .A2(n3317), .ZN(n3367) );
  NAND2_X1 U3342 ( .A1(n3368), .A2(n3369), .ZN(n3317) );
  NAND2_X1 U3343 ( .A1(n3238), .A2(n3370), .ZN(n3369) );
  NAND2_X1 U3344 ( .A1(n3235), .A2(n3237), .ZN(n3370) );
  NOR2_X1 U3345 ( .A1(n3177), .A2(n2309), .ZN(n3238) );
  INV_X1 U3346 ( .A(n3371), .ZN(n3368) );
  NOR2_X1 U3347 ( .A1(n3235), .A2(n3237), .ZN(n3371) );
  NOR2_X1 U3348 ( .A1(n3372), .A2(n3373), .ZN(n3237) );
  NOR3_X1 U3349 ( .A1(n2422), .A2(n3374), .A3(n3177), .ZN(n3373) );
  NOR2_X1 U3350 ( .A1(n3312), .A2(n3311), .ZN(n3374) );
  INV_X1 U3351 ( .A(n3375), .ZN(n3372) );
  NAND2_X1 U3352 ( .A1(n3311), .A2(n3312), .ZN(n3375) );
  NAND2_X1 U3353 ( .A1(n3376), .A2(n3377), .ZN(n3312) );
  NAND3_X1 U3354 ( .A1(b_8_), .A2(n3378), .A3(a_7_), .ZN(n3377) );
  NAND2_X1 U3355 ( .A1(n3379), .A2(n3380), .ZN(n3378) );
  INV_X1 U3356 ( .A(n3308), .ZN(n3380) );
  INV_X1 U3357 ( .A(n3306), .ZN(n3379) );
  NAND2_X1 U3358 ( .A1(n3308), .A2(n3306), .ZN(n3376) );
  XNOR2_X1 U3359 ( .A(n3381), .B(n3382), .ZN(n3306) );
  XOR2_X1 U3360 ( .A(n3383), .B(n3384), .Z(n3382) );
  NOR2_X1 U3361 ( .A1(n3385), .A2(n3386), .ZN(n3308) );
  INV_X1 U3362 ( .A(n3387), .ZN(n3386) );
  NAND2_X1 U3363 ( .A1(n3303), .A2(n3388), .ZN(n3387) );
  NAND2_X1 U3364 ( .A1(n2265), .A2(n3305), .ZN(n3388) );
  XOR2_X1 U3365 ( .A(n3389), .B(n3390), .Z(n3303) );
  NAND2_X1 U3366 ( .A1(n3391), .A2(n3392), .ZN(n3389) );
  NOR2_X1 U3367 ( .A1(n3305), .A2(n2265), .ZN(n3385) );
  NOR2_X1 U3368 ( .A1(n3177), .A2(n2663), .ZN(n2265) );
  NAND2_X1 U3369 ( .A1(n3258), .A2(n3393), .ZN(n3305) );
  NAND2_X1 U3370 ( .A1(n3257), .A2(n3259), .ZN(n3393) );
  NAND2_X1 U3371 ( .A1(n3394), .A2(n3395), .ZN(n3259) );
  NAND2_X1 U3372 ( .A1(a_9_), .A2(b_8_), .ZN(n3395) );
  INV_X1 U3373 ( .A(n3396), .ZN(n3394) );
  XNOR2_X1 U3374 ( .A(n3397), .B(n3398), .ZN(n3257) );
  NAND2_X1 U3375 ( .A1(n3399), .A2(n3400), .ZN(n3397) );
  NAND2_X1 U3376 ( .A1(a_9_), .A2(n3396), .ZN(n3258) );
  NAND2_X1 U3377 ( .A1(n3266), .A2(n3401), .ZN(n3396) );
  NAND2_X1 U3378 ( .A1(n3265), .A2(n3267), .ZN(n3401) );
  NAND2_X1 U3379 ( .A1(n3402), .A2(n3403), .ZN(n3267) );
  NAND2_X1 U3380 ( .A1(a_10_), .A2(b_8_), .ZN(n3403) );
  INV_X1 U3381 ( .A(n3404), .ZN(n3402) );
  XNOR2_X1 U3382 ( .A(n3405), .B(n3406), .ZN(n3265) );
  XOR2_X1 U3383 ( .A(n3407), .B(n3408), .Z(n3405) );
  NAND2_X1 U3384 ( .A1(a_11_), .A2(b_7_), .ZN(n3407) );
  NAND2_X1 U3385 ( .A1(a_10_), .A2(n3404), .ZN(n3266) );
  NAND2_X1 U3386 ( .A1(n3409), .A2(n3410), .ZN(n3404) );
  NAND3_X1 U3387 ( .A1(b_8_), .A2(n3411), .A3(a_11_), .ZN(n3410) );
  NAND2_X1 U3388 ( .A1(n3273), .A2(n3275), .ZN(n3411) );
  INV_X1 U3389 ( .A(n3412), .ZN(n3409) );
  NOR2_X1 U3390 ( .A1(n3273), .A2(n3275), .ZN(n3412) );
  NOR2_X1 U3391 ( .A1(n3413), .A2(n3414), .ZN(n3275) );
  INV_X1 U3392 ( .A(n3415), .ZN(n3414) );
  NAND2_X1 U3393 ( .A1(n3301), .A2(n3416), .ZN(n3415) );
  NAND2_X1 U3394 ( .A1(n3302), .A2(n3300), .ZN(n3416) );
  NOR2_X1 U3395 ( .A1(n3177), .A2(n2211), .ZN(n3301) );
  NOR2_X1 U3396 ( .A1(n3300), .A2(n3302), .ZN(n3413) );
  NOR2_X1 U3397 ( .A1(n3417), .A2(n3418), .ZN(n3302) );
  INV_X1 U3398 ( .A(n3419), .ZN(n3418) );
  NAND2_X1 U3399 ( .A1(n3296), .A2(n3420), .ZN(n3419) );
  NAND2_X1 U3400 ( .A1(n3421), .A2(n3298), .ZN(n3420) );
  NOR2_X1 U3401 ( .A1(n3177), .A2(n2191), .ZN(n3296) );
  INV_X1 U3402 ( .A(b_8_), .ZN(n3177) );
  NOR2_X1 U3403 ( .A1(n3298), .A2(n3421), .ZN(n3417) );
  INV_X1 U3404 ( .A(n3297), .ZN(n3421) );
  NAND2_X1 U3405 ( .A1(n3422), .A2(n3423), .ZN(n3297) );
  NAND2_X1 U3406 ( .A1(b_6_), .A2(n3424), .ZN(n3423) );
  NAND2_X1 U3407 ( .A1(n2170), .A2(n3425), .ZN(n3424) );
  NAND2_X1 U3408 ( .A1(a_15_), .A2(n2282), .ZN(n3425) );
  NAND2_X1 U3409 ( .A1(b_7_), .A2(n3426), .ZN(n3422) );
  NAND2_X1 U3410 ( .A1(n2173), .A2(n3427), .ZN(n3426) );
  NAND2_X1 U3411 ( .A1(a_14_), .A2(n2421), .ZN(n3427) );
  NAND3_X1 U3412 ( .A1(b_8_), .A2(n2416), .A3(b_7_), .ZN(n3298) );
  XNOR2_X1 U3413 ( .A(n3428), .B(n3429), .ZN(n3300) );
  XNOR2_X1 U3414 ( .A(n3430), .B(n3431), .ZN(n3428) );
  XOR2_X1 U3415 ( .A(n3432), .B(n3433), .Z(n3273) );
  XNOR2_X1 U3416 ( .A(n3434), .B(n3435), .ZN(n3432) );
  XNOR2_X1 U3417 ( .A(n3436), .B(n3437), .ZN(n3311) );
  XOR2_X1 U3418 ( .A(n3438), .B(n2397), .Z(n3436) );
  XOR2_X1 U3419 ( .A(n3439), .B(n3440), .Z(n3235) );
  XOR2_X1 U3420 ( .A(n3441), .B(n3442), .Z(n3440) );
  NAND2_X1 U3421 ( .A1(b_7_), .A2(a_6_), .ZN(n3442) );
  XOR2_X1 U3422 ( .A(n3443), .B(n3444), .Z(n3315) );
  XNOR2_X1 U3423 ( .A(n3445), .B(n3446), .ZN(n3444) );
  NAND2_X1 U3424 ( .A1(b_7_), .A2(a_5_), .ZN(n3446) );
  XOR2_X1 U3425 ( .A(n3447), .B(n3448), .Z(n3327) );
  XNOR2_X1 U3426 ( .A(n3449), .B(n3450), .ZN(n3448) );
  NAND2_X1 U3427 ( .A1(a_2_), .A2(b_7_), .ZN(n3450) );
  XNOR2_X1 U3428 ( .A(n3451), .B(n3452), .ZN(n3330) );
  XNOR2_X1 U3429 ( .A(n3453), .B(n3454), .ZN(n3451) );
  NOR2_X1 U3430 ( .A1(n2282), .A2(n2427), .ZN(n3454) );
  XNOR2_X1 U3431 ( .A(n3455), .B(n3456), .ZN(n2134) );
  XNOR2_X1 U3432 ( .A(n3457), .B(n3458), .ZN(n3456) );
  NAND2_X1 U3433 ( .A1(a_0_), .A2(b_7_), .ZN(n3458) );
  NAND2_X1 U3434 ( .A1(n3459), .A2(n3337), .ZN(n2473) );
  NAND2_X1 U3435 ( .A1(n3460), .A2(n3461), .ZN(n3337) );
  NAND3_X1 U3436 ( .A1(b_7_), .A2(n3462), .A3(a_0_), .ZN(n3461) );
  NAND2_X1 U3437 ( .A1(n3457), .A2(n3455), .ZN(n3462) );
  INV_X1 U3438 ( .A(n3463), .ZN(n3460) );
  NOR2_X1 U3439 ( .A1(n3455), .A2(n3457), .ZN(n3463) );
  NOR2_X1 U3440 ( .A1(n3464), .A2(n3465), .ZN(n3457) );
  INV_X1 U3441 ( .A(n3466), .ZN(n3465) );
  NAND3_X1 U3442 ( .A1(b_7_), .A2(n3467), .A3(a_1_), .ZN(n3466) );
  NAND2_X1 U3443 ( .A1(n3453), .A2(n3452), .ZN(n3467) );
  NOR2_X1 U3444 ( .A1(n3452), .A2(n3453), .ZN(n3464) );
  NOR2_X1 U3445 ( .A1(n3468), .A2(n3469), .ZN(n3453) );
  INV_X1 U3446 ( .A(n3470), .ZN(n3469) );
  NAND3_X1 U3447 ( .A1(b_7_), .A2(n3471), .A3(a_2_), .ZN(n3470) );
  NAND2_X1 U3448 ( .A1(n3447), .A2(n3449), .ZN(n3471) );
  NOR2_X1 U3449 ( .A1(n3447), .A2(n3449), .ZN(n3468) );
  NOR2_X1 U3450 ( .A1(n3472), .A2(n3473), .ZN(n3449) );
  INV_X1 U3451 ( .A(n3474), .ZN(n3473) );
  NAND3_X1 U3452 ( .A1(b_7_), .A2(n3475), .A3(a_3_), .ZN(n3474) );
  NAND2_X1 U3453 ( .A1(n3354), .A2(n3353), .ZN(n3475) );
  NOR2_X1 U3454 ( .A1(n3353), .A2(n3354), .ZN(n3472) );
  NOR2_X1 U3455 ( .A1(n3476), .A2(n3477), .ZN(n3354) );
  INV_X1 U3456 ( .A(n3478), .ZN(n3477) );
  NAND3_X1 U3457 ( .A1(b_7_), .A2(n3479), .A3(a_4_), .ZN(n3478) );
  NAND2_X1 U3458 ( .A1(n3361), .A2(n3359), .ZN(n3479) );
  NOR2_X1 U3459 ( .A1(n3359), .A2(n3361), .ZN(n3476) );
  NOR2_X1 U3460 ( .A1(n3480), .A2(n3481), .ZN(n3361) );
  INV_X1 U3461 ( .A(n3482), .ZN(n3481) );
  NAND3_X1 U3462 ( .A1(a_5_), .A2(n3483), .A3(b_7_), .ZN(n3482) );
  NAND2_X1 U3463 ( .A1(n3445), .A2(n3443), .ZN(n3483) );
  NOR2_X1 U3464 ( .A1(n3443), .A2(n3445), .ZN(n3480) );
  NOR2_X1 U3465 ( .A1(n3484), .A2(n3485), .ZN(n3445) );
  INV_X1 U3466 ( .A(n3486), .ZN(n3485) );
  NAND3_X1 U3467 ( .A1(a_6_), .A2(n3487), .A3(b_7_), .ZN(n3486) );
  NAND2_X1 U3468 ( .A1(n3439), .A2(n3441), .ZN(n3487) );
  NOR2_X1 U3469 ( .A1(n3441), .A2(n3439), .ZN(n3484) );
  XOR2_X1 U3470 ( .A(n3488), .B(n3489), .Z(n3439) );
  XNOR2_X1 U3471 ( .A(n3490), .B(n3491), .ZN(n3489) );
  NAND2_X1 U3472 ( .A1(n3492), .A2(n3493), .ZN(n3441) );
  NAND2_X1 U3473 ( .A1(n3437), .A2(n3494), .ZN(n3493) );
  NAND2_X1 U3474 ( .A1(n2277), .A2(n3495), .ZN(n3494) );
  INV_X1 U3475 ( .A(n3438), .ZN(n3495) );
  INV_X1 U3476 ( .A(n2397), .ZN(n2277) );
  XOR2_X1 U3477 ( .A(n3496), .B(n3497), .Z(n3437) );
  XOR2_X1 U3478 ( .A(n3498), .B(n3499), .Z(n3497) );
  NAND2_X1 U3479 ( .A1(b_6_), .A2(a_8_), .ZN(n3499) );
  NAND2_X1 U3480 ( .A1(n3438), .A2(n2397), .ZN(n3492) );
  NAND2_X1 U3481 ( .A1(a_7_), .A2(b_7_), .ZN(n2397) );
  NOR2_X1 U3482 ( .A1(n3500), .A2(n3501), .ZN(n3438) );
  NOR2_X1 U3483 ( .A1(n3384), .A2(n3502), .ZN(n3501) );
  NOR2_X1 U3484 ( .A1(n3383), .A2(n3381), .ZN(n3502) );
  NAND2_X1 U3485 ( .A1(b_7_), .A2(a_8_), .ZN(n3384) );
  INV_X1 U3486 ( .A(n3503), .ZN(n3500) );
  NAND2_X1 U3487 ( .A1(n3381), .A2(n3383), .ZN(n3503) );
  NAND2_X1 U3488 ( .A1(n3391), .A2(n3504), .ZN(n3383) );
  NAND2_X1 U3489 ( .A1(n3390), .A2(n3392), .ZN(n3504) );
  NAND2_X1 U3490 ( .A1(n3505), .A2(n3506), .ZN(n3392) );
  NAND2_X1 U3491 ( .A1(a_9_), .A2(b_7_), .ZN(n3506) );
  INV_X1 U3492 ( .A(n3507), .ZN(n3505) );
  XNOR2_X1 U3493 ( .A(n3508), .B(n3509), .ZN(n3390) );
  NAND2_X1 U3494 ( .A1(n3510), .A2(n3511), .ZN(n3508) );
  NAND2_X1 U3495 ( .A1(a_9_), .A2(n3507), .ZN(n3391) );
  NAND2_X1 U3496 ( .A1(n3399), .A2(n3512), .ZN(n3507) );
  NAND2_X1 U3497 ( .A1(n3398), .A2(n3400), .ZN(n3512) );
  NAND2_X1 U3498 ( .A1(n3513), .A2(n3514), .ZN(n3400) );
  NAND2_X1 U3499 ( .A1(a_10_), .A2(b_7_), .ZN(n3514) );
  INV_X1 U3500 ( .A(n3515), .ZN(n3513) );
  XNOR2_X1 U3501 ( .A(n3516), .B(n3517), .ZN(n3398) );
  XOR2_X1 U3502 ( .A(n3518), .B(n3519), .Z(n3516) );
  NAND2_X1 U3503 ( .A1(a_11_), .A2(b_6_), .ZN(n3518) );
  NAND2_X1 U3504 ( .A1(a_10_), .A2(n3515), .ZN(n3399) );
  NAND2_X1 U3505 ( .A1(n3520), .A2(n3521), .ZN(n3515) );
  NAND3_X1 U3506 ( .A1(b_7_), .A2(n3522), .A3(a_11_), .ZN(n3521) );
  NAND2_X1 U3507 ( .A1(n3406), .A2(n3408), .ZN(n3522) );
  INV_X1 U3508 ( .A(n3523), .ZN(n3520) );
  NOR2_X1 U3509 ( .A1(n3406), .A2(n3408), .ZN(n3523) );
  NOR2_X1 U3510 ( .A1(n3524), .A2(n3525), .ZN(n3408) );
  INV_X1 U3511 ( .A(n3526), .ZN(n3525) );
  NAND2_X1 U3512 ( .A1(n3434), .A2(n3527), .ZN(n3526) );
  NAND2_X1 U3513 ( .A1(n3435), .A2(n3433), .ZN(n3527) );
  NOR2_X1 U3514 ( .A1(n2282), .A2(n2211), .ZN(n3434) );
  NOR2_X1 U3515 ( .A1(n3433), .A2(n3435), .ZN(n3524) );
  NOR2_X1 U3516 ( .A1(n3528), .A2(n3529), .ZN(n3435) );
  INV_X1 U3517 ( .A(n3530), .ZN(n3529) );
  NAND2_X1 U3518 ( .A1(n3429), .A2(n3531), .ZN(n3530) );
  NAND2_X1 U3519 ( .A1(n3532), .A2(n3431), .ZN(n3531) );
  NOR2_X1 U3520 ( .A1(n2282), .A2(n2191), .ZN(n3429) );
  INV_X1 U3521 ( .A(b_7_), .ZN(n2282) );
  NOR2_X1 U3522 ( .A1(n3431), .A2(n3532), .ZN(n3528) );
  INV_X1 U3523 ( .A(n3430), .ZN(n3532) );
  NAND2_X1 U3524 ( .A1(n3533), .A2(n3534), .ZN(n3430) );
  NAND2_X1 U3525 ( .A1(b_5_), .A2(n3535), .ZN(n3534) );
  NAND2_X1 U3526 ( .A1(n2170), .A2(n3536), .ZN(n3535) );
  NAND2_X1 U3527 ( .A1(a_15_), .A2(n2421), .ZN(n3536) );
  NAND2_X1 U3528 ( .A1(b_6_), .A2(n3537), .ZN(n3533) );
  NAND2_X1 U3529 ( .A1(n2173), .A2(n3538), .ZN(n3537) );
  NAND2_X1 U3530 ( .A1(a_14_), .A2(n2311), .ZN(n3538) );
  NAND3_X1 U3531 ( .A1(b_7_), .A2(n2416), .A3(b_6_), .ZN(n3431) );
  XNOR2_X1 U3532 ( .A(n3539), .B(n3540), .ZN(n3433) );
  XNOR2_X1 U3533 ( .A(n3541), .B(n3542), .ZN(n3539) );
  XOR2_X1 U3534 ( .A(n3543), .B(n3544), .Z(n3406) );
  XNOR2_X1 U3535 ( .A(n3545), .B(n3546), .ZN(n3543) );
  XNOR2_X1 U3536 ( .A(n3547), .B(n3548), .ZN(n3381) );
  NAND2_X1 U3537 ( .A1(n3549), .A2(n3550), .ZN(n3547) );
  XOR2_X1 U3538 ( .A(n3551), .B(n3552), .Z(n3443) );
  XNOR2_X1 U3539 ( .A(n3553), .B(n2294), .ZN(n3551) );
  XNOR2_X1 U3540 ( .A(n3554), .B(n3555), .ZN(n3359) );
  XOR2_X1 U3541 ( .A(n3556), .B(n3557), .Z(n3554) );
  XNOR2_X1 U3542 ( .A(n3558), .B(n3559), .ZN(n3353) );
  XOR2_X1 U3543 ( .A(n3560), .B(n3561), .Z(n3558) );
  XOR2_X1 U3544 ( .A(n3562), .B(n3563), .Z(n3447) );
  XNOR2_X1 U3545 ( .A(n3564), .B(n3565), .ZN(n3563) );
  XOR2_X1 U3546 ( .A(n3566), .B(n3567), .Z(n3452) );
  XNOR2_X1 U3547 ( .A(n3568), .B(n3569), .ZN(n3567) );
  XNOR2_X1 U3548 ( .A(n3570), .B(n3571), .ZN(n3455) );
  XOR2_X1 U3549 ( .A(n3572), .B(n3573), .Z(n3570) );
  XNOR2_X1 U3550 ( .A(n3339), .B(n3338), .ZN(n3459) );
  XNOR2_X1 U3551 ( .A(n3574), .B(n3575), .ZN(n3338) );
  XNOR2_X1 U3552 ( .A(n3576), .B(n2146), .ZN(n2137) );
  INV_X1 U3553 ( .A(n2141), .ZN(n2470) );
  NOR3_X1 U3554 ( .A1(n2146), .A2(n2145), .A3(n2472), .ZN(n2141) );
  NAND2_X1 U3555 ( .A1(n3577), .A2(n2469), .ZN(n2472) );
  NAND2_X1 U3556 ( .A1(n3578), .A2(n3579), .ZN(n3577) );
  INV_X1 U3557 ( .A(n3580), .ZN(n3579) );
  XNOR2_X1 U3558 ( .A(n3581), .B(n3582), .ZN(n3578) );
  INV_X1 U3559 ( .A(n3576), .ZN(n2145) );
  NAND2_X1 U3560 ( .A1(n3583), .A2(n3584), .ZN(n3576) );
  NAND2_X1 U3561 ( .A1(n3575), .A2(n3585), .ZN(n3584) );
  INV_X1 U3562 ( .A(n3586), .ZN(n3585) );
  NOR2_X1 U3563 ( .A1(n3574), .A2(n3339), .ZN(n3586) );
  NOR2_X1 U3564 ( .A1(n2433), .A2(n2421), .ZN(n3575) );
  NAND2_X1 U3565 ( .A1(n3339), .A2(n3574), .ZN(n3583) );
  NAND2_X1 U3566 ( .A1(n3587), .A2(n3588), .ZN(n3574) );
  NAND2_X1 U3567 ( .A1(n3573), .A2(n3589), .ZN(n3588) );
  INV_X1 U3568 ( .A(n3590), .ZN(n3589) );
  NOR2_X1 U3569 ( .A1(n3571), .A2(n3572), .ZN(n3590) );
  NOR2_X1 U3570 ( .A1(n2427), .A2(n2421), .ZN(n3573) );
  NAND2_X1 U3571 ( .A1(n3571), .A2(n3572), .ZN(n3587) );
  NAND2_X1 U3572 ( .A1(n3591), .A2(n3592), .ZN(n3572) );
  NAND2_X1 U3573 ( .A1(n3569), .A2(n3593), .ZN(n3592) );
  INV_X1 U3574 ( .A(n3594), .ZN(n3593) );
  NOR2_X1 U3575 ( .A1(n3566), .A2(n3568), .ZN(n3594) );
  NOR2_X1 U3576 ( .A1(n2426), .A2(n2421), .ZN(n3569) );
  NAND2_X1 U3577 ( .A1(n3566), .A2(n3568), .ZN(n3591) );
  NAND2_X1 U3578 ( .A1(n3595), .A2(n3596), .ZN(n3568) );
  NAND2_X1 U3579 ( .A1(n3565), .A2(n3597), .ZN(n3596) );
  INV_X1 U3580 ( .A(n3598), .ZN(n3597) );
  NOR2_X1 U3581 ( .A1(n3564), .A2(n3562), .ZN(n3598) );
  NOR2_X1 U3582 ( .A1(n2344), .A2(n2421), .ZN(n3565) );
  NAND2_X1 U3583 ( .A1(n3562), .A2(n3564), .ZN(n3595) );
  NAND2_X1 U3584 ( .A1(n3599), .A2(n3600), .ZN(n3564) );
  NAND2_X1 U3585 ( .A1(n3561), .A2(n3601), .ZN(n3600) );
  INV_X1 U3586 ( .A(n3602), .ZN(n3601) );
  NOR2_X1 U3587 ( .A1(n3559), .A2(n3560), .ZN(n3602) );
  NOR2_X1 U3588 ( .A1(n2424), .A2(n2421), .ZN(n3561) );
  NAND2_X1 U3589 ( .A1(n3559), .A2(n3560), .ZN(n3599) );
  NAND2_X1 U3590 ( .A1(n3603), .A2(n3604), .ZN(n3560) );
  NAND2_X1 U3591 ( .A1(n3557), .A2(n3605), .ZN(n3604) );
  NAND2_X1 U3592 ( .A1(n3555), .A2(n3556), .ZN(n3605) );
  NOR2_X1 U3593 ( .A1(n2421), .A2(n2309), .ZN(n3557) );
  INV_X1 U3594 ( .A(n3606), .ZN(n3603) );
  NOR2_X1 U3595 ( .A1(n3555), .A2(n3556), .ZN(n3606) );
  NAND2_X1 U3596 ( .A1(n3607), .A2(n3608), .ZN(n3556) );
  NAND2_X1 U3597 ( .A1(n3552), .A2(n3609), .ZN(n3608) );
  NAND2_X1 U3598 ( .A1(n3610), .A2(n3553), .ZN(n3609) );
  INV_X1 U3599 ( .A(n2294), .ZN(n3610) );
  XNOR2_X1 U3600 ( .A(n3611), .B(n3612), .ZN(n3552) );
  XNOR2_X1 U3601 ( .A(n3613), .B(n3614), .ZN(n3612) );
  NAND2_X1 U3602 ( .A1(a_7_), .A2(b_5_), .ZN(n3614) );
  NAND2_X1 U3603 ( .A1(n3615), .A2(n2294), .ZN(n3607) );
  NAND2_X1 U3604 ( .A1(b_6_), .A2(a_6_), .ZN(n2294) );
  INV_X1 U3605 ( .A(n3553), .ZN(n3615) );
  NAND2_X1 U3606 ( .A1(n3616), .A2(n3617), .ZN(n3553) );
  NAND2_X1 U3607 ( .A1(n3491), .A2(n3618), .ZN(n3617) );
  INV_X1 U3608 ( .A(n3619), .ZN(n3618) );
  NOR2_X1 U3609 ( .A1(n3490), .A2(n3488), .ZN(n3619) );
  NOR2_X1 U3610 ( .A1(n2280), .A2(n2421), .ZN(n3491) );
  NAND2_X1 U3611 ( .A1(n3488), .A2(n3490), .ZN(n3616) );
  NAND2_X1 U3612 ( .A1(n3620), .A2(n3621), .ZN(n3490) );
  INV_X1 U3613 ( .A(n3622), .ZN(n3621) );
  NOR3_X1 U3614 ( .A1(n2663), .A2(n3623), .A3(n2421), .ZN(n3622) );
  NOR2_X1 U3615 ( .A1(n3498), .A2(n3496), .ZN(n3623) );
  NAND2_X1 U3616 ( .A1(n3496), .A2(n3498), .ZN(n3620) );
  NAND2_X1 U3617 ( .A1(n3549), .A2(n3624), .ZN(n3498) );
  NAND2_X1 U3618 ( .A1(n3548), .A2(n3550), .ZN(n3624) );
  NAND2_X1 U3619 ( .A1(n3625), .A2(n3626), .ZN(n3550) );
  NAND2_X1 U3620 ( .A1(a_9_), .A2(b_6_), .ZN(n3626) );
  INV_X1 U3621 ( .A(n3627), .ZN(n3625) );
  XNOR2_X1 U3622 ( .A(n3628), .B(n3629), .ZN(n3548) );
  NAND2_X1 U3623 ( .A1(n3630), .A2(n3631), .ZN(n3628) );
  NAND2_X1 U3624 ( .A1(a_9_), .A2(n3627), .ZN(n3549) );
  NAND2_X1 U3625 ( .A1(n3510), .A2(n3632), .ZN(n3627) );
  NAND2_X1 U3626 ( .A1(n3509), .A2(n3511), .ZN(n3632) );
  NAND2_X1 U3627 ( .A1(n3633), .A2(n3634), .ZN(n3511) );
  NAND2_X1 U3628 ( .A1(a_10_), .A2(b_6_), .ZN(n3634) );
  INV_X1 U3629 ( .A(n3635), .ZN(n3633) );
  XNOR2_X1 U3630 ( .A(n3636), .B(n3637), .ZN(n3509) );
  XOR2_X1 U3631 ( .A(n3638), .B(n3639), .Z(n3636) );
  NAND2_X1 U3632 ( .A1(a_11_), .A2(b_5_), .ZN(n3638) );
  NAND2_X1 U3633 ( .A1(a_10_), .A2(n3635), .ZN(n3510) );
  NAND2_X1 U3634 ( .A1(n3640), .A2(n3641), .ZN(n3635) );
  NAND3_X1 U3635 ( .A1(b_6_), .A2(n3642), .A3(a_11_), .ZN(n3641) );
  NAND2_X1 U3636 ( .A1(n3517), .A2(n3519), .ZN(n3642) );
  INV_X1 U3637 ( .A(n3643), .ZN(n3640) );
  NOR2_X1 U3638 ( .A1(n3517), .A2(n3519), .ZN(n3643) );
  NOR2_X1 U3639 ( .A1(n3644), .A2(n3645), .ZN(n3519) );
  INV_X1 U3640 ( .A(n3646), .ZN(n3645) );
  NAND2_X1 U3641 ( .A1(n3545), .A2(n3647), .ZN(n3646) );
  NAND2_X1 U3642 ( .A1(n3546), .A2(n3544), .ZN(n3647) );
  NOR2_X1 U3643 ( .A1(n2421), .A2(n2211), .ZN(n3545) );
  NOR2_X1 U3644 ( .A1(n3544), .A2(n3546), .ZN(n3644) );
  NOR2_X1 U3645 ( .A1(n3648), .A2(n3649), .ZN(n3546) );
  INV_X1 U3646 ( .A(n3650), .ZN(n3649) );
  NAND2_X1 U3647 ( .A1(n3540), .A2(n3651), .ZN(n3650) );
  NAND2_X1 U3648 ( .A1(n3652), .A2(n3542), .ZN(n3651) );
  NOR2_X1 U3649 ( .A1(n2421), .A2(n2191), .ZN(n3540) );
  INV_X1 U3650 ( .A(b_6_), .ZN(n2421) );
  NOR2_X1 U3651 ( .A1(n3542), .A2(n3652), .ZN(n3648) );
  INV_X1 U3652 ( .A(n3541), .ZN(n3652) );
  NAND2_X1 U3653 ( .A1(n3653), .A2(n3654), .ZN(n3541) );
  NAND2_X1 U3654 ( .A1(b_4_), .A2(n3655), .ZN(n3654) );
  NAND2_X1 U3655 ( .A1(n2170), .A2(n3656), .ZN(n3655) );
  NAND2_X1 U3656 ( .A1(a_15_), .A2(n2311), .ZN(n3656) );
  NAND2_X1 U3657 ( .A1(b_5_), .A2(n3657), .ZN(n3653) );
  NAND2_X1 U3658 ( .A1(n2173), .A2(n3658), .ZN(n3657) );
  NAND2_X1 U3659 ( .A1(a_14_), .A2(n2423), .ZN(n3658) );
  NAND3_X1 U3660 ( .A1(b_6_), .A2(n2416), .A3(b_5_), .ZN(n3542) );
  XNOR2_X1 U3661 ( .A(n3659), .B(n3660), .ZN(n3544) );
  XNOR2_X1 U3662 ( .A(n3661), .B(n3662), .ZN(n3659) );
  XOR2_X1 U3663 ( .A(n3663), .B(n3664), .Z(n3517) );
  XNOR2_X1 U3664 ( .A(n3665), .B(n3666), .ZN(n3663) );
  XNOR2_X1 U3665 ( .A(n3667), .B(n3668), .ZN(n3496) );
  NAND2_X1 U3666 ( .A1(n3669), .A2(n3670), .ZN(n3667) );
  XNOR2_X1 U3667 ( .A(n3671), .B(n3672), .ZN(n3488) );
  XOR2_X1 U3668 ( .A(n3673), .B(n3674), .Z(n3672) );
  NAND2_X1 U3669 ( .A1(b_5_), .A2(a_8_), .ZN(n3674) );
  XNOR2_X1 U3670 ( .A(n3675), .B(n3676), .ZN(n3555) );
  XNOR2_X1 U3671 ( .A(n3677), .B(n3678), .ZN(n3676) );
  NAND2_X1 U3672 ( .A1(b_5_), .A2(a_6_), .ZN(n3678) );
  XOR2_X1 U3673 ( .A(n3679), .B(n3680), .Z(n3559) );
  XOR2_X1 U3674 ( .A(n3681), .B(n2307), .Z(n3679) );
  XNOR2_X1 U3675 ( .A(n3682), .B(n3683), .ZN(n3562) );
  XNOR2_X1 U3676 ( .A(n3684), .B(n3685), .ZN(n3682) );
  NOR2_X1 U3677 ( .A1(n2311), .A2(n2424), .ZN(n3685) );
  XNOR2_X1 U3678 ( .A(n3686), .B(n3687), .ZN(n3566) );
  XNOR2_X1 U3679 ( .A(n3688), .B(n3689), .ZN(n3686) );
  NOR2_X1 U3680 ( .A1(n2311), .A2(n2344), .ZN(n3689) );
  XNOR2_X1 U3681 ( .A(n3690), .B(n3691), .ZN(n3571) );
  XNOR2_X1 U3682 ( .A(n3692), .B(n3693), .ZN(n3690) );
  NOR2_X1 U3683 ( .A1(n2311), .A2(n2426), .ZN(n3693) );
  XNOR2_X1 U3684 ( .A(n3694), .B(n3695), .ZN(n3339) );
  XNOR2_X1 U3685 ( .A(n3696), .B(n3697), .ZN(n3694) );
  NOR2_X1 U3686 ( .A1(n2311), .A2(n2427), .ZN(n3697) );
  XOR2_X1 U3687 ( .A(n3698), .B(n3699), .Z(n2146) );
  XNOR2_X1 U3688 ( .A(n3700), .B(n3701), .ZN(n3698) );
  NOR2_X1 U3689 ( .A1(n2311), .A2(n2433), .ZN(n3701) );
  NAND2_X1 U3690 ( .A1(n3702), .A2(n3580), .ZN(n2469) );
  NAND2_X1 U3691 ( .A1(n3703), .A2(n3704), .ZN(n3580) );
  NAND3_X1 U3692 ( .A1(b_5_), .A2(n3705), .A3(a_0_), .ZN(n3704) );
  NAND2_X1 U3693 ( .A1(n3700), .A2(n3699), .ZN(n3705) );
  INV_X1 U3694 ( .A(n3706), .ZN(n3703) );
  NOR2_X1 U3695 ( .A1(n3699), .A2(n3700), .ZN(n3706) );
  NOR2_X1 U3696 ( .A1(n3707), .A2(n3708), .ZN(n3700) );
  INV_X1 U3697 ( .A(n3709), .ZN(n3708) );
  NAND3_X1 U3698 ( .A1(b_5_), .A2(n3710), .A3(a_1_), .ZN(n3709) );
  NAND2_X1 U3699 ( .A1(n3695), .A2(n3696), .ZN(n3710) );
  NOR2_X1 U3700 ( .A1(n3695), .A2(n3696), .ZN(n3707) );
  NOR2_X1 U3701 ( .A1(n3711), .A2(n3712), .ZN(n3696) );
  INV_X1 U3702 ( .A(n3713), .ZN(n3712) );
  NAND3_X1 U3703 ( .A1(b_5_), .A2(n3714), .A3(a_2_), .ZN(n3713) );
  NAND2_X1 U3704 ( .A1(n3692), .A2(n3691), .ZN(n3714) );
  NOR2_X1 U3705 ( .A1(n3691), .A2(n3692), .ZN(n3711) );
  NOR2_X1 U3706 ( .A1(n3715), .A2(n3716), .ZN(n3692) );
  INV_X1 U3707 ( .A(n3717), .ZN(n3716) );
  NAND3_X1 U3708 ( .A1(b_5_), .A2(n3718), .A3(a_3_), .ZN(n3717) );
  NAND2_X1 U3709 ( .A1(n3688), .A2(n3687), .ZN(n3718) );
  NOR2_X1 U3710 ( .A1(n3687), .A2(n3688), .ZN(n3715) );
  NOR2_X1 U3711 ( .A1(n3719), .A2(n3720), .ZN(n3688) );
  INV_X1 U3712 ( .A(n3721), .ZN(n3720) );
  NAND3_X1 U3713 ( .A1(b_5_), .A2(n3722), .A3(a_4_), .ZN(n3721) );
  NAND2_X1 U3714 ( .A1(n3683), .A2(n3684), .ZN(n3722) );
  NOR2_X1 U3715 ( .A1(n3683), .A2(n3684), .ZN(n3719) );
  NOR2_X1 U3716 ( .A1(n3723), .A2(n3724), .ZN(n3684) );
  INV_X1 U3717 ( .A(n3725), .ZN(n3724) );
  NAND2_X1 U3718 ( .A1(n3680), .A2(n3726), .ZN(n3725) );
  NAND2_X1 U3719 ( .A1(n3681), .A2(n2307), .ZN(n3726) );
  XNOR2_X1 U3720 ( .A(n3727), .B(n3728), .ZN(n3680) );
  XNOR2_X1 U3721 ( .A(n3729), .B(n3730), .ZN(n3727) );
  NOR2_X1 U3722 ( .A1(n2307), .A2(n3681), .ZN(n3723) );
  NOR2_X1 U3723 ( .A1(n3731), .A2(n3732), .ZN(n3681) );
  INV_X1 U3724 ( .A(n3733), .ZN(n3732) );
  NAND3_X1 U3725 ( .A1(a_6_), .A2(n3734), .A3(b_5_), .ZN(n3733) );
  NAND2_X1 U3726 ( .A1(n3675), .A2(n3677), .ZN(n3734) );
  NOR2_X1 U3727 ( .A1(n3675), .A2(n3677), .ZN(n3731) );
  NOR2_X1 U3728 ( .A1(n3735), .A2(n3736), .ZN(n3677) );
  INV_X1 U3729 ( .A(n3737), .ZN(n3736) );
  NAND3_X1 U3730 ( .A1(b_5_), .A2(n3738), .A3(a_7_), .ZN(n3737) );
  NAND2_X1 U3731 ( .A1(n3613), .A2(n3611), .ZN(n3738) );
  NOR2_X1 U3732 ( .A1(n3611), .A2(n3613), .ZN(n3735) );
  NOR2_X1 U3733 ( .A1(n3739), .A2(n3740), .ZN(n3613) );
  NOR3_X1 U3734 ( .A1(n2663), .A2(n3741), .A3(n2311), .ZN(n3740) );
  NOR2_X1 U3735 ( .A1(n3671), .A2(n3673), .ZN(n3741) );
  INV_X1 U3736 ( .A(n3742), .ZN(n3739) );
  NAND2_X1 U3737 ( .A1(n3671), .A2(n3673), .ZN(n3742) );
  NAND2_X1 U3738 ( .A1(n3669), .A2(n3743), .ZN(n3673) );
  NAND2_X1 U3739 ( .A1(n3668), .A2(n3670), .ZN(n3743) );
  NAND2_X1 U3740 ( .A1(n3744), .A2(n3745), .ZN(n3670) );
  NAND2_X1 U3741 ( .A1(a_9_), .A2(b_5_), .ZN(n3745) );
  INV_X1 U3742 ( .A(n3746), .ZN(n3744) );
  XOR2_X1 U3743 ( .A(n3747), .B(n3748), .Z(n3668) );
  XNOR2_X1 U3744 ( .A(n3749), .B(n3750), .ZN(n3748) );
  NAND2_X1 U3745 ( .A1(a_9_), .A2(n3746), .ZN(n3669) );
  NAND2_X1 U3746 ( .A1(n3630), .A2(n3751), .ZN(n3746) );
  NAND2_X1 U3747 ( .A1(n3629), .A2(n3631), .ZN(n3751) );
  NAND2_X1 U3748 ( .A1(n3752), .A2(n3753), .ZN(n3631) );
  NAND2_X1 U3749 ( .A1(a_10_), .A2(b_5_), .ZN(n3753) );
  INV_X1 U3750 ( .A(n3754), .ZN(n3752) );
  XNOR2_X1 U3751 ( .A(n3755), .B(n3756), .ZN(n3629) );
  XOR2_X1 U3752 ( .A(n3757), .B(n3758), .Z(n3755) );
  NAND2_X1 U3753 ( .A1(b_4_), .A2(a_11_), .ZN(n3757) );
  NAND2_X1 U3754 ( .A1(a_10_), .A2(n3754), .ZN(n3630) );
  NAND2_X1 U3755 ( .A1(n3759), .A2(n3760), .ZN(n3754) );
  NAND3_X1 U3756 ( .A1(b_5_), .A2(n3761), .A3(a_11_), .ZN(n3760) );
  NAND2_X1 U3757 ( .A1(n3637), .A2(n3639), .ZN(n3761) );
  INV_X1 U3758 ( .A(n3762), .ZN(n3759) );
  NOR2_X1 U3759 ( .A1(n3637), .A2(n3639), .ZN(n3762) );
  NOR2_X1 U3760 ( .A1(n3763), .A2(n3764), .ZN(n3639) );
  INV_X1 U3761 ( .A(n3765), .ZN(n3764) );
  NAND2_X1 U3762 ( .A1(n3665), .A2(n3766), .ZN(n3765) );
  NAND2_X1 U3763 ( .A1(n3666), .A2(n3664), .ZN(n3766) );
  NOR2_X1 U3764 ( .A1(n2311), .A2(n2211), .ZN(n3665) );
  NOR2_X1 U3765 ( .A1(n3664), .A2(n3666), .ZN(n3763) );
  NOR2_X1 U3766 ( .A1(n3767), .A2(n3768), .ZN(n3666) );
  INV_X1 U3767 ( .A(n3769), .ZN(n3768) );
  NAND2_X1 U3768 ( .A1(n3660), .A2(n3770), .ZN(n3769) );
  NAND2_X1 U3769 ( .A1(n3771), .A2(n3662), .ZN(n3770) );
  NOR2_X1 U3770 ( .A1(n2311), .A2(n2191), .ZN(n3660) );
  INV_X1 U3771 ( .A(b_5_), .ZN(n2311) );
  NOR2_X1 U3772 ( .A1(n3662), .A2(n3771), .ZN(n3767) );
  INV_X1 U3773 ( .A(n3661), .ZN(n3771) );
  NAND2_X1 U3774 ( .A1(n3772), .A2(n3773), .ZN(n3661) );
  NAND2_X1 U3775 ( .A1(b_3_), .A2(n3774), .ZN(n3773) );
  NAND2_X1 U3776 ( .A1(n2170), .A2(n3775), .ZN(n3774) );
  NAND2_X1 U3777 ( .A1(a_15_), .A2(n2423), .ZN(n3775) );
  NAND2_X1 U3778 ( .A1(b_4_), .A2(n3776), .ZN(n3772) );
  NAND2_X1 U3779 ( .A1(n2173), .A2(n3777), .ZN(n3776) );
  NAND2_X1 U3780 ( .A1(a_14_), .A2(n2346), .ZN(n3777) );
  NAND3_X1 U3781 ( .A1(b_5_), .A2(n2416), .A3(b_4_), .ZN(n3662) );
  XNOR2_X1 U3782 ( .A(n3778), .B(n3779), .ZN(n3664) );
  XNOR2_X1 U3783 ( .A(n3780), .B(n3781), .ZN(n3778) );
  XOR2_X1 U3784 ( .A(n3782), .B(n3783), .Z(n3637) );
  XNOR2_X1 U3785 ( .A(n3784), .B(n3785), .ZN(n3782) );
  XNOR2_X1 U3786 ( .A(n3786), .B(n3787), .ZN(n3671) );
  XNOR2_X1 U3787 ( .A(n3788), .B(n3789), .ZN(n3787) );
  XOR2_X1 U3788 ( .A(n3790), .B(n3791), .Z(n3611) );
  XNOR2_X1 U3789 ( .A(n3792), .B(n3793), .ZN(n3790) );
  XOR2_X1 U3790 ( .A(n3794), .B(n3795), .Z(n3675) );
  XNOR2_X1 U3791 ( .A(n3796), .B(n3797), .ZN(n3794) );
  NAND2_X1 U3792 ( .A1(b_5_), .A2(a_5_), .ZN(n2307) );
  XOR2_X1 U3793 ( .A(n3798), .B(n3799), .Z(n3683) );
  XNOR2_X1 U3794 ( .A(n3800), .B(n3801), .ZN(n3798) );
  XNOR2_X1 U3795 ( .A(n3802), .B(n3803), .ZN(n3687) );
  XOR2_X1 U3796 ( .A(n3804), .B(n2324), .Z(n3802) );
  XNOR2_X1 U3797 ( .A(n3805), .B(n3806), .ZN(n3691) );
  XOR2_X1 U3798 ( .A(n3807), .B(n3808), .Z(n3806) );
  XNOR2_X1 U3799 ( .A(n3809), .B(n3810), .ZN(n3695) );
  XNOR2_X1 U3800 ( .A(n3811), .B(n3812), .ZN(n3810) );
  XOR2_X1 U3801 ( .A(n3813), .B(n3814), .Z(n3699) );
  XNOR2_X1 U3802 ( .A(n3815), .B(n3816), .ZN(n3813) );
  XNOR2_X1 U3803 ( .A(n3817), .B(n3582), .ZN(n3702) );
  XNOR2_X1 U3804 ( .A(n3818), .B(n3819), .ZN(n3582) );
  XNOR2_X1 U3805 ( .A(n3820), .B(n2158), .ZN(n2149) );
  INV_X1 U3806 ( .A(n2153), .ZN(n2466) );
  NOR3_X1 U3807 ( .A1(n2158), .A2(n2157), .A3(n2468), .ZN(n2153) );
  NAND2_X1 U3808 ( .A1(n3821), .A2(n2465), .ZN(n2468) );
  NAND2_X1 U3809 ( .A1(n3822), .A2(n3823), .ZN(n3821) );
  XOR2_X1 U3810 ( .A(n3824), .B(n3825), .Z(n3823) );
  INV_X1 U3811 ( .A(n3826), .ZN(n3822) );
  INV_X1 U3812 ( .A(n3820), .ZN(n2157) );
  NAND2_X1 U3813 ( .A1(n3827), .A2(n3828), .ZN(n3820) );
  NAND2_X1 U3814 ( .A1(n3819), .A2(n3829), .ZN(n3828) );
  NAND2_X1 U3815 ( .A1(n3830), .A2(n3581), .ZN(n3829) );
  NOR2_X1 U3816 ( .A1(n2433), .A2(n2423), .ZN(n3819) );
  NAND2_X1 U3817 ( .A1(n3817), .A2(n3818), .ZN(n3827) );
  INV_X1 U3818 ( .A(n3830), .ZN(n3818) );
  NOR2_X1 U3819 ( .A1(n3831), .A2(n3832), .ZN(n3830) );
  INV_X1 U3820 ( .A(n3833), .ZN(n3832) );
  NAND2_X1 U3821 ( .A1(n3815), .A2(n3834), .ZN(n3833) );
  NAND2_X1 U3822 ( .A1(n3814), .A2(n3816), .ZN(n3834) );
  NOR2_X1 U3823 ( .A1(n2427), .A2(n2423), .ZN(n3815) );
  NOR2_X1 U3824 ( .A1(n3814), .A2(n3816), .ZN(n3831) );
  NOR2_X1 U3825 ( .A1(n3835), .A2(n3836), .ZN(n3816) );
  INV_X1 U3826 ( .A(n3837), .ZN(n3836) );
  NAND2_X1 U3827 ( .A1(n3812), .A2(n3838), .ZN(n3837) );
  NAND2_X1 U3828 ( .A1(n3839), .A2(n3809), .ZN(n3838) );
  NOR2_X1 U3829 ( .A1(n2426), .A2(n2423), .ZN(n3812) );
  NOR2_X1 U3830 ( .A1(n3809), .A2(n3839), .ZN(n3835) );
  INV_X1 U3831 ( .A(n3811), .ZN(n3839) );
  NAND2_X1 U3832 ( .A1(n3840), .A2(n3841), .ZN(n3811) );
  NAND2_X1 U3833 ( .A1(n3808), .A2(n3842), .ZN(n3841) );
  INV_X1 U3834 ( .A(n3843), .ZN(n3842) );
  NOR2_X1 U3835 ( .A1(n3805), .A2(n3807), .ZN(n3843) );
  NOR2_X1 U3836 ( .A1(n2344), .A2(n2423), .ZN(n3808) );
  NAND2_X1 U3837 ( .A1(n3805), .A2(n3807), .ZN(n3840) );
  NOR2_X1 U3838 ( .A1(n3844), .A2(n3845), .ZN(n3807) );
  NOR2_X1 U3839 ( .A1(n3803), .A2(n3846), .ZN(n3845) );
  NOR2_X1 U3840 ( .A1(n2324), .A2(n3804), .ZN(n3846) );
  XNOR2_X1 U3841 ( .A(n3847), .B(n3848), .ZN(n3803) );
  NAND2_X1 U3842 ( .A1(n3849), .A2(n3850), .ZN(n3847) );
  INV_X1 U3843 ( .A(n3851), .ZN(n3844) );
  NAND2_X1 U3844 ( .A1(n3804), .A2(n2324), .ZN(n3851) );
  NAND2_X1 U3845 ( .A1(a_4_), .A2(b_4_), .ZN(n2324) );
  NOR2_X1 U3846 ( .A1(n3852), .A2(n3853), .ZN(n3804) );
  INV_X1 U3847 ( .A(n3854), .ZN(n3853) );
  NAND2_X1 U3848 ( .A1(n3801), .A2(n3855), .ZN(n3854) );
  NAND2_X1 U3849 ( .A1(n3800), .A2(n3799), .ZN(n3855) );
  NOR2_X1 U3850 ( .A1(n2423), .A2(n2309), .ZN(n3801) );
  NOR2_X1 U3851 ( .A1(n3799), .A2(n3800), .ZN(n3852) );
  NOR2_X1 U3852 ( .A1(n3856), .A2(n3857), .ZN(n3800) );
  INV_X1 U3853 ( .A(n3858), .ZN(n3857) );
  NAND2_X1 U3854 ( .A1(n3730), .A2(n3859), .ZN(n3858) );
  NAND2_X1 U3855 ( .A1(n3728), .A2(n3729), .ZN(n3859) );
  NOR2_X1 U3856 ( .A1(n2423), .A2(n2422), .ZN(n3730) );
  NOR2_X1 U3857 ( .A1(n3728), .A2(n3729), .ZN(n3856) );
  NOR2_X1 U3858 ( .A1(n3860), .A2(n3861), .ZN(n3729) );
  INV_X1 U3859 ( .A(n3862), .ZN(n3861) );
  NAND2_X1 U3860 ( .A1(n3797), .A2(n3863), .ZN(n3862) );
  NAND2_X1 U3861 ( .A1(n3796), .A2(n3795), .ZN(n3863) );
  NOR2_X1 U3862 ( .A1(n2280), .A2(n2423), .ZN(n3797) );
  NOR2_X1 U3863 ( .A1(n3795), .A2(n3796), .ZN(n3860) );
  NOR2_X1 U3864 ( .A1(n3864), .A2(n3865), .ZN(n3796) );
  INV_X1 U3865 ( .A(n3866), .ZN(n3865) );
  NAND2_X1 U3866 ( .A1(n3793), .A2(n3867), .ZN(n3866) );
  NAND2_X1 U3867 ( .A1(n3791), .A2(n3792), .ZN(n3867) );
  NOR2_X1 U3868 ( .A1(n2423), .A2(n2663), .ZN(n3793) );
  NOR2_X1 U3869 ( .A1(n3791), .A2(n3792), .ZN(n3864) );
  NOR2_X1 U3870 ( .A1(n3868), .A2(n3869), .ZN(n3792) );
  INV_X1 U3871 ( .A(n3870), .ZN(n3869) );
  NAND2_X1 U3872 ( .A1(n3789), .A2(n3871), .ZN(n3870) );
  NAND2_X1 U3873 ( .A1(n3786), .A2(n3788), .ZN(n3871) );
  NOR2_X1 U3874 ( .A1(n2251), .A2(n2423), .ZN(n3789) );
  NOR2_X1 U3875 ( .A1(n3788), .A2(n3786), .ZN(n3868) );
  XOR2_X1 U3876 ( .A(n3872), .B(n3873), .Z(n3786) );
  NAND2_X1 U3877 ( .A1(n3874), .A2(n3875), .ZN(n3872) );
  NAND2_X1 U3878 ( .A1(n3876), .A2(n3877), .ZN(n3788) );
  NAND2_X1 U3879 ( .A1(n3747), .A2(n3878), .ZN(n3877) );
  INV_X1 U3880 ( .A(n3879), .ZN(n3878) );
  NOR2_X1 U3881 ( .A1(n3750), .A2(n3749), .ZN(n3879) );
  XOR2_X1 U3882 ( .A(n3880), .B(n3881), .Z(n3747) );
  XOR2_X1 U3883 ( .A(n3882), .B(n3883), .Z(n3880) );
  NAND2_X1 U3884 ( .A1(b_3_), .A2(a_11_), .ZN(n3882) );
  NAND2_X1 U3885 ( .A1(n3749), .A2(n3750), .ZN(n3876) );
  NAND2_X1 U3886 ( .A1(b_4_), .A2(a_10_), .ZN(n3750) );
  NOR2_X1 U3887 ( .A1(n3884), .A2(n3885), .ZN(n3749) );
  INV_X1 U3888 ( .A(n3886), .ZN(n3885) );
  NAND3_X1 U3889 ( .A1(a_11_), .A2(n3887), .A3(b_4_), .ZN(n3886) );
  NAND2_X1 U3890 ( .A1(n3756), .A2(n3758), .ZN(n3887) );
  NOR2_X1 U3891 ( .A1(n3756), .A2(n3758), .ZN(n3884) );
  NOR2_X1 U3892 ( .A1(n3888), .A2(n3889), .ZN(n3758) );
  INV_X1 U3893 ( .A(n3890), .ZN(n3889) );
  NAND2_X1 U3894 ( .A1(n3784), .A2(n3891), .ZN(n3890) );
  NAND2_X1 U3895 ( .A1(n3785), .A2(n3783), .ZN(n3891) );
  NOR2_X1 U3896 ( .A1(n2423), .A2(n2211), .ZN(n3784) );
  NOR2_X1 U3897 ( .A1(n3783), .A2(n3785), .ZN(n3888) );
  NOR2_X1 U3898 ( .A1(n3892), .A2(n3893), .ZN(n3785) );
  INV_X1 U3899 ( .A(n3894), .ZN(n3893) );
  NAND2_X1 U3900 ( .A1(n3779), .A2(n3895), .ZN(n3894) );
  NAND2_X1 U3901 ( .A1(n3896), .A2(n3781), .ZN(n3895) );
  NOR2_X1 U3902 ( .A1(n2423), .A2(n2191), .ZN(n3779) );
  INV_X1 U3903 ( .A(b_4_), .ZN(n2423) );
  NOR2_X1 U3904 ( .A1(n3781), .A2(n3896), .ZN(n3892) );
  INV_X1 U3905 ( .A(n3780), .ZN(n3896) );
  NAND2_X1 U3906 ( .A1(n3897), .A2(n3898), .ZN(n3780) );
  NAND2_X1 U3907 ( .A1(b_2_), .A2(n3899), .ZN(n3898) );
  NAND2_X1 U3908 ( .A1(n2170), .A2(n3900), .ZN(n3899) );
  NAND2_X1 U3909 ( .A1(a_15_), .A2(n2346), .ZN(n3900) );
  NAND2_X1 U3910 ( .A1(b_3_), .A2(n3901), .ZN(n3897) );
  NAND2_X1 U3911 ( .A1(n2173), .A2(n3902), .ZN(n3901) );
  NAND2_X1 U3912 ( .A1(a_14_), .A2(n2425), .ZN(n3902) );
  NAND3_X1 U3913 ( .A1(b_4_), .A2(n2416), .A3(b_3_), .ZN(n3781) );
  XNOR2_X1 U3914 ( .A(n3903), .B(n3904), .ZN(n3783) );
  XNOR2_X1 U3915 ( .A(n3905), .B(n3906), .ZN(n3903) );
  XOR2_X1 U3916 ( .A(n3907), .B(n3908), .Z(n3756) );
  XNOR2_X1 U3917 ( .A(n3909), .B(n3910), .ZN(n3907) );
  XOR2_X1 U3918 ( .A(n3911), .B(n3912), .Z(n3791) );
  NAND2_X1 U3919 ( .A1(n3913), .A2(n3914), .ZN(n3911) );
  XNOR2_X1 U3920 ( .A(n3915), .B(n3916), .ZN(n3795) );
  XOR2_X1 U3921 ( .A(n3917), .B(n3918), .Z(n3915) );
  NOR2_X1 U3922 ( .A1(n2663), .A2(n2346), .ZN(n3918) );
  XOR2_X1 U3923 ( .A(n3919), .B(n3920), .Z(n3728) );
  NAND2_X1 U3924 ( .A1(n3921), .A2(n3922), .ZN(n3919) );
  XNOR2_X1 U3925 ( .A(n3923), .B(n3924), .ZN(n3799) );
  XOR2_X1 U3926 ( .A(n3925), .B(n3926), .Z(n3923) );
  NOR2_X1 U3927 ( .A1(n2422), .A2(n2346), .ZN(n3926) );
  XOR2_X1 U3928 ( .A(n3927), .B(n3928), .Z(n3805) );
  XOR2_X1 U3929 ( .A(n3929), .B(n3930), .Z(n3927) );
  NOR2_X1 U3930 ( .A1(n2346), .A2(n2424), .ZN(n3930) );
  XOR2_X1 U3931 ( .A(n3931), .B(n3932), .Z(n3809) );
  XOR2_X1 U3932 ( .A(n2390), .B(n3933), .Z(n3931) );
  XNOR2_X1 U3933 ( .A(n3934), .B(n3935), .ZN(n3814) );
  XNOR2_X1 U3934 ( .A(n3936), .B(n3937), .ZN(n3934) );
  NAND2_X1 U3935 ( .A1(a_2_), .A2(b_3_), .ZN(n3936) );
  INV_X1 U3936 ( .A(n3581), .ZN(n3817) );
  XOR2_X1 U3937 ( .A(n3938), .B(n3939), .Z(n3581) );
  XNOR2_X1 U3938 ( .A(n3940), .B(n3941), .ZN(n3938) );
  NOR2_X1 U3939 ( .A1(n2346), .A2(n2427), .ZN(n3941) );
  XNOR2_X1 U3940 ( .A(n3942), .B(n3943), .ZN(n2158) );
  XNOR2_X1 U3941 ( .A(n3944), .B(n3945), .ZN(n3943) );
  NAND2_X1 U3942 ( .A1(a_0_), .A2(b_3_), .ZN(n3945) );
  NAND2_X1 U3943 ( .A1(n3946), .A2(n3826), .ZN(n2465) );
  NAND2_X1 U3944 ( .A1(n3947), .A2(n3948), .ZN(n3826) );
  NAND3_X1 U3945 ( .A1(b_3_), .A2(n3949), .A3(a_0_), .ZN(n3948) );
  NAND2_X1 U3946 ( .A1(n3944), .A2(n3942), .ZN(n3949) );
  INV_X1 U3947 ( .A(n3950), .ZN(n3947) );
  NOR2_X1 U3948 ( .A1(n3942), .A2(n3944), .ZN(n3950) );
  NOR2_X1 U3949 ( .A1(n3951), .A2(n3952), .ZN(n3944) );
  INV_X1 U3950 ( .A(n3953), .ZN(n3952) );
  NAND3_X1 U3951 ( .A1(b_3_), .A2(n3954), .A3(a_1_), .ZN(n3953) );
  NAND2_X1 U3952 ( .A1(n3939), .A2(n3940), .ZN(n3954) );
  NOR2_X1 U3953 ( .A1(n3939), .A2(n3940), .ZN(n3951) );
  NOR2_X1 U3954 ( .A1(n3955), .A2(n3956), .ZN(n3940) );
  INV_X1 U3955 ( .A(n3957), .ZN(n3956) );
  NAND3_X1 U3956 ( .A1(b_3_), .A2(n3958), .A3(a_2_), .ZN(n3957) );
  NAND2_X1 U3957 ( .A1(n3935), .A2(n3937), .ZN(n3958) );
  NOR2_X1 U3958 ( .A1(n3937), .A2(n3935), .ZN(n3955) );
  XOR2_X1 U3959 ( .A(n3959), .B(n3960), .Z(n3935) );
  XNOR2_X1 U3960 ( .A(n3961), .B(n3962), .ZN(n3959) );
  NAND2_X1 U3961 ( .A1(n3963), .A2(n3964), .ZN(n3937) );
  NAND2_X1 U3962 ( .A1(n3932), .A2(n3965), .ZN(n3964) );
  NAND2_X1 U3963 ( .A1(n2341), .A2(n3966), .ZN(n3965) );
  INV_X1 U3964 ( .A(n2390), .ZN(n2341) );
  XOR2_X1 U3965 ( .A(n3967), .B(n3968), .Z(n3932) );
  XNOR2_X1 U3966 ( .A(n3969), .B(n3970), .ZN(n3967) );
  NAND2_X1 U3967 ( .A1(n3933), .A2(n2390), .ZN(n3963) );
  NAND2_X1 U3968 ( .A1(a_3_), .A2(b_3_), .ZN(n2390) );
  INV_X1 U3969 ( .A(n3966), .ZN(n3933) );
  NAND2_X1 U3970 ( .A1(n3971), .A2(n3972), .ZN(n3966) );
  INV_X1 U3971 ( .A(n3973), .ZN(n3972) );
  NOR3_X1 U3972 ( .A1(n2346), .A2(n3974), .A3(n2424), .ZN(n3973) );
  NOR2_X1 U3973 ( .A1(n3928), .A2(n3929), .ZN(n3974) );
  NAND2_X1 U3974 ( .A1(n3928), .A2(n3929), .ZN(n3971) );
  NAND2_X1 U3975 ( .A1(n3849), .A2(n3975), .ZN(n3929) );
  NAND2_X1 U3976 ( .A1(n3848), .A2(n3850), .ZN(n3975) );
  NAND2_X1 U3977 ( .A1(n3976), .A2(n3977), .ZN(n3850) );
  NAND2_X1 U3978 ( .A1(b_3_), .A2(a_5_), .ZN(n3977) );
  INV_X1 U3979 ( .A(n3978), .ZN(n3976) );
  XNOR2_X1 U3980 ( .A(n3979), .B(n3980), .ZN(n3848) );
  XNOR2_X1 U3981 ( .A(n3981), .B(n3982), .ZN(n3979) );
  NAND2_X1 U3982 ( .A1(a_5_), .A2(n3978), .ZN(n3849) );
  NAND2_X1 U3983 ( .A1(n3983), .A2(n3984), .ZN(n3978) );
  NAND3_X1 U3984 ( .A1(a_6_), .A2(n3985), .A3(b_3_), .ZN(n3984) );
  INV_X1 U3985 ( .A(n3986), .ZN(n3985) );
  NOR2_X1 U3986 ( .A1(n3924), .A2(n3925), .ZN(n3986) );
  NAND2_X1 U3987 ( .A1(n3924), .A2(n3925), .ZN(n3983) );
  NAND2_X1 U3988 ( .A1(n3921), .A2(n3987), .ZN(n3925) );
  NAND2_X1 U3989 ( .A1(n3920), .A2(n3922), .ZN(n3987) );
  NAND2_X1 U3990 ( .A1(n3988), .A2(n3989), .ZN(n3922) );
  NAND2_X1 U3991 ( .A1(a_7_), .A2(b_3_), .ZN(n3989) );
  INV_X1 U3992 ( .A(n3990), .ZN(n3988) );
  XNOR2_X1 U3993 ( .A(n3991), .B(n3992), .ZN(n3920) );
  XNOR2_X1 U3994 ( .A(n3993), .B(n3994), .ZN(n3991) );
  NAND2_X1 U3995 ( .A1(a_7_), .A2(n3990), .ZN(n3921) );
  NAND2_X1 U3996 ( .A1(n3995), .A2(n3996), .ZN(n3990) );
  NAND3_X1 U3997 ( .A1(a_8_), .A2(n3997), .A3(b_3_), .ZN(n3996) );
  INV_X1 U3998 ( .A(n3998), .ZN(n3997) );
  NOR2_X1 U3999 ( .A1(n3916), .A2(n3917), .ZN(n3998) );
  NAND2_X1 U4000 ( .A1(n3916), .A2(n3917), .ZN(n3995) );
  NAND2_X1 U4001 ( .A1(n3913), .A2(n3999), .ZN(n3917) );
  NAND2_X1 U4002 ( .A1(n3912), .A2(n3914), .ZN(n3999) );
  NAND2_X1 U4003 ( .A1(n4000), .A2(n4001), .ZN(n3914) );
  NAND2_X1 U4004 ( .A1(b_3_), .A2(a_9_), .ZN(n4001) );
  INV_X1 U4005 ( .A(n4002), .ZN(n4000) );
  XNOR2_X1 U4006 ( .A(n4003), .B(n4004), .ZN(n3912) );
  XNOR2_X1 U4007 ( .A(n4005), .B(n4006), .ZN(n4003) );
  NAND2_X1 U4008 ( .A1(a_9_), .A2(n4002), .ZN(n3913) );
  NAND2_X1 U4009 ( .A1(n3874), .A2(n4007), .ZN(n4002) );
  NAND2_X1 U4010 ( .A1(n3873), .A2(n3875), .ZN(n4007) );
  NAND2_X1 U4011 ( .A1(n4008), .A2(n4009), .ZN(n3875) );
  NAND2_X1 U4012 ( .A1(b_3_), .A2(a_10_), .ZN(n4009) );
  INV_X1 U4013 ( .A(n4010), .ZN(n4008) );
  XNOR2_X1 U4014 ( .A(n4011), .B(n4012), .ZN(n3873) );
  XNOR2_X1 U4015 ( .A(n4013), .B(n4014), .ZN(n4012) );
  NAND2_X1 U4016 ( .A1(a_10_), .A2(n4010), .ZN(n3874) );
  NAND2_X1 U4017 ( .A1(n4015), .A2(n4016), .ZN(n4010) );
  NAND3_X1 U4018 ( .A1(a_11_), .A2(n4017), .A3(b_3_), .ZN(n4016) );
  NAND2_X1 U4019 ( .A1(n3883), .A2(n3881), .ZN(n4017) );
  INV_X1 U4020 ( .A(n4018), .ZN(n4015) );
  NOR2_X1 U4021 ( .A1(n3881), .A2(n3883), .ZN(n4018) );
  NOR2_X1 U4022 ( .A1(n4019), .A2(n4020), .ZN(n3883) );
  INV_X1 U4023 ( .A(n4021), .ZN(n4020) );
  NAND2_X1 U4024 ( .A1(n3909), .A2(n4022), .ZN(n4021) );
  NAND2_X1 U4025 ( .A1(n3910), .A2(n3908), .ZN(n4022) );
  NOR2_X1 U4026 ( .A1(n2346), .A2(n2211), .ZN(n3909) );
  NOR2_X1 U4027 ( .A1(n3908), .A2(n3910), .ZN(n4019) );
  NOR2_X1 U4028 ( .A1(n4023), .A2(n4024), .ZN(n3910) );
  INV_X1 U4029 ( .A(n4025), .ZN(n4024) );
  NAND2_X1 U4030 ( .A1(n3904), .A2(n4026), .ZN(n4025) );
  NAND2_X1 U4031 ( .A1(n4027), .A2(n3906), .ZN(n4026) );
  NOR2_X1 U4032 ( .A1(n2346), .A2(n2191), .ZN(n3904) );
  INV_X1 U4033 ( .A(b_3_), .ZN(n2346) );
  NOR2_X1 U4034 ( .A1(n3906), .A2(n4027), .ZN(n4023) );
  INV_X1 U4035 ( .A(n3905), .ZN(n4027) );
  NAND2_X1 U4036 ( .A1(n4028), .A2(n4029), .ZN(n3905) );
  NAND2_X1 U4037 ( .A1(b_1_), .A2(n4030), .ZN(n4029) );
  NAND2_X1 U4038 ( .A1(n2170), .A2(n4031), .ZN(n4030) );
  NAND2_X1 U4039 ( .A1(a_15_), .A2(n2425), .ZN(n4031) );
  NAND2_X1 U4040 ( .A1(b_2_), .A2(n4032), .ZN(n4028) );
  NAND2_X1 U4041 ( .A1(n2173), .A2(n4033), .ZN(n4032) );
  NAND2_X1 U4042 ( .A1(a_14_), .A2(n2375), .ZN(n4033) );
  NAND3_X1 U4043 ( .A1(b_3_), .A2(n2416), .A3(b_2_), .ZN(n3906) );
  XNOR2_X1 U4044 ( .A(n4034), .B(n4035), .ZN(n3908) );
  XNOR2_X1 U4045 ( .A(n4036), .B(n4037), .ZN(n4034) );
  XNOR2_X1 U4046 ( .A(n4038), .B(n4039), .ZN(n3881) );
  XOR2_X1 U4047 ( .A(n4040), .B(n4041), .Z(n4038) );
  XNOR2_X1 U4048 ( .A(n4042), .B(n4043), .ZN(n3916) );
  XNOR2_X1 U4049 ( .A(n4044), .B(n4045), .ZN(n4042) );
  XNOR2_X1 U4050 ( .A(n4046), .B(n4047), .ZN(n3924) );
  XNOR2_X1 U4051 ( .A(n4048), .B(n4049), .ZN(n4046) );
  XNOR2_X1 U4052 ( .A(n4050), .B(n4051), .ZN(n3928) );
  XNOR2_X1 U4053 ( .A(n4052), .B(n4053), .ZN(n4050) );
  XOR2_X1 U4054 ( .A(n4054), .B(n4055), .Z(n3939) );
  XOR2_X1 U4055 ( .A(n2358), .B(n4056), .Z(n4054) );
  XNOR2_X1 U4056 ( .A(n4057), .B(n4058), .ZN(n3942) );
  XNOR2_X1 U4057 ( .A(n4059), .B(n4060), .ZN(n4057) );
  NAND2_X1 U4058 ( .A1(a_1_), .A2(b_2_), .ZN(n4059) );
  XNOR2_X1 U4059 ( .A(n3824), .B(n3825), .ZN(n3946) );
  NAND2_X1 U4060 ( .A1(n4061), .A2(n4062), .ZN(n3824) );
  XOR2_X1 U4061 ( .A(n4063), .B(n4064), .Z(n2181) );
  INV_X1 U4062 ( .A(n4065), .ZN(n2334) );
  NAND2_X1 U4063 ( .A1(n4066), .A2(n4067), .ZN(n4065) );
  NAND2_X1 U4064 ( .A1(n4064), .A2(n4063), .ZN(n4067) );
  XOR2_X1 U4065 ( .A(n2387), .B(n4068), .Z(n4066) );
  INV_X1 U4066 ( .A(n4069), .ZN(n2333) );
  NAND4_X1 U4067 ( .A1(n2387), .A2(n4068), .A3(n4064), .A4(n4063), .ZN(n4069)
         );
  NAND2_X1 U4068 ( .A1(n4061), .A2(n4070), .ZN(n4063) );
  NAND2_X1 U4069 ( .A1(n3825), .A2(n4062), .ZN(n4070) );
  NAND2_X1 U4070 ( .A1(n4071), .A2(n4072), .ZN(n4062) );
  NAND2_X1 U4071 ( .A1(a_0_), .A2(b_2_), .ZN(n4072) );
  INV_X1 U4072 ( .A(n4073), .ZN(n4071) );
  XOR2_X1 U4073 ( .A(n4074), .B(n4075), .Z(n3825) );
  NOR2_X1 U4074 ( .A1(n4076), .A2(n2426), .ZN(n4075) );
  XOR2_X1 U4075 ( .A(n2371), .B(n4077), .Z(n4074) );
  NAND2_X1 U4076 ( .A1(a_0_), .A2(n4073), .ZN(n4061) );
  NAND2_X1 U4077 ( .A1(n4078), .A2(n4079), .ZN(n4073) );
  NAND3_X1 U4078 ( .A1(b_2_), .A2(n4080), .A3(a_1_), .ZN(n4079) );
  NAND2_X1 U4079 ( .A1(n4058), .A2(n4060), .ZN(n4080) );
  INV_X1 U4080 ( .A(n4081), .ZN(n4078) );
  NOR2_X1 U4081 ( .A1(n4058), .A2(n4060), .ZN(n4081) );
  NAND2_X1 U4082 ( .A1(n4082), .A2(n4083), .ZN(n4060) );
  NAND2_X1 U4083 ( .A1(n4055), .A2(n4084), .ZN(n4083) );
  INV_X1 U4084 ( .A(n4085), .ZN(n4084) );
  NOR2_X1 U4085 ( .A1(n2358), .A2(n4056), .ZN(n4085) );
  XNOR2_X1 U4086 ( .A(n4086), .B(n4087), .ZN(n4055) );
  NOR2_X1 U4087 ( .A1(n2375), .A2(n2344), .ZN(n4087) );
  XOR2_X1 U4088 ( .A(n4088), .B(n4089), .Z(n4086) );
  NAND2_X1 U4089 ( .A1(n4056), .A2(n2358), .ZN(n4082) );
  NAND2_X1 U4090 ( .A1(a_2_), .A2(b_2_), .ZN(n2358) );
  NOR2_X1 U4091 ( .A1(n4090), .A2(n4091), .ZN(n4056) );
  INV_X1 U4092 ( .A(n4092), .ZN(n4091) );
  NAND2_X1 U4093 ( .A1(n3962), .A2(n4093), .ZN(n4092) );
  NAND2_X1 U4094 ( .A1(n3961), .A2(n3960), .ZN(n4093) );
  NOR2_X1 U4095 ( .A1(n2344), .A2(n2425), .ZN(n3962) );
  INV_X1 U4096 ( .A(a_3_), .ZN(n2344) );
  NOR2_X1 U4097 ( .A1(n3960), .A2(n3961), .ZN(n4090) );
  NOR2_X1 U4098 ( .A1(n4094), .A2(n4095), .ZN(n3961) );
  INV_X1 U4099 ( .A(n4096), .ZN(n4095) );
  NAND2_X1 U4100 ( .A1(n3969), .A2(n4097), .ZN(n4096) );
  NAND2_X1 U4101 ( .A1(n3970), .A2(n3968), .ZN(n4097) );
  NOR2_X1 U4102 ( .A1(n2424), .A2(n2425), .ZN(n3969) );
  NOR2_X1 U4103 ( .A1(n3968), .A2(n3970), .ZN(n4094) );
  NOR2_X1 U4104 ( .A1(n4098), .A2(n4099), .ZN(n3970) );
  INV_X1 U4105 ( .A(n4100), .ZN(n4099) );
  NAND2_X1 U4106 ( .A1(n4053), .A2(n4101), .ZN(n4100) );
  NAND2_X1 U4107 ( .A1(n4052), .A2(n4051), .ZN(n4101) );
  NOR2_X1 U4108 ( .A1(n2425), .A2(n2309), .ZN(n4053) );
  NOR2_X1 U4109 ( .A1(n4051), .A2(n4052), .ZN(n4098) );
  NOR2_X1 U4110 ( .A1(n4102), .A2(n4103), .ZN(n4052) );
  INV_X1 U4111 ( .A(n4104), .ZN(n4103) );
  NAND2_X1 U4112 ( .A1(n3981), .A2(n4105), .ZN(n4104) );
  NAND2_X1 U4113 ( .A1(n3982), .A2(n3980), .ZN(n4105) );
  NOR2_X1 U4114 ( .A1(n2425), .A2(n2422), .ZN(n3981) );
  NOR2_X1 U4115 ( .A1(n3980), .A2(n3982), .ZN(n4102) );
  NOR2_X1 U4116 ( .A1(n4106), .A2(n4107), .ZN(n3982) );
  INV_X1 U4117 ( .A(n4108), .ZN(n4107) );
  NAND2_X1 U4118 ( .A1(n4049), .A2(n4109), .ZN(n4108) );
  NAND2_X1 U4119 ( .A1(n4048), .A2(n4047), .ZN(n4109) );
  NOR2_X1 U4120 ( .A1(n2280), .A2(n2425), .ZN(n4049) );
  NOR2_X1 U4121 ( .A1(n4047), .A2(n4048), .ZN(n4106) );
  NOR2_X1 U4122 ( .A1(n4110), .A2(n4111), .ZN(n4048) );
  INV_X1 U4123 ( .A(n4112), .ZN(n4111) );
  NAND2_X1 U4124 ( .A1(n3993), .A2(n4113), .ZN(n4112) );
  NAND2_X1 U4125 ( .A1(n3994), .A2(n3992), .ZN(n4113) );
  NOR2_X1 U4126 ( .A1(n2425), .A2(n2663), .ZN(n3993) );
  NOR2_X1 U4127 ( .A1(n3992), .A2(n3994), .ZN(n4110) );
  NOR2_X1 U4128 ( .A1(n4114), .A2(n4115), .ZN(n3994) );
  INV_X1 U4129 ( .A(n4116), .ZN(n4115) );
  NAND2_X1 U4130 ( .A1(n4045), .A2(n4117), .ZN(n4116) );
  NAND2_X1 U4131 ( .A1(n4044), .A2(n4043), .ZN(n4117) );
  NOR2_X1 U4132 ( .A1(n2425), .A2(n2251), .ZN(n4045) );
  NOR2_X1 U4133 ( .A1(n4043), .A2(n4044), .ZN(n4114) );
  NOR2_X1 U4134 ( .A1(n4118), .A2(n4119), .ZN(n4044) );
  INV_X1 U4135 ( .A(n4120), .ZN(n4119) );
  NAND2_X1 U4136 ( .A1(n4005), .A2(n4121), .ZN(n4120) );
  NAND2_X1 U4137 ( .A1(n4006), .A2(n4004), .ZN(n4121) );
  NOR2_X1 U4138 ( .A1(n2425), .A2(n2419), .ZN(n4005) );
  NOR2_X1 U4139 ( .A1(n4004), .A2(n4006), .ZN(n4118) );
  INV_X1 U4140 ( .A(n4122), .ZN(n4006) );
  NAND2_X1 U4141 ( .A1(n4123), .A2(n4124), .ZN(n4122) );
  NAND2_X1 U4142 ( .A1(n4014), .A2(n4125), .ZN(n4124) );
  INV_X1 U4143 ( .A(n4126), .ZN(n4125) );
  NOR2_X1 U4144 ( .A1(n4013), .A2(n4011), .ZN(n4126) );
  NOR2_X1 U4145 ( .A1(n2425), .A2(n2221), .ZN(n4014) );
  NAND2_X1 U4146 ( .A1(n4011), .A2(n4013), .ZN(n4123) );
  NAND2_X1 U4147 ( .A1(n4127), .A2(n4128), .ZN(n4013) );
  NAND2_X1 U4148 ( .A1(n4040), .A2(n4129), .ZN(n4128) );
  INV_X1 U4149 ( .A(n4130), .ZN(n4129) );
  NOR2_X1 U4150 ( .A1(n4039), .A2(n4041), .ZN(n4130) );
  NOR2_X1 U4151 ( .A1(n2425), .A2(n2211), .ZN(n4040) );
  NAND2_X1 U4152 ( .A1(n4039), .A2(n4041), .ZN(n4127) );
  NAND2_X1 U4153 ( .A1(n4131), .A2(n4132), .ZN(n4041) );
  NAND2_X1 U4154 ( .A1(n4035), .A2(n4133), .ZN(n4132) );
  NAND2_X1 U4155 ( .A1(n4134), .A2(n4037), .ZN(n4133) );
  INV_X1 U4156 ( .A(n4036), .ZN(n4134) );
  NOR2_X1 U4157 ( .A1(n2425), .A2(n2191), .ZN(n4035) );
  INV_X1 U4158 ( .A(b_2_), .ZN(n2425) );
  NAND2_X1 U4159 ( .A1(n4135), .A2(n4036), .ZN(n4131) );
  NAND2_X1 U4160 ( .A1(n4136), .A2(n4137), .ZN(n4036) );
  NAND2_X1 U4161 ( .A1(b_0_), .A2(n4138), .ZN(n4137) );
  NAND2_X1 U4162 ( .A1(n2170), .A2(n4139), .ZN(n4138) );
  NAND2_X1 U4163 ( .A1(a_15_), .A2(n2375), .ZN(n4139) );
  NAND2_X1 U4164 ( .A1(a_15_), .A2(n2415), .ZN(n2170) );
  NAND2_X1 U4165 ( .A1(b_1_), .A2(n4140), .ZN(n4136) );
  NAND2_X1 U4166 ( .A1(n2173), .A2(n4141), .ZN(n4140) );
  NAND2_X1 U4167 ( .A1(a_14_), .A2(n4076), .ZN(n4141) );
  NAND2_X1 U4168 ( .A1(a_14_), .A2(n4142), .ZN(n2173) );
  INV_X1 U4169 ( .A(n4037), .ZN(n4135) );
  NAND3_X1 U4170 ( .A1(b_2_), .A2(n2416), .A3(b_1_), .ZN(n4037) );
  XNOR2_X1 U4171 ( .A(n4143), .B(n4144), .ZN(n4039) );
  XNOR2_X1 U4172 ( .A(n4145), .B(n4146), .ZN(n4144) );
  NAND2_X1 U4173 ( .A1(b_0_), .A2(a_14_), .ZN(n4143) );
  XNOR2_X1 U4174 ( .A(n4147), .B(n4148), .ZN(n4011) );
  NAND2_X1 U4175 ( .A1(n4149), .A2(n4150), .ZN(n4147) );
  NAND2_X1 U4176 ( .A1(n4151), .A2(n4152), .ZN(n4150) );
  NAND2_X1 U4177 ( .A1(b_1_), .A2(a_12_), .ZN(n4151) );
  XNOR2_X1 U4178 ( .A(n4153), .B(n4154), .ZN(n4004) );
  XNOR2_X1 U4179 ( .A(n4155), .B(n4156), .ZN(n4154) );
  NAND2_X1 U4180 ( .A1(b_1_), .A2(a_11_), .ZN(n4153) );
  XNOR2_X1 U4181 ( .A(n4157), .B(n4158), .ZN(n4043) );
  XNOR2_X1 U4182 ( .A(n4159), .B(n4160), .ZN(n4158) );
  NAND2_X1 U4183 ( .A1(b_1_), .A2(a_10_), .ZN(n4157) );
  XNOR2_X1 U4184 ( .A(n4161), .B(n4162), .ZN(n3992) );
  NOR2_X1 U4185 ( .A1(n2251), .A2(n2375), .ZN(n4162) );
  INV_X1 U4186 ( .A(a_9_), .ZN(n2251) );
  XOR2_X1 U4187 ( .A(n4163), .B(n4164), .Z(n4161) );
  XNOR2_X1 U4188 ( .A(n4165), .B(n4166), .ZN(n4047) );
  XNOR2_X1 U4189 ( .A(n4167), .B(n4168), .ZN(n4166) );
  NAND2_X1 U4190 ( .A1(b_1_), .A2(a_8_), .ZN(n4165) );
  XNOR2_X1 U4191 ( .A(n4169), .B(n4170), .ZN(n3980) );
  NOR2_X1 U4192 ( .A1(n2375), .A2(n2280), .ZN(n4170) );
  INV_X1 U4193 ( .A(a_7_), .ZN(n2280) );
  XOR2_X1 U4194 ( .A(n4171), .B(n4172), .Z(n4169) );
  XNOR2_X1 U4195 ( .A(n4173), .B(n4174), .ZN(n4051) );
  XNOR2_X1 U4196 ( .A(n4175), .B(n4176), .ZN(n4174) );
  NAND2_X1 U4197 ( .A1(b_1_), .A2(a_6_), .ZN(n4173) );
  XNOR2_X1 U4198 ( .A(n4177), .B(n4178), .ZN(n3968) );
  NOR2_X1 U4199 ( .A1(n2309), .A2(n2375), .ZN(n4178) );
  INV_X1 U4200 ( .A(a_5_), .ZN(n2309) );
  XOR2_X1 U4201 ( .A(n4179), .B(n4180), .Z(n4177) );
  XNOR2_X1 U4202 ( .A(n4181), .B(n4182), .ZN(n3960) );
  XNOR2_X1 U4203 ( .A(n4183), .B(n4184), .ZN(n4182) );
  NAND2_X1 U4204 ( .A1(a_4_), .A2(b_1_), .ZN(n4181) );
  XNOR2_X1 U4205 ( .A(n4185), .B(n4186), .ZN(n4058) );
  XNOR2_X1 U4206 ( .A(n4187), .B(n4188), .ZN(n4186) );
  NAND2_X1 U4207 ( .A1(a_2_), .A2(b_1_), .ZN(n4185) );
  XOR2_X1 U4208 ( .A(n4189), .B(n4190), .Z(n4064) );
  XNOR2_X1 U4209 ( .A(n4191), .B(n4192), .ZN(n4190) );
  NAND2_X1 U4210 ( .A1(a_1_), .A2(b_0_), .ZN(n4189) );
  NOR2_X1 U4211 ( .A1(n2433), .A2(n4076), .ZN(n2387) );
  NOR2_X1 U4212 ( .A1(n4068), .A2(n2433), .ZN(n2463) );
  INV_X1 U4213 ( .A(a_0_), .ZN(n2433) );
  NOR2_X1 U4214 ( .A1(n4193), .A2(n4194), .ZN(n4068) );
  NOR3_X1 U4215 ( .A1(n4076), .A2(n4195), .A3(n2427), .ZN(n4194) );
  INV_X1 U4216 ( .A(a_1_), .ZN(n2427) );
  INV_X1 U4217 ( .A(n4196), .ZN(n4195) );
  NAND2_X1 U4218 ( .A1(n4192), .A2(n4191), .ZN(n4196) );
  NOR2_X1 U4219 ( .A1(n4191), .A2(n4192), .ZN(n4193) );
  NOR2_X1 U4220 ( .A1(n4197), .A2(n4198), .ZN(n4192) );
  NOR3_X1 U4221 ( .A1(n4076), .A2(n4199), .A3(n2426), .ZN(n4198) );
  INV_X1 U4222 ( .A(a_2_), .ZN(n2426) );
  INV_X1 U4223 ( .A(n4200), .ZN(n4199) );
  NAND2_X1 U4224 ( .A1(n4077), .A2(n2371), .ZN(n4200) );
  NOR2_X1 U4225 ( .A1(n2371), .A2(n4077), .ZN(n4197) );
  NOR2_X1 U4226 ( .A1(n4201), .A2(n4202), .ZN(n4077) );
  INV_X1 U4227 ( .A(n4203), .ZN(n4202) );
  NAND3_X1 U4228 ( .A1(b_1_), .A2(n4204), .A3(a_2_), .ZN(n4203) );
  NAND2_X1 U4229 ( .A1(n4188), .A2(n4187), .ZN(n4204) );
  NOR2_X1 U4230 ( .A1(n4187), .A2(n4188), .ZN(n4201) );
  NOR2_X1 U4231 ( .A1(n4205), .A2(n4206), .ZN(n4188) );
  INV_X1 U4232 ( .A(n4207), .ZN(n4206) );
  NAND3_X1 U4233 ( .A1(b_1_), .A2(n4208), .A3(a_3_), .ZN(n4207) );
  NAND2_X1 U4234 ( .A1(n4089), .A2(n4088), .ZN(n4208) );
  NOR2_X1 U4235 ( .A1(n4088), .A2(n4089), .ZN(n4205) );
  NOR2_X1 U4236 ( .A1(n4209), .A2(n4210), .ZN(n4089) );
  NOR3_X1 U4237 ( .A1(n2375), .A2(n4211), .A3(n2424), .ZN(n4210) );
  INV_X1 U4238 ( .A(a_4_), .ZN(n2424) );
  INV_X1 U4239 ( .A(n4212), .ZN(n4211) );
  NAND2_X1 U4240 ( .A1(n4184), .A2(n4183), .ZN(n4212) );
  NOR2_X1 U4241 ( .A1(n4183), .A2(n4184), .ZN(n4209) );
  NOR2_X1 U4242 ( .A1(n4213), .A2(n4214), .ZN(n4184) );
  INV_X1 U4243 ( .A(n4215), .ZN(n4214) );
  NAND3_X1 U4244 ( .A1(a_5_), .A2(n4216), .A3(b_1_), .ZN(n4215) );
  NAND2_X1 U4245 ( .A1(n4180), .A2(n4179), .ZN(n4216) );
  NOR2_X1 U4246 ( .A1(n4179), .A2(n4180), .ZN(n4213) );
  NOR2_X1 U4247 ( .A1(n4217), .A2(n4218), .ZN(n4180) );
  NOR3_X1 U4248 ( .A1(n2422), .A2(n4219), .A3(n2375), .ZN(n4218) );
  INV_X1 U4249 ( .A(n4220), .ZN(n4219) );
  NAND2_X1 U4250 ( .A1(n4176), .A2(n4175), .ZN(n4220) );
  INV_X1 U4251 ( .A(a_6_), .ZN(n2422) );
  NOR2_X1 U4252 ( .A1(n4175), .A2(n4176), .ZN(n4217) );
  NOR2_X1 U4253 ( .A1(n4221), .A2(n4222), .ZN(n4176) );
  INV_X1 U4254 ( .A(n4223), .ZN(n4222) );
  NAND3_X1 U4255 ( .A1(b_1_), .A2(n4224), .A3(a_7_), .ZN(n4223) );
  NAND2_X1 U4256 ( .A1(n4172), .A2(n4171), .ZN(n4224) );
  NOR2_X1 U4257 ( .A1(n4171), .A2(n4172), .ZN(n4221) );
  NOR2_X1 U4258 ( .A1(n4225), .A2(n4226), .ZN(n4172) );
  NOR3_X1 U4259 ( .A1(n2663), .A2(n4227), .A3(n2375), .ZN(n4226) );
  INV_X1 U4260 ( .A(n4228), .ZN(n4227) );
  NAND2_X1 U4261 ( .A1(n4168), .A2(n4167), .ZN(n4228) );
  INV_X1 U4262 ( .A(a_8_), .ZN(n2663) );
  NOR2_X1 U4263 ( .A1(n4167), .A2(n4168), .ZN(n4225) );
  NOR2_X1 U4264 ( .A1(n4229), .A2(n4230), .ZN(n4168) );
  INV_X1 U4265 ( .A(n4231), .ZN(n4230) );
  NAND3_X1 U4266 ( .A1(a_9_), .A2(n4232), .A3(b_1_), .ZN(n4231) );
  NAND2_X1 U4267 ( .A1(n4164), .A2(n4163), .ZN(n4232) );
  NOR2_X1 U4268 ( .A1(n4163), .A2(n4164), .ZN(n4229) );
  NOR2_X1 U4269 ( .A1(n4233), .A2(n4234), .ZN(n4164) );
  NOR3_X1 U4270 ( .A1(n2419), .A2(n4235), .A3(n2375), .ZN(n4234) );
  NOR2_X1 U4271 ( .A1(n4160), .A2(n4159), .ZN(n4235) );
  INV_X1 U4272 ( .A(a_10_), .ZN(n2419) );
  INV_X1 U4273 ( .A(n4236), .ZN(n4233) );
  NAND2_X1 U4274 ( .A1(n4159), .A2(n4160), .ZN(n4236) );
  NAND2_X1 U4275 ( .A1(n4237), .A2(n4238), .ZN(n4160) );
  NAND3_X1 U4276 ( .A1(a_11_), .A2(n4239), .A3(b_1_), .ZN(n4238) );
  NAND2_X1 U4277 ( .A1(n4156), .A2(n4155), .ZN(n4239) );
  INV_X1 U4278 ( .A(n4240), .ZN(n4155) );
  INV_X1 U4279 ( .A(n4241), .ZN(n4156) );
  NAND2_X1 U4280 ( .A1(n4240), .A2(n4241), .ZN(n4237) );
  NAND2_X1 U4281 ( .A1(n4149), .A2(n4242), .ZN(n4241) );
  NAND2_X1 U4282 ( .A1(n4243), .A2(n4148), .ZN(n4242) );
  NAND2_X1 U4283 ( .A1(n4146), .A2(n4244), .ZN(n4148) );
  NAND3_X1 U4284 ( .A1(b_0_), .A2(a_14_), .A3(n4145), .ZN(n4244) );
  NOR2_X1 U4285 ( .A1(n2375), .A2(n2191), .ZN(n4145) );
  INV_X1 U4286 ( .A(a_13_), .ZN(n2191) );
  INV_X1 U4287 ( .A(b_1_), .ZN(n2375) );
  NAND3_X1 U4288 ( .A1(b_1_), .A2(n2416), .A3(b_0_), .ZN(n4146) );
  INV_X1 U4289 ( .A(a_14_), .ZN(n2415) );
  INV_X1 U4290 ( .A(a_15_), .ZN(n4142) );
  NAND2_X1 U4291 ( .A1(n4152), .A2(n2211), .ZN(n4243) );
  NAND3_X1 U4292 ( .A1(b_1_), .A2(a_12_), .A3(n4245), .ZN(n4149) );
  INV_X1 U4293 ( .A(n4152), .ZN(n4245) );
  NAND2_X1 U4294 ( .A1(b_0_), .A2(a_13_), .ZN(n4152) );
  NOR2_X1 U4295 ( .A1(n4076), .A2(n2211), .ZN(n4240) );
  INV_X1 U4296 ( .A(a_12_), .ZN(n2211) );
  NOR2_X1 U4297 ( .A1(n4076), .A2(n2221), .ZN(n4159) );
  INV_X1 U4298 ( .A(a_11_), .ZN(n2221) );
  INV_X1 U4299 ( .A(b_0_), .ZN(n4076) );
  NAND2_X1 U4300 ( .A1(b_0_), .A2(a_10_), .ZN(n4163) );
  NAND2_X1 U4301 ( .A1(b_0_), .A2(a_9_), .ZN(n4167) );
  NAND2_X1 U4302 ( .A1(b_0_), .A2(a_8_), .ZN(n4171) );
  NAND2_X1 U4303 ( .A1(b_0_), .A2(a_7_), .ZN(n4175) );
  NAND2_X1 U4304 ( .A1(b_0_), .A2(a_6_), .ZN(n4179) );
  NAND2_X1 U4305 ( .A1(b_0_), .A2(a_5_), .ZN(n4183) );
  NAND2_X1 U4306 ( .A1(a_4_), .A2(b_0_), .ZN(n4088) );
  NAND2_X1 U4307 ( .A1(a_3_), .A2(b_0_), .ZN(n4187) );
  NAND2_X1 U4308 ( .A1(a_1_), .A2(b_1_), .ZN(n2371) );
  NAND2_X1 U4309 ( .A1(a_0_), .A2(b_1_), .ZN(n4191) );
endmodule

