module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270,
         WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278,
         DFF_167_n1, WX1280, DFF_168_n1, WX1282, DFF_169_n1, WX1284, WX1286,
         DFF_171_n1, WX1288, DFF_172_n1, WX1290, DFF_173_n1, WX1292,
         DFF_174_n1, WX1294, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1778, n8702, n8701, n8700, n8699, n8696, n8695, n8694,
         n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684,
         n8683, n8682, n8681, n8680, n8677, n8676, n8675, n8674, n8673, n8672,
         n8671, WX1839, n8670, WX1937, n8669, WX1939, n8668, WX1941, n8667,
         WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949, n8663, WX1951,
         n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959, n8657, WX1961,
         n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653, WX1969, WX1970,
         WX1971, WX1972, WX1973, WX1974, WX1975, WX1976, WX1977, WX1978,
         WX1979, WX1980, WX1981, WX1982, WX1983, WX1984, WX1985, WX1986,
         WX1987, WX1988, WX1989, WX1990, WX1991, WX1993, WX1994, WX1995,
         WX1996, WX1997, WX1998, WX1999, WX2000, WX2001, WX2002, WX2003,
         WX2004, WX2005, WX2006, WX2007, WX2008, WX2009, WX2010, WX2011,
         WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018, WX2019,
         WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026, WX2027,
         WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, WX2035, WX2036, n3783,
         WX2037, WX2038, WX2039, WX2040, WX2041, WX2042, WX2043, WX2044, n3775,
         WX2045, WX2046, WX2047, WX2048, WX2049, WX2050, WX2051, WX2052,
         WX2053, WX2054, WX2055, WX2056, n3763, WX2057, WX2058, WX2059, WX2060,
         WX2061, WX2062, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069,
         WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076, WX2077,
         WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084, WX2085,
         WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092, WX2093,
         WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101, WX2102,
         WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109, WX2110,
         WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117, WX2118,
         WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125, WX2126,
         WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133, WX2134,
         WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142, WX2143,
         WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150, WX2151,
         WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158, WX2159,
         WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166, WX2167,
         WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175, WX2176,
         WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183, WX2184,
         WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191, WX2192,
         WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563,
         WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571,
         WX2573, DFF_360_n1, WX2575, DFF_361_n1, WX2577, WX2579, DFF_363_n1,
         WX2581, DFF_364_n1, WX2583, DFF_365_n1, WX2585, DFF_366_n1, WX2587,
         WX2589, DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, DFF_379_n1, WX2613, DFF_380_n1, WX2615,
         DFF_381_n1, WX2617, DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644,
         n8643, n8642, n8641, n8640, n8639, n8638, n8637, n8636, n8635, n8632,
         n8631, n8630, n8629, n8628, n8627, n8626, n8625, n8624, n8623, n8622,
         n8621, n8620, n8619, n8618, n8617, n8616, n8613, WX3132, n8612,
         WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238,
         n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603,
         WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256,
         n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266,
         WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274,
         WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282,
         WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290,
         WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299,
         WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307,
         WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315,
         WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323,
         WX3324, WX3325, WX3326, WX3327, WX3328, WX3329, WX3330, WX3331,
         WX3332, WX3334, WX3335, WX3336, WX3337, WX3338, WX3339, WX3340,
         WX3341, n3739, WX3342, WX3343, WX3344, WX3345, n3735, WX3346, WX3347,
         WX3348, WX3349, WX3350, WX3351, WX3352, WX3353, WX3354, WX3355,
         WX3356, WX3357, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363,
         WX3364, WX3365, WX3366, WX3367, WX3368, WX3370, WX3371, WX3372,
         WX3373, WX3374, WX3375, WX3376, WX3377, WX3378, WX3379, WX3380,
         WX3381, WX3382, WX3383, WX3384, WX3385, WX3386, WX3387, WX3388,
         WX3389, WX3390, WX3391, WX3392, WX3393, WX3394, WX3395, WX3396,
         WX3397, WX3398, WX3399, WX3400, WX3401, WX3402, WX3403, WX3404,
         WX3406, WX3407, WX3408, WX3409, WX3410, WX3411, WX3412, WX3413,
         WX3414, WX3415, WX3416, WX3417, WX3418, WX3419, WX3420, WX3421,
         WX3422, WX3423, WX3424, WX3425, WX3426, WX3427, WX3428, WX3429,
         WX3430, WX3431, WX3432, WX3433, WX3434, WX3435, WX3436, WX3437,
         WX3438, WX3440, WX3441, WX3442, WX3443, WX3444, WX3445, WX3446,
         WX3447, WX3448, WX3449, WX3450, WX3451, WX3452, WX3453, WX3454,
         WX3455, WX3456, WX3457, WX3458, WX3459, WX3460, WX3461, WX3462,
         WX3463, WX3464, WX3465, WX3466, WX3467, WX3468, WX3469, WX3470,
         WX3471, WX3472, WX3474, WX3475, WX3476, WX3477, WX3478, WX3479,
         WX3480, WX3481, WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1,
         WX3852, DFF_545_n1, WX3854, DFF_546_n1, WX3856, WX3858, DFF_548_n1,
         WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864, DFF_551_n1, WX3866,
         DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872, DFF_555_n1, WX3874,
         DFF_556_n1, WX3876, DFF_557_n1, WX3878, DFF_558_n1, WX3880, WX3882,
         DFF_560_n1, WX3884, DFF_561_n1, WX3886, DFF_562_n1, WX3888,
         DFF_563_n1, WX3890, DFF_564_n1, WX3892, DFF_565_n1, WX3894,
         DFF_566_n1, WX3896, DFF_567_n1, WX3898, DFF_568_n1, WX3900,
         DFF_569_n1, WX3902, DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908,
         DFF_573_n1, WX3910, DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586,
         n8585, n8584, n8583, n8582, n8581, n8580, n8579, n8578, n8577, n8576,
         n8573, n8572, n8571, n8570, n8569, n8568, n8567, n8566, n8565, n8564,
         n8563, n8562, n8561, n8560, n8559, n8558, n8555, WX4425, n8554,
         WX4523, n8553, WX4525, n8552, WX4527, n8551, WX4529, n8550, WX4531,
         n8549, WX4533, n8548, WX4535, n8547, WX4537, n8546, WX4539, n8545,
         WX4541, n8544, WX4543, n8543, WX4545, n8542, WX4547, n8541, WX4549,
         n8540, WX4551, WX4553, n8537, WX4555, WX4556, WX4557, WX4558, WX4559,
         WX4560, WX4561, WX4562, WX4563, WX4564, WX4565, WX4566, WX4567,
         WX4568, WX4569, WX4570, WX4571, WX4572, WX4573, WX4574, WX4575,
         WX4576, WX4577, WX4578, WX4579, WX4580, WX4581, WX4582, WX4583,
         WX4584, WX4585, WX4587, WX4588, WX4589, WX4590, WX4591, WX4592,
         WX4593, WX4594, WX4595, WX4596, WX4597, WX4598, WX4599, WX4600,
         WX4601, WX4602, WX4603, WX4604, WX4605, WX4606, WX4607, WX4608,
         WX4609, WX4610, WX4611, WX4612, WX4613, WX4614, WX4615, WX4616,
         WX4617, WX4618, WX4619, WX4621, WX4622, WX4623, WX4624, n3717, WX4625,
         WX4626, WX4627, WX4628, n3713, WX4629, WX4630, WX4631, WX4632, WX4633,
         WX4634, WX4635, WX4636, WX4637, WX4638, WX4639, WX4640, WX4641,
         WX4642, WX4643, WX4644, WX4645, WX4646, WX4647, WX4648, WX4649,
         WX4650, n3691, WX4651, WX4652, WX4653, WX4655, WX4656, WX4657, WX4658,
         WX4659, WX4660, WX4661, WX4662, WX4663, WX4664, WX4665, WX4666,
         WX4667, WX4668, WX4669, WX4670, WX4671, WX4672, WX4673, WX4674,
         WX4675, WX4676, WX4677, WX4678, WX4679, WX4680, WX4681, WX4682,
         WX4683, WX4684, WX4685, WX4686, WX4687, WX4689, WX4690, WX4691,
         WX4692, WX4693, WX4694, WX4695, WX4696, WX4697, WX4698, WX4699,
         WX4700, WX4701, WX4702, WX4703, WX4704, WX4705, WX4706, WX4707,
         WX4708, WX4709, WX4710, WX4711, WX4712, WX4713, WX4714, WX4715,
         WX4716, WX4717, WX4718, WX4719, WX4720, WX4721, WX4723, WX4724,
         WX4725, WX4726, WX4727, WX4728, WX4729, WX4730, WX4731, WX4732,
         WX4733, WX4734, WX4735, WX4736, WX4737, WX4738, WX4739, WX4740,
         WX4741, WX4742, WX4743, WX4744, WX4745, WX4746, WX4747, WX4748,
         WX4749, WX4750, WX4751, WX4752, WX4753, WX4754, WX4755, WX4757,
         WX4758, WX4759, WX4760, WX4761, WX4762, WX4763, WX4764, WX4765,
         WX4766, WX4767, WX4768, WX4769, WX4770, WX4771, WX4772, WX4773,
         WX4774, WX4775, WX4776, WX4777, WX4778, WX5143, DFF_736_n1, WX5145,
         DFF_737_n1, WX5147, DFF_738_n1, WX5149, WX5151, DFF_740_n1, WX5153,
         WX5155, DFF_742_n1, WX5157, DFF_743_n1, WX5159, DFF_744_n1, WX5161,
         DFF_745_n1, WX5163, WX5165, DFF_747_n1, WX5167, DFF_748_n1, WX5169,
         DFF_749_n1, WX5171, DFF_750_n1, WX5173, WX5175, DFF_752_n1, WX5177,
         DFF_753_n1, WX5179, DFF_754_n1, WX5181, DFF_755_n1, WX5183,
         DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191,
         DFF_760_n1, WX5193, DFF_761_n1, WX5195, DFF_762_n1, WX5197,
         DFF_763_n1, WX5199, DFF_764_n1, WX5201, DFF_765_n1, WX5203,
         DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528, n8527, n8526, n8525,
         n8524, n8523, n8520, n8519, n8518, n8517, n8516, n8515, n8514, n8513,
         n8512, n8511, n8510, n8509, n8508, n8507, n8506, n8505, n8502, n8501,
         n8500, n8499, n8498, n8497, WX5718, n8496, WX5816, n8495, WX5818,
         n8494, WX5820, n8493, WX5822, n8492, WX5824, n8491, WX5826, n8490,
         WX5828, n8489, WX5830, n8488, WX5832, n8487, WX5834, WX5836, n8484,
         WX5838, n8483, WX5840, n8482, WX5842, n8481, WX5844, n8480, WX5846,
         n8479, WX5848, WX5849, WX5850, WX5851, WX5852, WX5853, WX5854, WX5855,
         WX5856, WX5857, WX5858, WX5859, WX5860, WX5861, WX5862, WX5863,
         WX5864, WX5865, WX5866, WX5867, WX5868, WX5870, WX5871, WX5872,
         WX5873, WX5874, WX5875, WX5876, WX5877, WX5878, WX5879, WX5880,
         WX5881, WX5882, WX5883, WX5884, WX5885, WX5886, WX5887, WX5888,
         WX5889, WX5890, WX5891, WX5892, WX5893, WX5894, WX5895, WX5896,
         WX5897, WX5898, WX5899, WX5900, WX5901, WX5902, WX5904, WX5905,
         WX5906, WX5907, WX5908, WX5909, WX5910, WX5911, WX5912, WX5913,
         WX5914, WX5915, WX5916, WX5917, WX5918, WX5919, WX5920, WX5921,
         WX5922, WX5923, WX5924, WX5925, WX5926, WX5927, WX5928, WX5929,
         WX5930, WX5931, WX5932, WX5933, n3669, WX5934, WX5935, WX5936, WX5938,
         WX5939, WX5940, WX5941, n3661, WX5942, WX5943, WX5944, WX5945, WX5946,
         WX5947, WX5948, WX5949, WX5950, WX5951, WX5952, WX5953, WX5954,
         WX5955, WX5956, WX5957, WX5958, WX5959, WX5960, WX5961, WX5962,
         WX5963, WX5964, WX5965, WX5966, WX5967, WX5968, WX5969, WX5970,
         WX5972, WX5973, WX5974, WX5975, WX5976, WX5977, WX5978, WX5979,
         WX5980, WX5981, WX5982, WX5983, WX5984, WX5985, WX5986, WX5987,
         WX5988, WX5989, WX5990, WX5991, WX5992, WX5993, WX5994, WX5995,
         WX5996, WX5997, WX5998, WX5999, WX6000, WX6001, WX6002, WX6003,
         WX6004, WX6006, WX6007, WX6008, WX6009, WX6010, WX6011, WX6012,
         WX6013, WX6014, WX6015, WX6016, WX6017, WX6018, WX6019, WX6020,
         WX6021, WX6022, WX6023, WX6024, WX6025, WX6026, WX6027, WX6028,
         WX6029, WX6030, WX6031, WX6032, WX6033, WX6034, WX6035, WX6036,
         WX6037, WX6038, WX6040, WX6041, WX6042, WX6043, WX6044, WX6045,
         WX6046, WX6047, WX6048, WX6049, WX6050, WX6051, WX6052, WX6053,
         WX6054, WX6055, WX6056, WX6057, WX6058, WX6059, WX6060, WX6061,
         WX6062, WX6063, WX6064, WX6065, WX6066, WX6067, WX6068, WX6069,
         WX6070, WX6071, WX6436, WX6438, DFF_929_n1, WX6440, DFF_930_n1,
         WX6442, WX6444, DFF_932_n1, WX6446, DFF_933_n1, WX6448, DFF_934_n1,
         WX6450, DFF_935_n1, WX6452, DFF_936_n1, WX6454, DFF_937_n1, WX6456,
         WX6458, DFF_939_n1, WX6460, DFF_940_n1, WX6462, DFF_941_n1, WX6464,
         DFF_942_n1, WX6466, WX6468, DFF_944_n1, WX6470, WX6472, DFF_946_n1,
         WX6474, DFF_947_n1, WX6476, DFF_948_n1, WX6478, DFF_949_n1, WX6480,
         DFF_950_n1, WX6482, DFF_951_n1, WX6484, DFF_952_n1, WX6486,
         DFF_953_n1, WX6488, DFF_954_n1, WX6490, DFF_955_n1, WX6492,
         DFF_956_n1, WX6494, DFF_957_n1, WX6496, DFF_958_n1, WX6498,
         DFF_959_n1, WX6950, n8470, n8467, n8466, n8465, n8464, n8463, n8462,
         n8461, n8460, n8459, n8458, n8457, n8456, n8455, n8454, n8453, n8452,
         n8449, n8448, n8447, n8446, n8445, n8444, n8443, n8442, n8441, n8440,
         n8439, WX7011, n8438, WX7109, n8437, WX7111, n8436, WX7113, n8435,
         WX7115, n8434, WX7117, WX7119, n8431, WX7121, n8430, WX7123, n8429,
         WX7125, n8428, WX7127, n8427, WX7129, n8426, WX7131, n8425, WX7133,
         n8424, WX7135, n8423, WX7137, n8422, WX7139, n8421, WX7141, WX7142,
         WX7143, WX7144, WX7145, WX7146, WX7147, WX7148, WX7149, WX7150,
         WX7151, WX7153, WX7154, WX7155, WX7156, WX7157, WX7158, WX7159,
         WX7160, WX7161, WX7162, WX7163, WX7164, WX7165, WX7166, WX7167,
         WX7168, WX7169, WX7170, WX7171, WX7172, WX7173, WX7174, WX7175,
         WX7176, WX7177, WX7178, WX7179, WX7180, WX7181, WX7182, WX7183,
         WX7184, WX7185, WX7187, WX7188, WX7189, WX7190, WX7191, WX7192,
         WX7193, WX7194, WX7195, WX7196, WX7197, WX7198, WX7199, WX7200,
         WX7201, WX7202, WX7203, WX7204, WX7205, WX7206, WX7207, WX7208,
         WX7209, WX7210, WX7211, WX7212, WX7213, WX7214, WX7215, WX7216, n3647,
         WX7217, WX7218, WX7219, WX7221, WX7222, WX7223, WX7224, n3639, WX7225,
         WX7226, WX7227, WX7228, n3635, WX7229, WX7230, WX7231, WX7232, WX7233,
         WX7234, WX7235, WX7236, WX7237, WX7238, WX7239, WX7240, WX7241,
         WX7242, WX7243, WX7244, WX7245, WX7246, WX7247, WX7248, WX7249,
         WX7250, WX7251, WX7252, WX7253, WX7255, WX7256, WX7257, WX7258,
         WX7259, WX7260, WX7261, WX7262, WX7263, WX7264, WX7265, WX7266,
         WX7267, WX7268, WX7269, WX7270, WX7271, WX7272, WX7273, WX7274,
         WX7275, WX7276, WX7277, WX7278, WX7279, WX7280, WX7281, WX7282,
         WX7283, WX7284, WX7285, WX7286, WX7287, WX7289, WX7290, WX7291,
         WX7292, WX7293, WX7294, WX7295, WX7296, WX7297, WX7298, WX7299,
         WX7300, WX7301, WX7302, WX7303, WX7304, WX7305, WX7306, WX7307,
         WX7308, WX7309, WX7310, WX7311, WX7312, WX7313, WX7314, WX7315,
         WX7316, WX7317, WX7318, WX7319, WX7320, WX7321, WX7323, WX7324,
         WX7325, WX7326, WX7327, WX7328, WX7329, WX7330, WX7331, WX7332,
         WX7333, WX7334, WX7335, WX7336, WX7337, WX7338, WX7339, WX7340,
         WX7341, WX7342, WX7343, WX7344, WX7345, WX7346, WX7347, WX7348,
         WX7349, WX7350, WX7351, WX7352, WX7353, WX7354, WX7355, WX7357,
         WX7358, WX7359, WX7360, WX7361, WX7362, WX7363, WX7364, WX7729,
         DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1, WX7735, WX7737,
         DFF_1124_n1, WX7739, DFF_1125_n1, WX7741, DFF_1126_n1, WX7743,
         DFF_1127_n1, WX7745, DFF_1128_n1, WX7747, DFF_1129_n1, WX7749, WX7751,
         DFF_1131_n1, WX7753, WX7755, DFF_1133_n1, WX7757, DFF_1134_n1, WX7759,
         WX7761, DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, DFF_1140_n1, WX7771, DFF_1141_n1, WX7773,
         DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n8410, n8409, n8408, n8407, n8406, n8405, n8404, n8403, n8402,
         n8401, n8400, n8399, n8396, n8395, n8394, n8393, n8392, n8391, n8390,
         n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381, WX8304,
         WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410,
         n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370,
         WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428,
         n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438,
         WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445, WX8446,
         WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453, WX8454,
         WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461, WX8462,
         WX8463, WX8464, WX8465, WX8466, WX8467, WX8468, WX8470, WX8471,
         WX8472, WX8473, WX8474, WX8475, WX8476, WX8477, WX8478, WX8479,
         WX8480, WX8481, WX8482, WX8483, WX8484, WX8485, WX8486, WX8487,
         WX8488, WX8489, WX8490, WX8491, WX8492, WX8493, WX8494, WX8495,
         WX8496, WX8497, WX8498, WX8499, n3625, WX8500, WX8501, WX8502, WX8504,
         WX8505, WX8506, WX8507, n3617, WX8508, WX8509, WX8510, WX8511, n3613,
         WX8512, WX8513, WX8514, WX8515, WX8516, WX8517, WX8518, WX8519,
         WX8520, WX8521, WX8522, WX8523, WX8524, WX8525, WX8526, WX8527,
         WX8528, WX8529, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535,
         WX8536, WX8538, WX8539, WX8540, WX8541, WX8542, WX8543, WX8544,
         WX8545, WX8546, WX8547, WX8548, WX8549, WX8550, WX8551, WX8552,
         WX8553, WX8554, WX8555, WX8556, WX8557, WX8558, WX8559, WX8560,
         WX8561, WX8562, WX8563, WX8564, WX8565, WX8566, WX8567, WX8568,
         WX8569, WX8570, WX8572, WX8573, WX8574, WX8575, WX8576, WX8577,
         WX8578, WX8579, WX8580, WX8581, WX8582, WX8583, WX8584, WX8585,
         WX8586, WX8587, WX8588, WX8589, WX8590, WX8591, WX8592, WX8593,
         WX8594, WX8595, WX8596, WX8597, WX8598, WX8599, WX8600, WX8601,
         WX8602, WX8603, WX8604, WX8606, WX8607, WX8608, WX8609, WX8610,
         WX8611, WX8612, WX8613, WX8614, WX8615, WX8616, WX8617, WX8618,
         WX8619, WX8620, WX8621, WX8622, WX8623, WX8624, WX8625, WX8626,
         WX8627, WX8628, WX8629, WX8630, WX8631, WX8632, WX8633, WX8634,
         WX8635, WX8636, WX8637, WX8638, WX8640, WX8641, WX8642, WX8643,
         WX8644, WX8645, WX8646, WX8647, WX8648, WX8649, WX8650, WX8651,
         WX8652, WX8653, WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1,
         WX9024, DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, WX9030, DFF_1316_n1,
         WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038, DFF_1320_n1,
         WX9040, DFF_1321_n1, WX9042, WX9044, DFF_1323_n1, WX9046, DFF_1324_n1,
         WX9048, DFF_1325_n1, WX9050, DFF_1326_n1, WX9052, WX9054, DFF_1328_n1,
         WX9056, DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350,
         n8349, n8348, n8347, n8346, n8343, n8342, n8341, n8340, n8339, n8338,
         n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328,
         n8325, n8324, n8323, n8322, WX9597, n8321, WX9695, n8320, WX9697,
         n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705, n8315,
         WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311, WX9715,
         n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305, WX9725,
         n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733, WX9734,
         WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741, WX9742,
         WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749, WX9750,
         WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758, WX9759,
         WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766, WX9767,
         WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774, WX9775,
         WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782, WX9783,
         WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791, WX9792,
         WX9793, WX9794, n3591, WX9795, WX9796, WX9797, WX9798, WX9799, WX9800,
         WX9801, WX9802, WX9803, WX9804, WX9805, WX9806, WX9807, WX9808,
         WX9809, WX9810, WX9811, WX9812, WX9813, WX9814, WX9815, WX9816, n3569,
         WX9817, WX9818, WX9819, WX9821, WX9822, WX9823, WX9824, WX9825,
         WX9826, WX9827, WX9828, WX9829, WX9830, WX9831, WX9832, WX9833,
         WX9834, WX9835, WX9836, WX9837, WX9838, WX9839, WX9840, WX9841,
         WX9842, WX9843, WX9844, WX9845, WX9846, WX9847, WX9848, WX9849,
         WX9850, WX9851, WX9852, WX9853, WX9855, WX9856, WX9857, WX9858,
         WX9859, WX9860, WX9861, WX9862, WX9863, WX9864, WX9865, WX9866,
         WX9867, WX9868, WX9869, WX9870, WX9871, WX9872, WX9873, WX9874,
         WX9875, WX9876, WX9877, WX9878, WX9879, WX9880, WX9881, WX9882,
         WX9883, WX9884, WX9885, WX9886, WX9887, WX9889, WX9890, WX9891,
         WX9892, WX9893, WX9894, WX9895, WX9896, WX9897, WX9898, WX9899,
         WX9900, WX9901, WX9902, WX9903, WX9904, WX9905, WX9906, WX9907,
         WX9908, WX9909, WX9910, WX9911, WX9912, WX9913, WX9914, WX9915,
         WX9916, WX9917, WX9918, WX9919, WX9920, WX9921, WX9923, WX9924,
         WX9925, WX9926, WX9927, WX9928, WX9929, WX9930, WX9931, WX9932,
         WX9933, WX9934, WX9935, WX9936, WX9937, WX9938, WX9939, WX9940,
         WX9941, WX9942, WX9943, WX9944, WX9945, WX9946, WX9947, WX9948,
         WX9949, WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319,
         WX10321, WX10323, DFF_1508_n1, WX10325, DFF_1509_n1, WX10327,
         DFF_1510_n1, WX10329, DFF_1511_n1, WX10331, DFF_1512_n1, WX10333,
         DFF_1513_n1, WX10335, WX10337, DFF_1515_n1, WX10339, DFF_1516_n1,
         WX10341, DFF_1517_n1, WX10343, DFF_1518_n1, WX10345, DFF_1519_n1,
         WX10347, DFF_1520_n1, WX10349, DFF_1521_n1, WX10351, DFF_1522_n1,
         WX10353, WX10355, DFF_1524_n1, WX10357, DFF_1525_n1, WX10359,
         DFF_1526_n1, WX10361, DFF_1527_n1, WX10363, DFF_1528_n1, WX10365,
         DFF_1529_n1, WX10367, DFF_1530_n1, WX10369, DFF_1531_n1, WX10371,
         DFF_1532_n1, WX10373, DFF_1533_n1, WX10375, DFF_1534_n1, WX10377,
         DFF_1535_n1, WX10829, n8295, n8294, n8293, n8290, n8289, n8288, n8287,
         n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279, n8278, n8277,
         n8276, n8275, n8272, n8271, n8270, n8269, n8268, n8267, n8266, n8265,
         n8264, WX10890, n8263, WX10988, n8262, WX10990, n8261, WX10992, n8260,
         WX10994, n8259, WX10996, n8258, WX10998, n8257, WX11000, WX11002,
         n8254, WX11004, n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250,
         WX11012, n8249, WX11014, n8248, WX11016, n8247, WX11018, n8246,
         WX11020, WX11021, WX11022, WX11023, WX11024, WX11025, WX11026,
         WX11027, WX11028, WX11029, WX11030, WX11031, WX11032, WX11033,
         WX11034, WX11036, WX11037, WX11038, WX11039, WX11040, WX11041,
         WX11042, WX11043, WX11044, WX11045, WX11046, WX11047, WX11048,
         WX11049, WX11050, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, WX11086, WX11087, WX11088, WX11089, WX11090, WX11091,
         WX11092, WX11093, WX11094, WX11095, WX11096, WX11097, WX11098,
         WX11099, n3547, WX11100, WX11101, WX11102, WX11104, WX11105, WX11106,
         WX11107, n3539, WX11108, WX11109, WX11110, WX11111, n3535, WX11112,
         WX11113, WX11114, WX11115, WX11116, WX11117, WX11118, WX11119,
         WX11120, WX11121, WX11122, WX11123, WX11124, WX11125, WX11126,
         WX11127, WX11128, WX11129, WX11130, WX11131, WX11132, WX11133,
         WX11134, WX11135, WX11136, WX11138, WX11139, WX11140, WX11141,
         WX11142, WX11143, WX11144, WX11145, WX11146, WX11147, WX11148,
         WX11149, WX11150, WX11151, WX11152, WX11153, WX11154, WX11155,
         WX11156, WX11157, WX11158, WX11159, WX11160, WX11161, WX11162,
         WX11163, WX11164, WX11165, WX11166, WX11167, WX11168, WX11169,
         WX11170, WX11172, WX11173, WX11174, WX11175, WX11176, WX11177,
         WX11178, WX11179, WX11180, WX11181, WX11182, WX11183, WX11184,
         WX11185, WX11186, WX11187, WX11188, WX11189, WX11190, WX11191,
         WX11192, WX11193, WX11194, WX11195, WX11196, WX11197, WX11198,
         WX11199, WX11200, WX11201, WX11202, WX11203, WX11204, WX11206,
         WX11207, WX11208, WX11209, WX11210, WX11211, WX11212, WX11213,
         WX11214, WX11215, WX11216, WX11217, WX11218, WX11219, WX11220,
         WX11221, WX11222, WX11223, WX11224, WX11225, WX11226, WX11227,
         WX11228, WX11229, WX11230, WX11231, WX11232, WX11233, WX11234,
         WX11235, WX11236, WX11237, WX11238, WX11240, WX11241, WX11242,
         WX11243, WX11608, DFF_1696_n1, WX11610, DFF_1697_n1, WX11612,
         DFF_1698_n1, WX11614, WX11616, DFF_1700_n1, WX11618, DFF_1701_n1,
         WX11620, DFF_1702_n1, WX11622, DFF_1703_n1, WX11624, DFF_1704_n1,
         WX11626, DFF_1705_n1, WX11628, WX11630, DFF_1707_n1, WX11632,
         DFF_1708_n1, WX11634, DFF_1709_n1, WX11636, WX11638, WX11640,
         DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, DFF_1714_n1, WX11646,
         DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1, WX11652,
         DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1, WX11658,
         DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1, WX11664,
         DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1, WX11670,
         n2245, n2153, n3278, n2152, n2148, Tj_Trigger, Tj_OUT1, Tj_OUT2,
         Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8,
         Tj_OUT5678, test_se_NOT, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n2182, n2183, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7863, n7864, n7866, n7867, n7868, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7887, n7888, n7889, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7938, n7939, n7941, n7942, n7943, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7958, n7959, n7961, n7962, n7963, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7978, n7979, n7981,
         n7982, n7983, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8031, n8032, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8052, n8053, n8054, n8055, n8056,
         n8057, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8094, n8095, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8255, n8256, n8273, n8274, n8291, n8292, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8308, n8309, n8326, n8327, n8344, n8345,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8379, n8380,
         n8397, n8398, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8432, n8450, n8451, n8468, n8469, n8471, n8472, n8473, n8475,
         n8476, n8477, n8478, n8485, n8486, n8503, n8504, n8521, n8522, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8538, n8539, n8556,
         n8557, n8574, n8575, n8587, n8588, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8614, n8615, n8633, n8634, n8645, n8646, n8647, n8649,
         n8650, n8651, n8652, n8659, n8660, n8678, n8679, n8697, n8698, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, U3558_n1, U3871_n1,
         U3991_n1, U5716_n1, U5717_n1, U5718_n1, U5719_n1, U5720_n1, U5721_n1,
         U5722_n1, U5723_n1, U5724_n1, U5725_n1, U5726_n1, U5727_n1, U5728_n1,
         U5729_n1, U5730_n1, U5731_n1, U5732_n1, U5733_n1, U5734_n1, U5735_n1,
         U5736_n1, U5737_n1, U5738_n1, U5739_n1, U5740_n1, U5741_n1, U5742_n1,
         U5743_n1, U5744_n1, U5745_n1, U5746_n1, U5747_n1, U5748_n1, U5749_n1,
         U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1,
         U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1,
         U5764_n1, U5765_n1, U5766_n1, U5767_n1, U5768_n1, U5769_n1, U5770_n1,
         U5771_n1, U5772_n1, U5773_n1, U5774_n1, U5775_n1, U5776_n1, U5777_n1,
         U5778_n1, U5779_n1, U5780_n1, U5781_n1, U5782_n1, U5783_n1, U5784_n1,
         U5785_n1, U5786_n1, U5787_n1, U5788_n1, U5789_n1, U5790_n1, U5791_n1,
         U5792_n1, U5793_n1, U5794_n1, U5795_n1, U5796_n1, U5797_n1, U5798_n1,
         U5799_n1, U5800_n1, U5801_n1, U5802_n1, U5803_n1, U5804_n1, U5805_n1,
         U5806_n1, U5807_n1, U5808_n1, U5809_n1, U5810_n1, U5811_n1, U5812_n1,
         U5813_n1, U5814_n1, U5815_n1, U5816_n1, U5817_n1, U5818_n1, U5819_n1,
         U5820_n1, U5821_n1, U5822_n1, U5823_n1, U5824_n1, U5825_n1, U5826_n1,
         U5827_n1, U5828_n1, U5829_n1, U5830_n1, U5831_n1, U5832_n1, U5833_n1,
         U5834_n1, U5835_n1, U5836_n1, U5837_n1, U5838_n1, U5839_n1, U5840_n1,
         U5841_n1, U5842_n1, U5843_n1, U5844_n1, U5845_n1, U5846_n1, U5847_n1,
         U5848_n1, U5849_n1, U5850_n1, U5851_n1, U5852_n1, U5853_n1, U5854_n1,
         U5855_n1, U5856_n1, U5857_n1, U5858_n1, U5859_n1, U5860_n1, U5861_n1,
         U5862_n1, U5863_n1, U5864_n1, U5865_n1, U5866_n1, U5867_n1, U5868_n1,
         U5869_n1, U5870_n1, U5871_n1, U5872_n1, U5873_n1, U5874_n1, U5875_n1,
         U5876_n1, U5877_n1, U5878_n1, U5879_n1, U5880_n1, U5881_n1, U5882_n1,
         U5883_n1, U5884_n1, U5885_n1, U5886_n1, U5887_n1, U5888_n1, U5889_n1,
         U5890_n1, U5891_n1, U5892_n1, U5893_n1, U5894_n1, U5895_n1, U5896_n1,
         U5897_n1, U5898_n1, U5899_n1, U5900_n1, U5901_n1, U5902_n1, U5903_n1,
         U5904_n1, U5905_n1, U5906_n1, U5907_n1, U5908_n1, U5909_n1, U5910_n1,
         U5911_n1, U5912_n1, U5913_n1, U5914_n1, U5915_n1, U5916_n1, U5917_n1,
         U5918_n1, U5919_n1, U5920_n1, U5921_n1, U5922_n1, U5923_n1, U5924_n1,
         U5925_n1, U5926_n1, U5927_n1, U5928_n1, U5929_n1, U5930_n1, U5931_n1,
         U5932_n1, U5933_n1, U5934_n1, U5935_n1, U5936_n1, U5937_n1, U5938_n1,
         U5939_n1, U5940_n1, U5941_n1, U5942_n1, U5943_n1, U5944_n1, U5945_n1,
         U5946_n1, U5947_n1, U5948_n1, U5949_n1, U5950_n1, U5951_n1, U5952_n1,
         U5953_n1, U5954_n1, U5955_n1, U5956_n1, U5957_n1, U5958_n1, U5959_n1,
         U5960_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1,
         U5967_n1, U5968_n1, U5969_n1, U5970_n1, U5971_n1, U5972_n1, U5973_n1,
         U5974_n1, U5975_n1, U5976_n1, U5977_n1, U5978_n1, U5979_n1, U5980_n1,
         U5981_n1, U5982_n1, U5983_n1, U5984_n1, U5985_n1, U5986_n1, U5987_n1,
         U5988_n1, U5989_n1, U5990_n1, U5991_n1, U5992_n1, U5993_n1, U5994_n1,
         U5995_n1, U5996_n1, U5997_n1, U5998_n1, U5999_n1, U6000_n1, U6001_n1,
         U6002_n1, U6003_n1, U6004_n1, U6005_n1, U6006_n1, U6007_n1, U6008_n1,
         U6009_n1, U6010_n1, U6011_n1, U6012_n1, U6013_n1, U6014_n1, U6015_n1,
         U6016_n1, U6017_n1, U6018_n1, U6019_n1, U6020_n1, U6021_n1, U6022_n1,
         U6023_n1, U6024_n1, U6025_n1, U6026_n1, U6027_n1, U6028_n1, U6029_n1,
         U6030_n1, U6031_n1, U6032_n1, U6033_n1, U6034_n1, U6035_n1, U6036_n1,
         U6037_n1, U6038_n1, U6039_n1, U6040_n1, U6041_n1, U6042_n1, U6043_n1,
         U6044_n1, U6045_n1, U6046_n1, U6047_n1, U6048_n1, U6049_n1, U6050_n1,
         U6051_n1, U6052_n1, U6053_n1, U6054_n1, U6055_n1, U6056_n1, U6057_n1,
         U6058_n1, U6059_n1, U6060_n1, U6061_n1, U6062_n1, U6063_n1, U6064_n1,
         U6065_n1, U6066_n1, U6067_n1, U6068_n1, U6069_n1, U6070_n1, U6071_n1,
         U6072_n1, U6073_n1, U6074_n1, U6075_n1, U6076_n1, U6077_n1, U6078_n1,
         U6079_n1, U6080_n1, U6081_n1, U6082_n1, U6083_n1, U6084_n1, U6085_n1,
         U6086_n1, U6087_n1, U6088_n1, U6089_n1, U6090_n1, U6091_n1, U6092_n1,
         U6093_n1, U6094_n1, U6095_n1, U6096_n1, U6097_n1, U6098_n1, U6099_n1,
         U6100_n1, U6101_n1, U6102_n1, U6103_n1, U6104_n1, U6105_n1, U6106_n1,
         U6107_n1, U6108_n1, U6109_n1, U6110_n1, U6111_n1, U6112_n1, U6113_n1,
         U6114_n1, U6115_n1, U6116_n1, U6117_n1, U6118_n1, U6119_n1, U6120_n1,
         U6121_n1, U6122_n1, U6123_n1, U6124_n1, U6125_n1, U6126_n1, U6127_n1,
         U6128_n1, U6129_n1, U6130_n1, U6131_n1, U6132_n1, U6133_n1, U6134_n1,
         U6135_n1, U6136_n1, U6137_n1, U6138_n1, U6139_n1, U6140_n1, U6141_n1,
         U6142_n1, U6143_n1, U6144_n1, U6145_n1, U6146_n1, U6147_n1, U6148_n1,
         U6149_n1, U6150_n1, U6151_n1, U6152_n1, U6153_n1, U6154_n1, U6155_n1,
         U6156_n1, U6157_n1, U6158_n1, U6159_n1, U6160_n1, U6161_n1, U6162_n1,
         U6163_n1, U6164_n1, U6165_n1, U6166_n1, U6167_n1, U6168_n1, U6169_n1,
         U6170_n1, U6171_n1, U6172_n1, U6173_n1, U6174_n1, U6175_n1, U6176_n1,
         U6177_n1, U6178_n1, U6179_n1, U6180_n1, U6181_n1, U6182_n1, U6183_n1,
         U6184_n1, U6185_n1, U6186_n1, U6187_n1, U6188_n1, U6189_n1, U6190_n1,
         U6191_n1, U6192_n1, U6193_n1, U6194_n1, U6195_n1, U6196_n1, U6197_n1,
         U6198_n1, U6199_n1, U6200_n1, U6201_n1, U6202_n1, U6203_n1, U6204_n1,
         U6205_n1, U6206_n1, U6207_n1, U6208_n1, U6209_n1, U6210_n1, U6211_n1,
         U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1,
         U6219_n1, U6220_n1, U6221_n1, U6222_n1, U6223_n1, U6224_n1, U6225_n1,
         U6226_n1, U6227_n1, U6228_n1, U6229_n1, U6230_n1, U6231_n1, U6232_n1,
         U6233_n1, U6234_n1, U6235_n1, U6236_n1, U6237_n1, U6238_n1, U6239_n1,
         U6240_n1, U6241_n1, U6242_n1, U6243_n1, U6244_n1, U6245_n1, U6246_n1,
         U6247_n1, U6248_n1, U6249_n1, U6250_n1, U6251_n1, U6252_n1, U6253_n1,
         U6254_n1, U6255_n1, U6256_n1, U6257_n1, U6258_n1, U6259_n1, U6260_n1,
         U6261_n1, U6262_n1, U6263_n1, U6264_n1, U6265_n1, U6266_n1, U6267_n1,
         U6268_n1, U6269_n1, U6270_n1, U6271_n1, U6272_n1, U6273_n1, U6274_n1,
         U6275_n1, U6276_n1, U6277_n1, U6278_n1, U6279_n1, U6280_n1, U6281_n1,
         U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1,
         U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6293_n1, U6294_n1, U6295_n1,
         U6296_n1, U6297_n1, U6298_n1, U6299_n1, U6300_n1, U6301_n1, U6302_n1,
         U6303_n1, U6304_n1, U6305_n1, U6306_n1, U6307_n1, U6308_n1, U6309_n1,
         U6310_n1, U6311_n1, U6312_n1, U6313_n1, U6314_n1, U6315_n1, U6316_n1,
         U6317_n1, U6318_n1, U6319_n1, U6320_n1, U6321_n1, U6322_n1, U6323_n1,
         U6324_n1, U6325_n1, U6326_n1, U6327_n1, U6328_n1, U6329_n1, U6330_n1,
         U6331_n1, U6332_n1, U6333_n1, U6334_n1, U6335_n1, U6336_n1, U6337_n1,
         U6338_n1, U6339_n1, U6340_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1,
         U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1,
         U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1,
         U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1,
         U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1,
         U6373_n1, U6374_n1, U6375_n1, U6376_n1, U6377_n1, U6378_n1, U6379_n1,
         U6380_n1, U6381_n1, U6382_n1, U6383_n1, U6384_n1, U6385_n1, U6386_n1,
         U6387_n1, U6388_n1, U6389_n1, U6390_n1, U6391_n1, U6392_n1, U6393_n1,
         U6394_n1, U6395_n1, U6396_n1, U6397_n1, U6398_n1, U6399_n1, U6400_n1,
         U6401_n1, U6402_n1, U6403_n1, U6404_n1, U6405_n1, U6406_n1, U6407_n1,
         U6408_n1, U6409_n1, U6410_n1, U6411_n1, U6412_n1, U6413_n1, U6414_n1,
         U6415_n1, U6416_n1, U6417_n1, U6418_n1, U6419_n1, U6420_n1, U6421_n1,
         U6422_n1, U6423_n1, U6424_n1, U6425_n1, U6426_n1, U6427_n1, U6428_n1,
         U6429_n1, U6430_n1, U6431_n1, U6432_n1, U6433_n1, U6434_n1, U6435_n1,
         U6436_n1, U6437_n1, U6438_n1, U6439_n1, U6440_n1, U6441_n1, U6442_n1,
         U6443_n1, U6444_n1, U6445_n1, U6446_n1, U6447_n1, U6448_n1, U6449_n1,
         U6450_n1, U6451_n1, U6452_n1, U6453_n1, U6454_n1, U6455_n1, U6456_n1,
         U6457_n1, U6458_n1, U6459_n1, U6460_n1, U6461_n1, U6462_n1, U6463_n1,
         U6464_n1, U6465_n1, U6466_n1, U6467_n1, U6468_n1, U6469_n1, U6470_n1,
         U6471_n1, U6472_n1, U6473_n1, U6474_n1, U6475_n1, U6476_n1, U6477_n1,
         U6478_n1, U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n9625), .CLK(n9771), .Q(
        WX485) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n9620), .CLK(n9773), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n9620), .CLK(n9773), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n9621), .CLK(n9773), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n9621), .CLK(n9773), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n9621), .CLK(n9773), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n9621), .CLK(n9773), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n9621), .CLK(n9773), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n9621), .CLK(n9773), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n9622), .CLK(n9772), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n9622), .CLK(n9772), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n9622), .CLK(n9772), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n9622), .CLK(n9772), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n9622), .CLK(n9772), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n9622), .CLK(n9772), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n9623), .CLK(n9772), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n9623), .CLK(n9772), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n9623), .CLK(n9772), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n9623), .CLK(n9772), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n9623), .CLK(n9772), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n9623), .CLK(n9772), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n9624), .CLK(n9771), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n9624), .CLK(n9771), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n9624), .CLK(n9771), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n9624), .CLK(n9771), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n9624), .CLK(n9771), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n9624), .CLK(n9771), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n9625), .CLK(n9771), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n9625), .CLK(n9771), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n9625), .CLK(n9771), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n9625), .CLK(n9771), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n9625), .CLK(n9771), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n9620), .CLK(n9773), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n9620), .CLK(n9773), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n9620), .CLK(n9773), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n9620), .CLK(n9773), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n9619), .CLK(n9774), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n9619), .CLK(n9774), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n9619), .CLK(n9774), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n9618), .CLK(n9774), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n9618), .CLK(n9774), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n9618), .CLK(n9774), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n9617), .CLK(n9775), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n9617), .CLK(n9775), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n9617), .CLK(n9775), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n9616), .CLK(n9775), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n9616), .CLK(n9775), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n9615), .CLK(n9776), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n9615), .CLK(n9776), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n9614), .CLK(n9776), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n9613), .CLK(n9777), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n9613), .CLK(n9777), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n9612), .CLK(n9777), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n9611), .CLK(n9778), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n9610), .CLK(n9778), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n9610), .CLK(n9778), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n9609), .CLK(n9779), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n9609), .CLK(n9779), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n9608), .CLK(n9779), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n9607), .CLK(n9780), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n9607), .CLK(n9780), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n9606), .CLK(n9780), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n9605), .CLK(n9781), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n9605), .CLK(n9781), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n9604), .CLK(n9781), .Q(
        WX709), .QN(n8773) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n9603), .CLK(n9782), .Q(
        WX711), .QN(n8678) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n9603), .CLK(n9782), .Q(
        WX713), .QN(n8710) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n9619), .CLK(n9774), .Q(
        WX715), .QN(n8719) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n9619), .CLK(n9774), .Q(
        WX717), .QN(n8725) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n9619), .CLK(n9774), .Q(
        WX719), .QN(n8728) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n9618), .CLK(n9774), .Q(
        WX721), .QN(n8737) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n9618), .CLK(n9774), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n9618), .CLK(n9774), .Q(
        WX725), .QN(n8748) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n9617), .CLK(n9775), .Q(
        WX727), .QN(n8760) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n9617), .CLK(n9775), .Q(
        WX729), .QN(n8766) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n9617), .CLK(n9775), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n9616), .CLK(n9775), .Q(
        WX733), .QN(n8707) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n9616), .CLK(n9775), .Q(
        WX735), .QN(n8722) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n9615), .CLK(n9776), .Q(
        WX737), .QN(n8734) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n9615), .CLK(n9776), .Q(
        WX739), .QN(n8749) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n9614), .CLK(n9776), .Q(
        WX741), .QN(n8763) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n9614), .CLK(n9776), .Q(
        WX743), .QN(n8778) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n9613), .CLK(n9777), .Q(
        WX745), .QN(n8713) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n9612), .CLK(n9777), .Q(
        WX747), .QN(n8740) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n9612), .CLK(n9777), .Q(
        WX749), .QN(n8786) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n9611), .CLK(n9778), .Q(
        WX751), .QN(n8731) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n9611), .CLK(n9778), .Q(
        WX753), .QN(n8741) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n9610), .CLK(n9778), .Q(
        WX755), .QN(n8753) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n9609), .CLK(n9779), .Q(
        WX757), .QN(n8781) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n9608), .CLK(n9779), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n9608), .CLK(n9779), .Q(
        WX761), .QN(n8756) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n9607), .CLK(n9780), .Q(
        WX763), .QN(n8759) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n9606), .CLK(n9780), .Q(
        WX765), .QN(n8704) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n9606), .CLK(n9780), .Q(
        WX767), .QN(n8779) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n9605), .CLK(n9781), .Q(
        WX769), .QN(n8715) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n9604), .CLK(n9781), .Q(
        WX771), .QN(n8787) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n9604), .CLK(n9781), .Q(
        WX773), .QN(n8774) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n9603), .CLK(n9782), .Q(
        WX775), .QN(n8679) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n9603), .CLK(n9782), .Q(
        WX777), .QN(n8708) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n9602), .CLK(n9782), .Q(
        WX779), .QN(n8717) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n9602), .CLK(n9782), .Q(
        WX781), .QN(n8723) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n9602), .CLK(n9782), .Q(
        WX783), .QN(n8726) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n9601), .CLK(n9783), .Q(
        WX785), .QN(n8735) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n9601), .CLK(n9783), .Q(
        WX787), .QN(n8744) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n9601), .CLK(n9783), .Q(
        WX789), .QN(n8746) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n9600), .CLK(n9783), .Q(
        WX791), .QN(n8761) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n9600), .CLK(n9783), .Q(
        WX793), .QN(n8767) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n9600), .CLK(n9783), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n9616), .CLK(n9775), 
        .Q(WX797), .QN(n8705) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n9616), .CLK(n9775), .Q(
        WX799), .QN(n8720) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n9615), .CLK(n9776), .Q(
        WX801), .QN(n8732) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n9615), .CLK(n9776), .Q(
        WX803), .QN(n8750) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n9614), .CLK(n9776), .Q(
        WX805), .QN(n8764) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n9614), .CLK(n9776), .Q(
        WX807), .QN(n8776) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n9613), .CLK(n9777), .Q(
        WX809), .QN(n8711) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n9612), .CLK(n9777), .Q(
        WX811), .QN(n8738) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n9612), .CLK(n9777), .Q(
        WX813), .QN(n8784) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n9611), .CLK(n9778), .Q(
        WX815), .QN(n8729) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n9610), .CLK(n9778), .Q(
        WX817), .QN(n8742) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n9610), .CLK(n9778), .Q(
        WX819), .QN(n8751) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n9609), .CLK(n9779), .Q(
        WX821), .QN(n8782) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n9608), .CLK(n9779), .Q(
        WX823), .QN(n8769) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n9608), .CLK(n9779), .Q(
        WX825), .QN(n8754) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n9607), .CLK(n9780), .Q(
        WX827), .QN(n8757) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n9606), .CLK(n9780), .Q(
        WX829), .QN(n8698) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n9606), .CLK(n9780), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n9605), .CLK(n9781), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n9604), .CLK(n9781), .Q(
        WX835), .QN(n8788) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n9604), .CLK(n9781), .Q(
        WX837), .QN(n8775) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n9603), .CLK(n9782), .Q(
        WX839), .QN(n8697) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n9603), .CLK(n9782), .Q(
        WX841), .QN(n8709) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n9602), .CLK(n9782), .Q(
        WX843), .QN(n8718) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n9602), .CLK(n9782), .Q(
        WX845), .QN(n8724) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n9602), .CLK(n9782), .Q(
        WX847), .QN(n8727) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n9601), .CLK(n9783), .Q(
        WX849), .QN(n8736) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n9601), .CLK(n9783), .Q(
        WX851), .QN(n8745) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n9601), .CLK(n9783), .Q(
        WX853), .QN(n8747) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n9600), .CLK(n9783), .Q(
        WX855), .QN(n8762) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n9600), .CLK(n9783), .Q(
        WX857), .QN(n8768) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n9600), .CLK(n9783), .Q(
        WX859), .QN(n8771) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n9599), .CLK(n9784), .Q(
        WX861), .QN(n8706) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n9599), .CLK(n9784), .Q(
        WX863), .QN(n8721) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n9599), .CLK(n9784), .Q(
        WX865), .QN(n8733) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n9599), .CLK(n9784), .Q(
        test_so8), .QN(n8798) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n9614), .CLK(n9776), 
        .Q(WX869), .QN(n8765) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n9613), .CLK(n9777), .Q(
        WX871), .QN(n8777) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n9613), .CLK(n9777), .Q(
        WX873), .QN(n8712) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n9612), .CLK(n9777), .Q(
        WX875), .QN(n8739) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n9611), .CLK(n9778), .Q(
        WX877), .QN(n8785) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n9611), .CLK(n9778), .Q(
        WX879), .QN(n8730) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n9610), .CLK(n9778), .Q(
        WX881), .QN(n8743) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n9609), .CLK(n9779), .Q(
        WX883), .QN(n8752) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n9609), .CLK(n9779), .Q(
        WX885), .QN(n8783) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n9608), .CLK(n9779), .Q(
        WX887), .QN(n8770) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n9607), .CLK(n9780), .Q(
        WX889), .QN(n8755) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n9607), .CLK(n9780), .Q(
        WX891), .QN(n8758) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n9606), .CLK(n9780), .Q(
        WX893), .QN(n8703) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n9605), .CLK(n9781), .Q(
        WX895) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n9605), .CLK(n9781), .Q(
        WX897), .QN(n8714) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n9604), .CLK(n9781), .Q(
        WX899), .QN(n8789) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n9341), .CLK(n9913), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n9341), .CLK(n9913), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n9340), .CLK(n9913), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n9339), .CLK(n9914), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n9339), .CLK(n9914), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n9339), .CLK(n9914), 
        .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n9339), .CLK(n9914), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n9339), .CLK(n9914), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n9339), .CLK(n9914), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n9338), .CLK(n9914), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n9338), .CLK(n9914), .Q(CRC_OUT_9_15) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n9338), .CLK(n9914), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n9338), .CLK(n9914), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n9338), .CLK(n9914), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n9338), .CLK(n9914), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n9599), .CLK(n9784), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n9599), .CLK(n9784), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n9598), .CLK(n9784), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n9597), .CLK(n9785), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n9597), .CLK(n9785), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n9597), .CLK(n9785), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n9597), .CLK(n9785), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n250), .SI(CRC_OUT_9_31), .SE(n9597), .CLK(n9785), 
        .Q(WX1778) );
  SDFFX1 DFF_193_Q_reg ( .D(n251), .SI(WX1778), .SE(n9592), .CLK(n9787), .Q(
        n8702), .QN(n9031) );
  SDFFX1 DFF_194_Q_reg ( .D(n252), .SI(n8702), .SE(n9592), .CLK(n9787), .Q(
        n8701), .QN(n9030) );
  SDFFX1 DFF_195_Q_reg ( .D(n253), .SI(n8701), .SE(n9592), .CLK(n9787), .Q(
        n8700), .QN(n9029) );
  SDFFX1 DFF_196_Q_reg ( .D(n254), .SI(n8700), .SE(n9592), .CLK(n9787), .Q(
        n8699), .QN(n9028) );
  SDFFX1 DFF_197_Q_reg ( .D(n255), .SI(n8699), .SE(n9592), .CLK(n9787), .Q(
        test_so11), .QN(n9074) );
  SDFFX1 DFF_198_Q_reg ( .D(n256), .SI(test_si12), .SE(n9592), .CLK(n9787), 
        .Q(n8696), .QN(n9027) );
  SDFFX1 DFF_199_Q_reg ( .D(n257), .SI(n8696), .SE(n9593), .CLK(n9787), .Q(
        n8695), .QN(n9026) );
  SDFFX1 DFF_200_Q_reg ( .D(n258), .SI(n8695), .SE(n9593), .CLK(n9787), .Q(
        n8694), .QN(n9025) );
  SDFFX1 DFF_201_Q_reg ( .D(n259), .SI(n8694), .SE(n9593), .CLK(n9787), .Q(
        n8693), .QN(n9024) );
  SDFFX1 DFF_202_Q_reg ( .D(n260), .SI(n8693), .SE(n9593), .CLK(n9787), .Q(
        n8692), .QN(n9023) );
  SDFFX1 DFF_203_Q_reg ( .D(n261), .SI(n8692), .SE(n9593), .CLK(n9787), .Q(
        n8691), .QN(n9022) );
  SDFFX1 DFF_204_Q_reg ( .D(n262), .SI(n8691), .SE(n9593), .CLK(n9787), .Q(
        n8690), .QN(n9021) );
  SDFFX1 DFF_205_Q_reg ( .D(n263), .SI(n8690), .SE(n9594), .CLK(n9786), .Q(
        n8689), .QN(n9020) );
  SDFFX1 DFF_206_Q_reg ( .D(n264), .SI(n8689), .SE(n9594), .CLK(n9786), .Q(
        n8688), .QN(n9019) );
  SDFFX1 DFF_207_Q_reg ( .D(n265), .SI(n8688), .SE(n9594), .CLK(n9786), .Q(
        n8687), .QN(n9018) );
  SDFFX1 DFF_208_Q_reg ( .D(n266), .SI(n8687), .SE(n9594), .CLK(n9786), .Q(
        n8686), .QN(n9017) );
  SDFFX1 DFF_209_Q_reg ( .D(n267), .SI(n8686), .SE(n9594), .CLK(n9786), .Q(
        n8685), .QN(n9016) );
  SDFFX1 DFF_210_Q_reg ( .D(n268), .SI(n8685), .SE(n9594), .CLK(n9786), .Q(
        n8684), .QN(n9015) );
  SDFFX1 DFF_211_Q_reg ( .D(n269), .SI(n8684), .SE(n9595), .CLK(n9786), .Q(
        n8683), .QN(n9014) );
  SDFFX1 DFF_212_Q_reg ( .D(n270), .SI(n8683), .SE(n9595), .CLK(n9786), .Q(
        n8682), .QN(n9013) );
  SDFFX1 DFF_213_Q_reg ( .D(n271), .SI(n8682), .SE(n9595), .CLK(n9786), .Q(
        n8681), .QN(n9012) );
  SDFFX1 DFF_214_Q_reg ( .D(n272), .SI(n8681), .SE(n9595), .CLK(n9786), .Q(
        n8680), .QN(n9011) );
  SDFFX1 DFF_215_Q_reg ( .D(n273), .SI(n8680), .SE(n9595), .CLK(n9786), .Q(
        test_so12), .QN(n9073) );
  SDFFX1 DFF_216_Q_reg ( .D(n274), .SI(test_si13), .SE(n9595), .CLK(n9786), 
        .Q(n8677), .QN(n9010) );
  SDFFX1 DFF_217_Q_reg ( .D(n275), .SI(n8677), .SE(n9596), .CLK(n9785), .Q(
        n8676), .QN(n9009) );
  SDFFX1 DFF_218_Q_reg ( .D(n276), .SI(n8676), .SE(n9596), .CLK(n9785), .Q(
        n8675), .QN(n9008) );
  SDFFX1 DFF_219_Q_reg ( .D(n277), .SI(n8675), .SE(n9596), .CLK(n9785), .Q(
        n8674), .QN(n9007) );
  SDFFX1 DFF_220_Q_reg ( .D(n278), .SI(n8674), .SE(n9596), .CLK(n9785), .Q(
        n8673), .QN(n9006) );
  SDFFX1 DFF_221_Q_reg ( .D(n279), .SI(n8673), .SE(n9596), .CLK(n9785), .Q(
        n8672), .QN(n9005) );
  SDFFX1 DFF_222_Q_reg ( .D(n280), .SI(n8672), .SE(n9596), .CLK(n9785), .Q(
        n8671), .QN(n9004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n9597), .CLK(n9785), .Q(
        n8670), .QN(n9003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n9591), .CLK(n9788), .Q(
        n8669), .QN(n16307) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n9591), .CLK(n9788), .Q(
        n8668), .QN(n16308) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n9590), .CLK(n9788), .Q(
        n8667), .QN(n16309) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n9590), .CLK(n9788), .Q(
        n8666), .QN(n16310) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n9589), .CLK(n9789), .Q(
        n8665), .QN(n16311) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n9588), .CLK(n9789), .Q(
        n8664), .QN(n16312) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n9588), .CLK(n9789), .Q(
        n8663), .QN(n16313) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n9587), .CLK(n9790), .Q(
        n8662), .QN(n16314) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n9587), .CLK(n9790), .Q(
        n8661), .QN(n16315) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n9341), .CLK(n9913), .Q(
        test_so13), .QN(n8825) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n9585), .CLK(n9791), 
        .Q(n8658), .QN(n16316) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n9585), .CLK(n9791), .Q(
        n8657), .QN(n16317) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n9584), .CLK(n9791), .Q(
        n8656), .QN(n16318) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n9584), .CLK(n9791), .Q(
        n8655), .QN(n16319) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n9583), .CLK(n9792), .Q(
        n8654), .QN(n16320) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n9582), .CLK(n9792), .Q(
        n8653), .QN(n16321) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n9582), .CLK(n9792), .Q(
        WX1970), .QN(n8094) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n9581), .CLK(n9793), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n9580), .CLK(n9793), .Q(
        WX1974), .QN(n8091) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n9580), .CLK(n9793), .Q(
        WX1976), .QN(n8089) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n9579), .CLK(n9794), .Q(
        WX1978), .QN(n8087) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n9578), .CLK(n9794), .Q(
        WX1980), .QN(n8085) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n9578), .CLK(n9794), .Q(
        WX1982), .QN(n8083) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n9577), .CLK(n9795), .Q(
        WX1984), .QN(n8081) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n9576), .CLK(n9795), .Q(
        WX1986), .QN(n8079) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n9576), .CLK(n9795), .Q(
        WX1988), .QN(n8077) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n9575), .CLK(n9796), .Q(
        WX1990), .QN(n8075) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n9574), .CLK(n9796), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n9573), .CLK(n9797), 
        .Q(WX1994), .QN(n8072) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n9573), .CLK(n9797), .Q(
        WX1996), .QN(n8070) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n9572), .CLK(n9797), .Q(
        WX1998), .QN(n8068) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n9572), .CLK(n9797), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n9591), .CLK(n9788), .Q(
        WX2002), .QN(n7626) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n9591), .CLK(n9788), .Q(
        WX2004), .QN(n7852) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n9590), .CLK(n9788), .Q(
        WX2006), .QN(n7850) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n9590), .CLK(n9788), .Q(
        WX2008), .QN(n7848) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n9589), .CLK(n9789), .Q(
        WX2010), .QN(n7846) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n9589), .CLK(n9789), .Q(
        WX2012), .QN(n7844) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n9588), .CLK(n9789), .Q(
        WX2014), .QN(n7842) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n9587), .CLK(n9790), .Q(
        WX2016), .QN(n7840) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n9587), .CLK(n9790), .Q(
        WX2018), .QN(n7838) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n9586), .CLK(n9790), .Q(
        WX2020), .QN(n7836) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n9586), .CLK(n9790), .Q(
        WX2022), .QN(n7834) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n9585), .CLK(n9791), .Q(
        WX2024), .QN(n7832) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n9584), .CLK(n9791), .Q(
        WX2026), .QN(n7830) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n9583), .CLK(n9792), .Q(
        test_so15), .QN(n8815) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n9582), .CLK(n9792), 
        .Q(WX2030), .QN(n7827) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n9582), .CLK(n9792), .Q(
        WX2032), .QN(n7825) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n9581), .CLK(n9793), .Q(
        WX2034) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n9581), .CLK(n9793), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n9580), .CLK(n9793), .Q(
        WX2038) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n9579), .CLK(n9794), .Q(
        WX2040) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n9579), .CLK(n9794), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n9578), .CLK(n9794), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n9577), .CLK(n9795), .Q(
        WX2046) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n9577), .CLK(n9795), .Q(
        WX2048) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n9576), .CLK(n9795), .Q(
        WX2050) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n9575), .CLK(n9796), .Q(
        WX2052) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n9575), .CLK(n9796), .Q(
        WX2054) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n9574), .CLK(n9796), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n9574), .CLK(n9796), .Q(
        WX2058) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n9573), .CLK(n9797), .Q(
        WX2060) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n9572), .CLK(n9797), .Q(
        WX2062) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n9571), .CLK(n9798), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n9591), .CLK(n9788), 
        .Q(WX2066), .QN(n7627) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n9591), .CLK(n9788), .Q(
        WX2068), .QN(n7853) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n9590), .CLK(n9788), .Q(
        WX2070), .QN(n7851) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n9590), .CLK(n9788), .Q(
        WX2072), .QN(n7849) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n9589), .CLK(n9789), .Q(
        WX2074), .QN(n7847) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n9589), .CLK(n9789), .Q(
        WX2076), .QN(n7845) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n9588), .CLK(n9789), .Q(
        WX2078), .QN(n7843) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n9587), .CLK(n9790), .Q(
        WX2080), .QN(n7841) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n9586), .CLK(n9790), .Q(
        WX2082), .QN(n7839) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n9586), .CLK(n9790), .Q(
        WX2084), .QN(n7837) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n9585), .CLK(n9791), .Q(
        WX2086), .QN(n7835) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n9585), .CLK(n9791), .Q(
        WX2088), .QN(n7833) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n9584), .CLK(n9791), .Q(
        WX2090), .QN(n7831) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n9583), .CLK(n9792), .Q(
        WX2092), .QN(n7829) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n9583), .CLK(n9792), .Q(
        WX2094), .QN(n7828) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n9582), .CLK(n9792), .Q(
        WX2096), .QN(n7826) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n9581), .CLK(n9793), .Q(
        WX2098), .QN(n8095) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n9581), .CLK(n9793), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n9580), .CLK(n9793), 
        .Q(WX2102), .QN(n8092) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n9579), .CLK(n9794), .Q(
        WX2104), .QN(n8090) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n9579), .CLK(n9794), .Q(
        WX2106), .QN(n8088) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n9578), .CLK(n9794), .Q(
        WX2108), .QN(n8086) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n9577), .CLK(n9795), .Q(
        WX2110), .QN(n8084) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n9577), .CLK(n9795), .Q(
        WX2112), .QN(n8082) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n9576), .CLK(n9795), .Q(
        WX2114), .QN(n8080) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n9575), .CLK(n9796), .Q(
        WX2116), .QN(n8078) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n9575), .CLK(n9796), .Q(
        WX2118), .QN(n8076) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n9574), .CLK(n9796), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n9573), .CLK(n9797), .Q(
        WX2122), .QN(n8073) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n9573), .CLK(n9797), .Q(
        WX2124), .QN(n8071) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n9572), .CLK(n9797), .Q(
        WX2126), .QN(n8069) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n9571), .CLK(n9798), .Q(
        WX2128), .QN(n8067) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n9571), .CLK(n9798), .Q(
        WX2130), .QN(n8574) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n9571), .CLK(n9798), .Q(
        WX2132), .QN(n8575) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n9571), .CLK(n9798), .Q(
        WX2134), .QN(n8587) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n9570), .CLK(n9798), .Q(
        test_so18), .QN(n8803) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n9589), .CLK(n9789), 
        .Q(WX2138), .QN(n8588) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n9588), .CLK(n9789), .Q(
        WX2140) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n9588), .CLK(n9789), .Q(
        WX2142), .QN(n8590) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n9587), .CLK(n9790), .Q(
        WX2144), .QN(n8591) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n9586), .CLK(n9790), .Q(
        WX2146), .QN(n8592) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n9586), .CLK(n9790), .Q(
        WX2148), .QN(n8593) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n9585), .CLK(n9791), .Q(
        WX2150), .QN(n8594) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n9584), .CLK(n9791), .Q(
        WX2152), .QN(n8595) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n9584), .CLK(n9791), .Q(
        WX2154), .QN(n8596) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n9583), .CLK(n9792), .Q(
        WX2156), .QN(n8614) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n9583), .CLK(n9792), .Q(
        WX2158), .QN(n8615) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n9582), .CLK(n9792), .Q(
        WX2160), .QN(n8123) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n9581), .CLK(n9793), .Q(
        WX2162), .QN(n8633) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n9580), .CLK(n9793), .Q(
        WX2164), .QN(n8634) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n9580), .CLK(n9793), .Q(
        WX2166), .QN(n8645) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n9579), .CLK(n9794), .Q(
        WX2168), .QN(n8646) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n9578), .CLK(n9794), .Q(
        WX2170), .QN(n8124) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n9578), .CLK(n9794), .Q(
        test_so19), .QN(n8793) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n9577), .CLK(n9795), 
        .Q(WX2174), .QN(n8647) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n9576), .CLK(n9795), .Q(
        WX2176) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n9576), .CLK(n9795), .Q(
        WX2178), .QN(n8649) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n9575), .CLK(n9796), .Q(
        WX2180), .QN(n8650) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n9574), .CLK(n9796), .Q(
        WX2182), .QN(n8651) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n9574), .CLK(n9796), .Q(
        WX2184), .QN(n8125) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n9573), .CLK(n9797), .Q(
        WX2186), .QN(n8652) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n9572), .CLK(n9797), .Q(
        WX2188), .QN(n8659) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n9572), .CLK(n9797), .Q(
        WX2190), .QN(n8660) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n9571), .CLK(n9798), .Q(
        WX2192), .QN(n8133) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n9346), .CLK(n9910), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n9346), .CLK(n9910), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n9346), .CLK(n9910), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n9346), .CLK(n9910), 
        .Q(CRC_OUT_8_3) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n9345), .CLK(n9911), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n9345), .CLK(n9911), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n9345), .CLK(n9911), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n9345), .CLK(n9911), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n9345), .CLK(n9911), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n9345), .CLK(n9911), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n9344), .CLK(n9911), 
        .Q(CRC_OUT_8_10) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n9344), .CLK(n9911), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n9344), .CLK(n9911), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n9344), .CLK(n9911), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n9344), .CLK(n9911), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n9344), .CLK(n9911), .Q(CRC_OUT_8_15) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n9343), .CLK(n9912), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n9342), .CLK(n9912), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n9342), .CLK(n9912), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n9342), .CLK(n9912), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n9342), .CLK(n9912), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n9342), .CLK(n9912), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n9342), .CLK(n9912), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n9341), .CLK(n9913), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n9341), .CLK(n9913), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n9341), .CLK(n9913), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n9570), .CLK(n9798), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n491), .SI(CRC_OUT_8_31), .SE(n9570), .CLK(n9798), 
        .Q(WX3071) );
  SDFFX1 DFF_385_Q_reg ( .D(n492), .SI(WX3071), .SE(n9565), .CLK(n9801), .Q(
        n8644), .QN(n9002) );
  SDFFX1 DFF_386_Q_reg ( .D(n493), .SI(n8644), .SE(n9565), .CLK(n9801), .Q(
        n8643), .QN(n9001) );
  SDFFX1 DFF_387_Q_reg ( .D(n494), .SI(n8643), .SE(n9565), .CLK(n9801), .Q(
        n8642), .QN(n9000) );
  SDFFX1 DFF_388_Q_reg ( .D(n495), .SI(n8642), .SE(n9565), .CLK(n9801), .Q(
        n8641), .QN(n8999) );
  SDFFX1 DFF_389_Q_reg ( .D(n496), .SI(n8641), .SE(n9566), .CLK(n9800), .Q(
        n8640), .QN(n8998) );
  SDFFX1 DFF_390_Q_reg ( .D(n497), .SI(n8640), .SE(n9566), .CLK(n9800), .Q(
        n8639), .QN(n8997) );
  SDFFX1 DFF_391_Q_reg ( .D(n498), .SI(n8639), .SE(n9566), .CLK(n9800), .Q(
        n8638), .QN(n8996) );
  SDFFX1 DFF_392_Q_reg ( .D(n499), .SI(n8638), .SE(n9566), .CLK(n9800), .Q(
        n8637), .QN(n8995) );
  SDFFX1 DFF_393_Q_reg ( .D(n500), .SI(n8637), .SE(n9566), .CLK(n9800), .Q(
        n8636), .QN(n8994) );
  SDFFX1 DFF_394_Q_reg ( .D(n501), .SI(n8636), .SE(n9566), .CLK(n9800), .Q(
        n8635), .QN(n8993) );
  SDFFX1 DFF_395_Q_reg ( .D(n502), .SI(n8635), .SE(n9567), .CLK(n9800), .Q(
        test_so22), .QN(n9072) );
  SDFFX1 DFF_396_Q_reg ( .D(n503), .SI(test_si23), .SE(n9567), .CLK(n9800), 
        .Q(n8632), .QN(n8992) );
  SDFFX1 DFF_397_Q_reg ( .D(n504), .SI(n8632), .SE(n9567), .CLK(n9800), .Q(
        n8631), .QN(n8991) );
  SDFFX1 DFF_398_Q_reg ( .D(n505), .SI(n8631), .SE(n9567), .CLK(n9800), .Q(
        n8630), .QN(n8990) );
  SDFFX1 DFF_399_Q_reg ( .D(n506), .SI(n8630), .SE(n9567), .CLK(n9800), .Q(
        n8629), .QN(n8989) );
  SDFFX1 DFF_400_Q_reg ( .D(n510), .SI(n8629), .SE(n9567), .CLK(n9800), .Q(
        n8628), .QN(n8988) );
  SDFFX1 DFF_401_Q_reg ( .D(n511), .SI(n8628), .SE(n9568), .CLK(n9799), .Q(
        n8627), .QN(n8987) );
  SDFFX1 DFF_402_Q_reg ( .D(n512), .SI(n8627), .SE(n9568), .CLK(n9799), .Q(
        n8626), .QN(n8986) );
  SDFFX1 DFF_403_Q_reg ( .D(n513), .SI(n8626), .SE(n9568), .CLK(n9799), .Q(
        n8625), .QN(n8985) );
  SDFFX1 DFF_404_Q_reg ( .D(n514), .SI(n8625), .SE(n9568), .CLK(n9799), .Q(
        n8624), .QN(n8984) );
  SDFFX1 DFF_405_Q_reg ( .D(n515), .SI(n8624), .SE(n9568), .CLK(n9799), .Q(
        n8623), .QN(n8983) );
  SDFFX1 DFF_406_Q_reg ( .D(n516), .SI(n8623), .SE(n9568), .CLK(n9799), .Q(
        n8622), .QN(n8982) );
  SDFFX1 DFF_407_Q_reg ( .D(n517), .SI(n8622), .SE(n9569), .CLK(n9799), .Q(
        n8621), .QN(n8981) );
  SDFFX1 DFF_408_Q_reg ( .D(n518), .SI(n8621), .SE(n9569), .CLK(n9799), .Q(
        n8620), .QN(n8980) );
  SDFFX1 DFF_409_Q_reg ( .D(n519), .SI(n8620), .SE(n9569), .CLK(n9799), .Q(
        n8619), .QN(n8979) );
  SDFFX1 DFF_410_Q_reg ( .D(n520), .SI(n8619), .SE(n9569), .CLK(n9799), .Q(
        n8618), .QN(n8978) );
  SDFFX1 DFF_411_Q_reg ( .D(n521), .SI(n8618), .SE(n9569), .CLK(n9799), .Q(
        n8617), .QN(n8977) );
  SDFFX1 DFF_412_Q_reg ( .D(n522), .SI(n8617), .SE(n9569), .CLK(n9799), .Q(
        n8616), .QN(n8976) );
  SDFFX1 DFF_413_Q_reg ( .D(n523), .SI(n8616), .SE(n9570), .CLK(n9798), .Q(
        test_so23), .QN(n9071) );
  SDFFX1 DFF_414_Q_reg ( .D(n524), .SI(test_si24), .SE(n9570), .CLK(n9798), 
        .Q(n8613), .QN(n8975) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n9570), .CLK(n9798), .Q(
        n8612), .QN(n8974) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n9565), .CLK(n9801), .Q(
        n8611), .QN(n16322) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n9564), .CLK(n9801), .Q(
        n8610), .QN(n16323) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n9564), .CLK(n9801), .Q(
        n8609), .QN(n16324) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n9564), .CLK(n9801), .Q(
        n8608), .QN(n16325) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n9563), .CLK(n9802), .Q(
        n8607), .QN(n16326) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n9563), .CLK(n9802), .Q(
        n8606), .QN(n16327) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n9563), .CLK(n9802), .Q(
        n8605), .QN(n16328) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n9562), .CLK(n9802), .Q(
        n8604), .QN(n16329) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n9562), .CLK(n9802), .Q(
        n8603), .QN(n16330) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n9561), .CLK(n9803), .Q(
        n8602), .QN(n16331) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n9561), .CLK(n9803), .Q(
        n8601), .QN(n16332) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n9559), .CLK(n9804), .Q(
        n8600), .QN(n16333) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n9559), .CLK(n9804), .Q(
        n8599), .QN(n16334) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n9558), .CLK(n9804), .Q(
        n8598), .QN(n16335) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n9558), .CLK(n9804), .Q(
        n8597), .QN(n16336) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n9557), .CLK(n9805), .Q(
        test_so24), .QN(n8824) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n9555), .CLK(n9806), 
        .Q(WX3263), .QN(n8064) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n9554), .CLK(n9806), .Q(
        WX3265), .QN(n8062) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n9553), .CLK(n9807), .Q(
        WX3267), .QN(n8060) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n9553), .CLK(n9807), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n9552), .CLK(n9807), .Q(
        WX3271), .QN(n8056) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n9551), .CLK(n9808), .Q(
        WX3273), .QN(n8054) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n9551), .CLK(n9808), .Q(
        WX3275), .QN(n8052) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n9550), .CLK(n9808), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n9549), .CLK(n9809), .Q(
        WX3279), .QN(n8049) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n9549), .CLK(n9809), .Q(
        WX3281), .QN(n8047) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n9548), .CLK(n9809), .Q(
        WX3283), .QN(n8045) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n9547), .CLK(n9810), .Q(
        WX3285), .QN(n8043) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n9547), .CLK(n9810), .Q(
        WX3287), .QN(n8041) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n9546), .CLK(n9810), .Q(
        WX3289), .QN(n8039) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n9545), .CLK(n9811), .Q(
        WX3291), .QN(n8037) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n9545), .CLK(n9811), .Q(
        WX3293), .QN(n8035) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n9565), .CLK(n9801), .Q(
        WX3295), .QN(n7624) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n9564), .CLK(n9801), .Q(
        test_so25), .QN(n8817) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n9564), .CLK(n9801), 
        .Q(WX3299), .QN(n7822) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n9564), .CLK(n9801), .Q(
        WX3301), .QN(n7820) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n9563), .CLK(n9802), .Q(
        WX3303), .QN(n7818) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n9563), .CLK(n9802), .Q(
        WX3305), .QN(n7817) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n9563), .CLK(n9802), .Q(
        WX3307), .QN(n7815) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n9562), .CLK(n9802), .Q(
        WX3309), .QN(n7813) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n9562), .CLK(n9802), .Q(
        WX3311), .QN(n7811) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n9561), .CLK(n9803), .Q(
        WX3313), .QN(n7809) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n9560), .CLK(n9803), .Q(
        WX3315), .QN(n7807) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n9560), .CLK(n9803), .Q(
        WX3317), .QN(n7805) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n9559), .CLK(n9804), .Q(
        WX3319), .QN(n7803) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n9559), .CLK(n9804), .Q(
        WX3321), .QN(n7801) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n9558), .CLK(n9804), .Q(
        WX3323), .QN(n7799) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n9557), .CLK(n9805), .Q(
        WX3325), .QN(n7797) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n9554), .CLK(n9806), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n9554), .CLK(n9806), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n9553), .CLK(n9807), .Q(
        WX3331) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n9552), .CLK(n9807), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n9552), .CLK(n9807), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n9551), .CLK(n9808), .Q(
        WX3337) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n9550), .CLK(n9808), .Q(
        WX3339) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n9550), .CLK(n9808), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n9549), .CLK(n9809), .Q(
        WX3343) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n9548), .CLK(n9809), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n9548), .CLK(n9809), .Q(
        WX3347) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n9547), .CLK(n9810), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n9546), .CLK(n9810), .Q(
        WX3351) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n9546), .CLK(n9810), .Q(
        WX3353) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n9545), .CLK(n9811), .Q(
        WX3355) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n9544), .CLK(n9811), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n9544), .CLK(n9811), .Q(
        WX3359), .QN(n7625) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n9544), .CLK(n9811), .Q(
        WX3361), .QN(n7824) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n9543), .CLK(n9812), .Q(
        WX3363), .QN(n7823) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n9543), .CLK(n9812), .Q(
        WX3365), .QN(n7821) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n9543), .CLK(n9812), .Q(
        WX3367), .QN(n7819) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n9542), .CLK(n9812), .Q(
        test_so27), .QN(n8816) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n9562), .CLK(n9802), 
        .Q(WX3371), .QN(n7816) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n9562), .CLK(n9802), .Q(
        WX3373), .QN(n7814) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n9561), .CLK(n9803), .Q(
        WX3375), .QN(n7812) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n9561), .CLK(n9803), .Q(
        WX3377), .QN(n7810) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n9560), .CLK(n9803), .Q(
        WX3379), .QN(n7808) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n9560), .CLK(n9803), .Q(
        WX3381), .QN(n7806) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n9559), .CLK(n9804), .Q(
        WX3383), .QN(n7804) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n9558), .CLK(n9804), .Q(
        WX3385), .QN(n7802) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n9558), .CLK(n9804), .Q(
        WX3387), .QN(n7800) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n9557), .CLK(n9805), .Q(
        WX3389), .QN(n7798) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n9554), .CLK(n9806), .Q(
        WX3391), .QN(n8065) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n9554), .CLK(n9806), .Q(
        WX3393), .QN(n8063) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n9553), .CLK(n9807), .Q(
        WX3395), .QN(n8061) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n9552), .CLK(n9807), .Q(
        WX3397), .QN(n8059) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n9552), .CLK(n9807), .Q(
        WX3399), .QN(n8057) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n9551), .CLK(n9808), .Q(
        WX3401), .QN(n8055) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n9550), .CLK(n9808), .Q(
        WX3403), .QN(n8053) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n9550), .CLK(n9808), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n9549), .CLK(n9809), 
        .Q(WX3407), .QN(n8050) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n9548), .CLK(n9809), .Q(
        WX3409), .QN(n8048) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n9548), .CLK(n9809), .Q(
        WX3411), .QN(n8046) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n9547), .CLK(n9810), .Q(
        WX3413), .QN(n8044) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n9546), .CLK(n9810), .Q(
        WX3415), .QN(n8042) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n9546), .CLK(n9810), .Q(
        WX3417), .QN(n8040) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n9545), .CLK(n9811), .Q(
        WX3419), .QN(n8038) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n9544), .CLK(n9811), .Q(
        WX3421), .QN(n8036) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n9544), .CLK(n9811), .Q(
        WX3423), .QN(n8471) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n9543), .CLK(n9812), .Q(
        WX3425), .QN(n8472) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n9543), .CLK(n9812), .Q(
        WX3427), .QN(n8473) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n9543), .CLK(n9812), .Q(
        WX3429) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n9542), .CLK(n9812), .Q(
        WX3431), .QN(n8475) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n9542), .CLK(n9812), .Q(
        WX3433), .QN(n8476) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n9542), .CLK(n9812), .Q(
        WX3435), .QN(n8477) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n9542), .CLK(n9812), .Q(
        WX3437), .QN(n8478) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n9542), .CLK(n9812), .Q(
        test_so29), .QN(n8802) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n9561), .CLK(n9803), 
        .Q(WX3441), .QN(n8485) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n9560), .CLK(n9803), .Q(
        WX3443), .QN(n8486) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n9560), .CLK(n9803), .Q(
        WX3445), .QN(n8503) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n9559), .CLK(n9804), .Q(
        WX3447), .QN(n8504) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n9558), .CLK(n9804), .Q(
        WX3449), .QN(n8521) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n9557), .CLK(n9805), .Q(
        WX3451), .QN(n8522) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n9557), .CLK(n9805), .Q(
        WX3453), .QN(n8120) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n9554), .CLK(n9806), .Q(
        WX3455), .QN(n8529) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n9553), .CLK(n9807), .Q(
        WX3457), .QN(n8530) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n9553), .CLK(n9807), .Q(
        WX3459), .QN(n8531) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n9552), .CLK(n9807), .Q(
        WX3461), .QN(n8532) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n9551), .CLK(n9808), .Q(
        WX3463) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n9551), .CLK(n9808), .Q(
        WX3465), .QN(n8533) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n9550), .CLK(n9808), .Q(
        WX3467), .QN(n8534) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n9549), .CLK(n9809), .Q(
        WX3469), .QN(n8535) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n9549), .CLK(n9809), .Q(
        WX3471), .QN(n8536) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n9548), .CLK(n9809), .Q(
        test_so30), .QN(n8792) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n9547), .CLK(n9810), 
        .Q(WX3475), .QN(n8538) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n9547), .CLK(n9810), .Q(
        WX3477), .QN(n8122) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n9546), .CLK(n9810), .Q(
        WX3479), .QN(n8539) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n9545), .CLK(n9811), .Q(
        WX3481), .QN(n8556) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n9545), .CLK(n9811), .Q(
        WX3483), .QN(n8557) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n9544), .CLK(n9811), .Q(
        WX3485), .QN(n8132) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n9350), .CLK(n9908), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n9350), .CLK(n9908), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n9350), .CLK(n9908), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n9350), .CLK(n9908), 
        .Q(CRC_OUT_7_3) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n9350), .CLK(n9908), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n9350), .CLK(n9908), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n9349), .CLK(n9909), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n9349), .CLK(n9909), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n9349), .CLK(n9909), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n9349), .CLK(n9909), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n9349), .CLK(n9909), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n9349), .CLK(n9909), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_15) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n9348), .CLK(n9909), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n9347), .CLK(n9910), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n9346), .CLK(n9910), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n9346), .CLK(n9910), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n9541), .CLK(n9813), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n9541), .CLK(n9813), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n9541), .CLK(n9813), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n9541), .CLK(n9813), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n9541), .CLK(n9813), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n9541), .CLK(n9813), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n735), .SI(CRC_OUT_7_31), .SE(n9540), .CLK(n9813), 
        .Q(WX4364) );
  SDFFX1 DFF_577_Q_reg ( .D(n736), .SI(WX4364), .SE(n9535), .CLK(n9816), .Q(
        n8586), .QN(n8973) );
  SDFFX1 DFF_578_Q_reg ( .D(n737), .SI(n8586), .SE(n9535), .CLK(n9816), .Q(
        n8585), .QN(n8972) );
  SDFFX1 DFF_579_Q_reg ( .D(n738), .SI(n8585), .SE(n9536), .CLK(n9815), .Q(
        n8584), .QN(n8971) );
  SDFFX1 DFF_580_Q_reg ( .D(n739), .SI(n8584), .SE(n9536), .CLK(n9815), .Q(
        n8583), .QN(n8970) );
  SDFFX1 DFF_581_Q_reg ( .D(n740), .SI(n8583), .SE(n9536), .CLK(n9815), .Q(
        n8582), .QN(n8969) );
  SDFFX1 DFF_582_Q_reg ( .D(n741), .SI(n8582), .SE(n9536), .CLK(n9815), .Q(
        n8581), .QN(n8968) );
  SDFFX1 DFF_583_Q_reg ( .D(n742), .SI(n8581), .SE(n9536), .CLK(n9815), .Q(
        n8580), .QN(n8967) );
  SDFFX1 DFF_584_Q_reg ( .D(n743), .SI(n8580), .SE(n9536), .CLK(n9815), .Q(
        n8579), .QN(n8966) );
  SDFFX1 DFF_585_Q_reg ( .D(n744), .SI(n8579), .SE(n9537), .CLK(n9815), .Q(
        n8578), .QN(n8965) );
  SDFFX1 DFF_586_Q_reg ( .D(n745), .SI(n8578), .SE(n9537), .CLK(n9815), .Q(
        n8577), .QN(n8964) );
  SDFFX1 DFF_587_Q_reg ( .D(n746), .SI(n8577), .SE(n9537), .CLK(n9815), .Q(
        n8576), .QN(n8963) );
  SDFFX1 DFF_588_Q_reg ( .D(n747), .SI(n8576), .SE(n9537), .CLK(n9815), .Q(
        test_so33), .QN(n9070) );
  SDFFX1 DFF_589_Q_reg ( .D(n748), .SI(test_si34), .SE(n9537), .CLK(n9815), 
        .Q(n8573), .QN(n8962) );
  SDFFX1 DFF_590_Q_reg ( .D(n749), .SI(n8573), .SE(n9537), .CLK(n9815), .Q(
        n8572), .QN(n8961) );
  SDFFX1 DFF_591_Q_reg ( .D(n750), .SI(n8572), .SE(n9538), .CLK(n9814), .Q(
        n8571), .QN(n8960) );
  SDFFX1 DFF_592_Q_reg ( .D(n751), .SI(n8571), .SE(n9538), .CLK(n9814), .Q(
        n8570), .QN(n8959) );
  SDFFX1 DFF_593_Q_reg ( .D(n752), .SI(n8570), .SE(n9538), .CLK(n9814), .Q(
        n8569), .QN(n8958) );
  SDFFX1 DFF_594_Q_reg ( .D(n753), .SI(n8569), .SE(n9538), .CLK(n9814), .Q(
        n8568), .QN(n8957) );
  SDFFX1 DFF_595_Q_reg ( .D(n754), .SI(n8568), .SE(n9538), .CLK(n9814), .Q(
        n8567), .QN(n8956) );
  SDFFX1 DFF_596_Q_reg ( .D(n755), .SI(n8567), .SE(n9538), .CLK(n9814), .Q(
        n8566), .QN(n8955) );
  SDFFX1 DFF_597_Q_reg ( .D(n756), .SI(n8566), .SE(n9539), .CLK(n9814), .Q(
        n8565), .QN(n8954) );
  SDFFX1 DFF_598_Q_reg ( .D(n757), .SI(n8565), .SE(n9539), .CLK(n9814), .Q(
        n8564), .QN(n8953) );
  SDFFX1 DFF_599_Q_reg ( .D(n758), .SI(n8564), .SE(n9539), .CLK(n9814), .Q(
        n8563), .QN(n8952) );
  SDFFX1 DFF_600_Q_reg ( .D(n759), .SI(n8563), .SE(n9539), .CLK(n9814), .Q(
        n8562), .QN(n8951) );
  SDFFX1 DFF_601_Q_reg ( .D(n760), .SI(n8562), .SE(n9539), .CLK(n9814), .Q(
        n8561), .QN(n8950) );
  SDFFX1 DFF_602_Q_reg ( .D(n761), .SI(n8561), .SE(n9539), .CLK(n9814), .Q(
        n8560), .QN(n8949) );
  SDFFX1 DFF_603_Q_reg ( .D(n762), .SI(n8560), .SE(n9540), .CLK(n9813), .Q(
        n8559), .QN(n8948) );
  SDFFX1 DFF_604_Q_reg ( .D(n763), .SI(n8559), .SE(n9540), .CLK(n9813), .Q(
        n8558), .QN(n8947) );
  SDFFX1 DFF_605_Q_reg ( .D(n764), .SI(n8558), .SE(n9540), .CLK(n9813), .Q(
        test_so34), .QN(n9069) );
  SDFFX1 DFF_606_Q_reg ( .D(n765), .SI(test_si35), .SE(n9540), .CLK(n9813), 
        .Q(n8555), .QN(n8946) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n9540), .CLK(n9813), .Q(
        n8554), .QN(n8945) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n9535), .CLK(n9816), .Q(
        n8553), .QN(n16337) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n9535), .CLK(n9816), .Q(
        n8552), .QN(n16338) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n9534), .CLK(n9816), .Q(
        n8551), .QN(n16339) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n9534), .CLK(n9816), .Q(
        n8550), .QN(n16340) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n9533), .CLK(n9817), .Q(
        n8549), .QN(n16341) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n9532), .CLK(n9817), .Q(
        n8548), .QN(n16342) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n9532), .CLK(n9817), .Q(
        n8547), .QN(n16343) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n9531), .CLK(n9818), .Q(
        n8546), .QN(n16344) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n9531), .CLK(n9818), .Q(
        n8545), .QN(n16345) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n9530), .CLK(n9818), .Q(
        n8544), .QN(n16346) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n9529), .CLK(n9819), .Q(
        n8543), .QN(n16347) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n9528), .CLK(n9819), .Q(
        n8542), .QN(n16348) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n9528), .CLK(n9819), .Q(
        n8541), .QN(n16349) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n9351), .CLK(n9908), .Q(
        n8540), .QN(n16350) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n9556), .CLK(n9805), .Q(
        test_so35), .QN(n8823) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n9555), .CLK(n9806), 
        .Q(n8537), .QN(n16351) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n9555), .CLK(n9806), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n9526), .CLK(n9820), .Q(
        WX4558), .QN(n8031) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n9525), .CLK(n9821), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n9525), .CLK(n9821), .Q(
        WX4562), .QN(n8028) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n9524), .CLK(n9821), .Q(
        WX4564), .QN(n8026) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n9523), .CLK(n9822), .Q(
        WX4566), .QN(n8024) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n9523), .CLK(n9822), .Q(
        WX4568), .QN(n8022) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n9522), .CLK(n9822), .Q(
        WX4570), .QN(n8020) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n9521), .CLK(n9823), .Q(
        WX4572), .QN(n8018) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n9521), .CLK(n9823), .Q(
        WX4574), .QN(n8016) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n9520), .CLK(n9823), .Q(
        WX4576), .QN(n8014) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n9519), .CLK(n9824), .Q(
        WX4578), .QN(n8012) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n9519), .CLK(n9824), .Q(
        WX4580), .QN(n8010) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n9518), .CLK(n9824), .Q(
        WX4582), .QN(n8008) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n9517), .CLK(n9825), .Q(
        WX4584), .QN(n8006) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n9517), .CLK(n9825), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n9535), .CLK(n9816), 
        .Q(WX4588), .QN(n7622) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n9535), .CLK(n9816), .Q(
        WX4590), .QN(n7796) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n9534), .CLK(n9816), .Q(
        WX4592), .QN(n7794) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n9534), .CLK(n9816), .Q(
        WX4594), .QN(n7792) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n9533), .CLK(n9817), .Q(
        WX4596), .QN(n7790) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n9533), .CLK(n9817), .Q(
        WX4598), .QN(n7788) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n9532), .CLK(n9817), .Q(
        WX4600), .QN(n7786) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n9531), .CLK(n9818), .Q(
        WX4602), .QN(n7784) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n9531), .CLK(n9818), .Q(
        WX4604), .QN(n7782) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n9530), .CLK(n9818), .Q(
        WX4606), .QN(n7780) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n9529), .CLK(n9819), .Q(
        WX4608), .QN(n7778) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n9529), .CLK(n9819), .Q(
        WX4610), .QN(n7776) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n9528), .CLK(n9819), .Q(
        WX4612), .QN(n7774) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n9527), .CLK(n9820), .Q(
        WX4614), .QN(n7772) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n9555), .CLK(n9806), .Q(
        WX4616), .QN(n7770) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n9555), .CLK(n9806), .Q(
        WX4618), .QN(n7768) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n9555), .CLK(n9806), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n9525), .CLK(n9821), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n9525), .CLK(n9821), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n9524), .CLK(n9821), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n9524), .CLK(n9821), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n9523), .CLK(n9822), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n9522), .CLK(n9822), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n9522), .CLK(n9822), .Q(
        WX4634) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n9521), .CLK(n9823), .Q(
        WX4636) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n9520), .CLK(n9823), .Q(
        WX4638) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n9520), .CLK(n9823), .Q(
        WX4640) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n9519), .CLK(n9824), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n9518), .CLK(n9824), .Q(
        WX4644) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n9518), .CLK(n9824), .Q(
        WX4646) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n9517), .CLK(n9825), .Q(
        WX4648) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n9516), .CLK(n9825), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n9516), .CLK(n9825), .Q(
        WX4652), .QN(n7623) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n9516), .CLK(n9825), .Q(
        test_so38), .QN(n8814) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n9534), .CLK(n9816), 
        .Q(WX4656), .QN(n7795) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n9534), .CLK(n9816), .Q(
        WX4658), .QN(n7793) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n9533), .CLK(n9817), .Q(
        WX4660), .QN(n7791) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n9533), .CLK(n9817), .Q(
        WX4662), .QN(n7789) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n9532), .CLK(n9817), .Q(
        WX4664), .QN(n7787) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n9531), .CLK(n9818), .Q(
        WX4666), .QN(n7785) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n9530), .CLK(n9818), .Q(
        WX4668), .QN(n7783) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n9530), .CLK(n9818), .Q(
        WX4670), .QN(n7781) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n9529), .CLK(n9819), .Q(
        WX4672), .QN(n7779) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n9529), .CLK(n9819), .Q(
        WX4674), .QN(n7777) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n9528), .CLK(n9819), .Q(
        WX4676), .QN(n7775) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n9527), .CLK(n9820), .Q(
        WX4678), .QN(n7773) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n9527), .CLK(n9820), .Q(
        WX4680), .QN(n7771) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n9527), .CLK(n9820), .Q(
        WX4682), .QN(n7769) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n9526), .CLK(n9820), .Q(
        WX4684), .QN(n8034) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n9526), .CLK(n9820), .Q(
        WX4686), .QN(n8032) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n9525), .CLK(n9821), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n9524), .CLK(n9821), 
        .Q(WX4690), .QN(n8029) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n9524), .CLK(n9821), .Q(
        WX4692), .QN(n8027) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n9523), .CLK(n9822), .Q(
        WX4694), .QN(n8025) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n9522), .CLK(n9822), .Q(
        WX4696), .QN(n8023) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n9522), .CLK(n9822), .Q(
        WX4698), .QN(n8021) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n9521), .CLK(n9823), .Q(
        WX4700), .QN(n8019) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n9520), .CLK(n9823), .Q(
        WX4702), .QN(n8017) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n9520), .CLK(n9823), .Q(
        WX4704), .QN(n8015) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n9519), .CLK(n9824), .Q(
        WX4706), .QN(n8013) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n9518), .CLK(n9824), .Q(
        WX4708), .QN(n8011) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n9518), .CLK(n9824), .Q(
        WX4710), .QN(n8009) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n9517), .CLK(n9825), .Q(
        WX4712), .QN(n8007) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n9516), .CLK(n9825), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n9516), .CLK(n9825), .Q(
        WX4716), .QN(n8355) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n9515), .CLK(n9826), .Q(
        WX4718), .QN(n8356) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n9515), .CLK(n9826), .Q(
        WX4720), .QN(n8357) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n9515), .CLK(n9826), .Q(
        test_so40), .QN(n8801) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n9533), .CLK(n9817), 
        .Q(WX4724), .QN(n8358) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n9532), .CLK(n9817), .Q(
        WX4726), .QN(n8359) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n9532), .CLK(n9817), .Q(
        WX4728), .QN(n8360) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n9531), .CLK(n9818), .Q(
        WX4730), .QN(n8361) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n9530), .CLK(n9818), .Q(
        WX4732) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n9530), .CLK(n9818), .Q(
        WX4734), .QN(n8379) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n9529), .CLK(n9819), .Q(
        WX4736), .QN(n8380) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n9528), .CLK(n9819), .Q(
        WX4738), .QN(n8397) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n9528), .CLK(n9819), .Q(
        WX4740), .QN(n8398) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n9527), .CLK(n9820), .Q(
        WX4742), .QN(n8412) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n9527), .CLK(n9820), .Q(
        WX4744), .QN(n8413) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n9526), .CLK(n9820), .Q(
        WX4746), .QN(n8118) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n9526), .CLK(n9820), .Q(
        WX4748), .QN(n8414) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n9526), .CLK(n9820), .Q(
        WX4750), .QN(n8415) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n9525), .CLK(n9821), .Q(
        WX4752), .QN(n8416) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n9524), .CLK(n9821), .Q(
        WX4754), .QN(n8417) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n9523), .CLK(n9822), .Q(
        test_so41), .QN(n8797) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n9523), .CLK(n9822), 
        .Q(WX4758), .QN(n8418) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n9522), .CLK(n9822), .Q(
        WX4760), .QN(n8419) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n9521), .CLK(n9823), .Q(
        WX4762), .QN(n8420) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n9521), .CLK(n9823), .Q(
        WX4764), .QN(n8432) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n9520), .CLK(n9823), .Q(
        WX4766) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n9519), .CLK(n9824), .Q(
        WX4768), .QN(n8450) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n9519), .CLK(n9824), .Q(
        WX4770), .QN(n8119) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n9518), .CLK(n9824), .Q(
        WX4772), .QN(n8451) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n9517), .CLK(n9825), .Q(
        WX4774), .QN(n8468) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n9517), .CLK(n9825), .Q(
        WX4776), .QN(n8469) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n9516), .CLK(n9825), .Q(
        WX4778), .QN(n8131) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n9356), .CLK(n9905), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n9355), .CLK(n9906), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n9355), .CLK(n9906), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n9355), .CLK(n9906), 
        .Q(CRC_OUT_6_3) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n9355), .CLK(n9906), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n9355), .CLK(n9906), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n9355), .CLK(n9906), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n9354), .CLK(n9906), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n9354), .CLK(n9906), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n9354), .CLK(n9906), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n9354), .CLK(n9906), 
        .Q(CRC_OUT_6_10) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n9354), .CLK(n9906), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n9354), .CLK(n9906), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_15) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n9353), .CLK(n9907), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n9352), .CLK(n9907), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n9352), .CLK(n9907), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n9352), .CLK(n9907), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n9352), .CLK(n9907), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n9352), .CLK(n9907), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n9352), .CLK(n9907), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n9351), .CLK(n9908), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n9351), .CLK(n9908), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n9351), .CLK(n9908), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n9351), .CLK(n9908), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n9351), .CLK(n9908), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n9515), .CLK(n9826), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n9515), .CLK(n9826), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n976), .SI(CRC_OUT_6_31), .SE(n9515), .CLK(n9826), 
        .Q(WX5657) );
  SDFFX1 DFF_769_Q_reg ( .D(n977), .SI(WX5657), .SE(n9509), .CLK(n9829), .Q(
        n8528), .QN(n8944) );
  SDFFX1 DFF_770_Q_reg ( .D(n978), .SI(n8528), .SE(n9510), .CLK(n9828), .Q(
        n8527), .QN(n8943) );
  SDFFX1 DFF_771_Q_reg ( .D(n979), .SI(n8527), .SE(n9510), .CLK(n9828), .Q(
        n8526), .QN(n8942) );
  SDFFX1 DFF_772_Q_reg ( .D(n980), .SI(n8526), .SE(n9510), .CLK(n9828), .Q(
        n8525), .QN(n8941) );
  SDFFX1 DFF_773_Q_reg ( .D(n981), .SI(n8525), .SE(n9510), .CLK(n9828), .Q(
        n8524), .QN(n8940) );
  SDFFX1 DFF_774_Q_reg ( .D(n982), .SI(n8524), .SE(n9510), .CLK(n9828), .Q(
        n8523), .QN(n8939) );
  SDFFX1 DFF_775_Q_reg ( .D(n983), .SI(n8523), .SE(n9510), .CLK(n9828), .Q(
        test_so44), .QN(n9068) );
  SDFFX1 DFF_776_Q_reg ( .D(n984), .SI(test_si45), .SE(n9511), .CLK(n9828), 
        .Q(n8520), .QN(n8938) );
  SDFFX1 DFF_777_Q_reg ( .D(n985), .SI(n8520), .SE(n9511), .CLK(n9828), .Q(
        n8519), .QN(n8937) );
  SDFFX1 DFF_778_Q_reg ( .D(n986), .SI(n8519), .SE(n9511), .CLK(n9828), .Q(
        n8518), .QN(n8936) );
  SDFFX1 DFF_779_Q_reg ( .D(n987), .SI(n8518), .SE(n9511), .CLK(n9828), .Q(
        n8517), .QN(n8935) );
  SDFFX1 DFF_780_Q_reg ( .D(n988), .SI(n8517), .SE(n9511), .CLK(n9828), .Q(
        n8516), .QN(n8934) );
  SDFFX1 DFF_781_Q_reg ( .D(n989), .SI(n8516), .SE(n9511), .CLK(n9828), .Q(
        n8515), .QN(n8933) );
  SDFFX1 DFF_782_Q_reg ( .D(n990), .SI(n8515), .SE(n9512), .CLK(n9827), .Q(
        n8514), .QN(n8932) );
  SDFFX1 DFF_783_Q_reg ( .D(n991), .SI(n8514), .SE(n9512), .CLK(n9827), .Q(
        n8513), .QN(n8931) );
  SDFFX1 DFF_784_Q_reg ( .D(n992), .SI(n8513), .SE(n9512), .CLK(n9827), .Q(
        n8512), .QN(n8930) );
  SDFFX1 DFF_785_Q_reg ( .D(n993), .SI(n8512), .SE(n9512), .CLK(n9827), .Q(
        n8511), .QN(n8929) );
  SDFFX1 DFF_786_Q_reg ( .D(n994), .SI(n8511), .SE(n9512), .CLK(n9827), .Q(
        n8510), .QN(n8928) );
  SDFFX1 DFF_787_Q_reg ( .D(n995), .SI(n8510), .SE(n9512), .CLK(n9827), .Q(
        n8509), .QN(n8927) );
  SDFFX1 DFF_788_Q_reg ( .D(n996), .SI(n8509), .SE(n9513), .CLK(n9827), .Q(
        n8508), .QN(n8926) );
  SDFFX1 DFF_789_Q_reg ( .D(n997), .SI(n8508), .SE(n9513), .CLK(n9827), .Q(
        n8507), .QN(n8925) );
  SDFFX1 DFF_790_Q_reg ( .D(n998), .SI(n8507), .SE(n9513), .CLK(n9827), .Q(
        n8506), .QN(n8924) );
  SDFFX1 DFF_791_Q_reg ( .D(n999), .SI(n8506), .SE(n9513), .CLK(n9827), .Q(
        n8505), .QN(n8923) );
  SDFFX1 DFF_792_Q_reg ( .D(n1000), .SI(n8505), .SE(n9513), .CLK(n9827), .Q(
        test_so45), .QN(n9067) );
  SDFFX1 DFF_793_Q_reg ( .D(n1001), .SI(test_si46), .SE(n9513), .CLK(n9827), 
        .Q(n8502), .QN(n8922) );
  SDFFX1 DFF_794_Q_reg ( .D(n1002), .SI(n8502), .SE(n9514), .CLK(n9826), .Q(
        n8501), .QN(n8921) );
  SDFFX1 DFF_795_Q_reg ( .D(n1003), .SI(n8501), .SE(n9514), .CLK(n9826), .Q(
        n8500), .QN(n8920) );
  SDFFX1 DFF_796_Q_reg ( .D(n1004), .SI(n8500), .SE(n9514), .CLK(n9826), .Q(
        n8499), .QN(n8919) );
  SDFFX1 DFF_797_Q_reg ( .D(n1005), .SI(n8499), .SE(n9514), .CLK(n9826), .Q(
        n8498), .QN(n8918) );
  SDFFX1 DFF_798_Q_reg ( .D(n1006), .SI(n8498), .SE(n9514), .CLK(n9826), .Q(
        n8497), .QN(n8917) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n9514), .CLK(n9826), .Q(
        n8496), .QN(n8916) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n9509), .CLK(n9829), .Q(
        n8495), .QN(n16352) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n9509), .CLK(n9829), .Q(
        n8494), .QN(n16353) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n9509), .CLK(n9829), .Q(
        n8493), .QN(n16354) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n9508), .CLK(n9829), .Q(
        n8492), .QN(n16355) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n9508), .CLK(n9829), .Q(
        n8491), .QN(n16356) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n9507), .CLK(n9830), .Q(
        n8490), .QN(n16357) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n9507), .CLK(n9830), .Q(
        n8489), .QN(n16358) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n9507), .CLK(n9830), .Q(
        n8488), .QN(n16359) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n9507), .CLK(n9830), .Q(
        n8487), .QN(n16360) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n9356), .CLK(n9905), .Q(
        test_so46), .QN(n8822) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n9506), .CLK(n9830), 
        .Q(n8484), .QN(n16361) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n9506), .CLK(n9830), .Q(
        n8483), .QN(n16362) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n9505), .CLK(n9831), .Q(
        n8482), .QN(n16363) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n9356), .CLK(n9905), .Q(
        n8481), .QN(n16364) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n9556), .CLK(n9805), .Q(
        n8480), .QN(n16365) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n9504), .CLK(n9831), .Q(
        n8479), .QN(n16366) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n9504), .CLK(n9831), .Q(
        WX5849), .QN(n8003) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n9503), .CLK(n9832), .Q(
        WX5851), .QN(n8001) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n9502), .CLK(n9832), .Q(
        WX5853), .QN(n7999) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n9502), .CLK(n9832), .Q(
        WX5855), .QN(n7997) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n9501), .CLK(n9833), .Q(
        WX5857), .QN(n7995) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n9500), .CLK(n9833), .Q(
        WX5859), .QN(n7993) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n9500), .CLK(n9833), .Q(
        WX5861), .QN(n7991) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n9499), .CLK(n9834), .Q(
        WX5863), .QN(n7989) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n9498), .CLK(n9834), .Q(
        WX5865), .QN(n7987) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n9498), .CLK(n9834), .Q(
        WX5867), .QN(n7985) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n9497), .CLK(n9835), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n9496), .CLK(n9835), 
        .Q(WX5871), .QN(n7982) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n9496), .CLK(n9835), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n9495), .CLK(n9836), .Q(
        WX5875), .QN(n7978) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n9494), .CLK(n9836), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n9494), .CLK(n9836), .Q(
        WX5879), .QN(n7975) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n9509), .CLK(n9829), .Q(
        WX5881), .QN(n7620) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n9509), .CLK(n9829), .Q(
        WX5883), .QN(n7766) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n9508), .CLK(n9829), .Q(
        WX5885), .QN(n7764) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n9508), .CLK(n9829), .Q(
        WX5887), .QN(n7762) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n9508), .CLK(n9829), .Q(
        WX5889), .QN(n7760) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n9508), .CLK(n9829), .Q(
        WX5891), .QN(n7758) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n9507), .CLK(n9830), .Q(
        WX5893), .QN(n7756) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n9507), .CLK(n9830), .Q(
        WX5895), .QN(n7754) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n9506), .CLK(n9830), .Q(
        WX5897), .QN(n7752) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n9506), .CLK(n9830), .Q(
        WX5899), .QN(n7750) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n9506), .CLK(n9830), .Q(
        WX5901), .QN(n7748) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n9506), .CLK(n9830), .Q(
        test_so48), .QN(n8813) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n9505), .CLK(n9831), 
        .Q(WX5905), .QN(n7745) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n9505), .CLK(n9831), .Q(
        WX5907), .QN(n7744) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n9504), .CLK(n9831), .Q(
        WX5909), .QN(n7742) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n9504), .CLK(n9831), .Q(
        WX5911), .QN(n7740) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n9503), .CLK(n9832), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n9503), .CLK(n9832), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n9502), .CLK(n9832), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n9501), .CLK(n9833), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n9501), .CLK(n9833), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n9500), .CLK(n9833), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n9499), .CLK(n9834), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n9499), .CLK(n9834), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n9498), .CLK(n9834), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n9497), .CLK(n9835), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n9497), .CLK(n9835), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n9496), .CLK(n9835), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n9495), .CLK(n9836), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n9495), .CLK(n9836), 
        .Q(WX5939) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n9494), .CLK(n9836), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n9493), .CLK(n9837), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n9493), .CLK(n9837), .Q(
        WX5945), .QN(n7621) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n9493), .CLK(n9837), .Q(
        WX5947), .QN(n7767) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n9492), .CLK(n9837), .Q(
        WX5949), .QN(n7765) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n9492), .CLK(n9837), .Q(
        WX5951), .QN(n7763) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n9492), .CLK(n9837), .Q(
        WX5953), .QN(n7761) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n9491), .CLK(n9838), .Q(
        WX5955), .QN(n7759) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n9491), .CLK(n9838), .Q(
        WX5957), .QN(n7757) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n9491), .CLK(n9838), .Q(
        WX5959), .QN(n7755) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n9490), .CLK(n9838), .Q(
        WX5961), .QN(n7753) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n9490), .CLK(n9838), .Q(
        WX5963), .QN(n7751) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n9490), .CLK(n9838), .Q(
        WX5965), .QN(n7749) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n9505), .CLK(n9831), .Q(
        WX5967), .QN(n7747) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n9505), .CLK(n9831), .Q(
        WX5969), .QN(n7746) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n9505), .CLK(n9831), .Q(
        test_so50), .QN(n8812) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n9504), .CLK(n9831), 
        .Q(WX5973), .QN(n7743) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n9504), .CLK(n9831), .Q(
        WX5975), .QN(n7741) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n9503), .CLK(n9832), .Q(
        WX5977), .QN(n8004) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n9503), .CLK(n9832), .Q(
        WX5979), .QN(n8002) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n9502), .CLK(n9832), .Q(
        WX5981), .QN(n8000) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n9501), .CLK(n9833), .Q(
        WX5983), .QN(n7998) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n9501), .CLK(n9833), .Q(
        WX5985), .QN(n7996) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n9500), .CLK(n9833), .Q(
        WX5987), .QN(n7994) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n9499), .CLK(n9834), .Q(
        WX5989), .QN(n7992) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n9499), .CLK(n9834), .Q(
        WX5991), .QN(n7990) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n9498), .CLK(n9834), .Q(
        WX5993), .QN(n7988) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n9497), .CLK(n9835), .Q(
        WX5995), .QN(n7986) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n9497), .CLK(n9835), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n9496), .CLK(n9835), .Q(
        WX5999), .QN(n7983) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n9495), .CLK(n9836), .Q(
        WX6001), .QN(n7981) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n9495), .CLK(n9836), .Q(
        WX6003), .QN(n7979) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n9494), .CLK(n9836), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n9493), .CLK(n9837), 
        .Q(WX6007), .QN(n7976) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n9493), .CLK(n9837), .Q(
        WX6009), .QN(n8239) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n9492), .CLK(n9837), .Q(
        WX6011), .QN(n8240) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n9492), .CLK(n9837), .Q(
        WX6013), .QN(n8241) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n9492), .CLK(n9837), .Q(
        WX6015), .QN(n8242) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n9491), .CLK(n9838), .Q(
        WX6017), .QN(n8243) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n9491), .CLK(n9838), .Q(
        WX6019), .QN(n8244) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n9491), .CLK(n9838), .Q(
        WX6021), .QN(n8245) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n9490), .CLK(n9838), .Q(
        WX6023), .QN(n8255) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n9490), .CLK(n9838), .Q(
        WX6025), .QN(n8256) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n9490), .CLK(n9838), .Q(
        WX6027), .QN(n8273) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n9489), .CLK(n9839), .Q(
        WX6029), .QN(n8274) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n9489), .CLK(n9839), .Q(
        WX6031), .QN(n8291) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n9489), .CLK(n9839), .Q(
        WX6033), .QN(n8292) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n9489), .CLK(n9839), .Q(
        WX6035), .QN(n8296) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n9489), .CLK(n9839), .Q(
        WX6037), .QN(n8297) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n9489), .CLK(n9839), .Q(
        test_so52), .QN(n8827) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n9503), .CLK(n9832), 
        .Q(WX6041), .QN(n8298) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n9502), .CLK(n9832), .Q(
        WX6043), .QN(n8299) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n9502), .CLK(n9832), .Q(
        WX6045), .QN(n8300) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n9501), .CLK(n9833), .Q(
        WX6047), .QN(n8301) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n9500), .CLK(n9833), .Q(
        WX6049), .QN(n8116) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n9500), .CLK(n9833), .Q(
        WX6051), .QN(n8302) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n9499), .CLK(n9834), .Q(
        WX6053), .QN(n8303) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n9498), .CLK(n9834), .Q(
        WX6055), .QN(n8308) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n9498), .CLK(n9834), .Q(
        WX6057), .QN(n8309) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n9497), .CLK(n9835), .Q(
        WX6059), .QN(n8326) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n9496), .CLK(n9835), .Q(
        WX6061), .QN(n8327) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n9496), .CLK(n9835), .Q(
        WX6063), .QN(n8117) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n9495), .CLK(n9836), .Q(
        WX6065), .QN(n8344) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n9494), .CLK(n9836), .Q(
        WX6067), .QN(n8345) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n9494), .CLK(n9836), .Q(
        WX6069), .QN(n8354) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n9493), .CLK(n9837), .Q(
        WX6071), .QN(n8130) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n9359), .CLK(n9904), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n9359), .CLK(n9904), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n9359), .CLK(n9904), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n9359), .CLK(n9904), 
        .Q(CRC_OUT_5_3) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n9359), .CLK(n9904), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n9359), .CLK(n9904), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n9358), .CLK(n9904), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n9358), .CLK(n9904), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n9358), .CLK(n9904), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n9358), .CLK(n9904), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n9358), .CLK(n9904), 
        .Q(CRC_OUT_5_10) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n9358), .CLK(n9904), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n9357), .CLK(n9905), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n9357), .CLK(n9905), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n9357), .CLK(n9905), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n9357), .CLK(n9905), .Q(CRC_OUT_5_15) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n9357), .CLK(n9905), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n9357), .CLK(n9905), .Q(test_so54), .QN(n8828) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n9356), .CLK(n9905), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n9356), .CLK(n9905), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n9356), .CLK(n9905), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n9488), .CLK(n9839), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n9487), .CLK(n9840), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n9487), .CLK(n9840), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n9487), .CLK(n9840), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n9487), .CLK(n9840), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n9487), .CLK(n9840), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n1217), .SI(CRC_OUT_5_31), .SE(n9487), .CLK(n9840), 
        .Q(WX6950) );
  SDFFX1 DFF_961_Q_reg ( .D(n1218), .SI(WX6950), .SE(n9481), .CLK(n9843), .Q(
        n8470), .QN(n8915) );
  SDFFX1 DFF_962_Q_reg ( .D(n1219), .SI(n8470), .SE(n9482), .CLK(n9842), .Q(
        test_so55), .QN(n9066) );
  SDFFX1 DFF_963_Q_reg ( .D(n1220), .SI(test_si56), .SE(n9482), .CLK(n9842), 
        .Q(n8467), .QN(n8914) );
  SDFFX1 DFF_964_Q_reg ( .D(n1221), .SI(n8467), .SE(n9482), .CLK(n9842), .Q(
        n8466), .QN(n8913) );
  SDFFX1 DFF_965_Q_reg ( .D(n1222), .SI(n8466), .SE(n9482), .CLK(n9842), .Q(
        n8465), .QN(n8912) );
  SDFFX1 DFF_966_Q_reg ( .D(n1223), .SI(n8465), .SE(n9482), .CLK(n9842), .Q(
        n8464), .QN(n8911) );
  SDFFX1 DFF_967_Q_reg ( .D(n1224), .SI(n8464), .SE(n9482), .CLK(n9842), .Q(
        n8463), .QN(n8910) );
  SDFFX1 DFF_968_Q_reg ( .D(n1225), .SI(n8463), .SE(n9483), .CLK(n9842), .Q(
        n8462), .QN(n8909) );
  SDFFX1 DFF_969_Q_reg ( .D(n1226), .SI(n8462), .SE(n9483), .CLK(n9842), .Q(
        n8461), .QN(n8908) );
  SDFFX1 DFF_970_Q_reg ( .D(n1227), .SI(n8461), .SE(n9483), .CLK(n9842), .Q(
        n8460), .QN(n8907) );
  SDFFX1 DFF_971_Q_reg ( .D(n1228), .SI(n8460), .SE(n9483), .CLK(n9842), .Q(
        n8459), .QN(n8906) );
  SDFFX1 DFF_972_Q_reg ( .D(n1229), .SI(n8459), .SE(n9483), .CLK(n9842), .Q(
        n8458), .QN(n8905) );
  SDFFX1 DFF_973_Q_reg ( .D(n1230), .SI(n8458), .SE(n9483), .CLK(n9842), .Q(
        n8457), .QN(n8904) );
  SDFFX1 DFF_974_Q_reg ( .D(n1231), .SI(n8457), .SE(n9484), .CLK(n9841), .Q(
        n8456), .QN(n8903) );
  SDFFX1 DFF_975_Q_reg ( .D(n1232), .SI(n8456), .SE(n9484), .CLK(n9841), .Q(
        n8455), .QN(n8902) );
  SDFFX1 DFF_976_Q_reg ( .D(n1233), .SI(n8455), .SE(n9484), .CLK(n9841), .Q(
        n8454), .QN(n8901) );
  SDFFX1 DFF_977_Q_reg ( .D(n1234), .SI(n8454), .SE(n9484), .CLK(n9841), .Q(
        n8453), .QN(n8900) );
  SDFFX1 DFF_978_Q_reg ( .D(n1235), .SI(n8453), .SE(n9484), .CLK(n9841), .Q(
        n8452), .QN(n8899) );
  SDFFX1 DFF_979_Q_reg ( .D(n1236), .SI(n8452), .SE(n9484), .CLK(n9841), .Q(
        test_so56), .QN(n9065) );
  SDFFX1 DFF_980_Q_reg ( .D(n1237), .SI(test_si57), .SE(n9485), .CLK(n9841), 
        .Q(n8449), .QN(n8898) );
  SDFFX1 DFF_981_Q_reg ( .D(n1238), .SI(n8449), .SE(n9485), .CLK(n9841), .Q(
        n8448), .QN(n8897) );
  SDFFX1 DFF_982_Q_reg ( .D(n1239), .SI(n8448), .SE(n9485), .CLK(n9841), .Q(
        n8447), .QN(n8896) );
  SDFFX1 DFF_983_Q_reg ( .D(n1240), .SI(n8447), .SE(n9485), .CLK(n9841), .Q(
        n8446), .QN(n8895) );
  SDFFX1 DFF_984_Q_reg ( .D(n1241), .SI(n8446), .SE(n9485), .CLK(n9841), .Q(
        n8445), .QN(n8894) );
  SDFFX1 DFF_985_Q_reg ( .D(n508), .SI(n8445), .SE(n9485), .CLK(n9841), .Q(
        n8444), .QN(n8893) );
  SDFFX1 DFF_986_Q_reg ( .D(n1242), .SI(n8444), .SE(n9486), .CLK(n9840), .Q(
        n8443), .QN(n8892) );
  SDFFX1 DFF_987_Q_reg ( .D(n1243), .SI(n8443), .SE(n9486), .CLK(n9840), .Q(
        n8442), .QN(n8891) );
  SDFFX1 DFF_988_Q_reg ( .D(n1244), .SI(n8442), .SE(n9486), .CLK(n9840), .Q(
        n8441), .QN(n8890) );
  SDFFX1 DFF_989_Q_reg ( .D(n1245), .SI(n8441), .SE(n9486), .CLK(n9840), .Q(
        n8440), .QN(n8889) );
  SDFFX1 DFF_990_Q_reg ( .D(n1246), .SI(n8440), .SE(n9486), .CLK(n9840), .Q(
        n8439), .QN(n8888) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n9486), .CLK(n9840), .Q(
        n8438), .QN(n8887) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n9481), .CLK(n9843), .Q(
        n8437), .QN(n16367) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n9481), .CLK(n9843), .Q(
        n8436), .QN(n16368) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n9481), .CLK(n9843), .Q(
        n8435), .QN(n16369) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n9480), .CLK(n9843), .Q(
        n8434), .QN(n16370) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n9480), .CLK(n9843), .Q(
        test_so57), .QN(n8821) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n9479), .CLK(n9844), 
        .Q(n8431), .QN(n16371) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n9479), .CLK(n9844), .Q(
        n8430), .QN(n16372) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n9479), .CLK(n9844), .Q(
        n8429), .QN(n16373) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n9478), .CLK(n9844), .Q(
        n8428), .QN(n16374) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n9478), .CLK(n9844), .Q(
        n8427), .QN(n16375) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n9477), .CLK(n9845), .Q(
        n8426), .QN(n16376) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n9477), .CLK(n9845), .Q(
        n8425), .QN(n16377) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n9476), .CLK(n9845), .Q(
        n8424), .QN(n16378) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n9475), .CLK(n9846), .Q(
        n8423), .QN(n16379) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n9556), .CLK(n9805), .Q(
        n8422), .QN(n16380) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n9474), .CLK(n9846), .Q(
        n8421), .QN(n16381) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n9474), .CLK(n9846), .Q(
        WX7142), .QN(n7973) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n9473), .CLK(n9847), 
        .Q(WX7144), .QN(n7971) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n9472), .CLK(n9847), 
        .Q(WX7146), .QN(n7969) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n9472), .CLK(n9847), 
        .Q(WX7148), .QN(n7967) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n9471), .CLK(n9848), 
        .Q(WX7150), .QN(n7965) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n9470), .CLK(n9848), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n9469), .CLK(n9849), 
        .Q(WX7154), .QN(n7962) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n9469), .CLK(n9849), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n9468), .CLK(n9849), 
        .Q(WX7158), .QN(n7958) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n9468), .CLK(n9849), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n9467), .CLK(n9850), 
        .Q(WX7162), .QN(n7955) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n9466), .CLK(n9850), 
        .Q(WX7164), .QN(n7953) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n9466), .CLK(n9850), 
        .Q(WX7166), .QN(n7951) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n9465), .CLK(n9851), 
        .Q(WX7168), .QN(n7949) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n9464), .CLK(n9851), 
        .Q(WX7170), .QN(n7947) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n9464), .CLK(n9851), 
        .Q(WX7172), .QN(n7945) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n9481), .CLK(n9843), 
        .Q(WX7174), .QN(n7618) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n9481), .CLK(n9843), 
        .Q(WX7176), .QN(n7738) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n9480), .CLK(n9843), 
        .Q(WX7178), .QN(n7736) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n9480), .CLK(n9843), 
        .Q(WX7180), .QN(n7734) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n9480), .CLK(n9843), 
        .Q(WX7182), .QN(n7732) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n9480), .CLK(n9843), 
        .Q(WX7184), .QN(n7730) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n9479), .CLK(n9844), 
        .Q(test_so59), .QN(n8811) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n9478), .CLK(n9844), 
        .Q(WX7188), .QN(n7727) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n9478), .CLK(n9844), 
        .Q(WX7190), .QN(n7726) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n9478), .CLK(n9844), 
        .Q(WX7192), .QN(n7724) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n9477), .CLK(n9845), 
        .Q(WX7194), .QN(n7722) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n9477), .CLK(n9845), 
        .Q(WX7196), .QN(n7720) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n9476), .CLK(n9845), 
        .Q(WX7198), .QN(n7718) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n9475), .CLK(n9846), 
        .Q(WX7200), .QN(n7716) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n9475), .CLK(n9846), 
        .Q(WX7202), .QN(n7714) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n9474), .CLK(n9846), 
        .Q(WX7204), .QN(n7712) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n9473), .CLK(n9847), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n9473), .CLK(n9847), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n9472), .CLK(n9847), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n9471), .CLK(n9848), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n9471), .CLK(n9848), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n9470), .CLK(n9848), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n9470), .CLK(n9848), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n9469), .CLK(n9849), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n9468), .CLK(n9849), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n9467), .CLK(n9850), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n9467), .CLK(n9850), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n9466), .CLK(n9850), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n9465), .CLK(n9851), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n9465), .CLK(n9851), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n9464), .CLK(n9851), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n9463), .CLK(n9852), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n9463), .CLK(n9852), 
        .Q(WX7238), .QN(n7619) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n9463), .CLK(n9852), 
        .Q(WX7240), .QN(n7739) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n9462), .CLK(n9852), 
        .Q(WX7242), .QN(n7737) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n9462), .CLK(n9852), 
        .Q(WX7244), .QN(n7735) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n9462), .CLK(n9852), 
        .Q(WX7246), .QN(n7733) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n9461), .CLK(n9853), 
        .Q(WX7248), .QN(n7731) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n9479), .CLK(n9844), 
        .Q(WX7250), .QN(n7729) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n9479), .CLK(n9844), 
        .Q(WX7252), .QN(n7728) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n9478), .CLK(n9844), 
        .Q(test_so61), .QN(n8810) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n9477), .CLK(n9845), 
        .Q(WX7256), .QN(n7725) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n9477), .CLK(n9845), 
        .Q(WX7258), .QN(n7723) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n9476), .CLK(n9845), 
        .Q(WX7260), .QN(n7721) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n9476), .CLK(n9845), 
        .Q(WX7262), .QN(n7719) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n9475), .CLK(n9846), 
        .Q(WX7264), .QN(n7717) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n9475), .CLK(n9846), 
        .Q(WX7266), .QN(n7715) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n9474), .CLK(n9846), 
        .Q(WX7268), .QN(n7713) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n9473), .CLK(n9847), 
        .Q(WX7270), .QN(n7974) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n9473), .CLK(n9847), 
        .Q(WX7272), .QN(n7972) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n9472), .CLK(n9847), 
        .Q(WX7274), .QN(n7970) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n9471), .CLK(n9848), 
        .Q(WX7276), .QN(n7968) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n9471), .CLK(n9848), 
        .Q(WX7278), .QN(n7966) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n9470), .CLK(n9848), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n9469), .CLK(n9849), 
        .Q(WX7282), .QN(n7963) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n9469), .CLK(n9849), 
        .Q(WX7284), .QN(n7961) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n9468), .CLK(n9849), 
        .Q(WX7286), .QN(n7959) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n9467), .CLK(n9850), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n9467), .CLK(n9850), 
        .Q(WX7290), .QN(n7956) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n9466), .CLK(n9850), 
        .Q(WX7292), .QN(n7954) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n9465), .CLK(n9851), 
        .Q(WX7294), .QN(n7952) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n9465), .CLK(n9851), 
        .Q(WX7296), .QN(n7950) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n9464), .CLK(n9851), 
        .Q(WX7298), .QN(n7948) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n9463), .CLK(n9852), 
        .Q(WX7300), .QN(n7946) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n9463), .CLK(n9852), 
        .Q(WX7302), .QN(n8212) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n9462), .CLK(n9852), 
        .Q(WX7304) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n9462), .CLK(n9852), 
        .Q(WX7306), .QN(n8214) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n9462), .CLK(n9852), 
        .Q(WX7308), .QN(n8215) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n9461), .CLK(n9853), 
        .Q(WX7310), .QN(n8216) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n9461), .CLK(n9853), 
        .Q(WX7312), .QN(n8217) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n9461), .CLK(n9853), 
        .Q(WX7314), .QN(n8218) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n9461), .CLK(n9853), 
        .Q(WX7316), .QN(n8219) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n9461), .CLK(n9853), 
        .Q(WX7318), .QN(n8220) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n9460), .CLK(n9853), 
        .Q(WX7320), .QN(n8221) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n9460), .CLK(n9853), 
        .Q(test_so63), .QN(n8800) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n9476), .CLK(n9845), 
        .Q(WX7324), .QN(n8222) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n9476), .CLK(n9845), 
        .Q(WX7326), .QN(n8223) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n9475), .CLK(n9846), 
        .Q(WX7328), .QN(n8224) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n9474), .CLK(n9846), 
        .Q(WX7330), .QN(n8225) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n9474), .CLK(n9846), 
        .Q(WX7332), .QN(n8114) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n9473), .CLK(n9847), 
        .Q(WX7334), .QN(n8226) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n9472), .CLK(n9847), 
        .Q(WX7336), .QN(n8227) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n9472), .CLK(n9847), 
        .Q(WX7338) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n9471), .CLK(n9848), 
        .Q(WX7340), .QN(n8229) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n9470), .CLK(n9848), 
        .Q(WX7342), .QN(n8115) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n9470), .CLK(n9848), 
        .Q(WX7344), .QN(n8230) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n9469), .CLK(n9849), 
        .Q(WX7346), .QN(n8231) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n9468), .CLK(n9849), 
        .Q(WX7348), .QN(n8232) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n9468), .CLK(n9849), 
        .Q(WX7350), .QN(n8233) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n9467), .CLK(n9850), 
        .Q(WX7352), .QN(n8234) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n9466), .CLK(n9850), 
        .Q(WX7354), .QN(n8235) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n9466), .CLK(n9850), 
        .Q(test_so64), .QN(n8796) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n9465), .CLK(n9851), 
        .Q(WX7358), .QN(n8236) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n9464), .CLK(n9851), 
        .Q(WX7360), .QN(n8237) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n9464), .CLK(n9851), 
        .Q(WX7362), .QN(n8238) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n9463), .CLK(n9852), 
        .Q(WX7364), .QN(n8129) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n9364), .CLK(n9901), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n9364), .CLK(n9901), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_3) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n9363), .CLK(n9902), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n9362), .CLK(n9902), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n9362), .CLK(n9902), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n9362), .CLK(n9902), .Q(CRC_OUT_4_10) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n9362), .CLK(
        n9902), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n9362), .CLK(
        n9902), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n9362), .CLK(n9902), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_15) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n9361), .CLK(
        n9903), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n9360), .CLK(
        n9903), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n9460), .CLK(
        n9853), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n9460), .CLK(
        n9853), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n9460), .CLK(
        n9853), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n9460), .CLK(
        n9853), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n9459), .CLK(n9854), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n9459), .CLK(
        n9854), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n1457), .SI(CRC_OUT_4_31), .SE(n9459), .CLK(n9854), .Q(WX8243) );
  SDFFX1 DFF_1153_Q_reg ( .D(n1458), .SI(WX8243), .SE(n9459), .CLK(n9854), .Q(
        n8411), .QN(n8886) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1459), .SI(n8411), .SE(n9459), .CLK(n9854), .Q(
        n8410), .QN(n8885) );
  SDFFX1 DFF_1155_Q_reg ( .D(n1460), .SI(n8410), .SE(n9459), .CLK(n9854), .Q(
        n8409), .QN(n8884) );
  SDFFX1 DFF_1156_Q_reg ( .D(n1461), .SI(n8409), .SE(n9458), .CLK(n9854), .Q(
        n8408), .QN(n8883) );
  SDFFX1 DFF_1157_Q_reg ( .D(n1462), .SI(n8408), .SE(n9458), .CLK(n9854), .Q(
        n8407), .QN(n8882) );
  SDFFX1 DFF_1158_Q_reg ( .D(n1463), .SI(n8407), .SE(n9458), .CLK(n9854), .Q(
        n8406), .QN(n8881) );
  SDFFX1 DFF_1159_Q_reg ( .D(n1464), .SI(n8406), .SE(n9458), .CLK(n9854), .Q(
        n8405), .QN(n8880) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1465), .SI(n8405), .SE(n9458), .CLK(n9854), .Q(
        n8404), .QN(n8879) );
  SDFFX1 DFF_1161_Q_reg ( .D(n1466), .SI(n8404), .SE(n9458), .CLK(n9854), .Q(
        n8403), .QN(n8878) );
  SDFFX1 DFF_1162_Q_reg ( .D(n1467), .SI(n8403), .SE(n9457), .CLK(n9855), .Q(
        n8402), .QN(n8877) );
  SDFFX1 DFF_1163_Q_reg ( .D(n1468), .SI(n8402), .SE(n9457), .CLK(n9855), .Q(
        n8401), .QN(n8876) );
  SDFFX1 DFF_1164_Q_reg ( .D(n509), .SI(n8401), .SE(n9557), .CLK(n9805), .Q(
        n8400), .QN(n8875) );
  SDFFX1 DFF_1165_Q_reg ( .D(n1469), .SI(n8400), .SE(n9556), .CLK(n9805), .Q(
        n8399), .QN(n8874) );
  SDFFX1 DFF_1166_Q_reg ( .D(n1470), .SI(n8399), .SE(n9556), .CLK(n9805), .Q(
        test_so67), .QN(n9064) );
  SDFFX1 DFF_1167_Q_reg ( .D(n1471), .SI(test_si68), .SE(n9454), .CLK(n9856), 
        .Q(n8396), .QN(n8873) );
  SDFFX1 DFF_1168_Q_reg ( .D(n1472), .SI(n8396), .SE(n9455), .CLK(n9856), .Q(
        n8395), .QN(n8872) );
  SDFFX1 DFF_1169_Q_reg ( .D(n1473), .SI(n8395), .SE(n9455), .CLK(n9856), .Q(
        n8394), .QN(n8871) );
  SDFFX1 DFF_1170_Q_reg ( .D(n1474), .SI(n8394), .SE(n9455), .CLK(n9856), .Q(
        n8393), .QN(n8870) );
  SDFFX1 DFF_1171_Q_reg ( .D(n1475), .SI(n8393), .SE(n9455), .CLK(n9856), .Q(
        n8392), .QN(n8869) );
  SDFFX1 DFF_1172_Q_reg ( .D(n1476), .SI(n8392), .SE(n9455), .CLK(n9856), .Q(
        n8391), .QN(n8868) );
  SDFFX1 DFF_1173_Q_reg ( .D(n1477), .SI(n8391), .SE(n9455), .CLK(n9856), .Q(
        n8390), .QN(n8867) );
  SDFFX1 DFF_1174_Q_reg ( .D(n1478), .SI(n8390), .SE(n9456), .CLK(n9855), .Q(
        n8389), .QN(n8866) );
  SDFFX1 DFF_1175_Q_reg ( .D(n1479), .SI(n8389), .SE(n9456), .CLK(n9855), .Q(
        n8388), .QN(n8865) );
  SDFFX1 DFF_1176_Q_reg ( .D(n1480), .SI(n8388), .SE(n9456), .CLK(n9855), .Q(
        n8387), .QN(n8864) );
  SDFFX1 DFF_1177_Q_reg ( .D(n1481), .SI(n8387), .SE(n9456), .CLK(n9855), .Q(
        n8386), .QN(n8863) );
  SDFFX1 DFF_1178_Q_reg ( .D(n1482), .SI(n8386), .SE(n9456), .CLK(n9855), .Q(
        n8385), .QN(n8862) );
  SDFFX1 DFF_1179_Q_reg ( .D(n1483), .SI(n8385), .SE(n9456), .CLK(n9855), .Q(
        n8384), .QN(n8861) );
  SDFFX1 DFF_1180_Q_reg ( .D(n1484), .SI(n8384), .SE(n9457), .CLK(n9855), .Q(
        n8383), .QN(n8860) );
  SDFFX1 DFF_1181_Q_reg ( .D(n1485), .SI(n8383), .SE(n9457), .CLK(n9855), .Q(
        n8382), .QN(n8859) );
  SDFFX1 DFF_1182_Q_reg ( .D(n1486), .SI(n8382), .SE(n9457), .CLK(n9855), .Q(
        n8381), .QN(n8858) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n9457), .CLK(n9855), .Q(
        test_so68), .QN(n9063) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n9454), .CLK(n9856), 
        .Q(n8378), .QN(n16382) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n9454), .CLK(n9856), .Q(
        n8377), .QN(n16383) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n9454), .CLK(n9856), .Q(
        n8376), .QN(n16384) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n9453), .CLK(n9857), .Q(
        n8375), .QN(n16385) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n9453), .CLK(n9857), .Q(
        n8374), .QN(n16386) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n9452), .CLK(n9857), .Q(
        n8373), .QN(n16387) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n9452), .CLK(n9857), .Q(
        n8372), .QN(n16388) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n9451), .CLK(n9858), .Q(
        n8371), .QN(n16389) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n9451), .CLK(n9858), .Q(
        n8370), .QN(n16390) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n9449), .CLK(n9859), .Q(
        n8369), .QN(n16391) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n9449), .CLK(n9859), .Q(
        n8368), .QN(n16392) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n9448), .CLK(n9859), .Q(
        n8367), .QN(n16393) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n9448), .CLK(n9859), .Q(
        n8366), .QN(n16394) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n9364), .CLK(n9901), .Q(
        n8365), .QN(n16395) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n9556), .CLK(n9805), .Q(
        n8364), .QN(n16396) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n9446), .CLK(n9860), .Q(
        n8363), .QN(n16397) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n9446), .CLK(n9860), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n9444), .CLK(n9861), 
        .Q(WX8437), .QN(n7942) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n9444), .CLK(n9861), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n9444), .CLK(n9861), 
        .Q(WX8441), .QN(n7938) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n9443), .CLK(n9862), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n9442), .CLK(n9862), 
        .Q(WX8445), .QN(n7935) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n9442), .CLK(n9862), 
        .Q(WX8447), .QN(n7933) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n9441), .CLK(n9863), 
        .Q(WX8449), .QN(n7931) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n9440), .CLK(n9863), 
        .Q(WX8451), .QN(n7929) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n9440), .CLK(n9863), 
        .Q(WX8453), .QN(n7927) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n9439), .CLK(n9864), 
        .Q(WX8455), .QN(n7925) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n9438), .CLK(n9864), 
        .Q(WX8457), .QN(n7923) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n9438), .CLK(n9864), 
        .Q(WX8459), .QN(n7921) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n9437), .CLK(n9865), 
        .Q(WX8461), .QN(n7919) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n9436), .CLK(n9865), 
        .Q(WX8463), .QN(n7917) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n9436), .CLK(n9865), 
        .Q(WX8465), .QN(n7915) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n9454), .CLK(n9856), 
        .Q(WX8467), .QN(n7616) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n9454), .CLK(n9856), 
        .Q(test_so70), .QN(n8809) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n9453), .CLK(n9857), 
        .Q(WX8471), .QN(n7709) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n9453), .CLK(n9857), 
        .Q(WX8473), .QN(n7708) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n9453), .CLK(n9857), 
        .Q(WX8475), .QN(n7706) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n9452), .CLK(n9857), 
        .Q(WX8477), .QN(n7704) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n9452), .CLK(n9857), 
        .Q(WX8479), .QN(n7702) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n9451), .CLK(n9858), 
        .Q(WX8481), .QN(n7700) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n9450), .CLK(n9858), 
        .Q(WX8483), .QN(n7698) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n9450), .CLK(n9858), 
        .Q(WX8485), .QN(n7696) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n9449), .CLK(n9859), 
        .Q(WX8487), .QN(n7694) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n9449), .CLK(n9859), 
        .Q(WX8489), .QN(n7692) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n9448), .CLK(n9859), 
        .Q(WX8491), .QN(n7690) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n9447), .CLK(n9860), 
        .Q(WX8493), .QN(n7688) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n9447), .CLK(n9860), 
        .Q(WX8495), .QN(n7686) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n9446), .CLK(n9860), 
        .Q(WX8497), .QN(n7684) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n9445), .CLK(n9861), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n9445), .CLK(n9861), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n9444), .CLK(n9861), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n9443), .CLK(n9862), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n9443), .CLK(n9862), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n9442), .CLK(n9862), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n9441), .CLK(n9863), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n9441), .CLK(n9863), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n9440), .CLK(n9863), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n9439), .CLK(n9864), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n9439), .CLK(n9864), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n9438), .CLK(n9864), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n9437), .CLK(n9865), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n9437), .CLK(n9865), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n9436), .CLK(n9865), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n9435), .CLK(n9866), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n9435), .CLK(n9866), 
        .Q(WX8531), .QN(n7617) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n9435), .CLK(n9866), 
        .Q(WX8533), .QN(n7711) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n9434), .CLK(n9866), 
        .Q(WX8535), .QN(n7710) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n9434), .CLK(n9866), 
        .Q(test_so72), .QN(n8808) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n9453), .CLK(n9857), 
        .Q(WX8539), .QN(n7707) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n9452), .CLK(n9857), 
        .Q(WX8541), .QN(n7705) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n9452), .CLK(n9857), 
        .Q(WX8543), .QN(n7703) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n9451), .CLK(n9858), 
        .Q(WX8545), .QN(n7701) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n9450), .CLK(n9858), 
        .Q(WX8547), .QN(n7699) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n9450), .CLK(n9858), 
        .Q(WX8549), .QN(n7697) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n9449), .CLK(n9859), 
        .Q(WX8551), .QN(n7695) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n9448), .CLK(n9859), 
        .Q(WX8553), .QN(n7693) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n9448), .CLK(n9859), 
        .Q(WX8555), .QN(n7691) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n9447), .CLK(n9860), 
        .Q(WX8557), .QN(n7689) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n9447), .CLK(n9860), 
        .Q(WX8559), .QN(n7687) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n9446), .CLK(n9860), 
        .Q(WX8561), .QN(n7685) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n9445), .CLK(n9861), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n9445), .CLK(n9861), 
        .Q(WX8565), .QN(n7943) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n9444), .CLK(n9861), 
        .Q(WX8567), .QN(n7941) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n9443), .CLK(n9862), 
        .Q(WX8569), .QN(n7939) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n9443), .CLK(n9862), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n9442), .CLK(n9862), 
        .Q(WX8573), .QN(n7936) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n9441), .CLK(n9863), 
        .Q(WX8575), .QN(n7934) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n9441), .CLK(n9863), 
        .Q(WX8577), .QN(n7932) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n9440), .CLK(n9863), 
        .Q(WX8579), .QN(n7930) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n9439), .CLK(n9864), 
        .Q(WX8581), .QN(n7928) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n9439), .CLK(n9864), 
        .Q(WX8583), .QN(n7926) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n9438), .CLK(n9864), 
        .Q(WX8585), .QN(n7924) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n9437), .CLK(n9865), 
        .Q(WX8587), .QN(n7922) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n9437), .CLK(n9865), 
        .Q(WX8589), .QN(n7920) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n9436), .CLK(n9865), 
        .Q(WX8591), .QN(n7918) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n9435), .CLK(n9866), 
        .Q(WX8593), .QN(n7916) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n9435), .CLK(n9866), 
        .Q(WX8595), .QN(n8186) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n9434), .CLK(n9866), 
        .Q(WX8597), .QN(n8187) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n9434), .CLK(n9866), 
        .Q(WX8599), .QN(n8188) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n9434), .CLK(n9866), 
        .Q(WX8601), .QN(n8189) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n9434), .CLK(n9866), 
        .Q(WX8603), .QN(n8190) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n9433), .CLK(n9867), 
        .Q(test_so74), .QN(n8799) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n9451), .CLK(n9858), 
        .Q(WX8607) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n9451), .CLK(n9858), 
        .Q(WX8609), .QN(n8192) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n9450), .CLK(n9858), 
        .Q(WX8611), .QN(n8193) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n9450), .CLK(n9858), 
        .Q(WX8613), .QN(n8194) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n9449), .CLK(n9859), 
        .Q(WX8615), .QN(n8195) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n9448), .CLK(n9859), 
        .Q(WX8617), .QN(n8196) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n9447), .CLK(n9860), 
        .Q(WX8619), .QN(n8197) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n9447), .CLK(n9860), 
        .Q(WX8621), .QN(n8198) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n9446), .CLK(n9860), 
        .Q(WX8623), .QN(n8199) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n9446), .CLK(n9860), 
        .Q(WX8625), .QN(n8111) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n9445), .CLK(n9861), 
        .Q(WX8627), .QN(n8200) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n9445), .CLK(n9861), 
        .Q(WX8629), .QN(n8201) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n9444), .CLK(n9861), 
        .Q(WX8631), .QN(n8202) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n9443), .CLK(n9862), 
        .Q(WX8633), .QN(n8203) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n9442), .CLK(n9862), 
        .Q(WX8635), .QN(n8112) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n9442), .CLK(n9862), 
        .Q(WX8637), .QN(n8204) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n9441), .CLK(n9863), 
        .Q(test_so75), .QN(n8791) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n9440), .CLK(n9863), 
        .Q(WX8641) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n9440), .CLK(n9863), 
        .Q(WX8643), .QN(n8206) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n9439), .CLK(n9864), 
        .Q(WX8645), .QN(n8207) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n9438), .CLK(n9864), 
        .Q(WX8647), .QN(n8208) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n9438), .CLK(n9864), 
        .Q(WX8649), .QN(n8113) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n9437), .CLK(n9865), 
        .Q(WX8651), .QN(n8209) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n9436), .CLK(n9865), 
        .Q(WX8653), .QN(n8210) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n9436), .CLK(n9865), 
        .Q(WX8655), .QN(n8211) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n9435), .CLK(n9866), 
        .Q(WX8657), .QN(n8128) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n9369), .CLK(n9899), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_3) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n9368), .CLK(n9899), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n9367), .CLK(n9900), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n9367), .CLK(n9900), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n9367), .CLK(n9900), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n9367), .CLK(n9900), .Q(CRC_OUT_3_10) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n9367), .CLK(
        n9900), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n9367), .CLK(
        n9900), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_15) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n9366), .CLK(
        n9900), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n9365), .CLK(
        n9901), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n9365), .CLK(
        n9901), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n9365), .CLK(
        n9901), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n9365), .CLK(
        n9901), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n9365), .CLK(
        n9901), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n9365), .CLK(
        n9901), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n9364), .CLK(n9901), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n9364), .CLK(
        n9901), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n9364), .CLK(
        n9901), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n9433), .CLK(
        n9867), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n9433), .CLK(
        n9867), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n9433), .CLK(
        n9867), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n9433), .CLK(
        n9867), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n1698), .SI(CRC_OUT_3_31), .SE(n9433), .CLK(n9867), .Q(WX9536) );
  SDFFX1 DFF_1345_Q_reg ( .D(n1699), .SI(WX9536), .SE(n9427), .CLK(n9870), .Q(
        n8353), .QN(n8857) );
  SDFFX1 DFF_1346_Q_reg ( .D(n1700), .SI(n8353), .SE(n9428), .CLK(n9869), .Q(
        n8352), .QN(n8856) );
  SDFFX1 DFF_1347_Q_reg ( .D(n1701), .SI(n8352), .SE(n9428), .CLK(n9869), .Q(
        n8351), .QN(n8855) );
  SDFFX1 DFF_1348_Q_reg ( .D(n1702), .SI(n8351), .SE(n9428), .CLK(n9869), .Q(
        n8350), .QN(n8854) );
  SDFFX1 DFF_1349_Q_reg ( .D(n1703), .SI(n8350), .SE(n9428), .CLK(n9869), .Q(
        n8349), .QN(n8853) );
  SDFFX1 DFF_1350_Q_reg ( .D(n1704), .SI(n8349), .SE(n9428), .CLK(n9869), .Q(
        n8348), .QN(n8852) );
  SDFFX1 DFF_1351_Q_reg ( .D(n1705), .SI(n8348), .SE(n9428), .CLK(n9869), .Q(
        n8347), .QN(n8851) );
  SDFFX1 DFF_1352_Q_reg ( .D(n1706), .SI(n8347), .SE(n9429), .CLK(n9869), .Q(
        n8346), .QN(n8850) );
  SDFFX1 DFF_1353_Q_reg ( .D(n1707), .SI(n8346), .SE(n9429), .CLK(n9869), .Q(
        test_so78), .QN(n9062) );
  SDFFX1 DFF_1354_Q_reg ( .D(n1708), .SI(test_si79), .SE(n9429), .CLK(n9869), 
        .Q(n8343), .QN(n8849) );
  SDFFX1 DFF_1355_Q_reg ( .D(n1709), .SI(n8343), .SE(n9429), .CLK(n9869), .Q(
        n8342), .QN(n8848) );
  SDFFX1 DFF_1356_Q_reg ( .D(n1710), .SI(n8342), .SE(n9429), .CLK(n9869), .Q(
        n8341), .QN(n8847) );
  SDFFX1 DFF_1357_Q_reg ( .D(n1711), .SI(n8341), .SE(n9429), .CLK(n9869), .Q(
        n8340), .QN(n8846) );
  SDFFX1 DFF_1358_Q_reg ( .D(n1712), .SI(n8340), .SE(n9430), .CLK(n9868), .Q(
        n8339), .QN(n8845) );
  SDFFX1 DFF_1359_Q_reg ( .D(n1713), .SI(n8339), .SE(n9430), .CLK(n9868), .Q(
        n8338), .QN(n8844) );
  SDFFX1 DFF_1360_Q_reg ( .D(n1714), .SI(n8338), .SE(n9430), .CLK(n9868), .Q(
        n8337), .QN(n8843) );
  SDFFX1 DFF_1361_Q_reg ( .D(n1715), .SI(n8337), .SE(n9430), .CLK(n9868), .Q(
        n8336), .QN(n8842) );
  SDFFX1 DFF_1362_Q_reg ( .D(n1716), .SI(n8336), .SE(n9430), .CLK(n9868), .Q(
        n8335), .QN(n8841) );
  SDFFX1 DFF_1363_Q_reg ( .D(n1717), .SI(n8335), .SE(n9430), .CLK(n9868), .Q(
        n8334), .QN(n8840) );
  SDFFX1 DFF_1364_Q_reg ( .D(n1718), .SI(n8334), .SE(n9431), .CLK(n9868), .Q(
        n8333), .QN(n8839) );
  SDFFX1 DFF_1365_Q_reg ( .D(n1719), .SI(n8333), .SE(n9431), .CLK(n9868), .Q(
        n8332), .QN(n8838) );
  SDFFX1 DFF_1366_Q_reg ( .D(n1720), .SI(n8332), .SE(n9431), .CLK(n9868), .Q(
        n8331), .QN(n8837) );
  SDFFX1 DFF_1367_Q_reg ( .D(n1721), .SI(n8331), .SE(n9431), .CLK(n9868), .Q(
        n8330), .QN(n8836) );
  SDFFX1 DFF_1368_Q_reg ( .D(n1722), .SI(n8330), .SE(n9431), .CLK(n9868), .Q(
        n8329), .QN(n8835) );
  SDFFX1 DFF_1369_Q_reg ( .D(n1723), .SI(n8329), .SE(n9431), .CLK(n9868), .Q(
        n8328), .QN(n8834) );
  SDFFX1 DFF_1370_Q_reg ( .D(n1724), .SI(n8328), .SE(n9432), .CLK(n9867), .Q(
        test_so79), .QN(n9061) );
  SDFFX1 DFF_1371_Q_reg ( .D(n1725), .SI(test_si80), .SE(n9432), .CLK(n9867), 
        .Q(n8325), .QN(n8833) );
  SDFFX1 DFF_1372_Q_reg ( .D(n1726), .SI(n8325), .SE(n9432), .CLK(n9867), .Q(
        n8324), .QN(n8832) );
  SDFFX1 DFF_1373_Q_reg ( .D(n1727), .SI(n8324), .SE(n9432), .CLK(n9867), .Q(
        n8323), .QN(n8831) );
  SDFFX1 DFF_1374_Q_reg ( .D(n1728), .SI(n8323), .SE(n9432), .CLK(n9867), .Q(
        n8322), .QN(n8830) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n9432), .CLK(n9867), .Q(
        n8321), .QN(n8829) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n9427), .CLK(n9870), .Q(
        n8320), .QN(n16398) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n9427), .CLK(n9870), .Q(
        n8319), .QN(n16399) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n9427), .CLK(n9870), .Q(
        n8318), .QN(n16400) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n9426), .CLK(n9870), .Q(
        n8317), .QN(n16401) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n9426), .CLK(n9870), .Q(
        n8316), .QN(n16402) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n9425), .CLK(n9871), .Q(
        n8315), .QN(n16403) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n9425), .CLK(n9871), .Q(
        n8314), .QN(n16404) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n9425), .CLK(n9871), .Q(
        n8313), .QN(n16405) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n9425), .CLK(n9871), .Q(
        n8312), .QN(n16406) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n9424), .CLK(n9871), .Q(
        n8311), .QN(n16407) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n9424), .CLK(n9871), .Q(
        n8310), .QN(n16408) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n9369), .CLK(n9899), .Q(
        test_so80), .QN(n8820) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n9423), .CLK(n9872), 
        .Q(n8307), .QN(n16409) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n9423), .CLK(n9872), .Q(
        n8306), .QN(n16410) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n9422), .CLK(n9872), .Q(
        n8305), .QN(n16411) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n9422), .CLK(n9872), .Q(
        n8304), .QN(n16412) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n9422), .CLK(n9872), .Q(
        WX9728), .QN(n7913) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n9421), .CLK(n9873), 
        .Q(WX9730), .QN(n7911) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n9421), .CLK(n9873), 
        .Q(WX9732), .QN(n7909) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n9420), .CLK(n9873), 
        .Q(WX9734), .QN(n7907) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n9419), .CLK(n9874), 
        .Q(WX9736), .QN(n7905) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n9419), .CLK(n9874), 
        .Q(WX9738), .QN(n7903) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n9418), .CLK(n9874), 
        .Q(WX9740), .QN(n7901) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n9417), .CLK(n9875), 
        .Q(WX9742), .QN(n7899) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n9417), .CLK(n9875), 
        .Q(WX9744), .QN(n7897) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n9416), .CLK(n9875), 
        .Q(WX9746), .QN(n7895) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n9415), .CLK(n9876), 
        .Q(WX9748), .QN(n7893) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n9415), .CLK(n9876), 
        .Q(WX9750), .QN(n7891) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n9414), .CLK(n9876), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n9413), .CLK(n9877), 
        .Q(WX9754), .QN(n7888) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n9413), .CLK(n9877), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n9412), .CLK(n9877), 
        .Q(WX9758), .QN(n7884) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n9427), .CLK(n9870), 
        .Q(WX9760), .QN(n7614) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n9427), .CLK(n9870), 
        .Q(WX9762), .QN(n7682) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n9426), .CLK(n9870), 
        .Q(WX9764), .QN(n7680) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n9426), .CLK(n9870), 
        .Q(WX9766), .QN(n7678) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n9426), .CLK(n9870), 
        .Q(WX9768), .QN(n7676) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n9426), .CLK(n9870), 
        .Q(WX9770), .QN(n7674) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n9425), .CLK(n9871), 
        .Q(WX9772), .QN(n7672) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n9425), .CLK(n9871), 
        .Q(WX9774), .QN(n7670) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n9424), .CLK(n9871), 
        .Q(WX9776), .QN(n7668) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n9424), .CLK(n9871), 
        .Q(WX9778), .QN(n7666) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n9424), .CLK(n9871), 
        .Q(WX9780), .QN(n7664) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n9424), .CLK(n9871), 
        .Q(WX9782), .QN(n7662) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n9423), .CLK(n9872), 
        .Q(WX9784), .QN(n7660) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n9423), .CLK(n9872), 
        .Q(test_so82), .QN(n8807) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n9422), .CLK(n9872), 
        .Q(WX9788), .QN(n7657) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n9422), .CLK(n9872), 
        .Q(WX9790), .QN(n7656) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n9421), .CLK(n9873), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n9421), .CLK(n9873), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n9420), .CLK(n9873), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n9420), .CLK(n9873), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n9419), .CLK(n9874), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n9418), .CLK(n9874), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n9418), .CLK(n9874), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n9417), .CLK(n9875), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n9416), .CLK(n9875), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n9416), .CLK(n9875), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n9415), .CLK(n9876), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n9414), .CLK(n9876), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n9414), .CLK(n9876), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n9413), .CLK(n9877), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n9412), .CLK(n9877), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n9412), .CLK(n9877), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n9411), .CLK(n9878), 
        .Q(WX9824), .QN(n7615) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n9411), .CLK(n9878), 
        .Q(WX9826), .QN(n7683) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n9411), .CLK(n9878), 
        .Q(WX9828), .QN(n7681) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n9410), .CLK(n9878), 
        .Q(WX9830), .QN(n7679) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n9410), .CLK(n9878), 
        .Q(WX9832), .QN(n7677) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n9410), .CLK(n9878), 
        .Q(WX9834), .QN(n7675) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n9409), .CLK(n9879), 
        .Q(WX9836), .QN(n7673) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n9409), .CLK(n9879), 
        .Q(WX9838), .QN(n7671) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n9409), .CLK(n9879), 
        .Q(WX9840), .QN(n7669) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n9408), .CLK(n9879), 
        .Q(WX9842), .QN(n7667) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n9408), .CLK(n9879), 
        .Q(WX9844), .QN(n7665) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n9408), .CLK(n9879), 
        .Q(WX9846), .QN(n7663) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n9407), .CLK(n9880), 
        .Q(WX9848), .QN(n7661) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n9423), .CLK(n9872), 
        .Q(WX9850), .QN(n7659) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n9423), .CLK(n9872), 
        .Q(WX9852), .QN(n7658) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n9422), .CLK(n9872), 
        .Q(test_so84), .QN(n8806) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n9421), .CLK(n9873), 
        .Q(WX9856), .QN(n7914) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n9421), .CLK(n9873), 
        .Q(WX9858), .QN(n7912) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n9420), .CLK(n9873), 
        .Q(WX9860), .QN(n7910) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n9420), .CLK(n9873), 
        .Q(WX9862), .QN(n7908) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n9419), .CLK(n9874), 
        .Q(WX9864), .QN(n7906) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n9418), .CLK(n9874), 
        .Q(WX9866), .QN(n7904) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n9418), .CLK(n9874), 
        .Q(WX9868), .QN(n7902) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n9417), .CLK(n9875), 
        .Q(WX9870), .QN(n7900) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n9416), .CLK(n9875), 
        .Q(WX9872), .QN(n7898) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n9416), .CLK(n9875), 
        .Q(WX9874), .QN(n7896) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n9415), .CLK(n9876), 
        .Q(WX9876), .QN(n7894) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n9414), .CLK(n9876), 
        .Q(WX9878), .QN(n7892) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n9414), .CLK(n9876), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n9413), .CLK(n9877), 
        .Q(WX9882), .QN(n7889) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n9412), .CLK(n9877), 
        .Q(WX9884), .QN(n7887) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n9412), .CLK(n9877), 
        .Q(WX9886), .QN(n7885) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n9411), .CLK(n9878), 
        .Q(test_so85), .QN(n8805) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n9411), .CLK(n9878), 
        .Q(WX9890), .QN(n8160) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n9410), .CLK(n9878), 
        .Q(WX9892), .QN(n8161) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n9410), .CLK(n9878), 
        .Q(WX9894), .QN(n8162) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n9410), .CLK(n9878), 
        .Q(WX9896), .QN(n8163) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n9409), .CLK(n9879), 
        .Q(WX9898), .QN(n8164) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n9409), .CLK(n9879), 
        .Q(WX9900), .QN(n8165) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n9409), .CLK(n9879), 
        .Q(WX9902), .QN(n8166) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n9408), .CLK(n9879), 
        .Q(WX9904), .QN(n8167) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n9408), .CLK(n9879), 
        .Q(WX9906), .QN(n8168) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n9408), .CLK(n9879), 
        .Q(WX9908), .QN(n8169) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n9407), .CLK(n9880), 
        .Q(WX9910), .QN(n8170) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n9407), .CLK(n9880), 
        .Q(WX9912), .QN(n8171) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n9407), .CLK(n9880), 
        .Q(WX9914), .QN(n8172) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n9407), .CLK(n9880), 
        .Q(WX9916), .QN(n8173) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n9407), .CLK(n9880), 
        .Q(WX9918), .QN(n8108) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n9406), .CLK(n9880), 
        .Q(WX9920), .QN(n8174) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n9406), .CLK(n9880), 
        .Q(test_so86), .QN(n8795) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n9420), .CLK(n9873), 
        .Q(WX9924), .QN(n8175) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n9419), .CLK(n9874), 
        .Q(WX9926), .QN(n8176) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n9419), .CLK(n9874), 
        .Q(WX9928), .QN(n8109) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n9418), .CLK(n9874), 
        .Q(WX9930), .QN(n8177) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n9417), .CLK(n9875), 
        .Q(WX9932), .QN(n8178) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n9417), .CLK(n9875), 
        .Q(WX9934), .QN(n8179) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n9416), .CLK(n9875), 
        .Q(WX9936), .QN(n8180) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n9415), .CLK(n9876), 
        .Q(WX9938), .QN(n8181) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n9415), .CLK(n9876), 
        .Q(WX9940), .QN(n8182) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n9414), .CLK(n9876), 
        .Q(WX9942), .QN(n8110) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n9413), .CLK(n9877), 
        .Q(WX9944), .QN(n8183) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n9413), .CLK(n9877), 
        .Q(WX9946), .QN(n8184) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n9412), .CLK(n9877), 
        .Q(WX9948), .QN(n8185) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n9411), .CLK(n9878), 
        .Q(WX9950), .QN(n8127) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n9372), .CLK(n9897), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n9372), .CLK(
        n9897), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n9372), .CLK(
        n9897), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n9371), .CLK(n9898), 
        .Q(CRC_OUT_2_3) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n9371), .CLK(
        n9898), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n9371), .CLK(
        n9898), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n9371), .CLK(
        n9898), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n9371), .CLK(
        n9898), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n9371), .CLK(
        n9898), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_10) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n9370), .CLK(
        n9898), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n9369), .CLK(
        n9899), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n9369), .CLK(
        n9899), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n9369), .CLK(
        n9899), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n9369), .CLK(
        n9899), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n9406), .CLK(
        n9880), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n9406), .CLK(n9880), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n9406), .CLK(
        n9880), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n9406), .CLK(
        n9880), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n9405), .CLK(
        n9881), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n9404), .CLK(
        n9881), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n9404), .CLK(
        n9881), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n9404), .CLK(
        n9881), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n1939), .SI(CRC_OUT_2_31), .SE(n9404), .CLK(n9881), .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(n1940), .SI(WX10829), .SE(n9399), .CLK(n9884), 
        .Q(n8295), .QN(n9060) );
  SDFFX1 DFF_1538_Q_reg ( .D(n1941), .SI(n8295), .SE(n9399), .CLK(n9884), .Q(
        n8294), .QN(n9059) );
  SDFFX1 DFF_1539_Q_reg ( .D(n1942), .SI(n8294), .SE(n9399), .CLK(n9884), .Q(
        n8293), .QN(n9058) );
  SDFFX1 DFF_1540_Q_reg ( .D(n1943), .SI(n8293), .SE(n9399), .CLK(n9884), .Q(
        test_so89), .QN(n9076) );
  SDFFX1 DFF_1541_Q_reg ( .D(n1944), .SI(test_si90), .SE(n9399), .CLK(n9884), 
        .Q(n8290), .QN(n9057) );
  SDFFX1 DFF_1542_Q_reg ( .D(n1945), .SI(n8290), .SE(n9400), .CLK(n9883), .Q(
        n8289), .QN(n9056) );
  SDFFX1 DFF_1543_Q_reg ( .D(n1946), .SI(n8289), .SE(n9400), .CLK(n9883), .Q(
        n8288), .QN(n9055) );
  SDFFX1 DFF_1544_Q_reg ( .D(n1947), .SI(n8288), .SE(n9400), .CLK(n9883), .Q(
        n8287), .QN(n9054) );
  SDFFX1 DFF_1545_Q_reg ( .D(n1948), .SI(n8287), .SE(n9400), .CLK(n9883), .Q(
        n8286), .QN(n9053) );
  SDFFX1 DFF_1546_Q_reg ( .D(n1949), .SI(n8286), .SE(n9400), .CLK(n9883), .Q(
        n8285), .QN(n9052) );
  SDFFX1 DFF_1547_Q_reg ( .D(n1950), .SI(n8285), .SE(n9400), .CLK(n9883), .Q(
        n8284), .QN(n9051) );
  SDFFX1 DFF_1548_Q_reg ( .D(n1951), .SI(n8284), .SE(n9401), .CLK(n9883), .Q(
        n8283), .QN(n9050) );
  SDFFX1 DFF_1549_Q_reg ( .D(n1952), .SI(n8283), .SE(n9401), .CLK(n9883), .Q(
        n8282), .QN(n9049) );
  SDFFX1 DFF_1550_Q_reg ( .D(n1953), .SI(n8282), .SE(n9401), .CLK(n9883), .Q(
        n8281), .QN(n9048) );
  SDFFX1 DFF_1551_Q_reg ( .D(n1954), .SI(n8281), .SE(n9401), .CLK(n9883), .Q(
        n8280), .QN(n9047) );
  SDFFX1 DFF_1552_Q_reg ( .D(n1955), .SI(n8280), .SE(n9401), .CLK(n9883), .Q(
        n8279), .QN(n9046) );
  SDFFX1 DFF_1553_Q_reg ( .D(n1956), .SI(n8279), .SE(n9401), .CLK(n9883), .Q(
        n8278), .QN(n9045) );
  SDFFX1 DFF_1554_Q_reg ( .D(n1957), .SI(n8278), .SE(n9402), .CLK(n9882), .Q(
        n8277), .QN(n9044) );
  SDFFX1 DFF_1555_Q_reg ( .D(n1958), .SI(n8277), .SE(n9402), .CLK(n9882), .Q(
        n8276), .QN(n9043) );
  SDFFX1 DFF_1556_Q_reg ( .D(n1959), .SI(n8276), .SE(n9402), .CLK(n9882), .Q(
        n8275), .QN(n9042) );
  SDFFX1 DFF_1557_Q_reg ( .D(n1960), .SI(n8275), .SE(n9402), .CLK(n9882), .Q(
        test_so90), .QN(n9075) );
  SDFFX1 DFF_1558_Q_reg ( .D(n1961), .SI(test_si91), .SE(n9402), .CLK(n9882), 
        .Q(n8272), .QN(n9041) );
  SDFFX1 DFF_1559_Q_reg ( .D(n1962), .SI(n8272), .SE(n9402), .CLK(n9882), .Q(
        n8271), .QN(n9040) );
  SDFFX1 DFF_1560_Q_reg ( .D(n1963), .SI(n8271), .SE(n9403), .CLK(n9882), .Q(
        n8270), .QN(n9039) );
  SDFFX1 DFF_1561_Q_reg ( .D(n1964), .SI(n8270), .SE(n9403), .CLK(n9882), .Q(
        n8269), .QN(n9038) );
  SDFFX1 DFF_1562_Q_reg ( .D(n1965), .SI(n8269), .SE(n9403), .CLK(n9882), .Q(
        n8268), .QN(n9037) );
  SDFFX1 DFF_1563_Q_reg ( .D(n1966), .SI(n8268), .SE(n9403), .CLK(n9882), .Q(
        n8267), .QN(n9036) );
  SDFFX1 DFF_1564_Q_reg ( .D(n1967), .SI(n8267), .SE(n9403), .CLK(n9882), .Q(
        n8266), .QN(n9035) );
  SDFFX1 DFF_1565_Q_reg ( .D(n1968), .SI(n8266), .SE(n9403), .CLK(n9882), .Q(
        n8265), .QN(n9034) );
  SDFFX1 DFF_1566_Q_reg ( .D(n1969), .SI(n8265), .SE(n9404), .CLK(n9881), .Q(
        n8264), .QN(n9033) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n9404), .CLK(n9881), 
        .Q(n8263), .QN(n9032) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n9399), .CLK(n9884), 
        .Q(n8262), .QN(n16413) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n9398), .CLK(n9884), 
        .Q(n8261), .QN(n16414) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n9398), .CLK(n9884), 
        .Q(n8260), .QN(n16415) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n9397), .CLK(n9885), 
        .Q(n8259), .QN(n16416) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n9397), .CLK(n9885), 
        .Q(n8258), .QN(n16417) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n9397), .CLK(n9885), 
        .Q(n8257), .QN(n16418) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n9397), .CLK(n9885), 
        .Q(test_so91), .QN(n8826) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n9396), .CLK(n9885), 
        .Q(n8254), .QN(n16419) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n9396), .CLK(n9885), 
        .Q(n8253), .QN(n16420) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n9395), .CLK(n9886), 
        .Q(n8252), .QN(n16421) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n9395), .CLK(n9886), 
        .Q(n8251), .QN(n16422) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n9394), .CLK(n9886), 
        .Q(n8250), .QN(n16423) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n9394), .CLK(n9886), 
        .Q(n8249), .QN(n16424) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n9393), .CLK(n9887), 
        .Q(n8248), .QN(n16425) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n9392), .CLK(n9887), 
        .Q(n8247), .QN(n16426) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n9392), .CLK(n9887), 
        .Q(n8246), .QN(n16427) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n9391), .CLK(n9888), 
        .Q(WX11021), .QN(n7882) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n9391), .CLK(n9888), 
        .Q(WX11023), .QN(n7880) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n9390), .CLK(n9888), 
        .Q(WX11025), .QN(n7878) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n9389), .CLK(n9889), 
        .Q(WX11027), .QN(n7876) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n9389), .CLK(n9889), 
        .Q(WX11029), .QN(n7874) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n9388), .CLK(n9889), 
        .Q(WX11031), .QN(n7872) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n9387), .CLK(n9890), 
        .Q(WX11033), .QN(n7870) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n9387), .CLK(n9890), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n9386), .CLK(n9890), 
        .Q(WX11037), .QN(n7867) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n9385), .CLK(n9891), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n9385), .CLK(n9891), 
        .Q(WX11041), .QN(n7863) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n9384), .CLK(n9891), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n9383), .CLK(n9892), 
        .Q(WX11045), .QN(n7860) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n9383), .CLK(n9892), 
        .Q(WX11047), .QN(n7858) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n9382), .CLK(n9892), 
        .Q(WX11049), .QN(n7856) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n9381), .CLK(n9893), 
        .Q(WX11051), .QN(n7854) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n9398), .CLK(n9884), 
        .Q(WX11053), .QN(n7612) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n9398), .CLK(n9884), 
        .Q(WX11055), .QN(n7654) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n9398), .CLK(n9884), 
        .Q(WX11057), .QN(n7652) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n9398), .CLK(n9884), 
        .Q(WX11059), .QN(n7650) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n9397), .CLK(n9885), 
        .Q(WX11061), .QN(n7648) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n9397), .CLK(n9885), 
        .Q(WX11063), .QN(n7646) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n9396), .CLK(n9885), 
        .Q(WX11065), .QN(n7644) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n9396), .CLK(n9885), 
        .Q(WX11067), .QN(n7642) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n9396), .CLK(n9885), 
        .Q(test_so93), .QN(n8819) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n9395), .CLK(n9886), 
        .Q(WX11071), .QN(n7639) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n9395), .CLK(n9886), 
        .Q(WX11073), .QN(n7638) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n9394), .CLK(n9886), 
        .Q(WX11075), .QN(n7636) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n9394), .CLK(n9886), 
        .Q(WX11077), .QN(n7634) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n9393), .CLK(n9887), 
        .Q(WX11079), .QN(n7632) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n9393), .CLK(n9887), 
        .Q(WX11081), .QN(n7630) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n9392), .CLK(n9887), 
        .Q(WX11083), .QN(n7628) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n9391), .CLK(n9888), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n9391), .CLK(n9888), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n9390), .CLK(n9888), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n9389), .CLK(n9889), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n9389), .CLK(n9889), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n9388), .CLK(n9889), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n9387), .CLK(n9890), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n9387), .CLK(n9890), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n9386), .CLK(n9890), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n9385), .CLK(n9891), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n9385), .CLK(n9891), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n9384), .CLK(n9891), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n9383), .CLK(n9892), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n9383), .CLK(n9892), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n9382), .CLK(n9892), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n9381), .CLK(n9893), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n9381), .CLK(n9893), 
        .Q(WX11117), .QN(n7613) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n9380), .CLK(n9893), 
        .Q(WX11119), .QN(n7655) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n9380), .CLK(n9893), 
        .Q(WX11121), .QN(n7653) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n9380), .CLK(n9893), 
        .Q(WX11123), .QN(n7651) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n9379), .CLK(n9894), 
        .Q(WX11125), .QN(n7649) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n9379), .CLK(n9894), 
        .Q(WX11127), .QN(n7647) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n9379), .CLK(n9894), 
        .Q(WX11129), .QN(n7645) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n9378), .CLK(n9894), 
        .Q(WX11131), .QN(n7643) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n9396), .CLK(n9885), 
        .Q(WX11133), .QN(n7641) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n9395), .CLK(n9886), 
        .Q(WX11135), .QN(n7640) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n9395), .CLK(n9886), 
        .Q(test_so95), .QN(n8818) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n9394), .CLK(n9886), 
        .Q(WX11139), .QN(n7637) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n9394), .CLK(n9886), 
        .Q(WX11141), .QN(n7635) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n9393), .CLK(n9887), 
        .Q(WX11143), .QN(n7633) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n9393), .CLK(n9887), 
        .Q(WX11145), .QN(n7631) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n9392), .CLK(n9887), 
        .Q(WX11147), .QN(n7629) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n9391), .CLK(n9888), 
        .Q(WX11149), .QN(n7883) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n9390), .CLK(n9888), 
        .Q(WX11151), .QN(n7881) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n9390), .CLK(n9888), 
        .Q(WX11153), .QN(n7879) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n9389), .CLK(n9889), 
        .Q(WX11155), .QN(n7877) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n9388), .CLK(n9889), 
        .Q(WX11157), .QN(n7875) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n9388), .CLK(n9889), 
        .Q(WX11159), .QN(n7873) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n9387), .CLK(n9890), 
        .Q(WX11161), .QN(n7871) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n9386), .CLK(n9890), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n9386), .CLK(n9890), 
        .Q(WX11165), .QN(n7868) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n9385), .CLK(n9891), 
        .Q(WX11167), .QN(n7866) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n9384), .CLK(n9891), 
        .Q(WX11169), .QN(n7864) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n9384), .CLK(n9891), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n9383), .CLK(n9892), 
        .Q(WX11173), .QN(n7861) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n9382), .CLK(n9892), 
        .Q(WX11175), .QN(n7859) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n9382), .CLK(n9892), 
        .Q(WX11177), .QN(n7857) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n9381), .CLK(n9893), 
        .Q(WX11179), .QN(n7855) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n9381), .CLK(n9893), 
        .Q(WX11181), .QN(n8134) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n9380), .CLK(n9893), 
        .Q(WX11183), .QN(n8135) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n9380), .CLK(n9893), 
        .Q(WX11185), .QN(n8136) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n9380), .CLK(n9893), 
        .Q(WX11187), .QN(n8137) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n9379), .CLK(n9894), 
        .Q(WX11189), .QN(n8138) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n9379), .CLK(n9894), 
        .Q(WX11191), .QN(n8139) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n9379), .CLK(n9894), 
        .Q(WX11193), .QN(n8140) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n9378), .CLK(n9894), 
        .Q(WX11195), .QN(n8141) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n9378), .CLK(n9894), 
        .Q(WX11197), .QN(n8142) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n9378), .CLK(n9894), 
        .Q(WX11199), .QN(n8143) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n9378), .CLK(n9894), 
        .Q(WX11201), .QN(n8144) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n9378), .CLK(n9894), 
        .Q(WX11203), .QN(n8145) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n9377), .CLK(n9895), 
        .Q(test_so97), .QN(n8804) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n9393), .CLK(n9887), 
        .Q(WX11207), .QN(n8146) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n9392), .CLK(n9887), 
        .Q(WX11209), .QN(n8147) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n9392), .CLK(n9887), 
        .Q(WX11211), .QN(n8105) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n9391), .CLK(n9888), 
        .Q(WX11213) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n9390), .CLK(n9888), 
        .Q(WX11215), .QN(n8149) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n9390), .CLK(n9888), 
        .Q(WX11217), .QN(n8150) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n9389), .CLK(n9889), 
        .Q(WX11219), .QN(n8151) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n9388), .CLK(n9889), 
        .Q(WX11221), .QN(n8106) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n9388), .CLK(n9889), 
        .Q(WX11223), .QN(n8152) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n9387), .CLK(n9890), 
        .Q(WX11225), .QN(n8153) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n9386), .CLK(n9890), 
        .Q(WX11227), .QN(n8154) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n9386), .CLK(n9890), 
        .Q(WX11229), .QN(n8155) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n9385), .CLK(n9891), 
        .Q(WX11231), .QN(n8156) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n9384), .CLK(n9891), 
        .Q(WX11233), .QN(n8157) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n9384), .CLK(n9891), 
        .Q(WX11235), .QN(n8107) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n9383), .CLK(n9892), 
        .Q(WX11237), .QN(n8158) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n9382), .CLK(n9892), 
        .Q(test_so98), .QN(n8794) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n9382), .CLK(n9892), 
        .Q(WX11241), .QN(n8159) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n9381), .CLK(n9893), 
        .Q(WX11243), .QN(n8126) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n9376), .CLK(n9895), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n9376), .CLK(
        n9895), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n9376), .CLK(
        n9895), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_3) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n9375), .CLK(
        n9896), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n9374), .CLK(
        n9896), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n9374), .CLK(
        n9896), .Q(CRC_OUT_1_10) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n9374), .CLK(
        n9896), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n9374), .CLK(
        n9896), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n9374), .CLK(
        n9896), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n9374), .CLK(
        n9896), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n9373), .CLK(n9897), .Q(CRC_OUT_1_15) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n9373), .CLK(
        n9897), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n9373), .CLK(
        n9897), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n9373), .CLK(
        n9897), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n9373), .CLK(
        n9897), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n9373), .CLK(
        n9897), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n9372), .CLK(
        n9897), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n9372), .CLK(
        n9897), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n9372), .CLK(
        n9897), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n9377), .CLK(
        n9895), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n9377), .CLK(
        n9895), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n9377), .CLK(
        n9895), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n9377), .CLK(
        n9895), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n9377), .CLK(
        n9895), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n9376), .CLK(
        n9895), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n9376), .CLK(
        n9895), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n9376), .CLK(
        n9895), .Q(test_so100), .QN(n8790) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n510), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n522), .IN2(n514), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n1956), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  INVX0 TrojanINVtest_se ( .INP(n9755), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  INVX0 U8974 ( .INP(n10069), .ZN(n9077) );
  INVX0 U8975 ( .INP(n9077), .ZN(n9078) );
  INVX0 U8976 ( .INP(n9077), .ZN(n9079) );
  INVX0 U8977 ( .INP(n9077), .ZN(n9080) );
  INVX0 U8978 ( .INP(n10068), .ZN(n9081) );
  INVX0 U8979 ( .INP(n9081), .ZN(n9082) );
  INVX0 U8980 ( .INP(n9081), .ZN(n9083) );
  INVX0 U8981 ( .INP(n9081), .ZN(n9084) );
  NBUFFX2 U8982 ( .INP(n9260), .Z(n9155) );
  NBUFFX2 U8983 ( .INP(n9245), .Z(n9228) );
  NBUFFX2 U8984 ( .INP(n9245), .Z(n9229) );
  NBUFFX2 U8985 ( .INP(n9245), .Z(n9231) );
  NBUFFX2 U8986 ( .INP(n9245), .Z(n9230) );
  NBUFFX2 U8987 ( .INP(n9246), .Z(n9224) );
  NBUFFX2 U8988 ( .INP(n9245), .Z(n9232) );
  NBUFFX2 U8989 ( .INP(n9244), .Z(n9233) );
  NBUFFX2 U8990 ( .INP(n9244), .Z(n9234) );
  NBUFFX2 U8991 ( .INP(n9244), .Z(n9236) );
  NBUFFX2 U8992 ( .INP(n9244), .Z(n9237) );
  NBUFFX2 U8993 ( .INP(n9243), .Z(n9238) );
  NBUFFX2 U8994 ( .INP(n9243), .Z(n9239) );
  NBUFFX2 U8995 ( .INP(n9243), .Z(n9240) );
  NBUFFX2 U8996 ( .INP(n9243), .Z(n9241) );
  NBUFFX2 U8997 ( .INP(n9246), .Z(n9227) );
  NBUFFX2 U8998 ( .INP(n9246), .Z(n9226) );
  NBUFFX2 U8999 ( .INP(n9246), .Z(n9225) );
  NBUFFX2 U9000 ( .INP(n9244), .Z(n9235) );
  NBUFFX2 U9001 ( .INP(n9261), .Z(n9148) );
  NBUFFX2 U9002 ( .INP(n9261), .Z(n9152) );
  NBUFFX2 U9003 ( .INP(n9262), .Z(n9147) );
  NBUFFX2 U9004 ( .INP(n9262), .Z(n9146) );
  NBUFFX2 U9005 ( .INP(n9262), .Z(n9145) );
  NBUFFX2 U9006 ( .INP(n9262), .Z(n9144) );
  NBUFFX2 U9007 ( .INP(n9262), .Z(n9143) );
  NBUFFX2 U9008 ( .INP(n9263), .Z(n9142) );
  NBUFFX2 U9009 ( .INP(n9263), .Z(n9140) );
  NBUFFX2 U9010 ( .INP(n9263), .Z(n9139) );
  NBUFFX2 U9011 ( .INP(n9263), .Z(n9138) );
  NBUFFX2 U9012 ( .INP(n9263), .Z(n9141) );
  NBUFFX2 U9013 ( .INP(n9260), .Z(n9153) );
  NBUFFX2 U9014 ( .INP(n9260), .Z(n9154) );
  NBUFFX2 U9015 ( .INP(n9261), .Z(n9151) );
  NBUFFX2 U9016 ( .INP(n9261), .Z(n9150) );
  NBUFFX2 U9017 ( .INP(n9261), .Z(n9149) );
  NBUFFX2 U9018 ( .INP(n9259), .Z(n9158) );
  NBUFFX2 U9019 ( .INP(n9260), .Z(n9157) );
  NBUFFX2 U9020 ( .INP(n9260), .Z(n9156) );
  NBUFFX2 U9021 ( .INP(n9258), .Z(n9164) );
  NBUFFX2 U9022 ( .INP(n9258), .Z(n9163) );
  NBUFFX2 U9023 ( .INP(n9259), .Z(n9159) );
  NBUFFX2 U9024 ( .INP(n9259), .Z(n9160) );
  NBUFFX2 U9025 ( .INP(n9259), .Z(n9161) );
  NBUFFX2 U9026 ( .INP(n9259), .Z(n9162) );
  NBUFFX2 U9027 ( .INP(n9252), .Z(n9196) );
  NBUFFX2 U9028 ( .INP(n9252), .Z(n9197) );
  NBUFFX2 U9029 ( .INP(n9251), .Z(n9199) );
  NBUFFX2 U9030 ( .INP(n9251), .Z(n9200) );
  NBUFFX2 U9031 ( .INP(n9251), .Z(n9201) );
  NBUFFX2 U9032 ( .INP(n9251), .Z(n9202) );
  NBUFFX2 U9033 ( .INP(n9250), .Z(n9203) );
  NBUFFX2 U9034 ( .INP(n9255), .Z(n9181) );
  NBUFFX2 U9035 ( .INP(n9255), .Z(n9182) );
  NBUFFX2 U9036 ( .INP(n9254), .Z(n9183) );
  NBUFFX2 U9037 ( .INP(n9254), .Z(n9184) );
  NBUFFX2 U9038 ( .INP(n9254), .Z(n9185) );
  NBUFFX2 U9039 ( .INP(n9254), .Z(n9186) );
  NBUFFX2 U9040 ( .INP(n9254), .Z(n9187) );
  NBUFFX2 U9041 ( .INP(n9253), .Z(n9188) );
  NBUFFX2 U9042 ( .INP(n9253), .Z(n9189) );
  NBUFFX2 U9043 ( .INP(n9253), .Z(n9190) );
  NBUFFX2 U9044 ( .INP(n9253), .Z(n9191) );
  NBUFFX2 U9045 ( .INP(n9247), .Z(n9222) );
  NBUFFX2 U9046 ( .INP(n9246), .Z(n9223) );
  NBUFFX2 U9047 ( .INP(n9247), .Z(n9221) );
  NBUFFX2 U9048 ( .INP(n9247), .Z(n9220) );
  NBUFFX2 U9049 ( .INP(n9250), .Z(n9205) );
  NBUFFX2 U9050 ( .INP(n9250), .Z(n9206) );
  NBUFFX2 U9051 ( .INP(n9249), .Z(n9208) );
  NBUFFX2 U9052 ( .INP(n9249), .Z(n9209) );
  NBUFFX2 U9053 ( .INP(n9249), .Z(n9210) );
  NBUFFX2 U9054 ( .INP(n9249), .Z(n9211) );
  NBUFFX2 U9055 ( .INP(n9247), .Z(n9219) );
  NBUFFX2 U9056 ( .INP(n9247), .Z(n9218) );
  NBUFFX2 U9057 ( .INP(n9248), .Z(n9217) );
  NBUFFX2 U9058 ( .INP(n9248), .Z(n9216) );
  NBUFFX2 U9059 ( .INP(n9248), .Z(n9214) );
  NBUFFX2 U9060 ( .INP(n9248), .Z(n9213) );
  NBUFFX2 U9061 ( .INP(n9249), .Z(n9212) );
  NBUFFX2 U9062 ( .INP(n9248), .Z(n9215) );
  NBUFFX2 U9063 ( .INP(n9250), .Z(n9207) );
  NBUFFX2 U9064 ( .INP(n9252), .Z(n9195) );
  NBUFFX2 U9065 ( .INP(n9257), .Z(n9171) );
  NBUFFX2 U9066 ( .INP(n9257), .Z(n9170) );
  NBUFFX2 U9067 ( .INP(n9257), .Z(n9169) );
  NBUFFX2 U9068 ( .INP(n9258), .Z(n9167) );
  NBUFFX2 U9069 ( .INP(n9258), .Z(n9166) );
  NBUFFX2 U9070 ( .INP(n9257), .Z(n9168) );
  NBUFFX2 U9071 ( .INP(n9257), .Z(n9172) );
  NBUFFX2 U9072 ( .INP(n9256), .Z(n9173) );
  NBUFFX2 U9073 ( .INP(n9256), .Z(n9174) );
  NBUFFX2 U9074 ( .INP(n9256), .Z(n9175) );
  NBUFFX2 U9075 ( .INP(n9256), .Z(n9176) );
  NBUFFX2 U9076 ( .INP(n9256), .Z(n9177) );
  NBUFFX2 U9077 ( .INP(n9255), .Z(n9178) );
  NBUFFX2 U9078 ( .INP(n9255), .Z(n9179) );
  NBUFFX2 U9079 ( .INP(n9255), .Z(n9180) );
  NBUFFX2 U9080 ( .INP(n9250), .Z(n9204) );
  NBUFFX2 U9081 ( .INP(n9251), .Z(n9198) );
  NBUFFX2 U9082 ( .INP(n9253), .Z(n9192) );
  NBUFFX2 U9083 ( .INP(n9252), .Z(n9193) );
  NBUFFX2 U9084 ( .INP(n9252), .Z(n9194) );
  NBUFFX2 U9085 ( .INP(n9258), .Z(n9165) );
  NBUFFX2 U9086 ( .INP(n9265), .Z(n9273) );
  NBUFFX2 U9087 ( .INP(n9270), .Z(n9288) );
  NBUFFX2 U9088 ( .INP(n9265), .Z(n9274) );
  NBUFFX2 U9089 ( .INP(n9265), .Z(n9275) );
  NBUFFX2 U9090 ( .INP(n9266), .Z(n9276) );
  NBUFFX2 U9091 ( .INP(n9266), .Z(n9277) );
  NBUFFX2 U9092 ( .INP(n9267), .Z(n9281) );
  NBUFFX2 U9093 ( .INP(n9268), .Z(n9282) );
  NBUFFX2 U9094 ( .INP(n9268), .Z(n9283) );
  NBUFFX2 U9095 ( .INP(n9268), .Z(n9284) );
  NBUFFX2 U9096 ( .INP(n9269), .Z(n9285) );
  NBUFFX2 U9097 ( .INP(n9269), .Z(n9286) );
  NBUFFX2 U9098 ( .INP(n9269), .Z(n9287) );
  NBUFFX2 U9099 ( .INP(n9266), .Z(n9278) );
  NBUFFX2 U9100 ( .INP(n9267), .Z(n9279) );
  NBUFFX2 U9101 ( .INP(n9267), .Z(n9280) );
  NBUFFX2 U9102 ( .INP(n9316), .Z(n9314) );
  NBUFFX2 U9103 ( .INP(n9320), .Z(n9292) );
  NBUFFX2 U9104 ( .INP(n9320), .Z(n9293) );
  NBUFFX2 U9105 ( .INP(n9320), .Z(n9294) );
  NBUFFX2 U9106 ( .INP(n9320), .Z(n9295) );
  NBUFFX2 U9107 ( .INP(n9318), .Z(n9302) );
  NBUFFX2 U9108 ( .INP(n9318), .Z(n9304) );
  NBUFFX2 U9109 ( .INP(n9318), .Z(n9305) );
  NBUFFX2 U9110 ( .INP(n9317), .Z(n9306) );
  NBUFFX2 U9111 ( .INP(n9317), .Z(n9307) );
  NBUFFX2 U9112 ( .INP(n9317), .Z(n9308) );
  NBUFFX2 U9113 ( .INP(n9319), .Z(n9296) );
  NBUFFX2 U9114 ( .INP(n9319), .Z(n9297) );
  NBUFFX2 U9115 ( .INP(n9318), .Z(n9303) );
  NBUFFX2 U9116 ( .INP(n9319), .Z(n9298) );
  NBUFFX2 U9117 ( .INP(n9319), .Z(n9299) );
  NBUFFX2 U9118 ( .INP(n9319), .Z(n9300) );
  NBUFFX2 U9119 ( .INP(n9318), .Z(n9301) );
  NBUFFX2 U9120 ( .INP(n9317), .Z(n9310) );
  NBUFFX2 U9121 ( .INP(n9317), .Z(n9309) );
  NBUFFX2 U9122 ( .INP(n9316), .Z(n9311) );
  NBUFFX2 U9123 ( .INP(n9316), .Z(n9312) );
  NBUFFX2 U9124 ( .INP(n9316), .Z(n9313) );
  NBUFFX2 U9125 ( .INP(n9243), .Z(n9242) );
  NBUFFX2 U9126 ( .INP(n9316), .Z(n9315) );
  NBUFFX2 U9127 ( .INP(n9943), .Z(n9774) );
  NBUFFX2 U9128 ( .INP(n9943), .Z(n9772) );
  NBUFFX2 U9129 ( .INP(n9943), .Z(n9773) );
  NBUFFX2 U9130 ( .INP(n9943), .Z(n9771) );
  NBUFFX2 U9131 ( .INP(n9918), .Z(n9896) );
  NBUFFX2 U9132 ( .INP(n9918), .Z(n9895) );
  NBUFFX2 U9133 ( .INP(n9919), .Z(n9894) );
  NBUFFX2 U9134 ( .INP(n9919), .Z(n9893) );
  NBUFFX2 U9135 ( .INP(n9919), .Z(n9892) );
  NBUFFX2 U9136 ( .INP(n9919), .Z(n9891) );
  NBUFFX2 U9137 ( .INP(n9919), .Z(n9890) );
  NBUFFX2 U9138 ( .INP(n9920), .Z(n9889) );
  NBUFFX2 U9139 ( .INP(n9920), .Z(n9888) );
  NBUFFX2 U9140 ( .INP(n9920), .Z(n9887) );
  NBUFFX2 U9141 ( .INP(n9920), .Z(n9886) );
  NBUFFX2 U9142 ( .INP(n9920), .Z(n9885) );
  NBUFFX2 U9143 ( .INP(n9921), .Z(n9882) );
  NBUFFX2 U9144 ( .INP(n9921), .Z(n9883) );
  NBUFFX2 U9145 ( .INP(n9921), .Z(n9884) );
  NBUFFX2 U9146 ( .INP(n9921), .Z(n9881) );
  NBUFFX2 U9147 ( .INP(n9918), .Z(n9898) );
  NBUFFX2 U9148 ( .INP(n9918), .Z(n9897) );
  NBUFFX2 U9149 ( .INP(n9921), .Z(n9880) );
  NBUFFX2 U9150 ( .INP(n9922), .Z(n9879) );
  NBUFFX2 U9151 ( .INP(n9922), .Z(n9878) );
  NBUFFX2 U9152 ( .INP(n9922), .Z(n9877) );
  NBUFFX2 U9153 ( .INP(n9922), .Z(n9876) );
  NBUFFX2 U9154 ( .INP(n9922), .Z(n9875) );
  NBUFFX2 U9155 ( .INP(n9923), .Z(n9874) );
  NBUFFX2 U9156 ( .INP(n9923), .Z(n9873) );
  NBUFFX2 U9157 ( .INP(n9923), .Z(n9872) );
  NBUFFX2 U9158 ( .INP(n9923), .Z(n9871) );
  NBUFFX2 U9159 ( .INP(n9924), .Z(n9868) );
  NBUFFX2 U9160 ( .INP(n9924), .Z(n9869) );
  NBUFFX2 U9161 ( .INP(n9923), .Z(n9870) );
  NBUFFX2 U9162 ( .INP(n9917), .Z(n9900) );
  NBUFFX2 U9163 ( .INP(n9918), .Z(n9899) );
  NBUFFX2 U9164 ( .INP(n9924), .Z(n9867) );
  NBUFFX2 U9165 ( .INP(n9924), .Z(n9866) );
  NBUFFX2 U9166 ( .INP(n9924), .Z(n9865) );
  NBUFFX2 U9167 ( .INP(n9925), .Z(n9864) );
  NBUFFX2 U9168 ( .INP(n9925), .Z(n9863) );
  NBUFFX2 U9169 ( .INP(n9925), .Z(n9862) );
  NBUFFX2 U9170 ( .INP(n9925), .Z(n9861) );
  NBUFFX2 U9171 ( .INP(n9925), .Z(n9860) );
  NBUFFX2 U9172 ( .INP(n9926), .Z(n9859) );
  NBUFFX2 U9173 ( .INP(n9926), .Z(n9858) );
  NBUFFX2 U9174 ( .INP(n9926), .Z(n9857) );
  NBUFFX2 U9175 ( .INP(n9926), .Z(n9856) );
  NBUFFX2 U9176 ( .INP(n9926), .Z(n9855) );
  NBUFFX2 U9177 ( .INP(n9927), .Z(n9854) );
  NBUFFX2 U9178 ( .INP(n9917), .Z(n9903) );
  NBUFFX2 U9179 ( .INP(n9917), .Z(n9902) );
  NBUFFX2 U9180 ( .INP(n9917), .Z(n9901) );
  NBUFFX2 U9181 ( .INP(n9927), .Z(n9853) );
  NBUFFX2 U9182 ( .INP(n9927), .Z(n9852) );
  NBUFFX2 U9183 ( .INP(n9927), .Z(n9851) );
  NBUFFX2 U9184 ( .INP(n9927), .Z(n9850) );
  NBUFFX2 U9185 ( .INP(n9928), .Z(n9849) );
  NBUFFX2 U9186 ( .INP(n9928), .Z(n9848) );
  NBUFFX2 U9187 ( .INP(n9928), .Z(n9847) );
  NBUFFX2 U9188 ( .INP(n9928), .Z(n9846) );
  NBUFFX2 U9189 ( .INP(n9928), .Z(n9845) );
  NBUFFX2 U9190 ( .INP(n9929), .Z(n9844) );
  NBUFFX2 U9191 ( .INP(n9929), .Z(n9841) );
  NBUFFX2 U9192 ( .INP(n9929), .Z(n9842) );
  NBUFFX2 U9193 ( .INP(n9929), .Z(n9843) );
  NBUFFX2 U9194 ( .INP(n9929), .Z(n9840) );
  NBUFFX2 U9195 ( .INP(n9917), .Z(n9904) );
  NBUFFX2 U9196 ( .INP(n9930), .Z(n9839) );
  NBUFFX2 U9197 ( .INP(n9930), .Z(n9838) );
  NBUFFX2 U9198 ( .INP(n9930), .Z(n9837) );
  NBUFFX2 U9199 ( .INP(n9930), .Z(n9836) );
  NBUFFX2 U9200 ( .INP(n9930), .Z(n9835) );
  NBUFFX2 U9201 ( .INP(n9931), .Z(n9834) );
  NBUFFX2 U9202 ( .INP(n9931), .Z(n9833) );
  NBUFFX2 U9203 ( .INP(n9931), .Z(n9832) );
  NBUFFX2 U9204 ( .INP(n9931), .Z(n9831) );
  NBUFFX2 U9205 ( .INP(n9931), .Z(n9830) );
  NBUFFX2 U9206 ( .INP(n9932), .Z(n9827) );
  NBUFFX2 U9207 ( .INP(n9932), .Z(n9828) );
  NBUFFX2 U9208 ( .INP(n9932), .Z(n9829) );
  NBUFFX2 U9209 ( .INP(n9916), .Z(n9907) );
  NBUFFX2 U9210 ( .INP(n9916), .Z(n9906) );
  NBUFFX2 U9211 ( .INP(n9916), .Z(n9905) );
  NBUFFX2 U9212 ( .INP(n9932), .Z(n9826) );
  NBUFFX2 U9213 ( .INP(n9932), .Z(n9825) );
  NBUFFX2 U9214 ( .INP(n9933), .Z(n9824) );
  NBUFFX2 U9215 ( .INP(n9933), .Z(n9823) );
  NBUFFX2 U9216 ( .INP(n9933), .Z(n9822) );
  NBUFFX2 U9217 ( .INP(n9933), .Z(n9821) );
  NBUFFX2 U9218 ( .INP(n9933), .Z(n9820) );
  NBUFFX2 U9219 ( .INP(n9934), .Z(n9819) );
  NBUFFX2 U9220 ( .INP(n9934), .Z(n9818) );
  NBUFFX2 U9221 ( .INP(n9934), .Z(n9817) );
  NBUFFX2 U9222 ( .INP(n9935), .Z(n9814) );
  NBUFFX2 U9223 ( .INP(n9934), .Z(n9815) );
  NBUFFX2 U9224 ( .INP(n9934), .Z(n9816) );
  NBUFFX2 U9225 ( .INP(n9935), .Z(n9813) );
  NBUFFX2 U9226 ( .INP(n9916), .Z(n9909) );
  NBUFFX2 U9227 ( .INP(n9916), .Z(n9908) );
  NBUFFX2 U9228 ( .INP(n9935), .Z(n9812) );
  NBUFFX2 U9229 ( .INP(n9935), .Z(n9811) );
  NBUFFX2 U9230 ( .INP(n9935), .Z(n9810) );
  NBUFFX2 U9231 ( .INP(n9936), .Z(n9809) );
  NBUFFX2 U9232 ( .INP(n9936), .Z(n9808) );
  NBUFFX2 U9233 ( .INP(n9936), .Z(n9807) );
  NBUFFX2 U9234 ( .INP(n9936), .Z(n9806) );
  NBUFFX2 U9235 ( .INP(n9936), .Z(n9805) );
  NBUFFX2 U9236 ( .INP(n9937), .Z(n9804) );
  NBUFFX2 U9237 ( .INP(n9937), .Z(n9803) );
  NBUFFX2 U9238 ( .INP(n9937), .Z(n9802) );
  NBUFFX2 U9239 ( .INP(n9938), .Z(n9799) );
  NBUFFX2 U9240 ( .INP(n9937), .Z(n9800) );
  NBUFFX2 U9241 ( .INP(n9937), .Z(n9801) );
  NBUFFX2 U9242 ( .INP(n9915), .Z(n9912) );
  NBUFFX2 U9243 ( .INP(n9915), .Z(n9911) );
  NBUFFX2 U9244 ( .INP(n9915), .Z(n9910) );
  NBUFFX2 U9245 ( .INP(n9938), .Z(n9798) );
  NBUFFX2 U9246 ( .INP(n9938), .Z(n9797) );
  NBUFFX2 U9247 ( .INP(n9938), .Z(n9796) );
  NBUFFX2 U9248 ( .INP(n9938), .Z(n9795) );
  NBUFFX2 U9249 ( .INP(n9939), .Z(n9794) );
  NBUFFX2 U9250 ( .INP(n9939), .Z(n9793) );
  NBUFFX2 U9251 ( .INP(n9939), .Z(n9792) );
  NBUFFX2 U9252 ( .INP(n9939), .Z(n9791) );
  NBUFFX2 U9253 ( .INP(n9939), .Z(n9790) );
  NBUFFX2 U9254 ( .INP(n9940), .Z(n9789) );
  NBUFFX2 U9255 ( .INP(n9940), .Z(n9788) );
  NBUFFX2 U9256 ( .INP(n9940), .Z(n9786) );
  NBUFFX2 U9257 ( .INP(n9940), .Z(n9787) );
  NBUFFX2 U9258 ( .INP(n9940), .Z(n9785) );
  NBUFFX2 U9259 ( .INP(n9915), .Z(n9914) );
  NBUFFX2 U9260 ( .INP(n9915), .Z(n9913) );
  NBUFFX2 U9261 ( .INP(n9941), .Z(n9784) );
  NBUFFX2 U9262 ( .INP(n9941), .Z(n9783) );
  NBUFFX2 U9263 ( .INP(n9941), .Z(n9782) );
  NBUFFX2 U9264 ( .INP(n9941), .Z(n9781) );
  NBUFFX2 U9265 ( .INP(n9941), .Z(n9780) );
  NBUFFX2 U9266 ( .INP(n9942), .Z(n9779) );
  NBUFFX2 U9267 ( .INP(n9942), .Z(n9778) );
  NBUFFX2 U9268 ( .INP(n9942), .Z(n9777) );
  NBUFFX2 U9269 ( .INP(n9942), .Z(n9776) );
  NBUFFX2 U9270 ( .INP(n9942), .Z(n9775) );
  NBUFFX2 U9271 ( .INP(n9270), .Z(n9289) );
  NBUFFX2 U9272 ( .INP(n9264), .Z(n9137) );
  NBUFFX2 U9273 ( .INP(n9264), .Z(n9136) );
  NBUFFX2 U9274 ( .INP(n9272), .Z(n9265) );
  NBUFFX2 U9275 ( .INP(n9271), .Z(n9268) );
  NBUFFX2 U9276 ( .INP(n9271), .Z(n9269) );
  NBUFFX2 U9277 ( .INP(n9272), .Z(n9266) );
  NBUFFX2 U9278 ( .INP(n9272), .Z(n9267) );
  NBUFFX2 U9279 ( .INP(n9271), .Z(n9270) );
  NBUFFX2 U9280 ( .INP(n9113), .Z(n9117) );
  NBUFFX2 U9281 ( .INP(n9113), .Z(n9116) );
  NBUFFX2 U9282 ( .INP(n9113), .Z(n9118) );
  NBUFFX2 U9283 ( .INP(n9114), .Z(n9120) );
  NBUFFX2 U9284 ( .INP(n9114), .Z(n9119) );
  NBUFFX2 U9285 ( .INP(n9115), .Z(n9122) );
  NBUFFX2 U9286 ( .INP(n9115), .Z(n9123) );
  NBUFFX2 U9287 ( .INP(n9114), .Z(n9121) );
  NBUFFX2 U9288 ( .INP(n9085), .Z(n9092) );
  NBUFFX2 U9289 ( .INP(n9089), .Z(n9111) );
  NBUFFX2 U9290 ( .INP(n9089), .Z(n9110) );
  NBUFFX2 U9291 ( .INP(n9085), .Z(n9090) );
  NBUFFX2 U9292 ( .INP(n9085), .Z(n9091) );
  NBUFFX2 U9293 ( .INP(n9088), .Z(n9108) );
  NBUFFX2 U9294 ( .INP(n9088), .Z(n9106) );
  NBUFFX2 U9295 ( .INP(n9087), .Z(n9104) );
  NBUFFX2 U9296 ( .INP(n9087), .Z(n9103) );
  NBUFFX2 U9297 ( .INP(n9087), .Z(n9102) );
  NBUFFX2 U9298 ( .INP(n9087), .Z(n9101) );
  NBUFFX2 U9299 ( .INP(n9087), .Z(n9100) );
  NBUFFX2 U9300 ( .INP(n9086), .Z(n9099) );
  NBUFFX2 U9301 ( .INP(n9086), .Z(n9098) );
  NBUFFX2 U9302 ( .INP(n9086), .Z(n9097) );
  NBUFFX2 U9303 ( .INP(n9086), .Z(n9096) );
  NBUFFX2 U9304 ( .INP(n9088), .Z(n9107) );
  NBUFFX2 U9305 ( .INP(n9088), .Z(n9109) );
  NBUFFX2 U9306 ( .INP(n9088), .Z(n9105) );
  NBUFFX2 U9307 ( .INP(n9085), .Z(n9093) );
  NBUFFX2 U9308 ( .INP(n9085), .Z(n9094) );
  NBUFFX2 U9309 ( .INP(n9086), .Z(n9095) );
  NBUFFX2 U9310 ( .INP(n9115), .Z(n9124) );
  NBUFFX2 U9311 ( .INP(n9089), .Z(n9112) );
  NBUFFX2 U9312 ( .INP(n2148), .Z(n9271) );
  NBUFFX2 U9313 ( .INP(n2148), .Z(n9272) );
  NBUFFX2 U9314 ( .INP(n10633), .Z(n9115) );
  NBUFFX2 U9315 ( .INP(n10633), .Z(n9113) );
  NBUFFX2 U9316 ( .INP(n10633), .Z(n9114) );
  INVX0 U9317 ( .INP(n2153), .ZN(n9337) );
  NBUFFX2 U9318 ( .INP(n9958), .Z(n9085) );
  NBUFFX2 U9319 ( .INP(n9958), .Z(n9086) );
  NBUFFX2 U9320 ( .INP(n9958), .Z(n9087) );
  NBUFFX2 U9321 ( .INP(n9958), .Z(n9088) );
  NBUFFX2 U9322 ( .INP(n9958), .Z(n9089) );
  NBUFFX2 U9323 ( .INP(n9135), .Z(n9125) );
  NBUFFX2 U9324 ( .INP(n9135), .Z(n9126) );
  NBUFFX2 U9325 ( .INP(n9134), .Z(n9127) );
  NBUFFX2 U9326 ( .INP(n9134), .Z(n9128) );
  NBUFFX2 U9327 ( .INP(n9134), .Z(n9129) );
  NBUFFX2 U9328 ( .INP(n9133), .Z(n9130) );
  NBUFFX2 U9329 ( .INP(n9133), .Z(n9131) );
  NBUFFX2 U9330 ( .INP(n9133), .Z(n9132) );
  NBUFFX2 U9331 ( .INP(n2182), .Z(n9133) );
  NBUFFX2 U9332 ( .INP(n2182), .Z(n9134) );
  NBUFFX2 U9333 ( .INP(n2182), .Z(n9135) );
  NBUFFX2 U9334 ( .INP(n9125), .Z(n9243) );
  NBUFFX2 U9335 ( .INP(n9125), .Z(n9244) );
  NBUFFX2 U9336 ( .INP(n9125), .Z(n9245) );
  NBUFFX2 U9337 ( .INP(n9126), .Z(n9246) );
  NBUFFX2 U9338 ( .INP(n9126), .Z(n9247) );
  NBUFFX2 U9339 ( .INP(n9126), .Z(n9248) );
  NBUFFX2 U9340 ( .INP(n9127), .Z(n9249) );
  NBUFFX2 U9341 ( .INP(n9127), .Z(n9250) );
  NBUFFX2 U9342 ( .INP(n9127), .Z(n9251) );
  NBUFFX2 U9343 ( .INP(n9128), .Z(n9252) );
  NBUFFX2 U9344 ( .INP(n9128), .Z(n9253) );
  NBUFFX2 U9345 ( .INP(n9128), .Z(n9254) );
  NBUFFX2 U9346 ( .INP(n9129), .Z(n9255) );
  NBUFFX2 U9347 ( .INP(n9129), .Z(n9256) );
  NBUFFX2 U9348 ( .INP(n9129), .Z(n9257) );
  NBUFFX2 U9349 ( .INP(n9130), .Z(n9258) );
  NBUFFX2 U9350 ( .INP(n9130), .Z(n9259) );
  NBUFFX2 U9351 ( .INP(n9130), .Z(n9260) );
  NBUFFX2 U9352 ( .INP(n9131), .Z(n9261) );
  NBUFFX2 U9353 ( .INP(n9131), .Z(n9262) );
  NBUFFX2 U9354 ( .INP(n9131), .Z(n9263) );
  NBUFFX2 U9355 ( .INP(n9132), .Z(n9264) );
  NBUFFX2 U9356 ( .INP(n2152), .Z(n9290) );
  NBUFFX2 U9357 ( .INP(n2152), .Z(n9291) );
  NBUFFX2 U9358 ( .INP(n9290), .Z(n9316) );
  NBUFFX2 U9359 ( .INP(n9290), .Z(n9317) );
  NBUFFX2 U9360 ( .INP(n9290), .Z(n9318) );
  NBUFFX2 U9361 ( .INP(n9291), .Z(n9319) );
  NBUFFX2 U9362 ( .INP(n9291), .Z(n9320) );
  INVX0 U9363 ( .INP(n9337), .ZN(n9321) );
  INVX0 U9364 ( .INP(n9337), .ZN(n9322) );
  INVX0 U9365 ( .INP(n9337), .ZN(n9323) );
  INVX0 U9366 ( .INP(n9337), .ZN(n9324) );
  INVX0 U9367 ( .INP(n9337), .ZN(n9325) );
  INVX0 U9368 ( .INP(n9337), .ZN(n9326) );
  INVX0 U9369 ( .INP(n9337), .ZN(n9327) );
  INVX0 U9370 ( .INP(n9337), .ZN(n9328) );
  INVX0 U9371 ( .INP(n9337), .ZN(n9329) );
  INVX0 U9372 ( .INP(n9337), .ZN(n9330) );
  INVX0 U9373 ( .INP(n9337), .ZN(n9331) );
  INVX0 U9374 ( .INP(n9337), .ZN(n9332) );
  INVX0 U9375 ( .INP(n9337), .ZN(n9333) );
  INVX0 U9376 ( .INP(n9337), .ZN(n9334) );
  INVX0 U9377 ( .INP(n9337), .ZN(n9335) );
  INVX0 U9378 ( .INP(n9337), .ZN(n9336) );
  NBUFFX2 U9379 ( .INP(n9722), .Z(n9338) );
  NBUFFX2 U9380 ( .INP(n9721), .Z(n9339) );
  NBUFFX2 U9381 ( .INP(n9721), .Z(n9340) );
  NBUFFX2 U9382 ( .INP(n9721), .Z(n9341) );
  NBUFFX2 U9383 ( .INP(n9720), .Z(n9342) );
  NBUFFX2 U9384 ( .INP(n9720), .Z(n9343) );
  NBUFFX2 U9385 ( .INP(n9720), .Z(n9344) );
  NBUFFX2 U9386 ( .INP(n9719), .Z(n9345) );
  NBUFFX2 U9387 ( .INP(n9719), .Z(n9346) );
  NBUFFX2 U9388 ( .INP(n9719), .Z(n9347) );
  NBUFFX2 U9389 ( .INP(n9718), .Z(n9348) );
  NBUFFX2 U9390 ( .INP(n9718), .Z(n9349) );
  NBUFFX2 U9391 ( .INP(n9718), .Z(n9350) );
  NBUFFX2 U9392 ( .INP(n9717), .Z(n9351) );
  NBUFFX2 U9393 ( .INP(n9717), .Z(n9352) );
  NBUFFX2 U9394 ( .INP(n9717), .Z(n9353) );
  NBUFFX2 U9395 ( .INP(n9716), .Z(n9354) );
  NBUFFX2 U9396 ( .INP(n9716), .Z(n9355) );
  NBUFFX2 U9397 ( .INP(n9716), .Z(n9356) );
  NBUFFX2 U9398 ( .INP(n9715), .Z(n9357) );
  NBUFFX2 U9399 ( .INP(n9715), .Z(n9358) );
  NBUFFX2 U9400 ( .INP(n9715), .Z(n9359) );
  NBUFFX2 U9401 ( .INP(n9714), .Z(n9360) );
  NBUFFX2 U9402 ( .INP(n9714), .Z(n9361) );
  NBUFFX2 U9403 ( .INP(n9714), .Z(n9362) );
  NBUFFX2 U9404 ( .INP(n9713), .Z(n9363) );
  NBUFFX2 U9405 ( .INP(n9713), .Z(n9364) );
  NBUFFX2 U9406 ( .INP(n9713), .Z(n9365) );
  NBUFFX2 U9407 ( .INP(n9712), .Z(n9366) );
  NBUFFX2 U9408 ( .INP(n9712), .Z(n9367) );
  NBUFFX2 U9409 ( .INP(n9712), .Z(n9368) );
  NBUFFX2 U9410 ( .INP(n9711), .Z(n9369) );
  NBUFFX2 U9411 ( .INP(n9711), .Z(n9370) );
  NBUFFX2 U9412 ( .INP(n9711), .Z(n9371) );
  NBUFFX2 U9413 ( .INP(n9710), .Z(n9372) );
  NBUFFX2 U9414 ( .INP(n9710), .Z(n9373) );
  NBUFFX2 U9415 ( .INP(n9710), .Z(n9374) );
  NBUFFX2 U9416 ( .INP(n9709), .Z(n9375) );
  NBUFFX2 U9417 ( .INP(n9709), .Z(n9376) );
  NBUFFX2 U9418 ( .INP(n9709), .Z(n9377) );
  NBUFFX2 U9419 ( .INP(n9708), .Z(n9378) );
  NBUFFX2 U9420 ( .INP(n9708), .Z(n9379) );
  NBUFFX2 U9421 ( .INP(n9708), .Z(n9380) );
  NBUFFX2 U9422 ( .INP(n9707), .Z(n9381) );
  NBUFFX2 U9423 ( .INP(n9707), .Z(n9382) );
  NBUFFX2 U9424 ( .INP(n9707), .Z(n9383) );
  NBUFFX2 U9425 ( .INP(n9706), .Z(n9384) );
  NBUFFX2 U9426 ( .INP(n9706), .Z(n9385) );
  NBUFFX2 U9427 ( .INP(n9706), .Z(n9386) );
  NBUFFX2 U9428 ( .INP(n9705), .Z(n9387) );
  NBUFFX2 U9429 ( .INP(n9705), .Z(n9388) );
  NBUFFX2 U9430 ( .INP(n9705), .Z(n9389) );
  NBUFFX2 U9431 ( .INP(n9704), .Z(n9390) );
  NBUFFX2 U9432 ( .INP(n9704), .Z(n9391) );
  NBUFFX2 U9433 ( .INP(n9704), .Z(n9392) );
  NBUFFX2 U9434 ( .INP(n9703), .Z(n9393) );
  NBUFFX2 U9435 ( .INP(n9703), .Z(n9394) );
  NBUFFX2 U9436 ( .INP(n9703), .Z(n9395) );
  NBUFFX2 U9437 ( .INP(n9702), .Z(n9396) );
  NBUFFX2 U9438 ( .INP(n9702), .Z(n9397) );
  NBUFFX2 U9439 ( .INP(n9702), .Z(n9398) );
  NBUFFX2 U9440 ( .INP(n9701), .Z(n9399) );
  NBUFFX2 U9441 ( .INP(n9701), .Z(n9400) );
  NBUFFX2 U9442 ( .INP(n9701), .Z(n9401) );
  NBUFFX2 U9443 ( .INP(n9700), .Z(n9402) );
  NBUFFX2 U9444 ( .INP(n9700), .Z(n9403) );
  NBUFFX2 U9445 ( .INP(n9700), .Z(n9404) );
  NBUFFX2 U9446 ( .INP(n9699), .Z(n9405) );
  NBUFFX2 U9447 ( .INP(n9699), .Z(n9406) );
  NBUFFX2 U9448 ( .INP(n9699), .Z(n9407) );
  NBUFFX2 U9449 ( .INP(n9698), .Z(n9408) );
  NBUFFX2 U9450 ( .INP(n9698), .Z(n9409) );
  NBUFFX2 U9451 ( .INP(n9698), .Z(n9410) );
  NBUFFX2 U9452 ( .INP(n9697), .Z(n9411) );
  NBUFFX2 U9453 ( .INP(n9697), .Z(n9412) );
  NBUFFX2 U9454 ( .INP(n9697), .Z(n9413) );
  NBUFFX2 U9455 ( .INP(n9696), .Z(n9414) );
  NBUFFX2 U9456 ( .INP(n9696), .Z(n9415) );
  NBUFFX2 U9457 ( .INP(n9696), .Z(n9416) );
  NBUFFX2 U9458 ( .INP(n9695), .Z(n9417) );
  NBUFFX2 U9459 ( .INP(n9695), .Z(n9418) );
  NBUFFX2 U9460 ( .INP(n9695), .Z(n9419) );
  NBUFFX2 U9461 ( .INP(n9694), .Z(n9420) );
  NBUFFX2 U9462 ( .INP(n9694), .Z(n9421) );
  NBUFFX2 U9463 ( .INP(n9694), .Z(n9422) );
  NBUFFX2 U9464 ( .INP(n9693), .Z(n9423) );
  NBUFFX2 U9465 ( .INP(n9693), .Z(n9424) );
  NBUFFX2 U9466 ( .INP(n9693), .Z(n9425) );
  NBUFFX2 U9467 ( .INP(n9692), .Z(n9426) );
  NBUFFX2 U9468 ( .INP(n9692), .Z(n9427) );
  NBUFFX2 U9469 ( .INP(n9692), .Z(n9428) );
  NBUFFX2 U9470 ( .INP(n9691), .Z(n9429) );
  NBUFFX2 U9471 ( .INP(n9691), .Z(n9430) );
  NBUFFX2 U9472 ( .INP(n9691), .Z(n9431) );
  NBUFFX2 U9473 ( .INP(n9690), .Z(n9432) );
  NBUFFX2 U9474 ( .INP(n9690), .Z(n9433) );
  NBUFFX2 U9475 ( .INP(n9690), .Z(n9434) );
  NBUFFX2 U9476 ( .INP(n9689), .Z(n9435) );
  NBUFFX2 U9477 ( .INP(n9689), .Z(n9436) );
  NBUFFX2 U9478 ( .INP(n9689), .Z(n9437) );
  NBUFFX2 U9479 ( .INP(n9688), .Z(n9438) );
  NBUFFX2 U9480 ( .INP(n9688), .Z(n9439) );
  NBUFFX2 U9481 ( .INP(n9688), .Z(n9440) );
  NBUFFX2 U9482 ( .INP(n9687), .Z(n9441) );
  NBUFFX2 U9483 ( .INP(n9687), .Z(n9442) );
  NBUFFX2 U9484 ( .INP(n9687), .Z(n9443) );
  NBUFFX2 U9485 ( .INP(n9686), .Z(n9444) );
  NBUFFX2 U9486 ( .INP(n9686), .Z(n9445) );
  NBUFFX2 U9487 ( .INP(n9686), .Z(n9446) );
  NBUFFX2 U9488 ( .INP(n9685), .Z(n9447) );
  NBUFFX2 U9489 ( .INP(n9685), .Z(n9448) );
  NBUFFX2 U9490 ( .INP(n9685), .Z(n9449) );
  NBUFFX2 U9491 ( .INP(n9684), .Z(n9450) );
  NBUFFX2 U9492 ( .INP(n9684), .Z(n9451) );
  NBUFFX2 U9493 ( .INP(n9684), .Z(n9452) );
  NBUFFX2 U9494 ( .INP(n9683), .Z(n9453) );
  NBUFFX2 U9495 ( .INP(n9683), .Z(n9454) );
  NBUFFX2 U9496 ( .INP(n9683), .Z(n9455) );
  NBUFFX2 U9497 ( .INP(n9682), .Z(n9456) );
  NBUFFX2 U9498 ( .INP(n9682), .Z(n9457) );
  NBUFFX2 U9499 ( .INP(n9682), .Z(n9458) );
  NBUFFX2 U9500 ( .INP(n9681), .Z(n9459) );
  NBUFFX2 U9501 ( .INP(n9681), .Z(n9460) );
  NBUFFX2 U9502 ( .INP(n9681), .Z(n9461) );
  NBUFFX2 U9503 ( .INP(n9680), .Z(n9462) );
  NBUFFX2 U9504 ( .INP(n9680), .Z(n9463) );
  NBUFFX2 U9505 ( .INP(n9680), .Z(n9464) );
  NBUFFX2 U9506 ( .INP(n9679), .Z(n9465) );
  NBUFFX2 U9507 ( .INP(n9679), .Z(n9466) );
  NBUFFX2 U9508 ( .INP(n9679), .Z(n9467) );
  NBUFFX2 U9509 ( .INP(n9678), .Z(n9468) );
  NBUFFX2 U9510 ( .INP(n9678), .Z(n9469) );
  NBUFFX2 U9511 ( .INP(n9678), .Z(n9470) );
  NBUFFX2 U9512 ( .INP(n9677), .Z(n9471) );
  NBUFFX2 U9513 ( .INP(n9677), .Z(n9472) );
  NBUFFX2 U9514 ( .INP(n9677), .Z(n9473) );
  NBUFFX2 U9515 ( .INP(n9676), .Z(n9474) );
  NBUFFX2 U9516 ( .INP(n9676), .Z(n9475) );
  NBUFFX2 U9517 ( .INP(n9676), .Z(n9476) );
  NBUFFX2 U9518 ( .INP(n9675), .Z(n9477) );
  NBUFFX2 U9519 ( .INP(n9675), .Z(n9478) );
  NBUFFX2 U9520 ( .INP(n9675), .Z(n9479) );
  NBUFFX2 U9521 ( .INP(n9674), .Z(n9480) );
  NBUFFX2 U9522 ( .INP(n9674), .Z(n9481) );
  NBUFFX2 U9523 ( .INP(n9674), .Z(n9482) );
  NBUFFX2 U9524 ( .INP(n9673), .Z(n9483) );
  NBUFFX2 U9525 ( .INP(n9673), .Z(n9484) );
  NBUFFX2 U9526 ( .INP(n9673), .Z(n9485) );
  NBUFFX2 U9527 ( .INP(n9672), .Z(n9486) );
  NBUFFX2 U9528 ( .INP(n9672), .Z(n9487) );
  NBUFFX2 U9529 ( .INP(n9672), .Z(n9488) );
  NBUFFX2 U9530 ( .INP(n9671), .Z(n9489) );
  NBUFFX2 U9531 ( .INP(n9671), .Z(n9490) );
  NBUFFX2 U9532 ( .INP(n9671), .Z(n9491) );
  NBUFFX2 U9533 ( .INP(n9670), .Z(n9492) );
  NBUFFX2 U9534 ( .INP(n9670), .Z(n9493) );
  NBUFFX2 U9535 ( .INP(n9670), .Z(n9494) );
  NBUFFX2 U9536 ( .INP(n9669), .Z(n9495) );
  NBUFFX2 U9537 ( .INP(n9669), .Z(n9496) );
  NBUFFX2 U9538 ( .INP(n9669), .Z(n9497) );
  NBUFFX2 U9539 ( .INP(n9668), .Z(n9498) );
  NBUFFX2 U9540 ( .INP(n9668), .Z(n9499) );
  NBUFFX2 U9541 ( .INP(n9668), .Z(n9500) );
  NBUFFX2 U9542 ( .INP(n9667), .Z(n9501) );
  NBUFFX2 U9543 ( .INP(n9667), .Z(n9502) );
  NBUFFX2 U9544 ( .INP(n9667), .Z(n9503) );
  NBUFFX2 U9545 ( .INP(n9666), .Z(n9504) );
  NBUFFX2 U9546 ( .INP(n9666), .Z(n9505) );
  NBUFFX2 U9547 ( .INP(n9666), .Z(n9506) );
  NBUFFX2 U9548 ( .INP(n9665), .Z(n9507) );
  NBUFFX2 U9549 ( .INP(n9665), .Z(n9508) );
  NBUFFX2 U9550 ( .INP(n9665), .Z(n9509) );
  NBUFFX2 U9551 ( .INP(n9664), .Z(n9510) );
  NBUFFX2 U9552 ( .INP(n9664), .Z(n9511) );
  NBUFFX2 U9553 ( .INP(n9664), .Z(n9512) );
  NBUFFX2 U9554 ( .INP(n9663), .Z(n9513) );
  NBUFFX2 U9555 ( .INP(n9663), .Z(n9514) );
  NBUFFX2 U9556 ( .INP(n9663), .Z(n9515) );
  NBUFFX2 U9557 ( .INP(n9662), .Z(n9516) );
  NBUFFX2 U9558 ( .INP(n9662), .Z(n9517) );
  NBUFFX2 U9559 ( .INP(n9662), .Z(n9518) );
  NBUFFX2 U9560 ( .INP(n9661), .Z(n9519) );
  NBUFFX2 U9561 ( .INP(n9661), .Z(n9520) );
  NBUFFX2 U9562 ( .INP(n9661), .Z(n9521) );
  NBUFFX2 U9563 ( .INP(n9660), .Z(n9522) );
  NBUFFX2 U9564 ( .INP(n9660), .Z(n9523) );
  NBUFFX2 U9565 ( .INP(n9660), .Z(n9524) );
  NBUFFX2 U9566 ( .INP(n9659), .Z(n9525) );
  NBUFFX2 U9567 ( .INP(n9659), .Z(n9526) );
  NBUFFX2 U9568 ( .INP(n9659), .Z(n9527) );
  NBUFFX2 U9569 ( .INP(n9658), .Z(n9528) );
  NBUFFX2 U9570 ( .INP(n9658), .Z(n9529) );
  NBUFFX2 U9571 ( .INP(n9658), .Z(n9530) );
  NBUFFX2 U9572 ( .INP(n9657), .Z(n9531) );
  NBUFFX2 U9573 ( .INP(n9657), .Z(n9532) );
  NBUFFX2 U9574 ( .INP(n9657), .Z(n9533) );
  NBUFFX2 U9575 ( .INP(n9656), .Z(n9534) );
  NBUFFX2 U9576 ( .INP(n9656), .Z(n9535) );
  NBUFFX2 U9577 ( .INP(n9656), .Z(n9536) );
  NBUFFX2 U9578 ( .INP(n9655), .Z(n9537) );
  NBUFFX2 U9579 ( .INP(n9655), .Z(n9538) );
  NBUFFX2 U9580 ( .INP(n9655), .Z(n9539) );
  NBUFFX2 U9581 ( .INP(n9654), .Z(n9540) );
  NBUFFX2 U9582 ( .INP(n9654), .Z(n9541) );
  NBUFFX2 U9583 ( .INP(n9654), .Z(n9542) );
  NBUFFX2 U9584 ( .INP(n9653), .Z(n9543) );
  NBUFFX2 U9585 ( .INP(n9653), .Z(n9544) );
  NBUFFX2 U9586 ( .INP(n9653), .Z(n9545) );
  NBUFFX2 U9587 ( .INP(n9652), .Z(n9546) );
  NBUFFX2 U9588 ( .INP(n9652), .Z(n9547) );
  NBUFFX2 U9589 ( .INP(n9652), .Z(n9548) );
  NBUFFX2 U9590 ( .INP(n9651), .Z(n9549) );
  NBUFFX2 U9591 ( .INP(n9651), .Z(n9550) );
  NBUFFX2 U9592 ( .INP(n9651), .Z(n9551) );
  NBUFFX2 U9593 ( .INP(n9650), .Z(n9552) );
  NBUFFX2 U9594 ( .INP(n9650), .Z(n9553) );
  NBUFFX2 U9595 ( .INP(n9650), .Z(n9554) );
  NBUFFX2 U9596 ( .INP(n9649), .Z(n9555) );
  NBUFFX2 U9597 ( .INP(n9649), .Z(n9556) );
  NBUFFX2 U9598 ( .INP(n9649), .Z(n9557) );
  NBUFFX2 U9599 ( .INP(n9648), .Z(n9558) );
  NBUFFX2 U9600 ( .INP(n9648), .Z(n9559) );
  NBUFFX2 U9601 ( .INP(n9648), .Z(n9560) );
  NBUFFX2 U9602 ( .INP(n9647), .Z(n9561) );
  NBUFFX2 U9603 ( .INP(n9647), .Z(n9562) );
  NBUFFX2 U9604 ( .INP(n9647), .Z(n9563) );
  NBUFFX2 U9605 ( .INP(n9646), .Z(n9564) );
  NBUFFX2 U9606 ( .INP(n9646), .Z(n9565) );
  NBUFFX2 U9607 ( .INP(n9646), .Z(n9566) );
  NBUFFX2 U9608 ( .INP(n9645), .Z(n9567) );
  NBUFFX2 U9609 ( .INP(n9645), .Z(n9568) );
  NBUFFX2 U9610 ( .INP(n9645), .Z(n9569) );
  NBUFFX2 U9611 ( .INP(n9644), .Z(n9570) );
  NBUFFX2 U9612 ( .INP(n9644), .Z(n9571) );
  NBUFFX2 U9613 ( .INP(n9644), .Z(n9572) );
  NBUFFX2 U9614 ( .INP(n9643), .Z(n9573) );
  NBUFFX2 U9615 ( .INP(n9643), .Z(n9574) );
  NBUFFX2 U9616 ( .INP(n9643), .Z(n9575) );
  NBUFFX2 U9617 ( .INP(n9642), .Z(n9576) );
  NBUFFX2 U9618 ( .INP(n9642), .Z(n9577) );
  NBUFFX2 U9619 ( .INP(n9642), .Z(n9578) );
  NBUFFX2 U9620 ( .INP(n9641), .Z(n9579) );
  NBUFFX2 U9621 ( .INP(n9641), .Z(n9580) );
  NBUFFX2 U9622 ( .INP(n9641), .Z(n9581) );
  NBUFFX2 U9623 ( .INP(n9640), .Z(n9582) );
  NBUFFX2 U9624 ( .INP(n9640), .Z(n9583) );
  NBUFFX2 U9625 ( .INP(n9640), .Z(n9584) );
  NBUFFX2 U9626 ( .INP(n9639), .Z(n9585) );
  NBUFFX2 U9627 ( .INP(n9639), .Z(n9586) );
  NBUFFX2 U9628 ( .INP(n9639), .Z(n9587) );
  NBUFFX2 U9629 ( .INP(n9638), .Z(n9588) );
  NBUFFX2 U9630 ( .INP(n9638), .Z(n9589) );
  NBUFFX2 U9631 ( .INP(n9638), .Z(n9590) );
  NBUFFX2 U9632 ( .INP(n9637), .Z(n9591) );
  NBUFFX2 U9633 ( .INP(n9637), .Z(n9592) );
  NBUFFX2 U9634 ( .INP(n9637), .Z(n9593) );
  NBUFFX2 U9635 ( .INP(n9636), .Z(n9594) );
  NBUFFX2 U9636 ( .INP(n9636), .Z(n9595) );
  NBUFFX2 U9637 ( .INP(n9636), .Z(n9596) );
  NBUFFX2 U9638 ( .INP(n9635), .Z(n9597) );
  NBUFFX2 U9639 ( .INP(n9635), .Z(n9598) );
  NBUFFX2 U9640 ( .INP(n9635), .Z(n9599) );
  NBUFFX2 U9641 ( .INP(n9634), .Z(n9600) );
  NBUFFX2 U9642 ( .INP(n9634), .Z(n9601) );
  NBUFFX2 U9643 ( .INP(n9634), .Z(n9602) );
  NBUFFX2 U9644 ( .INP(n9633), .Z(n9603) );
  NBUFFX2 U9645 ( .INP(n9633), .Z(n9604) );
  NBUFFX2 U9646 ( .INP(n9633), .Z(n9605) );
  NBUFFX2 U9647 ( .INP(n9632), .Z(n9606) );
  NBUFFX2 U9648 ( .INP(n9632), .Z(n9607) );
  NBUFFX2 U9649 ( .INP(n9632), .Z(n9608) );
  NBUFFX2 U9650 ( .INP(n9631), .Z(n9609) );
  NBUFFX2 U9651 ( .INP(n9631), .Z(n9610) );
  NBUFFX2 U9652 ( .INP(n9631), .Z(n9611) );
  NBUFFX2 U9653 ( .INP(n9630), .Z(n9612) );
  NBUFFX2 U9654 ( .INP(n9630), .Z(n9613) );
  NBUFFX2 U9655 ( .INP(n9630), .Z(n9614) );
  NBUFFX2 U9656 ( .INP(n9629), .Z(n9615) );
  NBUFFX2 U9657 ( .INP(n9629), .Z(n9616) );
  NBUFFX2 U9658 ( .INP(n9629), .Z(n9617) );
  NBUFFX2 U9659 ( .INP(n9628), .Z(n9618) );
  NBUFFX2 U9660 ( .INP(n9628), .Z(n9619) );
  NBUFFX2 U9661 ( .INP(n9628), .Z(n9620) );
  NBUFFX2 U9662 ( .INP(n9627), .Z(n9621) );
  NBUFFX2 U9663 ( .INP(n9627), .Z(n9622) );
  NBUFFX2 U9664 ( .INP(n9627), .Z(n9623) );
  NBUFFX2 U9665 ( .INP(n9626), .Z(n9624) );
  NBUFFX2 U9666 ( .INP(n9626), .Z(n9625) );
  NBUFFX2 U9667 ( .INP(n9755), .Z(n9626) );
  NBUFFX2 U9668 ( .INP(n9754), .Z(n9627) );
  NBUFFX2 U9669 ( .INP(n9754), .Z(n9628) );
  NBUFFX2 U9670 ( .INP(n9754), .Z(n9629) );
  NBUFFX2 U9671 ( .INP(n9753), .Z(n9630) );
  NBUFFX2 U9672 ( .INP(n9753), .Z(n9631) );
  NBUFFX2 U9673 ( .INP(n9753), .Z(n9632) );
  NBUFFX2 U9674 ( .INP(n9752), .Z(n9633) );
  NBUFFX2 U9675 ( .INP(n9752), .Z(n9634) );
  NBUFFX2 U9676 ( .INP(n9752), .Z(n9635) );
  NBUFFX2 U9677 ( .INP(n9751), .Z(n9636) );
  NBUFFX2 U9678 ( .INP(n9751), .Z(n9637) );
  NBUFFX2 U9679 ( .INP(n9751), .Z(n9638) );
  NBUFFX2 U9680 ( .INP(n9750), .Z(n9639) );
  NBUFFX2 U9681 ( .INP(n9750), .Z(n9640) );
  NBUFFX2 U9682 ( .INP(n9750), .Z(n9641) );
  NBUFFX2 U9683 ( .INP(n9749), .Z(n9642) );
  NBUFFX2 U9684 ( .INP(n9749), .Z(n9643) );
  NBUFFX2 U9685 ( .INP(n9749), .Z(n9644) );
  NBUFFX2 U9686 ( .INP(n9748), .Z(n9645) );
  NBUFFX2 U9687 ( .INP(n9748), .Z(n9646) );
  NBUFFX2 U9688 ( .INP(n9748), .Z(n9647) );
  NBUFFX2 U9689 ( .INP(n9747), .Z(n9648) );
  NBUFFX2 U9690 ( .INP(n9747), .Z(n9649) );
  NBUFFX2 U9691 ( .INP(n9747), .Z(n9650) );
  NBUFFX2 U9692 ( .INP(n9746), .Z(n9651) );
  NBUFFX2 U9693 ( .INP(n9746), .Z(n9652) );
  NBUFFX2 U9694 ( .INP(n9746), .Z(n9653) );
  NBUFFX2 U9695 ( .INP(n9745), .Z(n9654) );
  NBUFFX2 U9696 ( .INP(n9745), .Z(n9655) );
  NBUFFX2 U9697 ( .INP(n9745), .Z(n9656) );
  NBUFFX2 U9698 ( .INP(n9744), .Z(n9657) );
  NBUFFX2 U9699 ( .INP(n9744), .Z(n9658) );
  NBUFFX2 U9700 ( .INP(n9744), .Z(n9659) );
  NBUFFX2 U9701 ( .INP(n9743), .Z(n9660) );
  NBUFFX2 U9702 ( .INP(n9743), .Z(n9661) );
  NBUFFX2 U9703 ( .INP(n9743), .Z(n9662) );
  NBUFFX2 U9704 ( .INP(n9742), .Z(n9663) );
  NBUFFX2 U9705 ( .INP(n9742), .Z(n9664) );
  NBUFFX2 U9706 ( .INP(n9742), .Z(n9665) );
  NBUFFX2 U9707 ( .INP(n9741), .Z(n9666) );
  NBUFFX2 U9708 ( .INP(n9741), .Z(n9667) );
  NBUFFX2 U9709 ( .INP(n9741), .Z(n9668) );
  NBUFFX2 U9710 ( .INP(n9740), .Z(n9669) );
  NBUFFX2 U9711 ( .INP(n9740), .Z(n9670) );
  NBUFFX2 U9712 ( .INP(n9740), .Z(n9671) );
  NBUFFX2 U9713 ( .INP(n9739), .Z(n9672) );
  NBUFFX2 U9714 ( .INP(n9739), .Z(n9673) );
  NBUFFX2 U9715 ( .INP(n9739), .Z(n9674) );
  NBUFFX2 U9716 ( .INP(n9738), .Z(n9675) );
  NBUFFX2 U9717 ( .INP(n9738), .Z(n9676) );
  NBUFFX2 U9718 ( .INP(n9738), .Z(n9677) );
  NBUFFX2 U9719 ( .INP(n9737), .Z(n9678) );
  NBUFFX2 U9720 ( .INP(n9737), .Z(n9679) );
  NBUFFX2 U9721 ( .INP(n9737), .Z(n9680) );
  NBUFFX2 U9722 ( .INP(n9736), .Z(n9681) );
  NBUFFX2 U9723 ( .INP(n9736), .Z(n9682) );
  NBUFFX2 U9724 ( .INP(n9736), .Z(n9683) );
  NBUFFX2 U9725 ( .INP(n9735), .Z(n9684) );
  NBUFFX2 U9726 ( .INP(n9735), .Z(n9685) );
  NBUFFX2 U9727 ( .INP(n9735), .Z(n9686) );
  NBUFFX2 U9728 ( .INP(n9734), .Z(n9687) );
  NBUFFX2 U9729 ( .INP(n9734), .Z(n9688) );
  NBUFFX2 U9730 ( .INP(n9734), .Z(n9689) );
  NBUFFX2 U9731 ( .INP(n9733), .Z(n9690) );
  NBUFFX2 U9732 ( .INP(n9733), .Z(n9691) );
  NBUFFX2 U9733 ( .INP(n9733), .Z(n9692) );
  NBUFFX2 U9734 ( .INP(n9732), .Z(n9693) );
  NBUFFX2 U9735 ( .INP(n9732), .Z(n9694) );
  NBUFFX2 U9736 ( .INP(n9732), .Z(n9695) );
  NBUFFX2 U9737 ( .INP(n9731), .Z(n9696) );
  NBUFFX2 U9738 ( .INP(n9731), .Z(n9697) );
  NBUFFX2 U9739 ( .INP(n9731), .Z(n9698) );
  NBUFFX2 U9740 ( .INP(n9730), .Z(n9699) );
  NBUFFX2 U9741 ( .INP(n9730), .Z(n9700) );
  NBUFFX2 U9742 ( .INP(n9730), .Z(n9701) );
  NBUFFX2 U9743 ( .INP(n9729), .Z(n9702) );
  NBUFFX2 U9744 ( .INP(n9729), .Z(n9703) );
  NBUFFX2 U9745 ( .INP(n9729), .Z(n9704) );
  NBUFFX2 U9746 ( .INP(n9728), .Z(n9705) );
  NBUFFX2 U9747 ( .INP(n9728), .Z(n9706) );
  NBUFFX2 U9748 ( .INP(n9728), .Z(n9707) );
  NBUFFX2 U9749 ( .INP(n9727), .Z(n9708) );
  NBUFFX2 U9750 ( .INP(n9727), .Z(n9709) );
  NBUFFX2 U9751 ( .INP(n9727), .Z(n9710) );
  NBUFFX2 U9752 ( .INP(n9726), .Z(n9711) );
  NBUFFX2 U9753 ( .INP(n9726), .Z(n9712) );
  NBUFFX2 U9754 ( .INP(n9726), .Z(n9713) );
  NBUFFX2 U9755 ( .INP(n9725), .Z(n9714) );
  NBUFFX2 U9756 ( .INP(n9725), .Z(n9715) );
  NBUFFX2 U9757 ( .INP(n9725), .Z(n9716) );
  NBUFFX2 U9758 ( .INP(n9724), .Z(n9717) );
  NBUFFX2 U9759 ( .INP(n9724), .Z(n9718) );
  NBUFFX2 U9760 ( .INP(n9724), .Z(n9719) );
  NBUFFX2 U9761 ( .INP(n9723), .Z(n9720) );
  NBUFFX2 U9762 ( .INP(n9723), .Z(n9721) );
  NBUFFX2 U9763 ( .INP(n9723), .Z(n9722) );
  NBUFFX2 U9764 ( .INP(n9766), .Z(n9723) );
  NBUFFX2 U9765 ( .INP(n9766), .Z(n9724) );
  NBUFFX2 U9766 ( .INP(n9766), .Z(n9725) );
  NBUFFX2 U9767 ( .INP(n9765), .Z(n9726) );
  NBUFFX2 U9768 ( .INP(n9765), .Z(n9727) );
  NBUFFX2 U9769 ( .INP(n9765), .Z(n9728) );
  NBUFFX2 U9770 ( .INP(n9764), .Z(n9729) );
  NBUFFX2 U9771 ( .INP(n9764), .Z(n9730) );
  NBUFFX2 U9772 ( .INP(n9764), .Z(n9731) );
  NBUFFX2 U9773 ( .INP(n9763), .Z(n9732) );
  NBUFFX2 U9774 ( .INP(n9763), .Z(n9733) );
  NBUFFX2 U9775 ( .INP(n9763), .Z(n9734) );
  NBUFFX2 U9776 ( .INP(n9762), .Z(n9735) );
  NBUFFX2 U9777 ( .INP(n9762), .Z(n9736) );
  NBUFFX2 U9778 ( .INP(n9762), .Z(n9737) );
  NBUFFX2 U9779 ( .INP(n9761), .Z(n9738) );
  NBUFFX2 U9780 ( .INP(n9761), .Z(n9739) );
  NBUFFX2 U9781 ( .INP(n9761), .Z(n9740) );
  NBUFFX2 U9782 ( .INP(n9760), .Z(n9741) );
  NBUFFX2 U9783 ( .INP(n9760), .Z(n9742) );
  NBUFFX2 U9784 ( .INP(n9760), .Z(n9743) );
  NBUFFX2 U9785 ( .INP(n9759), .Z(n9744) );
  NBUFFX2 U9786 ( .INP(n9759), .Z(n9745) );
  NBUFFX2 U9787 ( .INP(n9759), .Z(n9746) );
  NBUFFX2 U9788 ( .INP(n9758), .Z(n9747) );
  NBUFFX2 U9789 ( .INP(n9758), .Z(n9748) );
  NBUFFX2 U9790 ( .INP(n9758), .Z(n9749) );
  NBUFFX2 U9791 ( .INP(n9757), .Z(n9750) );
  NBUFFX2 U9792 ( .INP(n9757), .Z(n9751) );
  NBUFFX2 U9793 ( .INP(n9757), .Z(n9752) );
  NBUFFX2 U9794 ( .INP(n9756), .Z(n9753) );
  NBUFFX2 U9795 ( .INP(n9756), .Z(n9754) );
  NBUFFX2 U9796 ( .INP(n9756), .Z(n9755) );
  NBUFFX2 U9797 ( .INP(n9770), .Z(n9756) );
  NBUFFX2 U9798 ( .INP(n9770), .Z(n9757) );
  NBUFFX2 U9799 ( .INP(n9769), .Z(n9758) );
  NBUFFX2 U9800 ( .INP(n9769), .Z(n9759) );
  NBUFFX2 U9801 ( .INP(n9769), .Z(n9760) );
  NBUFFX2 U9802 ( .INP(n9768), .Z(n9761) );
  NBUFFX2 U9803 ( .INP(n9768), .Z(n9762) );
  NBUFFX2 U9804 ( .INP(n9768), .Z(n9763) );
  NBUFFX2 U9805 ( .INP(n9767), .Z(n9764) );
  NBUFFX2 U9806 ( .INP(n9767), .Z(n9765) );
  NBUFFX2 U9807 ( .INP(n9767), .Z(n9766) );
  NBUFFX2 U9808 ( .INP(test_se), .Z(n9767) );
  NBUFFX2 U9809 ( .INP(test_se), .Z(n9768) );
  NBUFFX2 U9810 ( .INP(test_se), .Z(n9769) );
  NBUFFX2 U9811 ( .INP(test_se), .Z(n9770) );
  NBUFFX2 U9812 ( .INP(n9953), .Z(n9915) );
  NBUFFX2 U9813 ( .INP(n9953), .Z(n9916) );
  NBUFFX2 U9814 ( .INP(n9952), .Z(n9917) );
  NBUFFX2 U9815 ( .INP(n9952), .Z(n9918) );
  NBUFFX2 U9816 ( .INP(n9952), .Z(n9919) );
  NBUFFX2 U9817 ( .INP(n9951), .Z(n9920) );
  NBUFFX2 U9818 ( .INP(n9951), .Z(n9921) );
  NBUFFX2 U9819 ( .INP(n9951), .Z(n9922) );
  NBUFFX2 U9820 ( .INP(n9950), .Z(n9923) );
  NBUFFX2 U9821 ( .INP(n9950), .Z(n9924) );
  NBUFFX2 U9822 ( .INP(n9950), .Z(n9925) );
  NBUFFX2 U9823 ( .INP(n9949), .Z(n9926) );
  NBUFFX2 U9824 ( .INP(n9949), .Z(n9927) );
  NBUFFX2 U9825 ( .INP(n9949), .Z(n9928) );
  NBUFFX2 U9826 ( .INP(n9948), .Z(n9929) );
  NBUFFX2 U9827 ( .INP(n9948), .Z(n9930) );
  NBUFFX2 U9828 ( .INP(n9948), .Z(n9931) );
  NBUFFX2 U9829 ( .INP(n9947), .Z(n9932) );
  NBUFFX2 U9830 ( .INP(n9947), .Z(n9933) );
  NBUFFX2 U9831 ( .INP(n9947), .Z(n9934) );
  NBUFFX2 U9832 ( .INP(n9946), .Z(n9935) );
  NBUFFX2 U9833 ( .INP(n9946), .Z(n9936) );
  NBUFFX2 U9834 ( .INP(n9946), .Z(n9937) );
  NBUFFX2 U9835 ( .INP(n9945), .Z(n9938) );
  NBUFFX2 U9836 ( .INP(n9945), .Z(n9939) );
  NBUFFX2 U9837 ( .INP(n9945), .Z(n9940) );
  NBUFFX2 U9838 ( .INP(n9944), .Z(n9941) );
  NBUFFX2 U9839 ( .INP(n9944), .Z(n9942) );
  NBUFFX2 U9840 ( .INP(n9944), .Z(n9943) );
  NBUFFX2 U9841 ( .INP(CK), .Z(n9944) );
  NBUFFX2 U9842 ( .INP(CK), .Z(n9945) );
  NBUFFX2 U9843 ( .INP(n9953), .Z(n9946) );
  NBUFFX2 U9844 ( .INP(CK), .Z(n9947) );
  NBUFFX2 U9845 ( .INP(n9949), .Z(n9948) );
  NBUFFX2 U9846 ( .INP(CK), .Z(n9949) );
  NBUFFX2 U9847 ( .INP(n9944), .Z(n9950) );
  NBUFFX2 U9848 ( .INP(n9945), .Z(n9951) );
  NBUFFX2 U9849 ( .INP(n9947), .Z(n9952) );
  NBUFFX2 U9850 ( .INP(n9784), .Z(n9953) );
  NOR2X0 U9851 ( .IN1(TM1), .IN2(n9159), .QN(n3278) );
  NOR2X0 U9852 ( .IN1(n16412), .IN2(n9159), .QN(WX9789) );
  NOR2X0 U9853 ( .IN1(n16411), .IN2(n9159), .QN(WX9787) );
  NOR2X0 U9854 ( .IN1(n16410), .IN2(n9159), .QN(WX9785) );
  NOR2X0 U9855 ( .IN1(n16409), .IN2(n9158), .QN(WX9783) );
  NOR2X0 U9856 ( .IN1(n9224), .IN2(n8820), .QN(WX9781) );
  NOR2X0 U9857 ( .IN1(n16408), .IN2(n9158), .QN(WX9779) );
  NOR2X0 U9858 ( .IN1(n16407), .IN2(n9158), .QN(WX9777) );
  NOR2X0 U9859 ( .IN1(n16406), .IN2(n9158), .QN(WX9775) );
  NOR2X0 U9860 ( .IN1(n16405), .IN2(n9158), .QN(WX9773) );
  NOR2X0 U9861 ( .IN1(n16404), .IN2(n9158), .QN(WX9771) );
  NOR2X0 U9862 ( .IN1(n16403), .IN2(n9157), .QN(WX9769) );
  NOR2X0 U9863 ( .IN1(n16402), .IN2(n9157), .QN(WX9767) );
  NOR2X0 U9864 ( .IN1(n16401), .IN2(n9157), .QN(WX9765) );
  NOR2X0 U9865 ( .IN1(n16400), .IN2(n9157), .QN(WX9763) );
  NOR2X0 U9866 ( .IN1(n16399), .IN2(n9157), .QN(WX9761) );
  NOR2X0 U9867 ( .IN1(n16398), .IN2(n9157), .QN(WX9759) );
  NAND4X0 U9868 ( .IN1(n9954), .IN2(n9955), .IN3(n9956), .IN4(n9957), .QN(
        WX9757) );
  NAND2X0 U9869 ( .IN1(n9101), .IN2(n9959), .QN(n9957) );
  NAND2X0 U9870 ( .IN1(n9323), .IN2(n9960), .QN(n9956) );
  NAND2X0 U9871 ( .IN1(n9273), .IN2(n1728), .QN(n9955) );
  NOR2X0 U9872 ( .IN1(n9234), .IN2(n8829), .QN(n1728) );
  NAND2X0 U9873 ( .IN1(n9292), .IN2(CRC_OUT_2_0), .QN(n9954) );
  NAND4X0 U9874 ( .IN1(n9961), .IN2(n9962), .IN3(n9963), .IN4(n9964), .QN(
        WX9755) );
  NAND3X0 U9875 ( .IN1(n9965), .IN2(n9966), .IN3(n9090), .QN(n9964) );
  NAND2X0 U9876 ( .IN1(n9332), .IN2(n9967), .QN(n9963) );
  NAND2X0 U9877 ( .IN1(n1727), .IN2(n9273), .QN(n9962) );
  NOR2X0 U9878 ( .IN1(n9234), .IN2(n8830), .QN(n1727) );
  NAND2X0 U9879 ( .IN1(n9309), .IN2(CRC_OUT_2_1), .QN(n9961) );
  NAND4X0 U9880 ( .IN1(n9968), .IN2(n9969), .IN3(n9970), .IN4(n9971), .QN(
        WX9753) );
  NAND3X0 U9881 ( .IN1(n9972), .IN2(n9973), .IN3(n9321), .QN(n9971) );
  NAND2X0 U9882 ( .IN1(n9101), .IN2(n9974), .QN(n9970) );
  NAND2X0 U9883 ( .IN1(n1726), .IN2(n9273), .QN(n9969) );
  NOR2X0 U9884 ( .IN1(n9234), .IN2(n8831), .QN(n1726) );
  NAND2X0 U9885 ( .IN1(test_so87), .IN2(n9315), .QN(n9968) );
  NAND4X0 U9886 ( .IN1(n9975), .IN2(n9976), .IN3(n9977), .IN4(n9978), .QN(
        WX9751) );
  NAND3X0 U9887 ( .IN1(n9979), .IN2(n9980), .IN3(n9090), .QN(n9978) );
  NAND2X0 U9888 ( .IN1(n9329), .IN2(n9981), .QN(n9977) );
  NAND2X0 U9889 ( .IN1(n1725), .IN2(n9273), .QN(n9976) );
  NOR2X0 U9890 ( .IN1(n9234), .IN2(n8832), .QN(n1725) );
  NAND2X0 U9891 ( .IN1(n9303), .IN2(CRC_OUT_2_3), .QN(n9975) );
  NAND4X0 U9892 ( .IN1(n9982), .IN2(n9983), .IN3(n9984), .IN4(n9985), .QN(
        WX9749) );
  NAND3X0 U9893 ( .IN1(n9986), .IN2(n9987), .IN3(n9321), .QN(n9985) );
  NAND2X0 U9894 ( .IN1(n9101), .IN2(n9988), .QN(n9984) );
  NAND2X0 U9895 ( .IN1(n1724), .IN2(n9273), .QN(n9983) );
  NOR2X0 U9896 ( .IN1(n9234), .IN2(n8833), .QN(n1724) );
  NAND2X0 U9897 ( .IN1(n9303), .IN2(CRC_OUT_2_4), .QN(n9982) );
  NAND4X0 U9898 ( .IN1(n9989), .IN2(n9990), .IN3(n9991), .IN4(n9992), .QN(
        WX9747) );
  NAND2X0 U9899 ( .IN1(n9101), .IN2(n9993), .QN(n9992) );
  NAND2X0 U9900 ( .IN1(n9329), .IN2(n9994), .QN(n9991) );
  NAND2X0 U9901 ( .IN1(n1723), .IN2(n9273), .QN(n9990) );
  NOR2X0 U9902 ( .IN1(n9061), .IN2(n9157), .QN(n1723) );
  NAND2X0 U9903 ( .IN1(n9303), .IN2(CRC_OUT_2_5), .QN(n9989) );
  NAND4X0 U9904 ( .IN1(n9995), .IN2(n9996), .IN3(n9997), .IN4(n9998), .QN(
        WX9745) );
  NAND3X0 U9905 ( .IN1(n9999), .IN2(n10000), .IN3(n9321), .QN(n9998) );
  NAND2X0 U9906 ( .IN1(n9101), .IN2(n10001), .QN(n9997) );
  NAND2X0 U9907 ( .IN1(n1722), .IN2(n9273), .QN(n9996) );
  NOR2X0 U9908 ( .IN1(n9234), .IN2(n8834), .QN(n1722) );
  NAND2X0 U9909 ( .IN1(n9303), .IN2(CRC_OUT_2_6), .QN(n9995) );
  NAND4X0 U9910 ( .IN1(n10002), .IN2(n10003), .IN3(n10004), .IN4(n10005), .QN(
        WX9743) );
  NAND2X0 U9911 ( .IN1(n9101), .IN2(n10006), .QN(n10005) );
  NAND2X0 U9912 ( .IN1(n9329), .IN2(n10007), .QN(n10004) );
  NAND2X0 U9913 ( .IN1(n1721), .IN2(n9273), .QN(n10003) );
  NOR2X0 U9914 ( .IN1(n9235), .IN2(n8835), .QN(n1721) );
  NAND2X0 U9915 ( .IN1(n9304), .IN2(CRC_OUT_2_7), .QN(n10002) );
  NAND4X0 U9916 ( .IN1(n10008), .IN2(n10009), .IN3(n10010), .IN4(n10011), .QN(
        WX9741) );
  NAND3X0 U9917 ( .IN1(n10012), .IN2(n10013), .IN3(n9321), .QN(n10011) );
  NAND2X0 U9918 ( .IN1(n9101), .IN2(n10014), .QN(n10010) );
  NAND2X0 U9919 ( .IN1(n1720), .IN2(n9273), .QN(n10009) );
  NOR2X0 U9920 ( .IN1(n9235), .IN2(n8836), .QN(n1720) );
  NAND2X0 U9921 ( .IN1(n9304), .IN2(CRC_OUT_2_8), .QN(n10008) );
  NAND4X0 U9922 ( .IN1(n10015), .IN2(n10016), .IN3(n10017), .IN4(n10018), .QN(
        WX9739) );
  NAND2X0 U9923 ( .IN1(n9101), .IN2(n10019), .QN(n10018) );
  NAND2X0 U9924 ( .IN1(n9329), .IN2(n10020), .QN(n10017) );
  NAND2X0 U9925 ( .IN1(n1719), .IN2(n9273), .QN(n10016) );
  NOR2X0 U9926 ( .IN1(n9235), .IN2(n8837), .QN(n1719) );
  NAND2X0 U9927 ( .IN1(n9304), .IN2(CRC_OUT_2_9), .QN(n10015) );
  NAND4X0 U9928 ( .IN1(n10021), .IN2(n10022), .IN3(n10023), .IN4(n10024), .QN(
        WX9737) );
  NAND2X0 U9929 ( .IN1(n9101), .IN2(n10025), .QN(n10024) );
  NAND2X0 U9930 ( .IN1(n9329), .IN2(n10026), .QN(n10023) );
  NAND2X0 U9931 ( .IN1(n1718), .IN2(n9273), .QN(n10022) );
  NOR2X0 U9932 ( .IN1(n9235), .IN2(n8838), .QN(n1718) );
  NAND2X0 U9933 ( .IN1(n9304), .IN2(CRC_OUT_2_10), .QN(n10021) );
  NAND4X0 U9934 ( .IN1(n10027), .IN2(n10028), .IN3(n10029), .IN4(n10030), .QN(
        WX9735) );
  NAND2X0 U9935 ( .IN1(n9101), .IN2(n10031), .QN(n10030) );
  NAND2X0 U9936 ( .IN1(n9329), .IN2(n10032), .QN(n10029) );
  NAND2X0 U9937 ( .IN1(n1717), .IN2(n9273), .QN(n10028) );
  NOR2X0 U9938 ( .IN1(n9235), .IN2(n8839), .QN(n1717) );
  NAND2X0 U9939 ( .IN1(n9304), .IN2(CRC_OUT_2_11), .QN(n10027) );
  NAND4X0 U9940 ( .IN1(n10033), .IN2(n10034), .IN3(n10035), .IN4(n10036), .QN(
        WX9733) );
  NAND2X0 U9941 ( .IN1(n9100), .IN2(n10037), .QN(n10036) );
  NAND2X0 U9942 ( .IN1(n9329), .IN2(n10038), .QN(n10035) );
  NAND2X0 U9943 ( .IN1(n1716), .IN2(n9273), .QN(n10034) );
  NOR2X0 U9944 ( .IN1(n9235), .IN2(n8840), .QN(n1716) );
  NAND2X0 U9945 ( .IN1(n9304), .IN2(CRC_OUT_2_12), .QN(n10033) );
  NAND4X0 U9946 ( .IN1(n10039), .IN2(n10040), .IN3(n10041), .IN4(n10042), .QN(
        WX9731) );
  NAND2X0 U9947 ( .IN1(n9100), .IN2(n10043), .QN(n10042) );
  NAND2X0 U9948 ( .IN1(n9329), .IN2(n10044), .QN(n10041) );
  NAND2X0 U9949 ( .IN1(n1715), .IN2(n9273), .QN(n10040) );
  NOR2X0 U9950 ( .IN1(n9235), .IN2(n8841), .QN(n1715) );
  NAND2X0 U9951 ( .IN1(n9304), .IN2(CRC_OUT_2_13), .QN(n10039) );
  NAND4X0 U9952 ( .IN1(n10045), .IN2(n10046), .IN3(n10047), .IN4(n10048), .QN(
        WX9729) );
  NAND3X0 U9953 ( .IN1(n10049), .IN2(n10050), .IN3(n9090), .QN(n10048) );
  NAND2X0 U9954 ( .IN1(n9329), .IN2(n10051), .QN(n10047) );
  NAND2X0 U9955 ( .IN1(n1714), .IN2(n9273), .QN(n10046) );
  NOR2X0 U9956 ( .IN1(n9235), .IN2(n8842), .QN(n1714) );
  NAND2X0 U9957 ( .IN1(n9304), .IN2(CRC_OUT_2_14), .QN(n10045) );
  NAND4X0 U9958 ( .IN1(n10052), .IN2(n10053), .IN3(n10054), .IN4(n10055), .QN(
        WX9727) );
  NAND2X0 U9959 ( .IN1(n9100), .IN2(n10056), .QN(n10055) );
  NAND2X0 U9960 ( .IN1(n9329), .IN2(n10057), .QN(n10054) );
  NAND2X0 U9961 ( .IN1(n1713), .IN2(n9273), .QN(n10053) );
  NOR2X0 U9962 ( .IN1(n9235), .IN2(n8843), .QN(n1713) );
  NAND2X0 U9963 ( .IN1(n9304), .IN2(CRC_OUT_2_15), .QN(n10052) );
  NAND4X0 U9964 ( .IN1(n10058), .IN2(n10059), .IN3(n10060), .IN4(n10061), .QN(
        WX9725) );
  NAND2X0 U9965 ( .IN1(n10062), .IN2(n10063), .QN(n10061) );
  NAND3X0 U9966 ( .IN1(n10064), .IN2(n10065), .IN3(n10066), .QN(n10062) );
  NAND2X0 U9967 ( .IN1(n9329), .IN2(n10067), .QN(n10066) );
  NAND2X0 U9968 ( .IN1(n9084), .IN2(n8246), .QN(n10065) );
  NAND2X0 U9969 ( .IN1(n9078), .IN2(n16427), .QN(n10064) );
  NAND2X0 U9970 ( .IN1(n10070), .IN2(n9111), .QN(n10060) );
  NAND2X0 U9971 ( .IN1(n1712), .IN2(n9274), .QN(n10059) );
  NOR2X0 U9972 ( .IN1(n9235), .IN2(n8844), .QN(n1712) );
  NAND2X0 U9973 ( .IN1(n9304), .IN2(CRC_OUT_2_16), .QN(n10058) );
  NAND4X0 U9974 ( .IN1(n10071), .IN2(n10072), .IN3(n10073), .IN4(n10074), .QN(
        WX9723) );
  NAND2X0 U9975 ( .IN1(n10075), .IN2(n10076), .QN(n10074) );
  NAND2X0 U9976 ( .IN1(n10077), .IN2(n10078), .QN(n10075) );
  NAND2X0 U9977 ( .IN1(n9100), .IN2(n10079), .QN(n10078) );
  NAND2X0 U9978 ( .IN1(n9100), .IN2(n8305), .QN(n10077) );
  NAND2X0 U9979 ( .IN1(n10080), .IN2(n10081), .QN(n10073) );
  NAND3X0 U9980 ( .IN1(n10082), .IN2(n10083), .IN3(n10084), .QN(n10080) );
  NAND2X0 U9981 ( .IN1(n9329), .IN2(n10085), .QN(n10084) );
  NAND2X0 U9982 ( .IN1(n9083), .IN2(n8247), .QN(n10083) );
  NAND2X0 U9983 ( .IN1(n16426), .IN2(n9080), .QN(n10082) );
  NAND2X0 U9984 ( .IN1(n1711), .IN2(n9274), .QN(n10072) );
  NOR2X0 U9985 ( .IN1(n9235), .IN2(n8845), .QN(n1711) );
  NAND2X0 U9986 ( .IN1(n9304), .IN2(CRC_OUT_2_17), .QN(n10071) );
  NAND4X0 U9987 ( .IN1(n10086), .IN2(n10087), .IN3(n10088), .IN4(n10089), .QN(
        WX9721) );
  NAND2X0 U9988 ( .IN1(n10090), .IN2(n10091), .QN(n10089) );
  NAND3X0 U9989 ( .IN1(n10092), .IN2(n10093), .IN3(n10094), .QN(n10090) );
  NAND2X0 U9990 ( .IN1(n9329), .IN2(n10095), .QN(n10094) );
  NAND2X0 U9991 ( .IN1(n9082), .IN2(n8248), .QN(n10093) );
  NAND2X0 U9992 ( .IN1(n16425), .IN2(n9079), .QN(n10092) );
  NAND2X0 U9993 ( .IN1(n10096), .IN2(n9111), .QN(n10088) );
  NAND2X0 U9994 ( .IN1(n1710), .IN2(n9274), .QN(n10087) );
  NOR2X0 U9995 ( .IN1(n9236), .IN2(n8846), .QN(n1710) );
  NAND2X0 U9996 ( .IN1(n9304), .IN2(CRC_OUT_2_18), .QN(n10086) );
  NAND4X0 U9997 ( .IN1(n10097), .IN2(n10098), .IN3(n10099), .IN4(n10100), .QN(
        WX9719) );
  NAND2X0 U9998 ( .IN1(n10101), .IN2(n10102), .QN(n10100) );
  NAND2X0 U9999 ( .IN1(n10103), .IN2(n10104), .QN(n10101) );
  NAND2X0 U10000 ( .IN1(n9100), .IN2(n10105), .QN(n10104) );
  NAND2X0 U10001 ( .IN1(n9100), .IN2(n8307), .QN(n10103) );
  NAND2X0 U10002 ( .IN1(n10106), .IN2(n9336), .QN(n10099) );
  NAND2X0 U10003 ( .IN1(n1709), .IN2(n9274), .QN(n10098) );
  NOR2X0 U10004 ( .IN1(n9239), .IN2(n8847), .QN(n1709) );
  NAND2X0 U10005 ( .IN1(test_so88), .IN2(n9314), .QN(n10097) );
  NAND4X0 U10006 ( .IN1(n10107), .IN2(n10108), .IN3(n10109), .IN4(n10110), 
        .QN(WX9717) );
  NAND2X0 U10007 ( .IN1(n10111), .IN2(n10112), .QN(n10110) );
  NAND2X0 U10008 ( .IN1(n10113), .IN2(n10114), .QN(n10111) );
  NAND2X0 U10009 ( .IN1(n9100), .IN2(n10115), .QN(n10114) );
  NAND2X0 U10010 ( .IN1(n8170), .IN2(n9111), .QN(n10113) );
  NAND2X0 U10011 ( .IN1(n10116), .IN2(n10117), .QN(n10109) );
  NAND3X0 U10012 ( .IN1(n10118), .IN2(n10119), .IN3(n10120), .QN(n10116) );
  NAND2X0 U10013 ( .IN1(n9329), .IN2(n10121), .QN(n10120) );
  NAND2X0 U10014 ( .IN1(n9082), .IN2(n8250), .QN(n10119) );
  NAND2X0 U10015 ( .IN1(n16423), .IN2(n9078), .QN(n10118) );
  NAND2X0 U10016 ( .IN1(n1708), .IN2(n9274), .QN(n10108) );
  NOR2X0 U10017 ( .IN1(n9240), .IN2(n8848), .QN(n1708) );
  NAND2X0 U10018 ( .IN1(n9305), .IN2(CRC_OUT_2_20), .QN(n10107) );
  NAND4X0 U10019 ( .IN1(n10122), .IN2(n10123), .IN3(n10124), .IN4(n10125), 
        .QN(WX9715) );
  NAND2X0 U10020 ( .IN1(n10126), .IN2(n10127), .QN(n10125) );
  NAND2X0 U10021 ( .IN1(n10128), .IN2(n10129), .QN(n10126) );
  NAND2X0 U10022 ( .IN1(n9100), .IN2(n10130), .QN(n10129) );
  NAND2X0 U10023 ( .IN1(n9100), .IN2(n8310), .QN(n10128) );
  NAND2X0 U10024 ( .IN1(n10131), .IN2(n9336), .QN(n10124) );
  NAND2X0 U10025 ( .IN1(n1707), .IN2(n9274), .QN(n10123) );
  NOR2X0 U10026 ( .IN1(n9240), .IN2(n8849), .QN(n1707) );
  NAND2X0 U10027 ( .IN1(n9305), .IN2(CRC_OUT_2_21), .QN(n10122) );
  NAND4X0 U10028 ( .IN1(n10132), .IN2(n10133), .IN3(n10134), .IN4(n10135), 
        .QN(WX9713) );
  NAND2X0 U10029 ( .IN1(n10136), .IN2(n10137), .QN(n10135) );
  NAND2X0 U10030 ( .IN1(n10138), .IN2(n10139), .QN(n10136) );
  NAND2X0 U10031 ( .IN1(n9100), .IN2(n10140), .QN(n10139) );
  NAND2X0 U10032 ( .IN1(n9100), .IN2(n8311), .QN(n10138) );
  NAND2X0 U10033 ( .IN1(n10141), .IN2(n10142), .QN(n10134) );
  NAND3X0 U10034 ( .IN1(n10143), .IN2(n10144), .IN3(n10145), .QN(n10141) );
  NAND2X0 U10035 ( .IN1(n9329), .IN2(n10146), .QN(n10145) );
  NAND2X0 U10036 ( .IN1(n9084), .IN2(n8252), .QN(n10144) );
  NAND2X0 U10037 ( .IN1(n16421), .IN2(n9078), .QN(n10143) );
  NAND2X0 U10038 ( .IN1(n1706), .IN2(n9274), .QN(n10133) );
  NOR2X0 U10039 ( .IN1(n9062), .IN2(n9156), .QN(n1706) );
  NAND2X0 U10040 ( .IN1(n9305), .IN2(CRC_OUT_2_22), .QN(n10132) );
  NAND4X0 U10041 ( .IN1(n10147), .IN2(n10148), .IN3(n10149), .IN4(n10150), 
        .QN(WX9711) );
  NAND2X0 U10042 ( .IN1(n10151), .IN2(n10152), .QN(n10150) );
  NAND2X0 U10043 ( .IN1(n10153), .IN2(n10154), .QN(n10151) );
  NAND2X0 U10044 ( .IN1(n9100), .IN2(n10155), .QN(n10154) );
  NAND2X0 U10045 ( .IN1(n9100), .IN2(n8312), .QN(n10153) );
  NAND2X0 U10046 ( .IN1(n10156), .IN2(n9336), .QN(n10149) );
  NAND2X0 U10047 ( .IN1(n1705), .IN2(n9274), .QN(n10148) );
  NOR2X0 U10048 ( .IN1(n9240), .IN2(n8850), .QN(n1705) );
  NAND2X0 U10049 ( .IN1(n9305), .IN2(CRC_OUT_2_23), .QN(n10147) );
  NAND4X0 U10050 ( .IN1(n10157), .IN2(n10158), .IN3(n10159), .IN4(n10160), 
        .QN(WX9709) );
  NAND2X0 U10051 ( .IN1(n10161), .IN2(n10162), .QN(n10160) );
  NAND2X0 U10052 ( .IN1(n10163), .IN2(n10164), .QN(n10161) );
  NAND2X0 U10053 ( .IN1(n9100), .IN2(n10165), .QN(n10164) );
  NAND2X0 U10054 ( .IN1(n9100), .IN2(n8313), .QN(n10163) );
  NAND2X0 U10055 ( .IN1(n10166), .IN2(n10167), .QN(n10159) );
  NAND3X0 U10056 ( .IN1(n10168), .IN2(n10169), .IN3(n10170), .QN(n10166) );
  NAND2X0 U10057 ( .IN1(n9329), .IN2(n10171), .QN(n10170) );
  NAND2X0 U10058 ( .IN1(n9083), .IN2(n8254), .QN(n10169) );
  NAND2X0 U10059 ( .IN1(n16419), .IN2(n9080), .QN(n10168) );
  NAND2X0 U10060 ( .IN1(n1704), .IN2(n9274), .QN(n10158) );
  NOR2X0 U10061 ( .IN1(n9240), .IN2(n8851), .QN(n1704) );
  NAND2X0 U10062 ( .IN1(n9305), .IN2(CRC_OUT_2_24), .QN(n10157) );
  NAND4X0 U10063 ( .IN1(n10172), .IN2(n10173), .IN3(n10174), .IN4(n10175), 
        .QN(WX9707) );
  NAND2X0 U10064 ( .IN1(n10176), .IN2(n10177), .QN(n10175) );
  NAND2X0 U10065 ( .IN1(n10178), .IN2(n10179), .QN(n10176) );
  NAND2X0 U10066 ( .IN1(n9100), .IN2(n10180), .QN(n10179) );
  NAND2X0 U10067 ( .IN1(n9100), .IN2(n8314), .QN(n10178) );
  NAND2X0 U10068 ( .IN1(n10181), .IN2(n10182), .QN(n10174) );
  NAND3X0 U10069 ( .IN1(n10183), .IN2(n10184), .IN3(n10185), .QN(n10181) );
  NAND2X0 U10070 ( .IN1(n9329), .IN2(n10186), .QN(n10185) );
  NAND2X0 U10071 ( .IN1(n10069), .IN2(WX11193), .QN(n10184) );
  NAND2X0 U10072 ( .IN1(n9082), .IN2(n8140), .QN(n10183) );
  NAND2X0 U10073 ( .IN1(n1703), .IN2(n9274), .QN(n10173) );
  NOR2X0 U10074 ( .IN1(n9240), .IN2(n8852), .QN(n1703) );
  NAND2X0 U10075 ( .IN1(n9305), .IN2(CRC_OUT_2_25), .QN(n10172) );
  NAND4X0 U10076 ( .IN1(n10187), .IN2(n10188), .IN3(n10189), .IN4(n10190), 
        .QN(WX9705) );
  NAND2X0 U10077 ( .IN1(n10191), .IN2(n10192), .QN(n10190) );
  NAND2X0 U10078 ( .IN1(n10193), .IN2(n10194), .QN(n10191) );
  NAND2X0 U10079 ( .IN1(n9099), .IN2(n10195), .QN(n10194) );
  NAND2X0 U10080 ( .IN1(n9099), .IN2(n8315), .QN(n10193) );
  NAND2X0 U10081 ( .IN1(n10196), .IN2(n10197), .QN(n10189) );
  NAND3X0 U10082 ( .IN1(n10198), .IN2(n10199), .IN3(n10200), .QN(n10196) );
  NAND2X0 U10083 ( .IN1(n9330), .IN2(n10201), .QN(n10200) );
  NAND2X0 U10084 ( .IN1(n10068), .IN2(n8257), .QN(n10199) );
  NAND2X0 U10085 ( .IN1(n16418), .IN2(n9079), .QN(n10198) );
  NAND2X0 U10086 ( .IN1(n1702), .IN2(n9274), .QN(n10188) );
  NOR2X0 U10087 ( .IN1(n9240), .IN2(n8853), .QN(n1702) );
  NAND2X0 U10088 ( .IN1(n9305), .IN2(CRC_OUT_2_26), .QN(n10187) );
  NAND4X0 U10089 ( .IN1(n10202), .IN2(n10203), .IN3(n10204), .IN4(n10205), 
        .QN(WX9703) );
  NAND2X0 U10090 ( .IN1(n10206), .IN2(n10207), .QN(n10205) );
  NAND2X0 U10091 ( .IN1(n10208), .IN2(n10209), .QN(n10206) );
  NAND2X0 U10092 ( .IN1(n9099), .IN2(n10210), .QN(n10209) );
  NAND2X0 U10093 ( .IN1(n9099), .IN2(n8316), .QN(n10208) );
  NAND2X0 U10094 ( .IN1(n10211), .IN2(n10212), .QN(n10204) );
  NAND3X0 U10095 ( .IN1(n10213), .IN2(n10214), .IN3(n10215), .QN(n10211) );
  NAND2X0 U10096 ( .IN1(n9330), .IN2(n10216), .QN(n10215) );
  NAND2X0 U10097 ( .IN1(n9084), .IN2(n8258), .QN(n10214) );
  NAND2X0 U10098 ( .IN1(n16417), .IN2(n9078), .QN(n10213) );
  NAND2X0 U10099 ( .IN1(n1701), .IN2(n9274), .QN(n10203) );
  NOR2X0 U10100 ( .IN1(n9240), .IN2(n8854), .QN(n1701) );
  NAND2X0 U10101 ( .IN1(n9305), .IN2(CRC_OUT_2_27), .QN(n10202) );
  NAND4X0 U10102 ( .IN1(n10217), .IN2(n10218), .IN3(n10219), .IN4(n10220), 
        .QN(WX9701) );
  NAND2X0 U10103 ( .IN1(n10221), .IN2(n10222), .QN(n10220) );
  NAND2X0 U10104 ( .IN1(n10223), .IN2(n10224), .QN(n10221) );
  NAND2X0 U10105 ( .IN1(n9099), .IN2(n10225), .QN(n10224) );
  NAND2X0 U10106 ( .IN1(n9099), .IN2(n8317), .QN(n10223) );
  NAND2X0 U10107 ( .IN1(n10226), .IN2(n10227), .QN(n10219) );
  NAND3X0 U10108 ( .IN1(n10228), .IN2(n10229), .IN3(n10230), .QN(n10226) );
  NAND2X0 U10109 ( .IN1(n9330), .IN2(n10231), .QN(n10230) );
  NAND2X0 U10110 ( .IN1(n9083), .IN2(n8259), .QN(n10229) );
  NAND2X0 U10111 ( .IN1(n16416), .IN2(n10069), .QN(n10228) );
  NAND2X0 U10112 ( .IN1(n1700), .IN2(n9274), .QN(n10218) );
  NOR2X0 U10113 ( .IN1(n9240), .IN2(n8855), .QN(n1700) );
  NAND2X0 U10114 ( .IN1(n9305), .IN2(CRC_OUT_2_28), .QN(n10217) );
  NAND4X0 U10115 ( .IN1(n10232), .IN2(n10233), .IN3(n10234), .IN4(n10235), 
        .QN(WX9699) );
  NAND2X0 U10116 ( .IN1(n10236), .IN2(n10237), .QN(n10235) );
  NAND2X0 U10117 ( .IN1(n10238), .IN2(n10239), .QN(n10236) );
  NAND2X0 U10118 ( .IN1(n9099), .IN2(n10240), .QN(n10239) );
  NAND2X0 U10119 ( .IN1(n9099), .IN2(n8318), .QN(n10238) );
  NAND2X0 U10120 ( .IN1(n10241), .IN2(n10242), .QN(n10234) );
  NAND3X0 U10121 ( .IN1(n10243), .IN2(n10244), .IN3(n10245), .QN(n10241) );
  NAND2X0 U10122 ( .IN1(n9330), .IN2(n10246), .QN(n10245) );
  NAND2X0 U10123 ( .IN1(n9082), .IN2(n8260), .QN(n10244) );
  NAND2X0 U10124 ( .IN1(n16415), .IN2(n9080), .QN(n10243) );
  NAND2X0 U10125 ( .IN1(n1699), .IN2(n9274), .QN(n10233) );
  NOR2X0 U10126 ( .IN1(n9241), .IN2(n8856), .QN(n1699) );
  NAND2X0 U10127 ( .IN1(n9305), .IN2(CRC_OUT_2_29), .QN(n10232) );
  NAND4X0 U10128 ( .IN1(n10247), .IN2(n10248), .IN3(n10249), .IN4(n10250), 
        .QN(WX9697) );
  NAND2X0 U10129 ( .IN1(n10251), .IN2(n10252), .QN(n10250) );
  NAND2X0 U10130 ( .IN1(n10253), .IN2(n10254), .QN(n10251) );
  NAND2X0 U10131 ( .IN1(n9099), .IN2(n10255), .QN(n10254) );
  NAND2X0 U10132 ( .IN1(n9099), .IN2(n8319), .QN(n10253) );
  NAND2X0 U10133 ( .IN1(n10256), .IN2(n10257), .QN(n10249) );
  NAND3X0 U10134 ( .IN1(n10258), .IN2(n10259), .IN3(n10260), .QN(n10256) );
  NAND2X0 U10135 ( .IN1(n9330), .IN2(n10261), .QN(n10260) );
  NAND2X0 U10136 ( .IN1(n10068), .IN2(n8261), .QN(n10259) );
  NAND2X0 U10137 ( .IN1(n16414), .IN2(n9079), .QN(n10258) );
  NAND2X0 U10138 ( .IN1(n1698), .IN2(n9274), .QN(n10248) );
  NOR2X0 U10139 ( .IN1(n9241), .IN2(n8857), .QN(n1698) );
  NAND2X0 U10140 ( .IN1(n9305), .IN2(CRC_OUT_2_30), .QN(n10247) );
  NAND4X0 U10141 ( .IN1(n10262), .IN2(n10263), .IN3(n10264), .IN4(n10265), 
        .QN(WX9695) );
  NAND2X0 U10142 ( .IN1(n10266), .IN2(n10267), .QN(n10265) );
  NAND3X0 U10143 ( .IN1(n10268), .IN2(n10269), .IN3(n10270), .QN(n10266) );
  NAND2X0 U10144 ( .IN1(n9330), .IN2(n10271), .QN(n10270) );
  NAND2X0 U10145 ( .IN1(n9084), .IN2(n8262), .QN(n10269) );
  NAND2X0 U10146 ( .IN1(n16413), .IN2(n9078), .QN(n10268) );
  NAND2X0 U10147 ( .IN1(n10272), .IN2(n9111), .QN(n10264) );
  NAND2X0 U10148 ( .IN1(n9305), .IN2(CRC_OUT_2_31), .QN(n10263) );
  NAND2X0 U10149 ( .IN1(n2245), .IN2(WX9536), .QN(n10262) );
  NOR2X0 U10150 ( .IN1(n9241), .IN2(WX9536), .QN(WX9597) );
  NOR3X0 U10151 ( .IN1(n9147), .IN2(n10273), .IN3(n10274), .QN(WX9084) );
  NOR2X0 U10152 ( .IN1(n8186), .IN2(CRC_OUT_3_30), .QN(n10274) );
  NOR2X0 U10153 ( .IN1(DFF_1342_n1), .IN2(WX8595), .QN(n10273) );
  NOR3X0 U10154 ( .IN1(n9147), .IN2(n10275), .IN3(n10276), .QN(WX9082) );
  NOR2X0 U10155 ( .IN1(n8187), .IN2(CRC_OUT_3_29), .QN(n10276) );
  NOR2X0 U10156 ( .IN1(DFF_1341_n1), .IN2(WX8597), .QN(n10275) );
  NOR3X0 U10157 ( .IN1(n9147), .IN2(n10277), .IN3(n10278), .QN(WX9080) );
  NOR2X0 U10158 ( .IN1(n8188), .IN2(CRC_OUT_3_28), .QN(n10278) );
  NOR2X0 U10159 ( .IN1(DFF_1340_n1), .IN2(WX8599), .QN(n10277) );
  NOR3X0 U10160 ( .IN1(n9147), .IN2(n10279), .IN3(n10280), .QN(WX9078) );
  NOR2X0 U10161 ( .IN1(n8189), .IN2(CRC_OUT_3_27), .QN(n10280) );
  NOR2X0 U10162 ( .IN1(DFF_1339_n1), .IN2(WX8601), .QN(n10279) );
  NOR3X0 U10163 ( .IN1(n9147), .IN2(n10281), .IN3(n10282), .QN(WX9076) );
  NOR2X0 U10164 ( .IN1(n8190), .IN2(CRC_OUT_3_26), .QN(n10282) );
  NOR2X0 U10165 ( .IN1(DFF_1338_n1), .IN2(WX8603), .QN(n10281) );
  NOR2X0 U10166 ( .IN1(n9241), .IN2(n10283), .QN(WX9074) );
  NOR2X0 U10167 ( .IN1(n10284), .IN2(n10285), .QN(n10283) );
  NOR2X0 U10168 ( .IN1(test_so74), .IN2(CRC_OUT_3_25), .QN(n10285) );
  NOR2X0 U10169 ( .IN1(DFF_1337_n1), .IN2(n8799), .QN(n10284) );
  NOR2X0 U10170 ( .IN1(n9241), .IN2(n10286), .QN(WX9072) );
  NOR2X0 U10171 ( .IN1(n10287), .IN2(n10288), .QN(n10286) );
  NOR2X0 U10172 ( .IN1(test_so77), .IN2(WX8607), .QN(n10288) );
  INVX0 U10173 ( .INP(n10289), .ZN(n10287) );
  NAND2X0 U10174 ( .IN1(WX8607), .IN2(test_so77), .QN(n10289) );
  NOR3X0 U10175 ( .IN1(n9146), .IN2(n10290), .IN3(n10291), .QN(WX9070) );
  NOR2X0 U10176 ( .IN1(n8192), .IN2(CRC_OUT_3_23), .QN(n10291) );
  NOR2X0 U10177 ( .IN1(DFF_1335_n1), .IN2(WX8609), .QN(n10290) );
  NOR3X0 U10178 ( .IN1(n9146), .IN2(n10292), .IN3(n10293), .QN(WX9068) );
  NOR2X0 U10179 ( .IN1(n8193), .IN2(CRC_OUT_3_22), .QN(n10293) );
  NOR2X0 U10180 ( .IN1(DFF_1334_n1), .IN2(WX8611), .QN(n10292) );
  NOR3X0 U10181 ( .IN1(n9146), .IN2(n10294), .IN3(n10295), .QN(WX9066) );
  NOR2X0 U10182 ( .IN1(n8194), .IN2(CRC_OUT_3_21), .QN(n10295) );
  NOR2X0 U10183 ( .IN1(DFF_1333_n1), .IN2(WX8613), .QN(n10294) );
  NOR3X0 U10184 ( .IN1(n9146), .IN2(n10296), .IN3(n10297), .QN(WX9064) );
  NOR2X0 U10185 ( .IN1(n8195), .IN2(CRC_OUT_3_20), .QN(n10297) );
  NOR2X0 U10186 ( .IN1(DFF_1332_n1), .IN2(WX8615), .QN(n10296) );
  NOR3X0 U10187 ( .IN1(n9146), .IN2(n10298), .IN3(n10299), .QN(WX9062) );
  NOR2X0 U10188 ( .IN1(n8196), .IN2(CRC_OUT_3_19), .QN(n10299) );
  NOR2X0 U10189 ( .IN1(DFF_1331_n1), .IN2(WX8617), .QN(n10298) );
  NOR3X0 U10190 ( .IN1(n9146), .IN2(n10300), .IN3(n10301), .QN(WX9060) );
  NOR2X0 U10191 ( .IN1(n8197), .IN2(CRC_OUT_3_18), .QN(n10301) );
  NOR2X0 U10192 ( .IN1(DFF_1330_n1), .IN2(WX8619), .QN(n10300) );
  NOR3X0 U10193 ( .IN1(n9146), .IN2(n10302), .IN3(n10303), .QN(WX9058) );
  NOR2X0 U10194 ( .IN1(n8198), .IN2(CRC_OUT_3_17), .QN(n10303) );
  NOR2X0 U10195 ( .IN1(DFF_1329_n1), .IN2(WX8621), .QN(n10302) );
  NOR3X0 U10196 ( .IN1(n9146), .IN2(n10304), .IN3(n10305), .QN(WX9056) );
  NOR2X0 U10197 ( .IN1(n8199), .IN2(CRC_OUT_3_16), .QN(n10305) );
  NOR2X0 U10198 ( .IN1(DFF_1328_n1), .IN2(WX8623), .QN(n10304) );
  NOR2X0 U10199 ( .IN1(n9226), .IN2(n10306), .QN(WX9054) );
  NOR2X0 U10200 ( .IN1(n10307), .IN2(n10308), .QN(n10306) );
  INVX0 U10201 ( .INP(n10309), .ZN(n10308) );
  NAND2X0 U10202 ( .IN1(CRC_OUT_3_15), .IN2(n10310), .QN(n10309) );
  NOR2X0 U10203 ( .IN1(n10310), .IN2(CRC_OUT_3_15), .QN(n10307) );
  NAND2X0 U10204 ( .IN1(n10311), .IN2(n10312), .QN(n10310) );
  NAND2X0 U10205 ( .IN1(n8111), .IN2(CRC_OUT_3_31), .QN(n10312) );
  NAND2X0 U10206 ( .IN1(DFF_1343_n1), .IN2(WX8625), .QN(n10311) );
  NOR3X0 U10207 ( .IN1(n9146), .IN2(n10313), .IN3(n10314), .QN(WX9052) );
  NOR2X0 U10208 ( .IN1(n8200), .IN2(CRC_OUT_3_14), .QN(n10314) );
  NOR2X0 U10209 ( .IN1(DFF_1326_n1), .IN2(WX8627), .QN(n10313) );
  NOR3X0 U10210 ( .IN1(n9146), .IN2(n10315), .IN3(n10316), .QN(WX9050) );
  NOR2X0 U10211 ( .IN1(n8201), .IN2(CRC_OUT_3_13), .QN(n10316) );
  NOR2X0 U10212 ( .IN1(DFF_1325_n1), .IN2(WX8629), .QN(n10315) );
  NOR3X0 U10213 ( .IN1(n9146), .IN2(n10317), .IN3(n10318), .QN(WX9048) );
  NOR2X0 U10214 ( .IN1(n8202), .IN2(CRC_OUT_3_12), .QN(n10318) );
  NOR2X0 U10215 ( .IN1(DFF_1324_n1), .IN2(WX8631), .QN(n10317) );
  NOR3X0 U10216 ( .IN1(n9146), .IN2(n10319), .IN3(n10320), .QN(WX9046) );
  NOR2X0 U10217 ( .IN1(n8203), .IN2(CRC_OUT_3_11), .QN(n10320) );
  NOR2X0 U10218 ( .IN1(DFF_1323_n1), .IN2(WX8633), .QN(n10319) );
  NOR2X0 U10219 ( .IN1(n9226), .IN2(n10321), .QN(WX9044) );
  NOR2X0 U10220 ( .IN1(n10322), .IN2(n10323), .QN(n10321) );
  INVX0 U10221 ( .INP(n10324), .ZN(n10323) );
  NAND2X0 U10222 ( .IN1(CRC_OUT_3_10), .IN2(n10325), .QN(n10324) );
  NOR2X0 U10223 ( .IN1(n10325), .IN2(CRC_OUT_3_10), .QN(n10322) );
  NAND2X0 U10224 ( .IN1(n10326), .IN2(n10327), .QN(n10325) );
  NAND2X0 U10225 ( .IN1(n8112), .IN2(CRC_OUT_3_31), .QN(n10327) );
  NAND2X0 U10226 ( .IN1(DFF_1343_n1), .IN2(WX8635), .QN(n10326) );
  NOR3X0 U10227 ( .IN1(n9145), .IN2(n10328), .IN3(n10329), .QN(WX9042) );
  NOR2X0 U10228 ( .IN1(n8204), .IN2(CRC_OUT_3_9), .QN(n10329) );
  NOR2X0 U10229 ( .IN1(DFF_1321_n1), .IN2(WX8637), .QN(n10328) );
  NOR2X0 U10230 ( .IN1(n9226), .IN2(n10330), .QN(WX9040) );
  NOR2X0 U10231 ( .IN1(n10331), .IN2(n10332), .QN(n10330) );
  NOR2X0 U10232 ( .IN1(test_so75), .IN2(CRC_OUT_3_8), .QN(n10332) );
  NOR2X0 U10233 ( .IN1(DFF_1320_n1), .IN2(n8791), .QN(n10331) );
  NOR2X0 U10234 ( .IN1(n9226), .IN2(n10333), .QN(WX9038) );
  NOR2X0 U10235 ( .IN1(n10334), .IN2(n10335), .QN(n10333) );
  NOR2X0 U10236 ( .IN1(test_so76), .IN2(WX8641), .QN(n10335) );
  INVX0 U10237 ( .INP(n10336), .ZN(n10334) );
  NAND2X0 U10238 ( .IN1(WX8641), .IN2(test_so76), .QN(n10336) );
  NOR3X0 U10239 ( .IN1(n9145), .IN2(n10337), .IN3(n10338), .QN(WX9036) );
  NOR2X0 U10240 ( .IN1(n8206), .IN2(CRC_OUT_3_6), .QN(n10338) );
  NOR2X0 U10241 ( .IN1(DFF_1318_n1), .IN2(WX8643), .QN(n10337) );
  NOR3X0 U10242 ( .IN1(n9145), .IN2(n10339), .IN3(n10340), .QN(WX9034) );
  NOR2X0 U10243 ( .IN1(n8207), .IN2(CRC_OUT_3_5), .QN(n10340) );
  NOR2X0 U10244 ( .IN1(DFF_1317_n1), .IN2(WX8645), .QN(n10339) );
  NOR3X0 U10245 ( .IN1(n9145), .IN2(n10341), .IN3(n10342), .QN(WX9032) );
  NOR2X0 U10246 ( .IN1(n8208), .IN2(CRC_OUT_3_4), .QN(n10342) );
  NOR2X0 U10247 ( .IN1(DFF_1316_n1), .IN2(WX8647), .QN(n10341) );
  NOR2X0 U10248 ( .IN1(n9226), .IN2(n10343), .QN(WX9030) );
  NOR2X0 U10249 ( .IN1(n10344), .IN2(n10345), .QN(n10343) );
  INVX0 U10250 ( .INP(n10346), .ZN(n10345) );
  NAND2X0 U10251 ( .IN1(CRC_OUT_3_3), .IN2(n10347), .QN(n10346) );
  NOR2X0 U10252 ( .IN1(n10347), .IN2(CRC_OUT_3_3), .QN(n10344) );
  NAND2X0 U10253 ( .IN1(n10348), .IN2(n10349), .QN(n10347) );
  NAND2X0 U10254 ( .IN1(n8113), .IN2(CRC_OUT_3_31), .QN(n10349) );
  NAND2X0 U10255 ( .IN1(DFF_1343_n1), .IN2(WX8649), .QN(n10348) );
  NOR3X0 U10256 ( .IN1(n9145), .IN2(n10350), .IN3(n10351), .QN(WX9028) );
  NOR2X0 U10257 ( .IN1(n8209), .IN2(CRC_OUT_3_2), .QN(n10351) );
  NOR2X0 U10258 ( .IN1(DFF_1314_n1), .IN2(WX8651), .QN(n10350) );
  NOR3X0 U10259 ( .IN1(n9145), .IN2(n10352), .IN3(n10353), .QN(WX9026) );
  NOR2X0 U10260 ( .IN1(n8210), .IN2(CRC_OUT_3_1), .QN(n10353) );
  NOR2X0 U10261 ( .IN1(DFF_1313_n1), .IN2(WX8653), .QN(n10352) );
  NOR3X0 U10262 ( .IN1(n9145), .IN2(n10354), .IN3(n10355), .QN(WX9024) );
  NOR2X0 U10263 ( .IN1(n8211), .IN2(CRC_OUT_3_0), .QN(n10355) );
  NOR2X0 U10264 ( .IN1(DFF_1312_n1), .IN2(WX8655), .QN(n10354) );
  NOR3X0 U10265 ( .IN1(n9145), .IN2(n10356), .IN3(n10357), .QN(WX9022) );
  NOR2X0 U10266 ( .IN1(n8128), .IN2(CRC_OUT_3_31), .QN(n10357) );
  NOR2X0 U10267 ( .IN1(DFF_1343_n1), .IN2(WX8657), .QN(n10356) );
  NOR2X0 U10268 ( .IN1(n16397), .IN2(n9155), .QN(WX8496) );
  NOR2X0 U10269 ( .IN1(n16396), .IN2(n9157), .QN(WX8494) );
  NOR2X0 U10270 ( .IN1(n16395), .IN2(n9156), .QN(WX8492) );
  NOR2X0 U10271 ( .IN1(n16394), .IN2(n9159), .QN(WX8490) );
  NOR2X0 U10272 ( .IN1(n16393), .IN2(n9155), .QN(WX8488) );
  NOR2X0 U10273 ( .IN1(n16392), .IN2(n9156), .QN(WX8486) );
  NOR2X0 U10274 ( .IN1(n16391), .IN2(n9156), .QN(WX8484) );
  NOR2X0 U10275 ( .IN1(n16390), .IN2(n9156), .QN(WX8482) );
  NOR2X0 U10276 ( .IN1(n16389), .IN2(n9156), .QN(WX8480) );
  NOR2X0 U10277 ( .IN1(n16388), .IN2(n9157), .QN(WX8478) );
  NOR2X0 U10278 ( .IN1(n16387), .IN2(n9156), .QN(WX8476) );
  NOR2X0 U10279 ( .IN1(n16386), .IN2(n9156), .QN(WX8474) );
  NOR2X0 U10280 ( .IN1(n16385), .IN2(n9157), .QN(WX8472) );
  NOR2X0 U10281 ( .IN1(n16384), .IN2(n9157), .QN(WX8470) );
  NOR2X0 U10282 ( .IN1(n16383), .IN2(n9156), .QN(WX8468) );
  NOR2X0 U10283 ( .IN1(n16382), .IN2(n9157), .QN(WX8466) );
  NAND4X0 U10284 ( .IN1(n10358), .IN2(n10359), .IN3(n10360), .IN4(n10361), 
        .QN(WX8464) );
  NAND2X0 U10285 ( .IN1(n9330), .IN2(n9959), .QN(n10361) );
  NAND2X0 U10286 ( .IN1(n10362), .IN2(n10363), .QN(n9959) );
  INVX0 U10287 ( .INP(n10364), .ZN(n10363) );
  NOR2X0 U10288 ( .IN1(n10365), .IN2(n10366), .QN(n10364) );
  NAND2X0 U10289 ( .IN1(n10366), .IN2(n10365), .QN(n10362) );
  NOR2X0 U10290 ( .IN1(n10367), .IN2(n10368), .QN(n10365) );
  NOR2X0 U10291 ( .IN1(WX9950), .IN2(n7885), .QN(n10368) );
  INVX0 U10292 ( .INP(n10369), .ZN(n10367) );
  NAND2X0 U10293 ( .IN1(n7885), .IN2(WX9950), .QN(n10369) );
  NAND2X0 U10294 ( .IN1(n10370), .IN2(n10371), .QN(n10366) );
  NAND2X0 U10295 ( .IN1(n7884), .IN2(WX9822), .QN(n10371) );
  INVX0 U10296 ( .INP(n10372), .ZN(n10370) );
  NOR2X0 U10297 ( .IN1(WX9822), .IN2(n7884), .QN(n10372) );
  NAND2X0 U10298 ( .IN1(n9099), .IN2(n10373), .QN(n10360) );
  NAND2X0 U10299 ( .IN1(n1486), .IN2(n9274), .QN(n10359) );
  NOR2X0 U10300 ( .IN1(n9063), .IN2(n9156), .QN(n1486) );
  NAND2X0 U10301 ( .IN1(n9306), .IN2(CRC_OUT_3_0), .QN(n10358) );
  NAND4X0 U10302 ( .IN1(n10374), .IN2(n10375), .IN3(n10376), .IN4(n10377), 
        .QN(WX8462) );
  NAND3X0 U10303 ( .IN1(n9965), .IN2(n9966), .IN3(n9322), .QN(n10377) );
  NAND3X0 U10304 ( .IN1(n10378), .IN2(n10379), .IN3(n10380), .QN(n9966) );
  INVX0 U10305 ( .INP(n10381), .ZN(n10380) );
  NAND2X0 U10306 ( .IN1(n10381), .IN2(n10382), .QN(n9965) );
  NAND2X0 U10307 ( .IN1(n10378), .IN2(n10379), .QN(n10382) );
  NAND2X0 U10308 ( .IN1(n8185), .IN2(WX9884), .QN(n10379) );
  NAND2X0 U10309 ( .IN1(n7887), .IN2(WX9948), .QN(n10378) );
  NOR2X0 U10310 ( .IN1(n10383), .IN2(n10384), .QN(n10381) );
  INVX0 U10311 ( .INP(n10385), .ZN(n10384) );
  NAND2X0 U10312 ( .IN1(test_so83), .IN2(WX9756), .QN(n10385) );
  NOR2X0 U10313 ( .IN1(WX9756), .IN2(test_so83), .QN(n10383) );
  NAND2X0 U10314 ( .IN1(n9099), .IN2(n10386), .QN(n10376) );
  NAND2X0 U10315 ( .IN1(n1485), .IN2(n9274), .QN(n10375) );
  NOR2X0 U10316 ( .IN1(n9227), .IN2(n8858), .QN(n1485) );
  NAND2X0 U10317 ( .IN1(n9306), .IN2(CRC_OUT_3_1), .QN(n10374) );
  NAND4X0 U10318 ( .IN1(n10387), .IN2(n10388), .IN3(n10389), .IN4(n10390), 
        .QN(WX8460) );
  NAND2X0 U10319 ( .IN1(n9330), .IN2(n9974), .QN(n10390) );
  NAND2X0 U10320 ( .IN1(n10391), .IN2(n10392), .QN(n9974) );
  INVX0 U10321 ( .INP(n10393), .ZN(n10392) );
  NOR2X0 U10322 ( .IN1(n10394), .IN2(n10395), .QN(n10393) );
  NAND2X0 U10323 ( .IN1(n10395), .IN2(n10394), .QN(n10391) );
  NOR2X0 U10324 ( .IN1(n10396), .IN2(n10397), .QN(n10394) );
  NOR2X0 U10325 ( .IN1(WX9946), .IN2(n7889), .QN(n10397) );
  INVX0 U10326 ( .INP(n10398), .ZN(n10396) );
  NAND2X0 U10327 ( .IN1(n7889), .IN2(WX9946), .QN(n10398) );
  NAND2X0 U10328 ( .IN1(n10399), .IN2(n10400), .QN(n10395) );
  NAND2X0 U10329 ( .IN1(n7888), .IN2(WX9818), .QN(n10400) );
  INVX0 U10330 ( .INP(n10401), .ZN(n10399) );
  NOR2X0 U10331 ( .IN1(WX9818), .IN2(n7888), .QN(n10401) );
  NAND2X0 U10332 ( .IN1(n9099), .IN2(n10402), .QN(n10389) );
  NAND2X0 U10333 ( .IN1(n1484), .IN2(n9275), .QN(n10388) );
  NOR2X0 U10334 ( .IN1(n9228), .IN2(n8859), .QN(n1484) );
  NAND2X0 U10335 ( .IN1(n9306), .IN2(CRC_OUT_3_2), .QN(n10387) );
  NAND4X0 U10336 ( .IN1(n10403), .IN2(n10404), .IN3(n10405), .IN4(n10406), 
        .QN(WX8458) );
  NAND3X0 U10337 ( .IN1(n9979), .IN2(n9980), .IN3(n9321), .QN(n10406) );
  NAND3X0 U10338 ( .IN1(n10407), .IN2(n10408), .IN3(n10409), .QN(n9980) );
  INVX0 U10339 ( .INP(n10410), .ZN(n10409) );
  NAND2X0 U10340 ( .IN1(n10410), .IN2(n10411), .QN(n9979) );
  NAND2X0 U10341 ( .IN1(n10407), .IN2(n10408), .QN(n10411) );
  NAND2X0 U10342 ( .IN1(n8183), .IN2(WX9816), .QN(n10408) );
  NAND2X0 U10343 ( .IN1(n3569), .IN2(WX9944), .QN(n10407) );
  NOR2X0 U10344 ( .IN1(n10412), .IN2(n10413), .QN(n10410) );
  INVX0 U10345 ( .INP(n10414), .ZN(n10413) );
  NAND2X0 U10346 ( .IN1(test_so81), .IN2(WX9880), .QN(n10414) );
  NOR2X0 U10347 ( .IN1(WX9880), .IN2(test_so81), .QN(n10412) );
  NAND2X0 U10348 ( .IN1(n9099), .IN2(n10415), .QN(n10405) );
  NAND2X0 U10349 ( .IN1(n1483), .IN2(n9275), .QN(n10404) );
  NOR2X0 U10350 ( .IN1(n9228), .IN2(n8860), .QN(n1483) );
  NAND2X0 U10351 ( .IN1(n9306), .IN2(CRC_OUT_3_3), .QN(n10403) );
  NAND4X0 U10352 ( .IN1(n10416), .IN2(n10417), .IN3(n10418), .IN4(n10419), 
        .QN(WX8456) );
  NAND2X0 U10353 ( .IN1(n9330), .IN2(n9988), .QN(n10419) );
  NAND2X0 U10354 ( .IN1(n10420), .IN2(n10421), .QN(n9988) );
  INVX0 U10355 ( .INP(n10422), .ZN(n10421) );
  NOR2X0 U10356 ( .IN1(n10423), .IN2(n10424), .QN(n10422) );
  NAND2X0 U10357 ( .IN1(n10424), .IN2(n10423), .QN(n10420) );
  NOR2X0 U10358 ( .IN1(n10425), .IN2(n10426), .QN(n10423) );
  NOR2X0 U10359 ( .IN1(WX9942), .IN2(n7892), .QN(n10426) );
  INVX0 U10360 ( .INP(n10427), .ZN(n10425) );
  NAND2X0 U10361 ( .IN1(n7892), .IN2(WX9942), .QN(n10427) );
  NAND2X0 U10362 ( .IN1(n10428), .IN2(n10429), .QN(n10424) );
  NAND2X0 U10363 ( .IN1(n7891), .IN2(WX9814), .QN(n10429) );
  INVX0 U10364 ( .INP(n10430), .ZN(n10428) );
  NOR2X0 U10365 ( .IN1(WX9814), .IN2(n7891), .QN(n10430) );
  NAND2X0 U10366 ( .IN1(n9099), .IN2(n10431), .QN(n10418) );
  NAND2X0 U10367 ( .IN1(n1482), .IN2(n9275), .QN(n10417) );
  NOR2X0 U10368 ( .IN1(n9228), .IN2(n8861), .QN(n1482) );
  NAND2X0 U10369 ( .IN1(n9306), .IN2(CRC_OUT_3_4), .QN(n10416) );
  NAND4X0 U10370 ( .IN1(n10432), .IN2(n10433), .IN3(n10434), .IN4(n10435), 
        .QN(WX8454) );
  NAND2X0 U10371 ( .IN1(n9330), .IN2(n9993), .QN(n10435) );
  NAND2X0 U10372 ( .IN1(n10436), .IN2(n10437), .QN(n9993) );
  INVX0 U10373 ( .INP(n10438), .ZN(n10437) );
  NOR2X0 U10374 ( .IN1(n10439), .IN2(n10440), .QN(n10438) );
  NAND2X0 U10375 ( .IN1(n10440), .IN2(n10439), .QN(n10436) );
  NOR2X0 U10376 ( .IN1(n10441), .IN2(n10442), .QN(n10439) );
  NOR2X0 U10377 ( .IN1(WX9940), .IN2(n7894), .QN(n10442) );
  INVX0 U10378 ( .INP(n10443), .ZN(n10441) );
  NAND2X0 U10379 ( .IN1(n7894), .IN2(WX9940), .QN(n10443) );
  NAND2X0 U10380 ( .IN1(n10444), .IN2(n10445), .QN(n10440) );
  NAND2X0 U10381 ( .IN1(n7893), .IN2(WX9812), .QN(n10445) );
  INVX0 U10382 ( .INP(n10446), .ZN(n10444) );
  NOR2X0 U10383 ( .IN1(WX9812), .IN2(n7893), .QN(n10446) );
  NAND2X0 U10384 ( .IN1(n9099), .IN2(n10447), .QN(n10434) );
  NAND2X0 U10385 ( .IN1(n1481), .IN2(n9275), .QN(n10433) );
  NOR2X0 U10386 ( .IN1(n9228), .IN2(n8862), .QN(n1481) );
  NAND2X0 U10387 ( .IN1(n9306), .IN2(CRC_OUT_3_5), .QN(n10432) );
  NAND4X0 U10388 ( .IN1(n10448), .IN2(n10449), .IN3(n10450), .IN4(n10451), 
        .QN(WX8452) );
  NAND2X0 U10389 ( .IN1(n9330), .IN2(n10001), .QN(n10451) );
  NAND2X0 U10390 ( .IN1(n10452), .IN2(n10453), .QN(n10001) );
  INVX0 U10391 ( .INP(n10454), .ZN(n10453) );
  NOR2X0 U10392 ( .IN1(n10455), .IN2(n10456), .QN(n10454) );
  NAND2X0 U10393 ( .IN1(n10456), .IN2(n10455), .QN(n10452) );
  NOR2X0 U10394 ( .IN1(n10457), .IN2(n10458), .QN(n10455) );
  NOR2X0 U10395 ( .IN1(WX9938), .IN2(n7896), .QN(n10458) );
  INVX0 U10396 ( .INP(n10459), .ZN(n10457) );
  NAND2X0 U10397 ( .IN1(n7896), .IN2(WX9938), .QN(n10459) );
  NAND2X0 U10398 ( .IN1(n10460), .IN2(n10461), .QN(n10456) );
  NAND2X0 U10399 ( .IN1(n7895), .IN2(WX9810), .QN(n10461) );
  INVX0 U10400 ( .INP(n10462), .ZN(n10460) );
  NOR2X0 U10401 ( .IN1(WX9810), .IN2(n7895), .QN(n10462) );
  NAND2X0 U10402 ( .IN1(n9099), .IN2(n10463), .QN(n10450) );
  NAND2X0 U10403 ( .IN1(n1480), .IN2(n9275), .QN(n10449) );
  NOR2X0 U10404 ( .IN1(n9228), .IN2(n8863), .QN(n1480) );
  NAND2X0 U10405 ( .IN1(n9306), .IN2(CRC_OUT_3_6), .QN(n10448) );
  NAND4X0 U10406 ( .IN1(n10464), .IN2(n10465), .IN3(n10466), .IN4(n10467), 
        .QN(WX8450) );
  NAND2X0 U10407 ( .IN1(n9330), .IN2(n10006), .QN(n10467) );
  NAND2X0 U10408 ( .IN1(n10468), .IN2(n10469), .QN(n10006) );
  INVX0 U10409 ( .INP(n10470), .ZN(n10469) );
  NOR2X0 U10410 ( .IN1(n10471), .IN2(n10472), .QN(n10470) );
  NAND2X0 U10411 ( .IN1(n10472), .IN2(n10471), .QN(n10468) );
  NOR2X0 U10412 ( .IN1(n10473), .IN2(n10474), .QN(n10471) );
  NOR2X0 U10413 ( .IN1(WX9936), .IN2(n7898), .QN(n10474) );
  INVX0 U10414 ( .INP(n10475), .ZN(n10473) );
  NAND2X0 U10415 ( .IN1(n7898), .IN2(WX9936), .QN(n10475) );
  NAND2X0 U10416 ( .IN1(n10476), .IN2(n10477), .QN(n10472) );
  NAND2X0 U10417 ( .IN1(n7897), .IN2(WX9808), .QN(n10477) );
  INVX0 U10418 ( .INP(n10478), .ZN(n10476) );
  NOR2X0 U10419 ( .IN1(WX9808), .IN2(n7897), .QN(n10478) );
  NAND2X0 U10420 ( .IN1(n9099), .IN2(n10479), .QN(n10466) );
  NAND2X0 U10421 ( .IN1(n1479), .IN2(n9275), .QN(n10465) );
  NOR2X0 U10422 ( .IN1(n9228), .IN2(n8864), .QN(n1479) );
  NAND2X0 U10423 ( .IN1(test_so76), .IN2(n9315), .QN(n10464) );
  NAND4X0 U10424 ( .IN1(n10480), .IN2(n10481), .IN3(n10482), .IN4(n10483), 
        .QN(WX8448) );
  NAND2X0 U10425 ( .IN1(n9330), .IN2(n10014), .QN(n10483) );
  NAND2X0 U10426 ( .IN1(n10484), .IN2(n10485), .QN(n10014) );
  INVX0 U10427 ( .INP(n10486), .ZN(n10485) );
  NOR2X0 U10428 ( .IN1(n10487), .IN2(n10488), .QN(n10486) );
  NAND2X0 U10429 ( .IN1(n10488), .IN2(n10487), .QN(n10484) );
  NOR2X0 U10430 ( .IN1(n10489), .IN2(n10490), .QN(n10487) );
  NOR2X0 U10431 ( .IN1(WX9934), .IN2(n7900), .QN(n10490) );
  INVX0 U10432 ( .INP(n10491), .ZN(n10489) );
  NAND2X0 U10433 ( .IN1(n7900), .IN2(WX9934), .QN(n10491) );
  NAND2X0 U10434 ( .IN1(n10492), .IN2(n10493), .QN(n10488) );
  NAND2X0 U10435 ( .IN1(n7899), .IN2(WX9806), .QN(n10493) );
  INVX0 U10436 ( .INP(n10494), .ZN(n10492) );
  NOR2X0 U10437 ( .IN1(WX9806), .IN2(n7899), .QN(n10494) );
  NAND2X0 U10438 ( .IN1(n9098), .IN2(n10495), .QN(n10482) );
  NAND2X0 U10439 ( .IN1(n1478), .IN2(n9275), .QN(n10481) );
  NOR2X0 U10440 ( .IN1(n9229), .IN2(n8865), .QN(n1478) );
  NAND2X0 U10441 ( .IN1(n9306), .IN2(CRC_OUT_3_8), .QN(n10480) );
  NAND4X0 U10442 ( .IN1(n10496), .IN2(n10497), .IN3(n10498), .IN4(n10499), 
        .QN(WX8446) );
  NAND3X0 U10443 ( .IN1(n10500), .IN2(n10501), .IN3(n9092), .QN(n10499) );
  NAND2X0 U10444 ( .IN1(n9330), .IN2(n10019), .QN(n10498) );
  NAND2X0 U10445 ( .IN1(n10502), .IN2(n10503), .QN(n10019) );
  INVX0 U10446 ( .INP(n10504), .ZN(n10503) );
  NOR2X0 U10447 ( .IN1(n10505), .IN2(n10506), .QN(n10504) );
  NAND2X0 U10448 ( .IN1(n10506), .IN2(n10505), .QN(n10502) );
  NOR2X0 U10449 ( .IN1(n10507), .IN2(n10508), .QN(n10505) );
  NOR2X0 U10450 ( .IN1(WX9932), .IN2(n7902), .QN(n10508) );
  INVX0 U10451 ( .INP(n10509), .ZN(n10507) );
  NAND2X0 U10452 ( .IN1(n7902), .IN2(WX9932), .QN(n10509) );
  NAND2X0 U10453 ( .IN1(n10510), .IN2(n10511), .QN(n10506) );
  NAND2X0 U10454 ( .IN1(n7901), .IN2(WX9804), .QN(n10511) );
  INVX0 U10455 ( .INP(n10512), .ZN(n10510) );
  NOR2X0 U10456 ( .IN1(WX9804), .IN2(n7901), .QN(n10512) );
  NAND2X0 U10457 ( .IN1(n1477), .IN2(n9275), .QN(n10497) );
  NOR2X0 U10458 ( .IN1(n9230), .IN2(n8866), .QN(n1477) );
  NAND2X0 U10459 ( .IN1(n9306), .IN2(CRC_OUT_3_9), .QN(n10496) );
  NAND4X0 U10460 ( .IN1(n10513), .IN2(n10514), .IN3(n10515), .IN4(n10516), 
        .QN(WX8444) );
  NAND2X0 U10461 ( .IN1(n9330), .IN2(n10025), .QN(n10516) );
  NAND2X0 U10462 ( .IN1(n10517), .IN2(n10518), .QN(n10025) );
  INVX0 U10463 ( .INP(n10519), .ZN(n10518) );
  NOR2X0 U10464 ( .IN1(n10520), .IN2(n10521), .QN(n10519) );
  NAND2X0 U10465 ( .IN1(n10521), .IN2(n10520), .QN(n10517) );
  NOR2X0 U10466 ( .IN1(n10522), .IN2(n10523), .QN(n10520) );
  NOR2X0 U10467 ( .IN1(WX9930), .IN2(n7904), .QN(n10523) );
  INVX0 U10468 ( .INP(n10524), .ZN(n10522) );
  NAND2X0 U10469 ( .IN1(n7904), .IN2(WX9930), .QN(n10524) );
  NAND2X0 U10470 ( .IN1(n10525), .IN2(n10526), .QN(n10521) );
  NAND2X0 U10471 ( .IN1(n7903), .IN2(WX9802), .QN(n10526) );
  INVX0 U10472 ( .INP(n10527), .ZN(n10525) );
  NOR2X0 U10473 ( .IN1(WX9802), .IN2(n7903), .QN(n10527) );
  NAND2X0 U10474 ( .IN1(n9098), .IN2(n10528), .QN(n10515) );
  NAND2X0 U10475 ( .IN1(n1476), .IN2(n9275), .QN(n10514) );
  NOR2X0 U10476 ( .IN1(n9230), .IN2(n8867), .QN(n1476) );
  NAND2X0 U10477 ( .IN1(n9306), .IN2(CRC_OUT_3_10), .QN(n10513) );
  NAND4X0 U10478 ( .IN1(n10529), .IN2(n10530), .IN3(n10531), .IN4(n10532), 
        .QN(WX8442) );
  NAND3X0 U10479 ( .IN1(n10533), .IN2(n10534), .IN3(n9091), .QN(n10532) );
  NAND2X0 U10480 ( .IN1(n9330), .IN2(n10031), .QN(n10531) );
  NAND2X0 U10481 ( .IN1(n10535), .IN2(n10536), .QN(n10031) );
  INVX0 U10482 ( .INP(n10537), .ZN(n10536) );
  NOR2X0 U10483 ( .IN1(n10538), .IN2(n10539), .QN(n10537) );
  NAND2X0 U10484 ( .IN1(n10539), .IN2(n10538), .QN(n10535) );
  NOR2X0 U10485 ( .IN1(n10540), .IN2(n10541), .QN(n10538) );
  NOR2X0 U10486 ( .IN1(WX9928), .IN2(n7906), .QN(n10541) );
  INVX0 U10487 ( .INP(n10542), .ZN(n10540) );
  NAND2X0 U10488 ( .IN1(n7906), .IN2(WX9928), .QN(n10542) );
  NAND2X0 U10489 ( .IN1(n10543), .IN2(n10544), .QN(n10539) );
  NAND2X0 U10490 ( .IN1(n7905), .IN2(WX9800), .QN(n10544) );
  INVX0 U10491 ( .INP(n10545), .ZN(n10543) );
  NOR2X0 U10492 ( .IN1(WX9800), .IN2(n7905), .QN(n10545) );
  NAND2X0 U10493 ( .IN1(n1475), .IN2(n9275), .QN(n10530) );
  NOR2X0 U10494 ( .IN1(n9230), .IN2(n8868), .QN(n1475) );
  NAND2X0 U10495 ( .IN1(n9306), .IN2(CRC_OUT_3_11), .QN(n10529) );
  NAND4X0 U10496 ( .IN1(n10546), .IN2(n10547), .IN3(n10548), .IN4(n10549), 
        .QN(WX8440) );
  NAND2X0 U10497 ( .IN1(n9330), .IN2(n10037), .QN(n10549) );
  NAND2X0 U10498 ( .IN1(n10550), .IN2(n10551), .QN(n10037) );
  INVX0 U10499 ( .INP(n10552), .ZN(n10551) );
  NOR2X0 U10500 ( .IN1(n10553), .IN2(n10554), .QN(n10552) );
  NAND2X0 U10501 ( .IN1(n10554), .IN2(n10553), .QN(n10550) );
  NOR2X0 U10502 ( .IN1(n10555), .IN2(n10556), .QN(n10553) );
  NOR2X0 U10503 ( .IN1(WX9926), .IN2(n7908), .QN(n10556) );
  INVX0 U10504 ( .INP(n10557), .ZN(n10555) );
  NAND2X0 U10505 ( .IN1(n7908), .IN2(WX9926), .QN(n10557) );
  NAND2X0 U10506 ( .IN1(n10558), .IN2(n10559), .QN(n10554) );
  NAND2X0 U10507 ( .IN1(n7907), .IN2(WX9798), .QN(n10559) );
  INVX0 U10508 ( .INP(n10560), .ZN(n10558) );
  NOR2X0 U10509 ( .IN1(WX9798), .IN2(n7907), .QN(n10560) );
  NAND2X0 U10510 ( .IN1(n9098), .IN2(n10561), .QN(n10548) );
  NAND2X0 U10511 ( .IN1(n1474), .IN2(n9275), .QN(n10547) );
  NOR2X0 U10512 ( .IN1(n9230), .IN2(n8869), .QN(n1474) );
  NAND2X0 U10513 ( .IN1(n9306), .IN2(CRC_OUT_3_12), .QN(n10546) );
  NAND4X0 U10514 ( .IN1(n10562), .IN2(n10563), .IN3(n10564), .IN4(n10565), 
        .QN(WX8438) );
  NAND3X0 U10515 ( .IN1(n10566), .IN2(n10567), .IN3(n9092), .QN(n10565) );
  NAND2X0 U10516 ( .IN1(n9330), .IN2(n10043), .QN(n10564) );
  NAND2X0 U10517 ( .IN1(n10568), .IN2(n10569), .QN(n10043) );
  INVX0 U10518 ( .INP(n10570), .ZN(n10569) );
  NOR2X0 U10519 ( .IN1(n10571), .IN2(n10572), .QN(n10570) );
  NAND2X0 U10520 ( .IN1(n10572), .IN2(n10571), .QN(n10568) );
  NOR2X0 U10521 ( .IN1(n10573), .IN2(n10574), .QN(n10571) );
  NOR2X0 U10522 ( .IN1(WX9924), .IN2(n7910), .QN(n10574) );
  INVX0 U10523 ( .INP(n10575), .ZN(n10573) );
  NAND2X0 U10524 ( .IN1(n7910), .IN2(WX9924), .QN(n10575) );
  NAND2X0 U10525 ( .IN1(n10576), .IN2(n10577), .QN(n10572) );
  NAND2X0 U10526 ( .IN1(n7909), .IN2(WX9796), .QN(n10577) );
  INVX0 U10527 ( .INP(n10578), .ZN(n10576) );
  NOR2X0 U10528 ( .IN1(WX9796), .IN2(n7909), .QN(n10578) );
  NAND2X0 U10529 ( .IN1(n1473), .IN2(n9275), .QN(n10563) );
  NOR2X0 U10530 ( .IN1(n9230), .IN2(n8870), .QN(n1473) );
  NAND2X0 U10531 ( .IN1(n9307), .IN2(CRC_OUT_3_13), .QN(n10562) );
  NAND4X0 U10532 ( .IN1(n10579), .IN2(n10580), .IN3(n10581), .IN4(n10582), 
        .QN(WX8436) );
  NAND3X0 U10533 ( .IN1(n10049), .IN2(n10050), .IN3(n9322), .QN(n10582) );
  NAND3X0 U10534 ( .IN1(n10583), .IN2(n10584), .IN3(n10585), .QN(n10050) );
  INVX0 U10535 ( .INP(n10586), .ZN(n10585) );
  NAND2X0 U10536 ( .IN1(n10586), .IN2(n10587), .QN(n10049) );
  NAND2X0 U10537 ( .IN1(n10583), .IN2(n10584), .QN(n10587) );
  NAND2X0 U10538 ( .IN1(n7912), .IN2(WX9794), .QN(n10584) );
  NAND2X0 U10539 ( .IN1(n3591), .IN2(WX9858), .QN(n10583) );
  NOR2X0 U10540 ( .IN1(n10588), .IN2(n10589), .QN(n10586) );
  NOR2X0 U10541 ( .IN1(n8795), .IN2(n7911), .QN(n10589) );
  INVX0 U10542 ( .INP(n10590), .ZN(n10588) );
  NAND2X0 U10543 ( .IN1(n7911), .IN2(n8795), .QN(n10590) );
  NAND2X0 U10544 ( .IN1(n9098), .IN2(n10591), .QN(n10581) );
  NAND2X0 U10545 ( .IN1(n1472), .IN2(n9275), .QN(n10580) );
  NOR2X0 U10546 ( .IN1(n9230), .IN2(n8871), .QN(n1472) );
  NAND2X0 U10547 ( .IN1(n9307), .IN2(CRC_OUT_3_14), .QN(n10579) );
  NAND4X0 U10548 ( .IN1(n10592), .IN2(n10593), .IN3(n10594), .IN4(n10595), 
        .QN(WX8434) );
  NAND3X0 U10549 ( .IN1(n10596), .IN2(n10597), .IN3(n9092), .QN(n10595) );
  NAND2X0 U10550 ( .IN1(n9331), .IN2(n10056), .QN(n10594) );
  NAND2X0 U10551 ( .IN1(n10598), .IN2(n10599), .QN(n10056) );
  INVX0 U10552 ( .INP(n10600), .ZN(n10599) );
  NOR2X0 U10553 ( .IN1(n10601), .IN2(n10602), .QN(n10600) );
  NAND2X0 U10554 ( .IN1(n10602), .IN2(n10601), .QN(n10598) );
  NOR2X0 U10555 ( .IN1(n10603), .IN2(n10604), .QN(n10601) );
  NOR2X0 U10556 ( .IN1(WX9920), .IN2(n7914), .QN(n10604) );
  INVX0 U10557 ( .INP(n10605), .ZN(n10603) );
  NAND2X0 U10558 ( .IN1(n7914), .IN2(WX9920), .QN(n10605) );
  NAND2X0 U10559 ( .IN1(n10606), .IN2(n10607), .QN(n10602) );
  NAND2X0 U10560 ( .IN1(n7913), .IN2(WX9792), .QN(n10607) );
  INVX0 U10561 ( .INP(n10608), .ZN(n10606) );
  NOR2X0 U10562 ( .IN1(WX9792), .IN2(n7913), .QN(n10608) );
  NAND2X0 U10563 ( .IN1(n1471), .IN2(n9275), .QN(n10593) );
  NOR2X0 U10564 ( .IN1(n9231), .IN2(n8872), .QN(n1471) );
  NAND2X0 U10565 ( .IN1(n9307), .IN2(CRC_OUT_3_15), .QN(n10592) );
  NAND4X0 U10566 ( .IN1(n10609), .IN2(n10610), .IN3(n10611), .IN4(n10612), 
        .QN(WX8432) );
  NAND2X0 U10567 ( .IN1(n10613), .IN2(n10614), .QN(n10612) );
  NAND2X0 U10568 ( .IN1(n10615), .IN2(n10616), .QN(n10613) );
  NAND2X0 U10569 ( .IN1(n9098), .IN2(n10617), .QN(n10616) );
  NAND2X0 U10570 ( .IN1(n9098), .IN2(n8363), .QN(n10615) );
  NAND2X0 U10571 ( .IN1(n10070), .IN2(n2153), .QN(n10611) );
  NOR2X0 U10572 ( .IN1(n10618), .IN2(n10619), .QN(n10070) );
  INVX0 U10573 ( .INP(n10620), .ZN(n10619) );
  NAND2X0 U10574 ( .IN1(n10621), .IN2(n10622), .QN(n10620) );
  NOR2X0 U10575 ( .IN1(n10622), .IN2(n10621), .QN(n10618) );
  NAND2X0 U10576 ( .IN1(n10623), .IN2(n10624), .QN(n10621) );
  NAND2X0 U10577 ( .IN1(n8108), .IN2(n10625), .QN(n10624) );
  INVX0 U10578 ( .INP(n10626), .ZN(n10625) );
  NAND2X0 U10579 ( .IN1(n10626), .IN2(WX9918), .QN(n10623) );
  NAND2X0 U10580 ( .IN1(n10627), .IN2(n10628), .QN(n10626) );
  INVX0 U10581 ( .INP(n10629), .ZN(n10628) );
  NOR2X0 U10582 ( .IN1(n8806), .IN2(n16412), .QN(n10629) );
  NAND2X0 U10583 ( .IN1(n16412), .IN2(n8806), .QN(n10627) );
  NOR2X0 U10584 ( .IN1(n10630), .IN2(n10631), .QN(n10622) );
  INVX0 U10585 ( .INP(n10632), .ZN(n10631) );
  NAND2X0 U10586 ( .IN1(n7656), .IN2(n9121), .QN(n10632) );
  NOR2X0 U10587 ( .IN1(n9116), .IN2(n7656), .QN(n10630) );
  NAND2X0 U10588 ( .IN1(n1470), .IN2(n9275), .QN(n10610) );
  NOR2X0 U10589 ( .IN1(n9231), .IN2(n8873), .QN(n1470) );
  NAND2X0 U10590 ( .IN1(n9307), .IN2(CRC_OUT_3_16), .QN(n10609) );
  NAND4X0 U10591 ( .IN1(n10634), .IN2(n10635), .IN3(n10636), .IN4(n10637), 
        .QN(WX8430) );
  NAND2X0 U10592 ( .IN1(n10638), .IN2(n10076), .QN(n10637) );
  NAND2X0 U10593 ( .IN1(n10639), .IN2(n10079), .QN(n10076) );
  NAND2X0 U10594 ( .IN1(n10640), .IN2(n10641), .QN(n10639) );
  NAND2X0 U10595 ( .IN1(n16411), .IN2(n9121), .QN(n10641) );
  NAND2X0 U10596 ( .IN1(TM1), .IN2(n8305), .QN(n10640) );
  NAND3X0 U10597 ( .IN1(n10642), .IN2(n10643), .IN3(n10644), .QN(n10638) );
  NAND2X0 U10598 ( .IN1(n9331), .IN2(n10079), .QN(n10644) );
  NAND2X0 U10599 ( .IN1(n10645), .IN2(n10646), .QN(n10079) );
  NAND2X0 U10600 ( .IN1(n7657), .IN2(n10647), .QN(n10646) );
  INVX0 U10601 ( .INP(n10648), .ZN(n10645) );
  NOR2X0 U10602 ( .IN1(n10647), .IN2(n7657), .QN(n10648) );
  NOR2X0 U10603 ( .IN1(n10649), .IN2(n10650), .QN(n10647) );
  NOR2X0 U10604 ( .IN1(WX9916), .IN2(n7658), .QN(n10650) );
  INVX0 U10605 ( .INP(n10651), .ZN(n10649) );
  NAND2X0 U10606 ( .IN1(n7658), .IN2(WX9916), .QN(n10651) );
  NAND2X0 U10607 ( .IN1(n9083), .IN2(n8305), .QN(n10643) );
  NAND2X0 U10608 ( .IN1(n16411), .IN2(n10069), .QN(n10642) );
  NAND2X0 U10609 ( .IN1(n10652), .IN2(n10653), .QN(n10636) );
  NAND2X0 U10610 ( .IN1(n10654), .IN2(n10655), .QN(n10652) );
  NAND2X0 U10611 ( .IN1(n9098), .IN2(n10656), .QN(n10655) );
  NAND2X0 U10612 ( .IN1(n9098), .IN2(n8364), .QN(n10654) );
  NAND2X0 U10613 ( .IN1(n1469), .IN2(n9275), .QN(n10635) );
  NOR2X0 U10614 ( .IN1(n9064), .IN2(n9156), .QN(n1469) );
  NAND2X0 U10615 ( .IN1(n9307), .IN2(CRC_OUT_3_17), .QN(n10634) );
  NAND4X0 U10616 ( .IN1(n10657), .IN2(n10658), .IN3(n10659), .IN4(n10660), 
        .QN(WX8428) );
  NAND2X0 U10617 ( .IN1(n10661), .IN2(n10662), .QN(n10660) );
  NAND2X0 U10618 ( .IN1(n10663), .IN2(n10664), .QN(n10661) );
  NAND2X0 U10619 ( .IN1(n9098), .IN2(n10665), .QN(n10664) );
  NAND2X0 U10620 ( .IN1(n9098), .IN2(n8365), .QN(n10663) );
  NAND2X0 U10621 ( .IN1(n10096), .IN2(n2153), .QN(n10659) );
  NOR2X0 U10622 ( .IN1(n10666), .IN2(n10667), .QN(n10096) );
  INVX0 U10623 ( .INP(n10668), .ZN(n10667) );
  NAND2X0 U10624 ( .IN1(n10669), .IN2(n10670), .QN(n10668) );
  NOR2X0 U10625 ( .IN1(n10670), .IN2(n10669), .QN(n10666) );
  NAND2X0 U10626 ( .IN1(n10671), .IN2(n10672), .QN(n10669) );
  NAND2X0 U10627 ( .IN1(n8172), .IN2(n10673), .QN(n10672) );
  INVX0 U10628 ( .INP(n10674), .ZN(n10673) );
  NAND2X0 U10629 ( .IN1(n10674), .IN2(WX9914), .QN(n10671) );
  NAND2X0 U10630 ( .IN1(n10675), .IN2(n10676), .QN(n10674) );
  INVX0 U10631 ( .INP(n10677), .ZN(n10676) );
  NOR2X0 U10632 ( .IN1(n8807), .IN2(n16410), .QN(n10677) );
  NAND2X0 U10633 ( .IN1(n16410), .IN2(n8807), .QN(n10675) );
  NOR2X0 U10634 ( .IN1(n10678), .IN2(n10679), .QN(n10670) );
  INVX0 U10635 ( .INP(n10680), .ZN(n10679) );
  NAND2X0 U10636 ( .IN1(n7659), .IN2(n9121), .QN(n10680) );
  NOR2X0 U10637 ( .IN1(n9116), .IN2(n7659), .QN(n10678) );
  NAND2X0 U10638 ( .IN1(n509), .IN2(n9275), .QN(n10658) );
  NOR2X0 U10639 ( .IN1(n10681), .IN2(n8874), .QN(n509) );
  NAND2X0 U10640 ( .IN1(n9307), .IN2(CRC_OUT_3_18), .QN(n10657) );
  NAND4X0 U10641 ( .IN1(n10682), .IN2(n10683), .IN3(n10684), .IN4(n10685), 
        .QN(WX8426) );
  NAND2X0 U10642 ( .IN1(n10686), .IN2(n10102), .QN(n10685) );
  NAND2X0 U10643 ( .IN1(n10687), .IN2(n10105), .QN(n10102) );
  NAND2X0 U10644 ( .IN1(n10688), .IN2(n10689), .QN(n10687) );
  NAND2X0 U10645 ( .IN1(n16409), .IN2(n9121), .QN(n10689) );
  NAND2X0 U10646 ( .IN1(TM1), .IN2(n8307), .QN(n10688) );
  NAND3X0 U10647 ( .IN1(n10690), .IN2(n10691), .IN3(n10692), .QN(n10686) );
  NAND2X0 U10648 ( .IN1(n9331), .IN2(n10105), .QN(n10692) );
  NAND2X0 U10649 ( .IN1(n10693), .IN2(n10694), .QN(n10105) );
  NAND2X0 U10650 ( .IN1(n7660), .IN2(n10695), .QN(n10694) );
  INVX0 U10651 ( .INP(n10696), .ZN(n10693) );
  NOR2X0 U10652 ( .IN1(n10695), .IN2(n7660), .QN(n10696) );
  NOR2X0 U10653 ( .IN1(n10697), .IN2(n10698), .QN(n10695) );
  NOR2X0 U10654 ( .IN1(WX9912), .IN2(n7661), .QN(n10698) );
  INVX0 U10655 ( .INP(n10699), .ZN(n10697) );
  NAND2X0 U10656 ( .IN1(n7661), .IN2(WX9912), .QN(n10699) );
  NAND2X0 U10657 ( .IN1(n9082), .IN2(n8307), .QN(n10691) );
  NAND2X0 U10658 ( .IN1(n16409), .IN2(n9080), .QN(n10690) );
  NAND2X0 U10659 ( .IN1(n10700), .IN2(n10701), .QN(n10684) );
  NAND2X0 U10660 ( .IN1(n10702), .IN2(n10703), .QN(n10700) );
  NAND2X0 U10661 ( .IN1(n9098), .IN2(n10704), .QN(n10703) );
  NAND2X0 U10662 ( .IN1(n9098), .IN2(n8366), .QN(n10702) );
  NAND2X0 U10663 ( .IN1(n1468), .IN2(n9276), .QN(n10683) );
  NOR2X0 U10664 ( .IN1(n9231), .IN2(n8875), .QN(n1468) );
  NAND2X0 U10665 ( .IN1(n9307), .IN2(CRC_OUT_3_19), .QN(n10682) );
  NAND4X0 U10666 ( .IN1(n10705), .IN2(n10706), .IN3(n10707), .IN4(n10708), 
        .QN(WX8424) );
  NAND2X0 U10667 ( .IN1(n10709), .IN2(n10112), .QN(n10708) );
  NAND3X0 U10668 ( .IN1(n10710), .IN2(n10711), .IN3(n10115), .QN(n10112) );
  NAND2X0 U10669 ( .IN1(n8170), .IN2(n9121), .QN(n10711) );
  NAND2X0 U10670 ( .IN1(TM1), .IN2(WX9910), .QN(n10710) );
  NAND3X0 U10671 ( .IN1(n10712), .IN2(n10713), .IN3(n10714), .QN(n10709) );
  NAND2X0 U10672 ( .IN1(n9331), .IN2(n10115), .QN(n10714) );
  NAND2X0 U10673 ( .IN1(n10715), .IN2(n10716), .QN(n10115) );
  NAND2X0 U10674 ( .IN1(n10717), .IN2(WX9846), .QN(n10716) );
  NAND2X0 U10675 ( .IN1(n10718), .IN2(n10719), .QN(n10717) );
  NAND3X0 U10676 ( .IN1(n10718), .IN2(n10719), .IN3(n7663), .QN(n10715) );
  NAND2X0 U10677 ( .IN1(test_so80), .IN2(WX9782), .QN(n10719) );
  NAND2X0 U10678 ( .IN1(n7662), .IN2(n8820), .QN(n10718) );
  NAND2X0 U10679 ( .IN1(n9080), .IN2(WX9910), .QN(n10713) );
  NAND2X0 U10680 ( .IN1(n10068), .IN2(n8170), .QN(n10712) );
  NAND2X0 U10681 ( .IN1(n10720), .IN2(n10721), .QN(n10707) );
  NAND2X0 U10682 ( .IN1(n10722), .IN2(n10723), .QN(n10720) );
  NAND2X0 U10683 ( .IN1(n9098), .IN2(n10724), .QN(n10723) );
  NAND2X0 U10684 ( .IN1(n9098), .IN2(n8367), .QN(n10722) );
  NAND2X0 U10685 ( .IN1(n1467), .IN2(n9276), .QN(n10706) );
  NOR2X0 U10686 ( .IN1(n9231), .IN2(n8876), .QN(n1467) );
  NAND2X0 U10687 ( .IN1(n9307), .IN2(CRC_OUT_3_20), .QN(n10705) );
  NAND4X0 U10688 ( .IN1(n10725), .IN2(n10726), .IN3(n10727), .IN4(n10728), 
        .QN(WX8422) );
  NAND2X0 U10689 ( .IN1(n10729), .IN2(n10127), .QN(n10728) );
  NAND2X0 U10690 ( .IN1(n10730), .IN2(n10130), .QN(n10127) );
  NAND2X0 U10691 ( .IN1(n10731), .IN2(n10732), .QN(n10730) );
  NAND2X0 U10692 ( .IN1(n16408), .IN2(n9121), .QN(n10732) );
  NAND2X0 U10693 ( .IN1(TM1), .IN2(n8310), .QN(n10731) );
  NAND3X0 U10694 ( .IN1(n10733), .IN2(n10734), .IN3(n10735), .QN(n10729) );
  NAND2X0 U10695 ( .IN1(n9331), .IN2(n10130), .QN(n10735) );
  NAND2X0 U10696 ( .IN1(n10736), .IN2(n10737), .QN(n10130) );
  NAND2X0 U10697 ( .IN1(n7664), .IN2(n10738), .QN(n10737) );
  INVX0 U10698 ( .INP(n10739), .ZN(n10736) );
  NOR2X0 U10699 ( .IN1(n10738), .IN2(n7664), .QN(n10739) );
  NOR2X0 U10700 ( .IN1(n10740), .IN2(n10741), .QN(n10738) );
  NOR2X0 U10701 ( .IN1(WX9908), .IN2(n7665), .QN(n10741) );
  INVX0 U10702 ( .INP(n10742), .ZN(n10740) );
  NAND2X0 U10703 ( .IN1(n7665), .IN2(WX9908), .QN(n10742) );
  NAND2X0 U10704 ( .IN1(n9084), .IN2(n8310), .QN(n10734) );
  NAND2X0 U10705 ( .IN1(n16408), .IN2(n9079), .QN(n10733) );
  NAND2X0 U10706 ( .IN1(n10743), .IN2(n10744), .QN(n10727) );
  NAND2X0 U10707 ( .IN1(n10745), .IN2(n10746), .QN(n10743) );
  NAND2X0 U10708 ( .IN1(n9098), .IN2(n10747), .QN(n10746) );
  NAND2X0 U10709 ( .IN1(n9098), .IN2(n8368), .QN(n10745) );
  NAND2X0 U10710 ( .IN1(n1466), .IN2(n9276), .QN(n10726) );
  NOR2X0 U10711 ( .IN1(n9231), .IN2(n8877), .QN(n1466) );
  NAND2X0 U10712 ( .IN1(n9307), .IN2(CRC_OUT_3_21), .QN(n10725) );
  NAND4X0 U10713 ( .IN1(n10748), .IN2(n10749), .IN3(n10750), .IN4(n10751), 
        .QN(WX8420) );
  NAND2X0 U10714 ( .IN1(n10752), .IN2(n10137), .QN(n10751) );
  NAND2X0 U10715 ( .IN1(n10753), .IN2(n10140), .QN(n10137) );
  NAND2X0 U10716 ( .IN1(n10754), .IN2(n10755), .QN(n10753) );
  NAND2X0 U10717 ( .IN1(n16407), .IN2(n9121), .QN(n10755) );
  NAND2X0 U10718 ( .IN1(TM1), .IN2(n8311), .QN(n10754) );
  NAND3X0 U10719 ( .IN1(n10756), .IN2(n10757), .IN3(n10758), .QN(n10752) );
  NAND2X0 U10720 ( .IN1(n9331), .IN2(n10140), .QN(n10758) );
  NAND2X0 U10721 ( .IN1(n10759), .IN2(n10760), .QN(n10140) );
  NAND2X0 U10722 ( .IN1(n7666), .IN2(n10761), .QN(n10760) );
  INVX0 U10723 ( .INP(n10762), .ZN(n10759) );
  NOR2X0 U10724 ( .IN1(n10761), .IN2(n7666), .QN(n10762) );
  NOR2X0 U10725 ( .IN1(n10763), .IN2(n10764), .QN(n10761) );
  NOR2X0 U10726 ( .IN1(WX9906), .IN2(n7667), .QN(n10764) );
  INVX0 U10727 ( .INP(n10765), .ZN(n10763) );
  NAND2X0 U10728 ( .IN1(n7667), .IN2(WX9906), .QN(n10765) );
  NAND2X0 U10729 ( .IN1(n9083), .IN2(n8311), .QN(n10757) );
  NAND2X0 U10730 ( .IN1(n16407), .IN2(n9078), .QN(n10756) );
  NAND2X0 U10731 ( .IN1(n10766), .IN2(n10767), .QN(n10750) );
  NAND2X0 U10732 ( .IN1(n10768), .IN2(n10769), .QN(n10766) );
  NAND2X0 U10733 ( .IN1(n9098), .IN2(n10770), .QN(n10769) );
  NAND2X0 U10734 ( .IN1(n9098), .IN2(n8369), .QN(n10768) );
  NAND2X0 U10735 ( .IN1(n1465), .IN2(n9276), .QN(n10749) );
  NOR2X0 U10736 ( .IN1(n9231), .IN2(n8878), .QN(n1465) );
  NAND2X0 U10737 ( .IN1(n9307), .IN2(CRC_OUT_3_22), .QN(n10748) );
  NAND4X0 U10738 ( .IN1(n10771), .IN2(n10772), .IN3(n10773), .IN4(n10774), 
        .QN(WX8418) );
  NAND2X0 U10739 ( .IN1(n10775), .IN2(n10152), .QN(n10774) );
  NAND2X0 U10740 ( .IN1(n10776), .IN2(n10155), .QN(n10152) );
  NAND2X0 U10741 ( .IN1(n10777), .IN2(n10778), .QN(n10776) );
  NAND2X0 U10742 ( .IN1(n16406), .IN2(n9120), .QN(n10778) );
  NAND2X0 U10743 ( .IN1(TM1), .IN2(n8312), .QN(n10777) );
  NAND3X0 U10744 ( .IN1(n10779), .IN2(n10780), .IN3(n10781), .QN(n10775) );
  NAND2X0 U10745 ( .IN1(n9331), .IN2(n10155), .QN(n10781) );
  NAND2X0 U10746 ( .IN1(n10782), .IN2(n10783), .QN(n10155) );
  NAND2X0 U10747 ( .IN1(n7668), .IN2(n10784), .QN(n10783) );
  INVX0 U10748 ( .INP(n10785), .ZN(n10782) );
  NOR2X0 U10749 ( .IN1(n10784), .IN2(n7668), .QN(n10785) );
  NOR2X0 U10750 ( .IN1(n10786), .IN2(n10787), .QN(n10784) );
  NOR2X0 U10751 ( .IN1(WX9904), .IN2(n7669), .QN(n10787) );
  INVX0 U10752 ( .INP(n10788), .ZN(n10786) );
  NAND2X0 U10753 ( .IN1(n7669), .IN2(WX9904), .QN(n10788) );
  NAND2X0 U10754 ( .IN1(n9082), .IN2(n8312), .QN(n10780) );
  NAND2X0 U10755 ( .IN1(n16406), .IN2(n10069), .QN(n10779) );
  NAND2X0 U10756 ( .IN1(n10789), .IN2(n10790), .QN(n10773) );
  NAND2X0 U10757 ( .IN1(n10791), .IN2(n10792), .QN(n10789) );
  NAND2X0 U10758 ( .IN1(n9097), .IN2(n10793), .QN(n10792) );
  NAND2X0 U10759 ( .IN1(n9097), .IN2(n8370), .QN(n10791) );
  NAND2X0 U10760 ( .IN1(n1464), .IN2(n9276), .QN(n10772) );
  NOR2X0 U10761 ( .IN1(n9231), .IN2(n8879), .QN(n1464) );
  NAND2X0 U10762 ( .IN1(n9307), .IN2(CRC_OUT_3_23), .QN(n10771) );
  NAND4X0 U10763 ( .IN1(n10794), .IN2(n10795), .IN3(n10796), .IN4(n10797), 
        .QN(WX8416) );
  NAND2X0 U10764 ( .IN1(n10798), .IN2(n10162), .QN(n10797) );
  NAND2X0 U10765 ( .IN1(n10799), .IN2(n10165), .QN(n10162) );
  NAND2X0 U10766 ( .IN1(n10800), .IN2(n10801), .QN(n10799) );
  NAND2X0 U10767 ( .IN1(n16405), .IN2(n9120), .QN(n10801) );
  NAND2X0 U10768 ( .IN1(TM1), .IN2(n8313), .QN(n10800) );
  NAND3X0 U10769 ( .IN1(n10802), .IN2(n10803), .IN3(n10804), .QN(n10798) );
  NAND2X0 U10770 ( .IN1(n9331), .IN2(n10165), .QN(n10804) );
  NAND2X0 U10771 ( .IN1(n10805), .IN2(n10806), .QN(n10165) );
  NAND2X0 U10772 ( .IN1(n7670), .IN2(n10807), .QN(n10806) );
  INVX0 U10773 ( .INP(n10808), .ZN(n10805) );
  NOR2X0 U10774 ( .IN1(n10807), .IN2(n7670), .QN(n10808) );
  NOR2X0 U10775 ( .IN1(n10809), .IN2(n10810), .QN(n10807) );
  NOR2X0 U10776 ( .IN1(WX9902), .IN2(n7671), .QN(n10810) );
  INVX0 U10777 ( .INP(n10811), .ZN(n10809) );
  NAND2X0 U10778 ( .IN1(n7671), .IN2(WX9902), .QN(n10811) );
  NAND2X0 U10779 ( .IN1(n10068), .IN2(n8313), .QN(n10803) );
  NAND2X0 U10780 ( .IN1(n16405), .IN2(n9080), .QN(n10802) );
  NAND2X0 U10781 ( .IN1(n10812), .IN2(n10813), .QN(n10796) );
  NAND2X0 U10782 ( .IN1(n10814), .IN2(n10815), .QN(n10812) );
  NAND2X0 U10783 ( .IN1(n9097), .IN2(n10816), .QN(n10815) );
  NAND2X0 U10784 ( .IN1(n9097), .IN2(n8371), .QN(n10814) );
  NAND2X0 U10785 ( .IN1(n1463), .IN2(n9276), .QN(n10795) );
  NOR2X0 U10786 ( .IN1(n9231), .IN2(n8880), .QN(n1463) );
  NAND2X0 U10787 ( .IN1(test_so77), .IN2(n9314), .QN(n10794) );
  NAND4X0 U10788 ( .IN1(n10817), .IN2(n10818), .IN3(n10819), .IN4(n10820), 
        .QN(WX8414) );
  NAND2X0 U10789 ( .IN1(n10821), .IN2(n10177), .QN(n10820) );
  NAND2X0 U10790 ( .IN1(n10822), .IN2(n10180), .QN(n10177) );
  NAND2X0 U10791 ( .IN1(n10823), .IN2(n10824), .QN(n10822) );
  NAND2X0 U10792 ( .IN1(n16404), .IN2(n9120), .QN(n10824) );
  NAND2X0 U10793 ( .IN1(TM1), .IN2(n8314), .QN(n10823) );
  NAND3X0 U10794 ( .IN1(n10825), .IN2(n10826), .IN3(n10827), .QN(n10821) );
  NAND2X0 U10795 ( .IN1(n9331), .IN2(n10180), .QN(n10827) );
  NAND2X0 U10796 ( .IN1(n10828), .IN2(n10829), .QN(n10180) );
  NAND2X0 U10797 ( .IN1(n7672), .IN2(n10830), .QN(n10829) );
  INVX0 U10798 ( .INP(n10831), .ZN(n10828) );
  NOR2X0 U10799 ( .IN1(n10830), .IN2(n7672), .QN(n10831) );
  NOR2X0 U10800 ( .IN1(n10832), .IN2(n10833), .QN(n10830) );
  NOR2X0 U10801 ( .IN1(WX9900), .IN2(n7673), .QN(n10833) );
  INVX0 U10802 ( .INP(n10834), .ZN(n10832) );
  NAND2X0 U10803 ( .IN1(n7673), .IN2(WX9900), .QN(n10834) );
  NAND2X0 U10804 ( .IN1(n9084), .IN2(n8314), .QN(n10826) );
  NAND2X0 U10805 ( .IN1(n16404), .IN2(n9079), .QN(n10825) );
  NAND2X0 U10806 ( .IN1(n10835), .IN2(n10836), .QN(n10819) );
  NAND2X0 U10807 ( .IN1(n10837), .IN2(n10838), .QN(n10835) );
  NAND2X0 U10808 ( .IN1(n9097), .IN2(n10839), .QN(n10838) );
  NAND2X0 U10809 ( .IN1(n9097), .IN2(n8372), .QN(n10837) );
  NAND2X0 U10810 ( .IN1(n1462), .IN2(n9276), .QN(n10818) );
  NOR2X0 U10811 ( .IN1(n9231), .IN2(n8881), .QN(n1462) );
  NAND2X0 U10812 ( .IN1(n9307), .IN2(CRC_OUT_3_25), .QN(n10817) );
  NAND4X0 U10813 ( .IN1(n10840), .IN2(n10841), .IN3(n10842), .IN4(n10843), 
        .QN(WX8412) );
  NAND2X0 U10814 ( .IN1(n10844), .IN2(n10192), .QN(n10843) );
  NAND2X0 U10815 ( .IN1(n10845), .IN2(n10195), .QN(n10192) );
  NAND2X0 U10816 ( .IN1(n10846), .IN2(n10847), .QN(n10845) );
  NAND2X0 U10817 ( .IN1(n16403), .IN2(n9120), .QN(n10847) );
  NAND2X0 U10818 ( .IN1(TM1), .IN2(n8315), .QN(n10846) );
  NAND3X0 U10819 ( .IN1(n10848), .IN2(n10849), .IN3(n10850), .QN(n10844) );
  NAND2X0 U10820 ( .IN1(n9331), .IN2(n10195), .QN(n10850) );
  NAND2X0 U10821 ( .IN1(n10851), .IN2(n10852), .QN(n10195) );
  NAND2X0 U10822 ( .IN1(n7674), .IN2(n10853), .QN(n10852) );
  INVX0 U10823 ( .INP(n10854), .ZN(n10851) );
  NOR2X0 U10824 ( .IN1(n10853), .IN2(n7674), .QN(n10854) );
  NOR2X0 U10825 ( .IN1(n10855), .IN2(n10856), .QN(n10853) );
  NOR2X0 U10826 ( .IN1(WX9898), .IN2(n7675), .QN(n10856) );
  INVX0 U10827 ( .INP(n10857), .ZN(n10855) );
  NAND2X0 U10828 ( .IN1(n7675), .IN2(WX9898), .QN(n10857) );
  NAND2X0 U10829 ( .IN1(n9083), .IN2(n8315), .QN(n10849) );
  NAND2X0 U10830 ( .IN1(n16403), .IN2(n9078), .QN(n10848) );
  NAND2X0 U10831 ( .IN1(n10858), .IN2(n9110), .QN(n10842) );
  NAND2X0 U10832 ( .IN1(n1461), .IN2(n9276), .QN(n10841) );
  NOR2X0 U10833 ( .IN1(n9232), .IN2(n8882), .QN(n1461) );
  NAND2X0 U10834 ( .IN1(n9308), .IN2(CRC_OUT_3_26), .QN(n10840) );
  NAND4X0 U10835 ( .IN1(n10859), .IN2(n10860), .IN3(n10861), .IN4(n10862), 
        .QN(WX8410) );
  NAND2X0 U10836 ( .IN1(n10863), .IN2(n10207), .QN(n10862) );
  NAND2X0 U10837 ( .IN1(n10864), .IN2(n10210), .QN(n10207) );
  NAND2X0 U10838 ( .IN1(n10865), .IN2(n10866), .QN(n10864) );
  NAND2X0 U10839 ( .IN1(n16402), .IN2(n9120), .QN(n10866) );
  NAND2X0 U10840 ( .IN1(TM1), .IN2(n8316), .QN(n10865) );
  NAND3X0 U10841 ( .IN1(n10867), .IN2(n10868), .IN3(n10869), .QN(n10863) );
  NAND2X0 U10842 ( .IN1(n9331), .IN2(n10210), .QN(n10869) );
  NAND2X0 U10843 ( .IN1(n10870), .IN2(n10871), .QN(n10210) );
  NAND2X0 U10844 ( .IN1(n7676), .IN2(n10872), .QN(n10871) );
  INVX0 U10845 ( .INP(n10873), .ZN(n10870) );
  NOR2X0 U10846 ( .IN1(n10872), .IN2(n7676), .QN(n10873) );
  NOR2X0 U10847 ( .IN1(n10874), .IN2(n10875), .QN(n10872) );
  NOR2X0 U10848 ( .IN1(WX9896), .IN2(n7677), .QN(n10875) );
  INVX0 U10849 ( .INP(n10876), .ZN(n10874) );
  NAND2X0 U10850 ( .IN1(n7677), .IN2(WX9896), .QN(n10876) );
  NAND2X0 U10851 ( .IN1(n9082), .IN2(n8316), .QN(n10868) );
  NAND2X0 U10852 ( .IN1(n16402), .IN2(n10069), .QN(n10867) );
  NAND2X0 U10853 ( .IN1(n10877), .IN2(n10878), .QN(n10861) );
  NAND2X0 U10854 ( .IN1(n10879), .IN2(n10880), .QN(n10877) );
  NAND2X0 U10855 ( .IN1(n9097), .IN2(n10881), .QN(n10880) );
  NAND2X0 U10856 ( .IN1(n9097), .IN2(n8374), .QN(n10879) );
  NAND2X0 U10857 ( .IN1(n1460), .IN2(n9276), .QN(n10860) );
  NOR2X0 U10858 ( .IN1(n9232), .IN2(n8883), .QN(n1460) );
  NAND2X0 U10859 ( .IN1(n9308), .IN2(CRC_OUT_3_27), .QN(n10859) );
  NAND4X0 U10860 ( .IN1(n10882), .IN2(n10883), .IN3(n10884), .IN4(n10885), 
        .QN(WX8408) );
  NAND2X0 U10861 ( .IN1(n10886), .IN2(n10222), .QN(n10885) );
  NAND2X0 U10862 ( .IN1(n10887), .IN2(n10225), .QN(n10222) );
  NAND2X0 U10863 ( .IN1(n10888), .IN2(n10889), .QN(n10887) );
  NAND2X0 U10864 ( .IN1(n16401), .IN2(n9120), .QN(n10889) );
  NAND2X0 U10865 ( .IN1(TM1), .IN2(n8317), .QN(n10888) );
  NAND3X0 U10866 ( .IN1(n10890), .IN2(n10891), .IN3(n10892), .QN(n10886) );
  NAND2X0 U10867 ( .IN1(n9331), .IN2(n10225), .QN(n10892) );
  NAND2X0 U10868 ( .IN1(n10893), .IN2(n10894), .QN(n10225) );
  NAND2X0 U10869 ( .IN1(n7678), .IN2(n10895), .QN(n10894) );
  INVX0 U10870 ( .INP(n10896), .ZN(n10893) );
  NOR2X0 U10871 ( .IN1(n10895), .IN2(n7678), .QN(n10896) );
  NOR2X0 U10872 ( .IN1(n10897), .IN2(n10898), .QN(n10895) );
  NOR2X0 U10873 ( .IN1(WX9894), .IN2(n7679), .QN(n10898) );
  INVX0 U10874 ( .INP(n10899), .ZN(n10897) );
  NAND2X0 U10875 ( .IN1(n7679), .IN2(WX9894), .QN(n10899) );
  NAND2X0 U10876 ( .IN1(n10068), .IN2(n8317), .QN(n10891) );
  NAND2X0 U10877 ( .IN1(n16401), .IN2(n9080), .QN(n10890) );
  NAND2X0 U10878 ( .IN1(n10900), .IN2(n9111), .QN(n10884) );
  NAND2X0 U10879 ( .IN1(n1459), .IN2(n9276), .QN(n10883) );
  NOR2X0 U10880 ( .IN1(n9232), .IN2(n8884), .QN(n1459) );
  NAND2X0 U10881 ( .IN1(n9308), .IN2(CRC_OUT_3_28), .QN(n10882) );
  NAND4X0 U10882 ( .IN1(n10901), .IN2(n10902), .IN3(n10903), .IN4(n10904), 
        .QN(WX8406) );
  NAND2X0 U10883 ( .IN1(n10905), .IN2(n10237), .QN(n10904) );
  NAND2X0 U10884 ( .IN1(n10906), .IN2(n10240), .QN(n10237) );
  NAND2X0 U10885 ( .IN1(n10907), .IN2(n10908), .QN(n10906) );
  NAND2X0 U10886 ( .IN1(n16400), .IN2(n9120), .QN(n10908) );
  NAND2X0 U10887 ( .IN1(TM1), .IN2(n8318), .QN(n10907) );
  NAND3X0 U10888 ( .IN1(n10909), .IN2(n10910), .IN3(n10911), .QN(n10905) );
  NAND2X0 U10889 ( .IN1(n9331), .IN2(n10240), .QN(n10911) );
  NAND2X0 U10890 ( .IN1(n10912), .IN2(n10913), .QN(n10240) );
  NAND2X0 U10891 ( .IN1(n7680), .IN2(n10914), .QN(n10913) );
  INVX0 U10892 ( .INP(n10915), .ZN(n10912) );
  NOR2X0 U10893 ( .IN1(n10914), .IN2(n7680), .QN(n10915) );
  NOR2X0 U10894 ( .IN1(n10916), .IN2(n10917), .QN(n10914) );
  NOR2X0 U10895 ( .IN1(WX9892), .IN2(n7681), .QN(n10917) );
  INVX0 U10896 ( .INP(n10918), .ZN(n10916) );
  NAND2X0 U10897 ( .IN1(n7681), .IN2(WX9892), .QN(n10918) );
  NAND2X0 U10898 ( .IN1(n9084), .IN2(n8318), .QN(n10910) );
  NAND2X0 U10899 ( .IN1(n16400), .IN2(n9079), .QN(n10909) );
  NAND2X0 U10900 ( .IN1(n10919), .IN2(n10920), .QN(n10903) );
  NAND2X0 U10901 ( .IN1(n10921), .IN2(n10922), .QN(n10919) );
  NAND2X0 U10902 ( .IN1(n9097), .IN2(n10923), .QN(n10922) );
  NAND2X0 U10903 ( .IN1(n9097), .IN2(n8376), .QN(n10921) );
  NAND2X0 U10904 ( .IN1(n1458), .IN2(n9276), .QN(n10902) );
  NOR2X0 U10905 ( .IN1(n9232), .IN2(n8885), .QN(n1458) );
  NAND2X0 U10906 ( .IN1(n9308), .IN2(CRC_OUT_3_29), .QN(n10901) );
  NAND4X0 U10907 ( .IN1(n10924), .IN2(n10925), .IN3(n10926), .IN4(n10927), 
        .QN(WX8404) );
  NAND2X0 U10908 ( .IN1(n10928), .IN2(n10252), .QN(n10927) );
  NAND2X0 U10909 ( .IN1(n10929), .IN2(n10255), .QN(n10252) );
  NAND2X0 U10910 ( .IN1(n10930), .IN2(n10931), .QN(n10929) );
  NAND2X0 U10911 ( .IN1(n16399), .IN2(n9120), .QN(n10931) );
  NAND2X0 U10912 ( .IN1(TM1), .IN2(n8319), .QN(n10930) );
  NAND3X0 U10913 ( .IN1(n10932), .IN2(n10933), .IN3(n10934), .QN(n10928) );
  NAND2X0 U10914 ( .IN1(n9331), .IN2(n10255), .QN(n10934) );
  NAND2X0 U10915 ( .IN1(n10935), .IN2(n10936), .QN(n10255) );
  NAND2X0 U10916 ( .IN1(n7682), .IN2(n10937), .QN(n10936) );
  INVX0 U10917 ( .INP(n10938), .ZN(n10935) );
  NOR2X0 U10918 ( .IN1(n10937), .IN2(n7682), .QN(n10938) );
  NOR2X0 U10919 ( .IN1(n10939), .IN2(n10940), .QN(n10937) );
  NOR2X0 U10920 ( .IN1(WX9890), .IN2(n7683), .QN(n10940) );
  INVX0 U10921 ( .INP(n10941), .ZN(n10939) );
  NAND2X0 U10922 ( .IN1(n7683), .IN2(WX9890), .QN(n10941) );
  NAND2X0 U10923 ( .IN1(n9083), .IN2(n8319), .QN(n10933) );
  NAND2X0 U10924 ( .IN1(n16399), .IN2(n9078), .QN(n10932) );
  NAND2X0 U10925 ( .IN1(n10942), .IN2(n9111), .QN(n10926) );
  NAND2X0 U10926 ( .IN1(n1457), .IN2(n9276), .QN(n10925) );
  NOR2X0 U10927 ( .IN1(n9232), .IN2(n8886), .QN(n1457) );
  NAND2X0 U10928 ( .IN1(n9308), .IN2(CRC_OUT_3_30), .QN(n10924) );
  NAND4X0 U10929 ( .IN1(n10943), .IN2(n10944), .IN3(n10945), .IN4(n10946), 
        .QN(WX8402) );
  NAND2X0 U10930 ( .IN1(n10947), .IN2(n10948), .QN(n10946) );
  NAND2X0 U10931 ( .IN1(n10949), .IN2(n10950), .QN(n10947) );
  NAND2X0 U10932 ( .IN1(n9097), .IN2(n10951), .QN(n10950) );
  NAND2X0 U10933 ( .IN1(n9097), .IN2(n8378), .QN(n10949) );
  NAND2X0 U10934 ( .IN1(n10272), .IN2(n9335), .QN(n10945) );
  NOR2X0 U10935 ( .IN1(n10952), .IN2(n10953), .QN(n10272) );
  INVX0 U10936 ( .INP(n10954), .ZN(n10953) );
  NAND2X0 U10937 ( .IN1(n10955), .IN2(n10956), .QN(n10954) );
  NOR2X0 U10938 ( .IN1(n10956), .IN2(n10955), .QN(n10952) );
  NAND2X0 U10939 ( .IN1(n10957), .IN2(n10958), .QN(n10955) );
  NAND2X0 U10940 ( .IN1(n10959), .IN2(WX9824), .QN(n10958) );
  NAND2X0 U10941 ( .IN1(n10960), .IN2(n10961), .QN(n10959) );
  NAND3X0 U10942 ( .IN1(n10960), .IN2(n10961), .IN3(n7615), .QN(n10957) );
  NAND2X0 U10943 ( .IN1(test_so85), .IN2(WX9760), .QN(n10961) );
  NAND2X0 U10944 ( .IN1(n7614), .IN2(n8805), .QN(n10960) );
  NOR2X0 U10945 ( .IN1(n10962), .IN2(n10963), .QN(n10956) );
  INVX0 U10946 ( .INP(n10964), .ZN(n10963) );
  NAND2X0 U10947 ( .IN1(n16398), .IN2(n9120), .QN(n10964) );
  NOR2X0 U10948 ( .IN1(n9117), .IN2(n16398), .QN(n10962) );
  NAND2X0 U10949 ( .IN1(n9308), .IN2(CRC_OUT_3_31), .QN(n10944) );
  NAND2X0 U10950 ( .IN1(n2245), .IN2(WX8243), .QN(n10943) );
  NOR2X0 U10951 ( .IN1(n9231), .IN2(WX8243), .QN(WX8304) );
  NOR3X0 U10952 ( .IN1(n9145), .IN2(n10965), .IN3(n10966), .QN(WX7791) );
  NOR2X0 U10953 ( .IN1(n8212), .IN2(CRC_OUT_4_30), .QN(n10966) );
  NOR2X0 U10954 ( .IN1(DFF_1150_n1), .IN2(WX7302), .QN(n10965) );
  NOR2X0 U10955 ( .IN1(n9231), .IN2(n10967), .QN(WX7789) );
  NOR2X0 U10956 ( .IN1(n10968), .IN2(n10969), .QN(n10967) );
  NOR2X0 U10957 ( .IN1(test_so66), .IN2(WX7304), .QN(n10969) );
  INVX0 U10958 ( .INP(n10970), .ZN(n10968) );
  NAND2X0 U10959 ( .IN1(WX7304), .IN2(test_so66), .QN(n10970) );
  NOR3X0 U10960 ( .IN1(n9145), .IN2(n10971), .IN3(n10972), .QN(WX7787) );
  NOR2X0 U10961 ( .IN1(n8214), .IN2(CRC_OUT_4_28), .QN(n10972) );
  NOR2X0 U10962 ( .IN1(DFF_1148_n1), .IN2(WX7306), .QN(n10971) );
  NOR3X0 U10963 ( .IN1(n9145), .IN2(n10973), .IN3(n10974), .QN(WX7785) );
  NOR2X0 U10964 ( .IN1(n8215), .IN2(CRC_OUT_4_27), .QN(n10974) );
  NOR2X0 U10965 ( .IN1(DFF_1147_n1), .IN2(WX7308), .QN(n10973) );
  NOR3X0 U10966 ( .IN1(n10681), .IN2(n10975), .IN3(n10976), .QN(WX7783) );
  NOR2X0 U10967 ( .IN1(n8216), .IN2(CRC_OUT_4_26), .QN(n10976) );
  NOR2X0 U10968 ( .IN1(DFF_1146_n1), .IN2(WX7310), .QN(n10975) );
  NOR3X0 U10969 ( .IN1(n9145), .IN2(n10977), .IN3(n10978), .QN(WX7781) );
  NOR2X0 U10970 ( .IN1(n8217), .IN2(CRC_OUT_4_25), .QN(n10978) );
  NOR2X0 U10971 ( .IN1(DFF_1145_n1), .IN2(WX7312), .QN(n10977) );
  NOR3X0 U10972 ( .IN1(n9144), .IN2(n10979), .IN3(n10980), .QN(WX7779) );
  NOR2X0 U10973 ( .IN1(n8218), .IN2(CRC_OUT_4_24), .QN(n10980) );
  NOR2X0 U10974 ( .IN1(DFF_1144_n1), .IN2(WX7314), .QN(n10979) );
  NOR3X0 U10975 ( .IN1(n9144), .IN2(n10981), .IN3(n10982), .QN(WX7777) );
  NOR2X0 U10976 ( .IN1(n8219), .IN2(CRC_OUT_4_23), .QN(n10982) );
  NOR2X0 U10977 ( .IN1(DFF_1143_n1), .IN2(WX7316), .QN(n10981) );
  NOR3X0 U10978 ( .IN1(n9144), .IN2(n10983), .IN3(n10984), .QN(WX7775) );
  NOR2X0 U10979 ( .IN1(n8220), .IN2(CRC_OUT_4_22), .QN(n10984) );
  NOR2X0 U10980 ( .IN1(DFF_1142_n1), .IN2(WX7318), .QN(n10983) );
  NOR3X0 U10981 ( .IN1(n9144), .IN2(n10985), .IN3(n10986), .QN(WX7773) );
  NOR2X0 U10982 ( .IN1(n8221), .IN2(CRC_OUT_4_21), .QN(n10986) );
  NOR2X0 U10983 ( .IN1(DFF_1141_n1), .IN2(WX7320), .QN(n10985) );
  NOR2X0 U10984 ( .IN1(n9231), .IN2(n10987), .QN(WX7771) );
  NOR2X0 U10985 ( .IN1(n10988), .IN2(n10989), .QN(n10987) );
  NOR2X0 U10986 ( .IN1(test_so63), .IN2(CRC_OUT_4_20), .QN(n10989) );
  NOR2X0 U10987 ( .IN1(DFF_1140_n1), .IN2(n8800), .QN(n10988) );
  NOR3X0 U10988 ( .IN1(n9144), .IN2(n10990), .IN3(n10991), .QN(WX7769) );
  NOR2X0 U10989 ( .IN1(n8222), .IN2(CRC_OUT_4_19), .QN(n10991) );
  NOR2X0 U10990 ( .IN1(DFF_1139_n1), .IN2(WX7324), .QN(n10990) );
  NOR3X0 U10991 ( .IN1(n9144), .IN2(n10992), .IN3(n10993), .QN(WX7767) );
  NOR2X0 U10992 ( .IN1(n8223), .IN2(CRC_OUT_4_18), .QN(n10993) );
  NOR2X0 U10993 ( .IN1(DFF_1138_n1), .IN2(WX7326), .QN(n10992) );
  NOR3X0 U10994 ( .IN1(n9144), .IN2(n10994), .IN3(n10995), .QN(WX7765) );
  NOR2X0 U10995 ( .IN1(n8224), .IN2(CRC_OUT_4_17), .QN(n10995) );
  NOR2X0 U10996 ( .IN1(DFF_1137_n1), .IN2(WX7328), .QN(n10994) );
  NOR3X0 U10997 ( .IN1(n9144), .IN2(n10996), .IN3(n10997), .QN(WX7763) );
  NOR2X0 U10998 ( .IN1(n8225), .IN2(CRC_OUT_4_16), .QN(n10997) );
  NOR2X0 U10999 ( .IN1(DFF_1136_n1), .IN2(WX7330), .QN(n10996) );
  NOR2X0 U11000 ( .IN1(n9230), .IN2(n10998), .QN(WX7761) );
  NOR2X0 U11001 ( .IN1(n10999), .IN2(n11000), .QN(n10998) );
  INVX0 U11002 ( .INP(n11001), .ZN(n11000) );
  NAND2X0 U11003 ( .IN1(CRC_OUT_4_15), .IN2(n11002), .QN(n11001) );
  NOR2X0 U11004 ( .IN1(n11002), .IN2(CRC_OUT_4_15), .QN(n10999) );
  NAND2X0 U11005 ( .IN1(n11003), .IN2(n11004), .QN(n11002) );
  NAND2X0 U11006 ( .IN1(n8114), .IN2(CRC_OUT_4_31), .QN(n11004) );
  NAND2X0 U11007 ( .IN1(DFF_1151_n1), .IN2(WX7332), .QN(n11003) );
  NOR3X0 U11008 ( .IN1(n9144), .IN2(n11005), .IN3(n11006), .QN(WX7759) );
  NOR2X0 U11009 ( .IN1(n8226), .IN2(CRC_OUT_4_14), .QN(n11006) );
  NOR2X0 U11010 ( .IN1(DFF_1134_n1), .IN2(WX7334), .QN(n11005) );
  NOR3X0 U11011 ( .IN1(n9144), .IN2(n11007), .IN3(n11008), .QN(WX7757) );
  NOR2X0 U11012 ( .IN1(n8227), .IN2(CRC_OUT_4_13), .QN(n11008) );
  NOR2X0 U11013 ( .IN1(DFF_1133_n1), .IN2(WX7336), .QN(n11007) );
  NOR2X0 U11014 ( .IN1(n9230), .IN2(n11009), .QN(WX7755) );
  NOR2X0 U11015 ( .IN1(n11010), .IN2(n11011), .QN(n11009) );
  NOR2X0 U11016 ( .IN1(test_so65), .IN2(WX7338), .QN(n11011) );
  INVX0 U11017 ( .INP(n11012), .ZN(n11010) );
  NAND2X0 U11018 ( .IN1(WX7338), .IN2(test_so65), .QN(n11012) );
  NOR3X0 U11019 ( .IN1(n9144), .IN2(n11013), .IN3(n11014), .QN(WX7753) );
  NOR2X0 U11020 ( .IN1(n8229), .IN2(CRC_OUT_4_11), .QN(n11014) );
  NOR2X0 U11021 ( .IN1(DFF_1131_n1), .IN2(WX7340), .QN(n11013) );
  NOR2X0 U11022 ( .IN1(n9230), .IN2(n11015), .QN(WX7751) );
  NOR2X0 U11023 ( .IN1(n11016), .IN2(n11017), .QN(n11015) );
  INVX0 U11024 ( .INP(n11018), .ZN(n11017) );
  NAND2X0 U11025 ( .IN1(CRC_OUT_4_10), .IN2(n11019), .QN(n11018) );
  NOR2X0 U11026 ( .IN1(n11019), .IN2(CRC_OUT_4_10), .QN(n11016) );
  NAND2X0 U11027 ( .IN1(n11020), .IN2(n11021), .QN(n11019) );
  NAND2X0 U11028 ( .IN1(n8115), .IN2(CRC_OUT_4_31), .QN(n11021) );
  NAND2X0 U11029 ( .IN1(DFF_1151_n1), .IN2(WX7342), .QN(n11020) );
  NOR3X0 U11030 ( .IN1(n9144), .IN2(n11022), .IN3(n11023), .QN(WX7749) );
  NOR2X0 U11031 ( .IN1(n8230), .IN2(CRC_OUT_4_9), .QN(n11023) );
  NOR2X0 U11032 ( .IN1(DFF_1129_n1), .IN2(WX7344), .QN(n11022) );
  NOR3X0 U11033 ( .IN1(n9143), .IN2(n11024), .IN3(n11025), .QN(WX7747) );
  NOR2X0 U11034 ( .IN1(n8231), .IN2(CRC_OUT_4_8), .QN(n11025) );
  NOR2X0 U11035 ( .IN1(DFF_1128_n1), .IN2(WX7346), .QN(n11024) );
  NOR3X0 U11036 ( .IN1(n9143), .IN2(n11026), .IN3(n11027), .QN(WX7745) );
  NOR2X0 U11037 ( .IN1(n8232), .IN2(CRC_OUT_4_7), .QN(n11027) );
  NOR2X0 U11038 ( .IN1(DFF_1127_n1), .IN2(WX7348), .QN(n11026) );
  NOR3X0 U11039 ( .IN1(n9143), .IN2(n11028), .IN3(n11029), .QN(WX7743) );
  NOR2X0 U11040 ( .IN1(n8233), .IN2(CRC_OUT_4_6), .QN(n11029) );
  NOR2X0 U11041 ( .IN1(DFF_1126_n1), .IN2(WX7350), .QN(n11028) );
  NOR3X0 U11042 ( .IN1(n9143), .IN2(n11030), .IN3(n11031), .QN(WX7741) );
  NOR2X0 U11043 ( .IN1(n8234), .IN2(CRC_OUT_4_5), .QN(n11031) );
  NOR2X0 U11044 ( .IN1(DFF_1125_n1), .IN2(WX7352), .QN(n11030) );
  NOR3X0 U11045 ( .IN1(n9143), .IN2(n11032), .IN3(n11033), .QN(WX7739) );
  NOR2X0 U11046 ( .IN1(n8235), .IN2(CRC_OUT_4_4), .QN(n11033) );
  NOR2X0 U11047 ( .IN1(DFF_1124_n1), .IN2(WX7354), .QN(n11032) );
  NOR3X0 U11048 ( .IN1(n9143), .IN2(n11034), .IN3(n11035), .QN(WX7737) );
  INVX0 U11049 ( .INP(n11036), .ZN(n11035) );
  NAND2X0 U11050 ( .IN1(CRC_OUT_4_3), .IN2(n11037), .QN(n11036) );
  NOR2X0 U11051 ( .IN1(n11037), .IN2(CRC_OUT_4_3), .QN(n11034) );
  NAND2X0 U11052 ( .IN1(n11038), .IN2(n11039), .QN(n11037) );
  NAND2X0 U11053 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .QN(n11039) );
  NAND2X0 U11054 ( .IN1(DFF_1151_n1), .IN2(n8796), .QN(n11038) );
  NOR3X0 U11055 ( .IN1(n9143), .IN2(n11040), .IN3(n11041), .QN(WX7735) );
  NOR2X0 U11056 ( .IN1(n8236), .IN2(CRC_OUT_4_2), .QN(n11041) );
  NOR2X0 U11057 ( .IN1(DFF_1122_n1), .IN2(WX7358), .QN(n11040) );
  NOR3X0 U11058 ( .IN1(n9143), .IN2(n11042), .IN3(n11043), .QN(WX7733) );
  NOR2X0 U11059 ( .IN1(n8237), .IN2(CRC_OUT_4_1), .QN(n11043) );
  NOR2X0 U11060 ( .IN1(DFF_1121_n1), .IN2(WX7360), .QN(n11042) );
  NOR3X0 U11061 ( .IN1(n9143), .IN2(n11044), .IN3(n11045), .QN(WX7731) );
  NOR2X0 U11062 ( .IN1(n8238), .IN2(CRC_OUT_4_0), .QN(n11045) );
  NOR2X0 U11063 ( .IN1(DFF_1120_n1), .IN2(WX7362), .QN(n11044) );
  NOR3X0 U11064 ( .IN1(n9143), .IN2(n11046), .IN3(n11047), .QN(WX7729) );
  NOR2X0 U11065 ( .IN1(n8129), .IN2(CRC_OUT_4_31), .QN(n11047) );
  NOR2X0 U11066 ( .IN1(DFF_1151_n1), .IN2(WX7364), .QN(n11046) );
  NOR2X0 U11067 ( .IN1(n16381), .IN2(n9164), .QN(WX7203) );
  NOR2X0 U11068 ( .IN1(n16380), .IN2(n9165), .QN(WX7201) );
  NOR2X0 U11069 ( .IN1(n16379), .IN2(n9164), .QN(WX7199) );
  NOR2X0 U11070 ( .IN1(n16378), .IN2(n9164), .QN(WX7197) );
  NOR2X0 U11071 ( .IN1(n16377), .IN2(n9164), .QN(WX7195) );
  NOR2X0 U11072 ( .IN1(n16376), .IN2(n9164), .QN(WX7193) );
  NOR2X0 U11073 ( .IN1(n16375), .IN2(n9164), .QN(WX7191) );
  NOR2X0 U11074 ( .IN1(n16374), .IN2(n9164), .QN(WX7189) );
  NOR2X0 U11075 ( .IN1(n16373), .IN2(n9164), .QN(WX7187) );
  NOR2X0 U11076 ( .IN1(n16372), .IN2(n9164), .QN(WX7185) );
  NOR2X0 U11077 ( .IN1(n16371), .IN2(n9164), .QN(WX7183) );
  NOR2X0 U11078 ( .IN1(n9227), .IN2(n8821), .QN(WX7181) );
  NOR2X0 U11079 ( .IN1(n16370), .IN2(n9164), .QN(WX7179) );
  NOR2X0 U11080 ( .IN1(n16369), .IN2(n9164), .QN(WX7177) );
  NOR2X0 U11081 ( .IN1(n16368), .IN2(n9164), .QN(WX7175) );
  NOR2X0 U11082 ( .IN1(n16367), .IN2(n9163), .QN(WX7173) );
  NAND4X0 U11083 ( .IN1(n11048), .IN2(n11049), .IN3(n11050), .IN4(n11051), 
        .QN(WX7171) );
  NAND2X0 U11084 ( .IN1(n9331), .IN2(n10373), .QN(n11051) );
  NAND2X0 U11085 ( .IN1(n11052), .IN2(n11053), .QN(n10373) );
  INVX0 U11086 ( .INP(n11054), .ZN(n11053) );
  NOR2X0 U11087 ( .IN1(n11055), .IN2(n11056), .QN(n11054) );
  NAND2X0 U11088 ( .IN1(n11056), .IN2(n11055), .QN(n11052) );
  NOR2X0 U11089 ( .IN1(n11057), .IN2(n11058), .QN(n11055) );
  NOR2X0 U11090 ( .IN1(WX8657), .IN2(n7916), .QN(n11058) );
  INVX0 U11091 ( .INP(n11059), .ZN(n11057) );
  NAND2X0 U11092 ( .IN1(n7916), .IN2(WX8657), .QN(n11059) );
  NAND2X0 U11093 ( .IN1(n11060), .IN2(n11061), .QN(n11056) );
  NAND2X0 U11094 ( .IN1(n7915), .IN2(WX8529), .QN(n11061) );
  INVX0 U11095 ( .INP(n11062), .ZN(n11060) );
  NOR2X0 U11096 ( .IN1(WX8529), .IN2(n7915), .QN(n11062) );
  NAND2X0 U11097 ( .IN1(n9097), .IN2(n11063), .QN(n11050) );
  NAND2X0 U11098 ( .IN1(n1246), .IN2(n9276), .QN(n11049) );
  NOR2X0 U11099 ( .IN1(n9227), .IN2(n8887), .QN(n1246) );
  NAND2X0 U11100 ( .IN1(n9308), .IN2(CRC_OUT_4_0), .QN(n11048) );
  NAND4X0 U11101 ( .IN1(n11064), .IN2(n11065), .IN3(n11066), .IN4(n11067), 
        .QN(WX7169) );
  NAND2X0 U11102 ( .IN1(n9331), .IN2(n10386), .QN(n11067) );
  NAND2X0 U11103 ( .IN1(n11068), .IN2(n11069), .QN(n10386) );
  INVX0 U11104 ( .INP(n11070), .ZN(n11069) );
  NOR2X0 U11105 ( .IN1(n11071), .IN2(n11072), .QN(n11070) );
  NAND2X0 U11106 ( .IN1(n11072), .IN2(n11071), .QN(n11068) );
  NOR2X0 U11107 ( .IN1(n11073), .IN2(n11074), .QN(n11071) );
  NOR2X0 U11108 ( .IN1(WX8655), .IN2(n7918), .QN(n11074) );
  INVX0 U11109 ( .INP(n11075), .ZN(n11073) );
  NAND2X0 U11110 ( .IN1(n7918), .IN2(WX8655), .QN(n11075) );
  NAND2X0 U11111 ( .IN1(n11076), .IN2(n11077), .QN(n11072) );
  NAND2X0 U11112 ( .IN1(n7917), .IN2(WX8527), .QN(n11077) );
  INVX0 U11113 ( .INP(n11078), .ZN(n11076) );
  NOR2X0 U11114 ( .IN1(WX8527), .IN2(n7917), .QN(n11078) );
  NAND2X0 U11115 ( .IN1(n9097), .IN2(n11079), .QN(n11066) );
  NAND2X0 U11116 ( .IN1(n1245), .IN2(n9276), .QN(n11065) );
  NOR2X0 U11117 ( .IN1(n9227), .IN2(n8888), .QN(n1245) );
  NAND2X0 U11118 ( .IN1(n9308), .IN2(CRC_OUT_4_1), .QN(n11064) );
  NAND4X0 U11119 ( .IN1(n11080), .IN2(n11081), .IN3(n11082), .IN4(n11083), 
        .QN(WX7167) );
  NAND2X0 U11120 ( .IN1(n9331), .IN2(n10402), .QN(n11083) );
  NAND2X0 U11121 ( .IN1(n11084), .IN2(n11085), .QN(n10402) );
  INVX0 U11122 ( .INP(n11086), .ZN(n11085) );
  NOR2X0 U11123 ( .IN1(n11087), .IN2(n11088), .QN(n11086) );
  NAND2X0 U11124 ( .IN1(n11088), .IN2(n11087), .QN(n11084) );
  NOR2X0 U11125 ( .IN1(n11089), .IN2(n11090), .QN(n11087) );
  NOR2X0 U11126 ( .IN1(WX8653), .IN2(n7920), .QN(n11090) );
  INVX0 U11127 ( .INP(n11091), .ZN(n11089) );
  NAND2X0 U11128 ( .IN1(n7920), .IN2(WX8653), .QN(n11091) );
  NAND2X0 U11129 ( .IN1(n11092), .IN2(n11093), .QN(n11088) );
  NAND2X0 U11130 ( .IN1(n7919), .IN2(WX8525), .QN(n11093) );
  INVX0 U11131 ( .INP(n11094), .ZN(n11092) );
  NOR2X0 U11132 ( .IN1(WX8525), .IN2(n7919), .QN(n11094) );
  NAND2X0 U11133 ( .IN1(n9097), .IN2(n11095), .QN(n11082) );
  NAND2X0 U11134 ( .IN1(n1244), .IN2(n9276), .QN(n11081) );
  NOR2X0 U11135 ( .IN1(n9227), .IN2(n8889), .QN(n1244) );
  NAND2X0 U11136 ( .IN1(n9308), .IN2(CRC_OUT_4_2), .QN(n11080) );
  NAND4X0 U11137 ( .IN1(n11096), .IN2(n11097), .IN3(n11098), .IN4(n11099), 
        .QN(WX7165) );
  NAND2X0 U11138 ( .IN1(n9331), .IN2(n10415), .QN(n11099) );
  NAND2X0 U11139 ( .IN1(n11100), .IN2(n11101), .QN(n10415) );
  INVX0 U11140 ( .INP(n11102), .ZN(n11101) );
  NOR2X0 U11141 ( .IN1(n11103), .IN2(n11104), .QN(n11102) );
  NAND2X0 U11142 ( .IN1(n11104), .IN2(n11103), .QN(n11100) );
  NOR2X0 U11143 ( .IN1(n11105), .IN2(n11106), .QN(n11103) );
  NOR2X0 U11144 ( .IN1(WX8651), .IN2(n7922), .QN(n11106) );
  INVX0 U11145 ( .INP(n11107), .ZN(n11105) );
  NAND2X0 U11146 ( .IN1(n7922), .IN2(WX8651), .QN(n11107) );
  NAND2X0 U11147 ( .IN1(n11108), .IN2(n11109), .QN(n11104) );
  NAND2X0 U11148 ( .IN1(n7921), .IN2(WX8523), .QN(n11109) );
  INVX0 U11149 ( .INP(n11110), .ZN(n11108) );
  NOR2X0 U11150 ( .IN1(WX8523), .IN2(n7921), .QN(n11110) );
  NAND2X0 U11151 ( .IN1(n9097), .IN2(n11111), .QN(n11098) );
  NAND2X0 U11152 ( .IN1(n1243), .IN2(n9276), .QN(n11097) );
  NOR2X0 U11153 ( .IN1(n9225), .IN2(n8890), .QN(n1243) );
  NAND2X0 U11154 ( .IN1(n9308), .IN2(CRC_OUT_4_3), .QN(n11096) );
  NAND4X0 U11155 ( .IN1(n11112), .IN2(n11113), .IN3(n11114), .IN4(n11115), 
        .QN(WX7163) );
  NAND3X0 U11156 ( .IN1(n11116), .IN2(n11117), .IN3(n9090), .QN(n11115) );
  NAND2X0 U11157 ( .IN1(n9332), .IN2(n10431), .QN(n11114) );
  NAND2X0 U11158 ( .IN1(n11118), .IN2(n11119), .QN(n10431) );
  INVX0 U11159 ( .INP(n11120), .ZN(n11119) );
  NOR2X0 U11160 ( .IN1(n11121), .IN2(n11122), .QN(n11120) );
  NAND2X0 U11161 ( .IN1(n11122), .IN2(n11121), .QN(n11118) );
  NOR2X0 U11162 ( .IN1(n11123), .IN2(n11124), .QN(n11121) );
  NOR2X0 U11163 ( .IN1(WX8649), .IN2(n7924), .QN(n11124) );
  INVX0 U11164 ( .INP(n11125), .ZN(n11123) );
  NAND2X0 U11165 ( .IN1(n7924), .IN2(WX8649), .QN(n11125) );
  NAND2X0 U11166 ( .IN1(n11126), .IN2(n11127), .QN(n11122) );
  NAND2X0 U11167 ( .IN1(n7923), .IN2(WX8521), .QN(n11127) );
  INVX0 U11168 ( .INP(n11128), .ZN(n11126) );
  NOR2X0 U11169 ( .IN1(WX8521), .IN2(n7923), .QN(n11128) );
  NAND2X0 U11170 ( .IN1(n1242), .IN2(n9276), .QN(n11113) );
  NOR2X0 U11171 ( .IN1(n9224), .IN2(n8891), .QN(n1242) );
  NAND2X0 U11172 ( .IN1(n9308), .IN2(CRC_OUT_4_4), .QN(n11112) );
  NAND4X0 U11173 ( .IN1(n11129), .IN2(n11130), .IN3(n11131), .IN4(n11132), 
        .QN(WX7161) );
  NAND2X0 U11174 ( .IN1(n9332), .IN2(n10447), .QN(n11132) );
  NAND2X0 U11175 ( .IN1(n11133), .IN2(n11134), .QN(n10447) );
  INVX0 U11176 ( .INP(n11135), .ZN(n11134) );
  NOR2X0 U11177 ( .IN1(n11136), .IN2(n11137), .QN(n11135) );
  NAND2X0 U11178 ( .IN1(n11137), .IN2(n11136), .QN(n11133) );
  NOR2X0 U11179 ( .IN1(n11138), .IN2(n11139), .QN(n11136) );
  NOR2X0 U11180 ( .IN1(WX8647), .IN2(n7926), .QN(n11139) );
  INVX0 U11181 ( .INP(n11140), .ZN(n11138) );
  NAND2X0 U11182 ( .IN1(n7926), .IN2(WX8647), .QN(n11140) );
  NAND2X0 U11183 ( .IN1(n11141), .IN2(n11142), .QN(n11137) );
  NAND2X0 U11184 ( .IN1(n7925), .IN2(WX8519), .QN(n11142) );
  INVX0 U11185 ( .INP(n11143), .ZN(n11141) );
  NOR2X0 U11186 ( .IN1(WX8519), .IN2(n7925), .QN(n11143) );
  NAND2X0 U11187 ( .IN1(n9097), .IN2(n11144), .QN(n11131) );
  NAND2X0 U11188 ( .IN1(n508), .IN2(n9277), .QN(n11130) );
  NOR2X0 U11189 ( .IN1(n10681), .IN2(n8892), .QN(n508) );
  NAND2X0 U11190 ( .IN1(n9308), .IN2(CRC_OUT_4_5), .QN(n11129) );
  NAND4X0 U11191 ( .IN1(n11145), .IN2(n11146), .IN3(n11147), .IN4(n11148), 
        .QN(WX7159) );
  NAND3X0 U11192 ( .IN1(n11149), .IN2(n11150), .IN3(n9090), .QN(n11148) );
  NAND2X0 U11193 ( .IN1(n9332), .IN2(n10463), .QN(n11147) );
  NAND2X0 U11194 ( .IN1(n11151), .IN2(n11152), .QN(n10463) );
  INVX0 U11195 ( .INP(n11153), .ZN(n11152) );
  NOR2X0 U11196 ( .IN1(n11154), .IN2(n11155), .QN(n11153) );
  NAND2X0 U11197 ( .IN1(n11155), .IN2(n11154), .QN(n11151) );
  NOR2X0 U11198 ( .IN1(n11156), .IN2(n11157), .QN(n11154) );
  NOR2X0 U11199 ( .IN1(WX8645), .IN2(n7928), .QN(n11157) );
  INVX0 U11200 ( .INP(n11158), .ZN(n11156) );
  NAND2X0 U11201 ( .IN1(n7928), .IN2(WX8645), .QN(n11158) );
  NAND2X0 U11202 ( .IN1(n11159), .IN2(n11160), .QN(n11155) );
  NAND2X0 U11203 ( .IN1(n7927), .IN2(WX8517), .QN(n11160) );
  INVX0 U11204 ( .INP(n11161), .ZN(n11159) );
  NOR2X0 U11205 ( .IN1(WX8517), .IN2(n7927), .QN(n11161) );
  NAND2X0 U11206 ( .IN1(n1241), .IN2(n9277), .QN(n11146) );
  NOR2X0 U11207 ( .IN1(n9224), .IN2(n8893), .QN(n1241) );
  NAND2X0 U11208 ( .IN1(n9309), .IN2(CRC_OUT_4_6), .QN(n11145) );
  NAND4X0 U11209 ( .IN1(n11162), .IN2(n11163), .IN3(n11164), .IN4(n11165), 
        .QN(WX7157) );
  NAND2X0 U11210 ( .IN1(n9332), .IN2(n10479), .QN(n11165) );
  NAND2X0 U11211 ( .IN1(n11166), .IN2(n11167), .QN(n10479) );
  INVX0 U11212 ( .INP(n11168), .ZN(n11167) );
  NOR2X0 U11213 ( .IN1(n11169), .IN2(n11170), .QN(n11168) );
  NAND2X0 U11214 ( .IN1(n11170), .IN2(n11169), .QN(n11166) );
  NOR2X0 U11215 ( .IN1(n11171), .IN2(n11172), .QN(n11169) );
  NOR2X0 U11216 ( .IN1(WX8643), .IN2(n7930), .QN(n11172) );
  INVX0 U11217 ( .INP(n11173), .ZN(n11171) );
  NAND2X0 U11218 ( .IN1(n7930), .IN2(WX8643), .QN(n11173) );
  NAND2X0 U11219 ( .IN1(n11174), .IN2(n11175), .QN(n11170) );
  NAND2X0 U11220 ( .IN1(n7929), .IN2(WX8515), .QN(n11175) );
  INVX0 U11221 ( .INP(n11176), .ZN(n11174) );
  NOR2X0 U11222 ( .IN1(WX8515), .IN2(n7929), .QN(n11176) );
  NAND2X0 U11223 ( .IN1(n9097), .IN2(n11177), .QN(n11164) );
  NAND2X0 U11224 ( .IN1(n1240), .IN2(n9277), .QN(n11163) );
  NOR2X0 U11225 ( .IN1(n9224), .IN2(n8894), .QN(n1240) );
  NAND2X0 U11226 ( .IN1(n9309), .IN2(CRC_OUT_4_7), .QN(n11162) );
  NAND4X0 U11227 ( .IN1(n11178), .IN2(n11179), .IN3(n11180), .IN4(n11181), 
        .QN(WX7155) );
  NAND3X0 U11228 ( .IN1(n11182), .IN2(n11183), .IN3(n9090), .QN(n11181) );
  NAND2X0 U11229 ( .IN1(n9332), .IN2(n10495), .QN(n11180) );
  NAND2X0 U11230 ( .IN1(n11184), .IN2(n11185), .QN(n10495) );
  INVX0 U11231 ( .INP(n11186), .ZN(n11185) );
  NOR2X0 U11232 ( .IN1(n11187), .IN2(n11188), .QN(n11186) );
  NAND2X0 U11233 ( .IN1(n11188), .IN2(n11187), .QN(n11184) );
  NOR2X0 U11234 ( .IN1(n11189), .IN2(n11190), .QN(n11187) );
  NOR2X0 U11235 ( .IN1(WX8641), .IN2(n7932), .QN(n11190) );
  INVX0 U11236 ( .INP(n11191), .ZN(n11189) );
  NAND2X0 U11237 ( .IN1(n7932), .IN2(WX8641), .QN(n11191) );
  NAND2X0 U11238 ( .IN1(n11192), .IN2(n11193), .QN(n11188) );
  NAND2X0 U11239 ( .IN1(n7931), .IN2(WX8513), .QN(n11193) );
  INVX0 U11240 ( .INP(n11194), .ZN(n11192) );
  NOR2X0 U11241 ( .IN1(WX8513), .IN2(n7931), .QN(n11194) );
  NAND2X0 U11242 ( .IN1(n1239), .IN2(n9277), .QN(n11179) );
  NOR2X0 U11243 ( .IN1(n9224), .IN2(n8895), .QN(n1239) );
  NAND2X0 U11244 ( .IN1(n9309), .IN2(CRC_OUT_4_8), .QN(n11178) );
  NAND4X0 U11245 ( .IN1(n11195), .IN2(n11196), .IN3(n11197), .IN4(n11198), 
        .QN(WX7153) );
  NAND3X0 U11246 ( .IN1(n10500), .IN2(n10501), .IN3(n9323), .QN(n11198) );
  NAND3X0 U11247 ( .IN1(n11199), .IN2(n11200), .IN3(n11201), .QN(n10501) );
  INVX0 U11248 ( .INP(n11202), .ZN(n11201) );
  NAND2X0 U11249 ( .IN1(n11202), .IN2(n11203), .QN(n10500) );
  NAND2X0 U11250 ( .IN1(n11199), .IN2(n11200), .QN(n11203) );
  NAND2X0 U11251 ( .IN1(n7934), .IN2(WX8511), .QN(n11200) );
  NAND2X0 U11252 ( .IN1(n3613), .IN2(WX8575), .QN(n11199) );
  NOR2X0 U11253 ( .IN1(n11204), .IN2(n11205), .QN(n11202) );
  NOR2X0 U11254 ( .IN1(n8791), .IN2(n7933), .QN(n11205) );
  INVX0 U11255 ( .INP(n11206), .ZN(n11204) );
  NAND2X0 U11256 ( .IN1(n7933), .IN2(n8791), .QN(n11206) );
  NAND2X0 U11257 ( .IN1(n9096), .IN2(n11207), .QN(n11197) );
  NAND2X0 U11258 ( .IN1(n1238), .IN2(n9277), .QN(n11196) );
  NOR2X0 U11259 ( .IN1(n9224), .IN2(n8896), .QN(n1238) );
  NAND2X0 U11260 ( .IN1(n9309), .IN2(CRC_OUT_4_9), .QN(n11195) );
  NAND4X0 U11261 ( .IN1(n11208), .IN2(n11209), .IN3(n11210), .IN4(n11211), 
        .QN(WX7151) );
  NAND3X0 U11262 ( .IN1(n11212), .IN2(n11213), .IN3(n9090), .QN(n11211) );
  NAND2X0 U11263 ( .IN1(n9332), .IN2(n10528), .QN(n11210) );
  NAND2X0 U11264 ( .IN1(n11214), .IN2(n11215), .QN(n10528) );
  INVX0 U11265 ( .INP(n11216), .ZN(n11215) );
  NOR2X0 U11266 ( .IN1(n11217), .IN2(n11218), .QN(n11216) );
  NAND2X0 U11267 ( .IN1(n11218), .IN2(n11217), .QN(n11214) );
  NOR2X0 U11268 ( .IN1(n11219), .IN2(n11220), .QN(n11217) );
  NOR2X0 U11269 ( .IN1(WX8637), .IN2(n7936), .QN(n11220) );
  INVX0 U11270 ( .INP(n11221), .ZN(n11219) );
  NAND2X0 U11271 ( .IN1(n7936), .IN2(WX8637), .QN(n11221) );
  NAND2X0 U11272 ( .IN1(n11222), .IN2(n11223), .QN(n11218) );
  NAND2X0 U11273 ( .IN1(n7935), .IN2(WX8509), .QN(n11223) );
  INVX0 U11274 ( .INP(n11224), .ZN(n11222) );
  NOR2X0 U11275 ( .IN1(WX8509), .IN2(n7935), .QN(n11224) );
  NAND2X0 U11276 ( .IN1(n1237), .IN2(n9277), .QN(n11209) );
  NOR2X0 U11277 ( .IN1(n9224), .IN2(n8897), .QN(n1237) );
  NAND2X0 U11278 ( .IN1(n9309), .IN2(CRC_OUT_4_10), .QN(n11208) );
  NAND4X0 U11279 ( .IN1(n11225), .IN2(n11226), .IN3(n11227), .IN4(n11228), 
        .QN(WX7149) );
  NAND3X0 U11280 ( .IN1(n10533), .IN2(n10534), .IN3(n9323), .QN(n11228) );
  NAND3X0 U11281 ( .IN1(n11229), .IN2(n11230), .IN3(n11231), .QN(n10534) );
  INVX0 U11282 ( .INP(n11232), .ZN(n11231) );
  NAND2X0 U11283 ( .IN1(n11232), .IN2(n11233), .QN(n10533) );
  NAND2X0 U11284 ( .IN1(n11229), .IN2(n11230), .QN(n11233) );
  NAND2X0 U11285 ( .IN1(n8112), .IN2(WX8507), .QN(n11230) );
  NAND2X0 U11286 ( .IN1(n3617), .IN2(WX8635), .QN(n11229) );
  NOR2X0 U11287 ( .IN1(n11234), .IN2(n11235), .QN(n11232) );
  INVX0 U11288 ( .INP(n11236), .ZN(n11235) );
  NAND2X0 U11289 ( .IN1(test_so73), .IN2(WX8443), .QN(n11236) );
  NOR2X0 U11290 ( .IN1(WX8443), .IN2(test_so73), .QN(n11234) );
  NAND2X0 U11291 ( .IN1(n9096), .IN2(n11237), .QN(n11227) );
  NAND2X0 U11292 ( .IN1(n1236), .IN2(n9277), .QN(n11226) );
  NOR2X0 U11293 ( .IN1(n9224), .IN2(n8898), .QN(n1236) );
  NAND2X0 U11294 ( .IN1(n9309), .IN2(CRC_OUT_4_11), .QN(n11225) );
  NAND4X0 U11295 ( .IN1(n11238), .IN2(n11239), .IN3(n11240), .IN4(n11241), 
        .QN(WX7147) );
  NAND2X0 U11296 ( .IN1(n9332), .IN2(n10561), .QN(n11241) );
  NAND2X0 U11297 ( .IN1(n11242), .IN2(n11243), .QN(n10561) );
  INVX0 U11298 ( .INP(n11244), .ZN(n11243) );
  NOR2X0 U11299 ( .IN1(n11245), .IN2(n11246), .QN(n11244) );
  NAND2X0 U11300 ( .IN1(n11246), .IN2(n11245), .QN(n11242) );
  NOR2X0 U11301 ( .IN1(n11247), .IN2(n11248), .QN(n11245) );
  NOR2X0 U11302 ( .IN1(WX8633), .IN2(n7939), .QN(n11248) );
  INVX0 U11303 ( .INP(n11249), .ZN(n11247) );
  NAND2X0 U11304 ( .IN1(n7939), .IN2(WX8633), .QN(n11249) );
  NAND2X0 U11305 ( .IN1(n11250), .IN2(n11251), .QN(n11246) );
  NAND2X0 U11306 ( .IN1(n7938), .IN2(WX8505), .QN(n11251) );
  INVX0 U11307 ( .INP(n11252), .ZN(n11250) );
  NOR2X0 U11308 ( .IN1(WX8505), .IN2(n7938), .QN(n11252) );
  NAND2X0 U11309 ( .IN1(n9096), .IN2(n11253), .QN(n11240) );
  NAND2X0 U11310 ( .IN1(n1235), .IN2(n9277), .QN(n11239) );
  NOR2X0 U11311 ( .IN1(n9065), .IN2(n9164), .QN(n1235) );
  NAND2X0 U11312 ( .IN1(test_so65), .IN2(n9314), .QN(n11238) );
  NAND4X0 U11313 ( .IN1(n11254), .IN2(n11255), .IN3(n11256), .IN4(n11257), 
        .QN(WX7145) );
  NAND3X0 U11314 ( .IN1(n10566), .IN2(n10567), .IN3(n9323), .QN(n11257) );
  NAND3X0 U11315 ( .IN1(n11258), .IN2(n11259), .IN3(n11260), .QN(n10567) );
  INVX0 U11316 ( .INP(n11261), .ZN(n11260) );
  NAND2X0 U11317 ( .IN1(n11261), .IN2(n11262), .QN(n10566) );
  NAND2X0 U11318 ( .IN1(n11258), .IN2(n11259), .QN(n11262) );
  NAND2X0 U11319 ( .IN1(n8202), .IN2(WX8567), .QN(n11259) );
  NAND2X0 U11320 ( .IN1(n7941), .IN2(WX8631), .QN(n11258) );
  NOR2X0 U11321 ( .IN1(n11263), .IN2(n11264), .QN(n11261) );
  INVX0 U11322 ( .INP(n11265), .ZN(n11264) );
  NAND2X0 U11323 ( .IN1(test_so71), .IN2(WX8439), .QN(n11265) );
  NOR2X0 U11324 ( .IN1(WX8439), .IN2(test_so71), .QN(n11263) );
  NAND2X0 U11325 ( .IN1(n9096), .IN2(n11266), .QN(n11256) );
  NAND2X0 U11326 ( .IN1(n1234), .IN2(n9277), .QN(n11255) );
  NOR2X0 U11327 ( .IN1(n9224), .IN2(n8899), .QN(n1234) );
  NAND2X0 U11328 ( .IN1(n9309), .IN2(CRC_OUT_4_13), .QN(n11254) );
  NAND4X0 U11329 ( .IN1(n11267), .IN2(n11268), .IN3(n11269), .IN4(n11270), 
        .QN(WX7143) );
  NAND2X0 U11330 ( .IN1(n9332), .IN2(n10591), .QN(n11270) );
  NAND2X0 U11331 ( .IN1(n11271), .IN2(n11272), .QN(n10591) );
  INVX0 U11332 ( .INP(n11273), .ZN(n11272) );
  NOR2X0 U11333 ( .IN1(n11274), .IN2(n11275), .QN(n11273) );
  NAND2X0 U11334 ( .IN1(n11275), .IN2(n11274), .QN(n11271) );
  NOR2X0 U11335 ( .IN1(n11276), .IN2(n11277), .QN(n11274) );
  NOR2X0 U11336 ( .IN1(WX8629), .IN2(n7943), .QN(n11277) );
  INVX0 U11337 ( .INP(n11278), .ZN(n11276) );
  NAND2X0 U11338 ( .IN1(n7943), .IN2(WX8629), .QN(n11278) );
  NAND2X0 U11339 ( .IN1(n11279), .IN2(n11280), .QN(n11275) );
  NAND2X0 U11340 ( .IN1(n7942), .IN2(WX8501), .QN(n11280) );
  INVX0 U11341 ( .INP(n11281), .ZN(n11279) );
  NOR2X0 U11342 ( .IN1(WX8501), .IN2(n7942), .QN(n11281) );
  NAND2X0 U11343 ( .IN1(n9096), .IN2(n11282), .QN(n11269) );
  NAND2X0 U11344 ( .IN1(n1233), .IN2(n9277), .QN(n11268) );
  NOR2X0 U11345 ( .IN1(n9224), .IN2(n8900), .QN(n1233) );
  NAND2X0 U11346 ( .IN1(n9309), .IN2(CRC_OUT_4_14), .QN(n11267) );
  NAND4X0 U11347 ( .IN1(n11283), .IN2(n11284), .IN3(n11285), .IN4(n11286), 
        .QN(WX7141) );
  NAND3X0 U11348 ( .IN1(n10596), .IN2(n10597), .IN3(n9322), .QN(n11286) );
  NAND3X0 U11349 ( .IN1(n11287), .IN2(n11288), .IN3(n11289), .QN(n10597) );
  INVX0 U11350 ( .INP(n11290), .ZN(n11289) );
  NAND2X0 U11351 ( .IN1(n11290), .IN2(n11291), .QN(n10596) );
  NAND2X0 U11352 ( .IN1(n11287), .IN2(n11288), .QN(n11291) );
  NAND2X0 U11353 ( .IN1(n8200), .IN2(WX8499), .QN(n11288) );
  NAND2X0 U11354 ( .IN1(n3625), .IN2(WX8627), .QN(n11287) );
  NOR2X0 U11355 ( .IN1(n11292), .IN2(n11293), .QN(n11290) );
  INVX0 U11356 ( .INP(n11294), .ZN(n11293) );
  NAND2X0 U11357 ( .IN1(test_so69), .IN2(WX8563), .QN(n11294) );
  NOR2X0 U11358 ( .IN1(WX8563), .IN2(test_so69), .QN(n11292) );
  NAND2X0 U11359 ( .IN1(n9094), .IN2(n11295), .QN(n11285) );
  NAND2X0 U11360 ( .IN1(n1232), .IN2(n9277), .QN(n11284) );
  NOR2X0 U11361 ( .IN1(n9224), .IN2(n8901), .QN(n1232) );
  NAND2X0 U11362 ( .IN1(n9309), .IN2(CRC_OUT_4_15), .QN(n11283) );
  NAND4X0 U11363 ( .IN1(n11296), .IN2(n11297), .IN3(n11298), .IN4(n11299), 
        .QN(WX7139) );
  NAND2X0 U11364 ( .IN1(n11300), .IN2(n10614), .QN(n11299) );
  NAND2X0 U11365 ( .IN1(n11301), .IN2(n10617), .QN(n10614) );
  NAND2X0 U11366 ( .IN1(n11302), .IN2(n11303), .QN(n11301) );
  NAND2X0 U11367 ( .IN1(n16397), .IN2(n9120), .QN(n11303) );
  NAND2X0 U11368 ( .IN1(TM1), .IN2(n8363), .QN(n11302) );
  NAND3X0 U11369 ( .IN1(n11304), .IN2(n11305), .IN3(n11306), .QN(n11300) );
  NAND2X0 U11370 ( .IN1(n9332), .IN2(n10617), .QN(n11306) );
  NAND2X0 U11371 ( .IN1(n11307), .IN2(n11308), .QN(n10617) );
  NAND2X0 U11372 ( .IN1(n7684), .IN2(n11309), .QN(n11308) );
  INVX0 U11373 ( .INP(n11310), .ZN(n11307) );
  NOR2X0 U11374 ( .IN1(n11309), .IN2(n7684), .QN(n11310) );
  NOR2X0 U11375 ( .IN1(n11311), .IN2(n11312), .QN(n11309) );
  NOR2X0 U11376 ( .IN1(WX8625), .IN2(n7685), .QN(n11312) );
  INVX0 U11377 ( .INP(n11313), .ZN(n11311) );
  NAND2X0 U11378 ( .IN1(n7685), .IN2(WX8625), .QN(n11313) );
  NAND2X0 U11379 ( .IN1(n9082), .IN2(n8363), .QN(n11305) );
  NAND2X0 U11380 ( .IN1(n16397), .IN2(n10069), .QN(n11304) );
  NAND2X0 U11381 ( .IN1(n11314), .IN2(n11315), .QN(n11298) );
  NAND2X0 U11382 ( .IN1(n11316), .IN2(n11317), .QN(n11314) );
  NAND2X0 U11383 ( .IN1(n9092), .IN2(n11318), .QN(n11317) );
  NAND2X0 U11384 ( .IN1(n9092), .IN2(n8421), .QN(n11316) );
  NAND2X0 U11385 ( .IN1(n1231), .IN2(n9277), .QN(n11297) );
  NOR2X0 U11386 ( .IN1(n9224), .IN2(n8902), .QN(n1231) );
  NAND2X0 U11387 ( .IN1(n9310), .IN2(CRC_OUT_4_16), .QN(n11296) );
  NAND4X0 U11388 ( .IN1(n11319), .IN2(n11320), .IN3(n11321), .IN4(n11322), 
        .QN(WX7137) );
  NAND2X0 U11389 ( .IN1(n11323), .IN2(n10653), .QN(n11322) );
  NAND2X0 U11390 ( .IN1(n11324), .IN2(n10656), .QN(n10653) );
  NAND2X0 U11391 ( .IN1(n11325), .IN2(n11326), .QN(n11324) );
  NAND2X0 U11392 ( .IN1(n16396), .IN2(n9120), .QN(n11326) );
  NAND2X0 U11393 ( .IN1(TM1), .IN2(n8364), .QN(n11325) );
  NAND3X0 U11394 ( .IN1(n11327), .IN2(n11328), .IN3(n11329), .QN(n11323) );
  NAND2X0 U11395 ( .IN1(n9332), .IN2(n10656), .QN(n11329) );
  NAND2X0 U11396 ( .IN1(n11330), .IN2(n11331), .QN(n10656) );
  NAND2X0 U11397 ( .IN1(n7686), .IN2(n11332), .QN(n11331) );
  INVX0 U11398 ( .INP(n11333), .ZN(n11330) );
  NOR2X0 U11399 ( .IN1(n11332), .IN2(n7686), .QN(n11333) );
  NOR2X0 U11400 ( .IN1(n11334), .IN2(n11335), .QN(n11332) );
  NOR2X0 U11401 ( .IN1(WX8623), .IN2(n7687), .QN(n11335) );
  INVX0 U11402 ( .INP(n11336), .ZN(n11334) );
  NAND2X0 U11403 ( .IN1(n7687), .IN2(WX8623), .QN(n11336) );
  NAND2X0 U11404 ( .IN1(n10068), .IN2(n8364), .QN(n11328) );
  NAND2X0 U11405 ( .IN1(n16396), .IN2(n9080), .QN(n11327) );
  NAND2X0 U11406 ( .IN1(n11337), .IN2(n11338), .QN(n11321) );
  NAND2X0 U11407 ( .IN1(n11339), .IN2(n11340), .QN(n11337) );
  NAND2X0 U11408 ( .IN1(n9092), .IN2(n11341), .QN(n11340) );
  NAND2X0 U11409 ( .IN1(n9093), .IN2(n8422), .QN(n11339) );
  NAND2X0 U11410 ( .IN1(n1230), .IN2(n9277), .QN(n11320) );
  NOR2X0 U11411 ( .IN1(n9224), .IN2(n8903), .QN(n1230) );
  NAND2X0 U11412 ( .IN1(n9310), .IN2(CRC_OUT_4_17), .QN(n11319) );
  NAND4X0 U11413 ( .IN1(n11342), .IN2(n11343), .IN3(n11344), .IN4(n11345), 
        .QN(WX7135) );
  NAND2X0 U11414 ( .IN1(n11346), .IN2(n10662), .QN(n11345) );
  NAND2X0 U11415 ( .IN1(n11347), .IN2(n10665), .QN(n10662) );
  NAND2X0 U11416 ( .IN1(n11348), .IN2(n11349), .QN(n11347) );
  NAND2X0 U11417 ( .IN1(n16395), .IN2(n9120), .QN(n11349) );
  NAND2X0 U11418 ( .IN1(TM1), .IN2(n8365), .QN(n11348) );
  NAND3X0 U11419 ( .IN1(n11350), .IN2(n11351), .IN3(n11352), .QN(n11346) );
  NAND2X0 U11420 ( .IN1(n9332), .IN2(n10665), .QN(n11352) );
  NAND2X0 U11421 ( .IN1(n11353), .IN2(n11354), .QN(n10665) );
  NAND2X0 U11422 ( .IN1(n7688), .IN2(n11355), .QN(n11354) );
  INVX0 U11423 ( .INP(n11356), .ZN(n11353) );
  NOR2X0 U11424 ( .IN1(n11355), .IN2(n7688), .QN(n11356) );
  NOR2X0 U11425 ( .IN1(n11357), .IN2(n11358), .QN(n11355) );
  NOR2X0 U11426 ( .IN1(WX8621), .IN2(n7689), .QN(n11358) );
  INVX0 U11427 ( .INP(n11359), .ZN(n11357) );
  NAND2X0 U11428 ( .IN1(n7689), .IN2(WX8621), .QN(n11359) );
  NAND2X0 U11429 ( .IN1(n9084), .IN2(n8365), .QN(n11351) );
  NAND2X0 U11430 ( .IN1(n16395), .IN2(n9079), .QN(n11350) );
  NAND2X0 U11431 ( .IN1(n11360), .IN2(n11361), .QN(n11344) );
  NAND2X0 U11432 ( .IN1(n11362), .IN2(n11363), .QN(n11360) );
  NAND2X0 U11433 ( .IN1(n9092), .IN2(n11364), .QN(n11363) );
  NAND2X0 U11434 ( .IN1(n9093), .IN2(n8423), .QN(n11362) );
  NAND2X0 U11435 ( .IN1(n1229), .IN2(n9277), .QN(n11343) );
  NOR2X0 U11436 ( .IN1(n9225), .IN2(n8904), .QN(n1229) );
  NAND2X0 U11437 ( .IN1(n9310), .IN2(CRC_OUT_4_18), .QN(n11342) );
  NAND4X0 U11438 ( .IN1(n11365), .IN2(n11366), .IN3(n11367), .IN4(n11368), 
        .QN(WX7133) );
  NAND2X0 U11439 ( .IN1(n11369), .IN2(n10701), .QN(n11368) );
  NAND2X0 U11440 ( .IN1(n11370), .IN2(n10704), .QN(n10701) );
  NAND2X0 U11441 ( .IN1(n11371), .IN2(n11372), .QN(n11370) );
  NAND2X0 U11442 ( .IN1(n16394), .IN2(n9120), .QN(n11372) );
  NAND2X0 U11443 ( .IN1(TM1), .IN2(n8366), .QN(n11371) );
  NAND3X0 U11444 ( .IN1(n11373), .IN2(n11374), .IN3(n11375), .QN(n11369) );
  NAND2X0 U11445 ( .IN1(n9332), .IN2(n10704), .QN(n11375) );
  NAND2X0 U11446 ( .IN1(n11376), .IN2(n11377), .QN(n10704) );
  NAND2X0 U11447 ( .IN1(n7690), .IN2(n11378), .QN(n11377) );
  INVX0 U11448 ( .INP(n11379), .ZN(n11376) );
  NOR2X0 U11449 ( .IN1(n11378), .IN2(n7690), .QN(n11379) );
  NOR2X0 U11450 ( .IN1(n11380), .IN2(n11381), .QN(n11378) );
  NOR2X0 U11451 ( .IN1(WX8619), .IN2(n7691), .QN(n11381) );
  INVX0 U11452 ( .INP(n11382), .ZN(n11380) );
  NAND2X0 U11453 ( .IN1(n7691), .IN2(WX8619), .QN(n11382) );
  NAND2X0 U11454 ( .IN1(n9083), .IN2(n8366), .QN(n11374) );
  NAND2X0 U11455 ( .IN1(n16394), .IN2(n9078), .QN(n11373) );
  NAND2X0 U11456 ( .IN1(n11383), .IN2(n11384), .QN(n11367) );
  NAND2X0 U11457 ( .IN1(n11385), .IN2(n11386), .QN(n11383) );
  NAND2X0 U11458 ( .IN1(n9092), .IN2(n11387), .QN(n11386) );
  NAND2X0 U11459 ( .IN1(n9093), .IN2(n8424), .QN(n11385) );
  NAND2X0 U11460 ( .IN1(n1228), .IN2(n9277), .QN(n11366) );
  NOR2X0 U11461 ( .IN1(n9225), .IN2(n8905), .QN(n1228) );
  NAND2X0 U11462 ( .IN1(n9309), .IN2(CRC_OUT_4_19), .QN(n11365) );
  NAND4X0 U11463 ( .IN1(n11388), .IN2(n11389), .IN3(n11390), .IN4(n11391), 
        .QN(WX7131) );
  NAND2X0 U11464 ( .IN1(n11392), .IN2(n10721), .QN(n11391) );
  NAND2X0 U11465 ( .IN1(n11393), .IN2(n10724), .QN(n10721) );
  NAND2X0 U11466 ( .IN1(n11394), .IN2(n11395), .QN(n11393) );
  NAND2X0 U11467 ( .IN1(n16393), .IN2(n9120), .QN(n11395) );
  NAND2X0 U11468 ( .IN1(TM1), .IN2(n8367), .QN(n11394) );
  NAND3X0 U11469 ( .IN1(n11396), .IN2(n11397), .IN3(n11398), .QN(n11392) );
  NAND2X0 U11470 ( .IN1(n9332), .IN2(n10724), .QN(n11398) );
  NAND2X0 U11471 ( .IN1(n11399), .IN2(n11400), .QN(n10724) );
  NAND2X0 U11472 ( .IN1(n7692), .IN2(n11401), .QN(n11400) );
  INVX0 U11473 ( .INP(n11402), .ZN(n11399) );
  NOR2X0 U11474 ( .IN1(n11401), .IN2(n7692), .QN(n11402) );
  NOR2X0 U11475 ( .IN1(n11403), .IN2(n11404), .QN(n11401) );
  NOR2X0 U11476 ( .IN1(WX8617), .IN2(n7693), .QN(n11404) );
  INVX0 U11477 ( .INP(n11405), .ZN(n11403) );
  NAND2X0 U11478 ( .IN1(n7693), .IN2(WX8617), .QN(n11405) );
  NAND2X0 U11479 ( .IN1(n9082), .IN2(n8367), .QN(n11397) );
  NAND2X0 U11480 ( .IN1(n16393), .IN2(n10069), .QN(n11396) );
  NAND2X0 U11481 ( .IN1(n11406), .IN2(n11407), .QN(n11390) );
  NAND2X0 U11482 ( .IN1(n11408), .IN2(n11409), .QN(n11406) );
  NAND2X0 U11483 ( .IN1(n9093), .IN2(n11410), .QN(n11409) );
  NAND2X0 U11484 ( .IN1(n9092), .IN2(n8425), .QN(n11408) );
  NAND2X0 U11485 ( .IN1(n1227), .IN2(n9277), .QN(n11389) );
  NOR2X0 U11486 ( .IN1(n9225), .IN2(n8906), .QN(n1227) );
  NAND2X0 U11487 ( .IN1(n9310), .IN2(CRC_OUT_4_20), .QN(n11388) );
  NAND4X0 U11488 ( .IN1(n11411), .IN2(n11412), .IN3(n11413), .IN4(n11414), 
        .QN(WX7129) );
  NAND2X0 U11489 ( .IN1(n11415), .IN2(n10744), .QN(n11414) );
  NAND2X0 U11490 ( .IN1(n11416), .IN2(n10747), .QN(n10744) );
  NAND2X0 U11491 ( .IN1(n11417), .IN2(n11418), .QN(n11416) );
  NAND2X0 U11492 ( .IN1(n16392), .IN2(n9120), .QN(n11418) );
  NAND2X0 U11493 ( .IN1(TM1), .IN2(n8368), .QN(n11417) );
  NAND3X0 U11494 ( .IN1(n11419), .IN2(n11420), .IN3(n11421), .QN(n11415) );
  NAND2X0 U11495 ( .IN1(n9332), .IN2(n10747), .QN(n11421) );
  NAND2X0 U11496 ( .IN1(n11422), .IN2(n11423), .QN(n10747) );
  NAND2X0 U11497 ( .IN1(n7694), .IN2(n11424), .QN(n11423) );
  INVX0 U11498 ( .INP(n11425), .ZN(n11422) );
  NOR2X0 U11499 ( .IN1(n11424), .IN2(n7694), .QN(n11425) );
  NOR2X0 U11500 ( .IN1(n11426), .IN2(n11427), .QN(n11424) );
  NOR2X0 U11501 ( .IN1(WX8615), .IN2(n7695), .QN(n11427) );
  INVX0 U11502 ( .INP(n11428), .ZN(n11426) );
  NAND2X0 U11503 ( .IN1(n7695), .IN2(WX8615), .QN(n11428) );
  NAND2X0 U11504 ( .IN1(n10068), .IN2(n8368), .QN(n11420) );
  NAND2X0 U11505 ( .IN1(n16392), .IN2(n9080), .QN(n11419) );
  NAND2X0 U11506 ( .IN1(n11429), .IN2(n9112), .QN(n11413) );
  NAND2X0 U11507 ( .IN1(n1226), .IN2(n9277), .QN(n11412) );
  NOR2X0 U11508 ( .IN1(n9225), .IN2(n8907), .QN(n1226) );
  NAND2X0 U11509 ( .IN1(n9310), .IN2(CRC_OUT_4_21), .QN(n11411) );
  NAND4X0 U11510 ( .IN1(n11430), .IN2(n11431), .IN3(n11432), .IN4(n11433), 
        .QN(WX7127) );
  NAND2X0 U11511 ( .IN1(n11434), .IN2(n10767), .QN(n11433) );
  NAND2X0 U11512 ( .IN1(n11435), .IN2(n10770), .QN(n10767) );
  NAND2X0 U11513 ( .IN1(n11436), .IN2(n11437), .QN(n11435) );
  NAND2X0 U11514 ( .IN1(n16391), .IN2(n9120), .QN(n11437) );
  NAND2X0 U11515 ( .IN1(TM1), .IN2(n8369), .QN(n11436) );
  NAND3X0 U11516 ( .IN1(n11438), .IN2(n11439), .IN3(n11440), .QN(n11434) );
  NAND2X0 U11517 ( .IN1(n9332), .IN2(n10770), .QN(n11440) );
  NAND2X0 U11518 ( .IN1(n11441), .IN2(n11442), .QN(n10770) );
  NAND2X0 U11519 ( .IN1(n7696), .IN2(n11443), .QN(n11442) );
  INVX0 U11520 ( .INP(n11444), .ZN(n11441) );
  NOR2X0 U11521 ( .IN1(n11443), .IN2(n7696), .QN(n11444) );
  NOR2X0 U11522 ( .IN1(n11445), .IN2(n11446), .QN(n11443) );
  NOR2X0 U11523 ( .IN1(WX8613), .IN2(n7697), .QN(n11446) );
  INVX0 U11524 ( .INP(n11447), .ZN(n11445) );
  NAND2X0 U11525 ( .IN1(n7697), .IN2(WX8613), .QN(n11447) );
  NAND2X0 U11526 ( .IN1(n9084), .IN2(n8369), .QN(n11439) );
  NAND2X0 U11527 ( .IN1(n16391), .IN2(n9079), .QN(n11438) );
  NAND2X0 U11528 ( .IN1(n11448), .IN2(n11449), .QN(n11432) );
  NAND2X0 U11529 ( .IN1(n11450), .IN2(n11451), .QN(n11448) );
  NAND2X0 U11530 ( .IN1(n9092), .IN2(n11452), .QN(n11451) );
  NAND2X0 U11531 ( .IN1(n9093), .IN2(n8427), .QN(n11450) );
  NAND2X0 U11532 ( .IN1(n1225), .IN2(n9278), .QN(n11431) );
  NOR2X0 U11533 ( .IN1(n9225), .IN2(n8908), .QN(n1225) );
  NAND2X0 U11534 ( .IN1(n9310), .IN2(CRC_OUT_4_22), .QN(n11430) );
  NAND4X0 U11535 ( .IN1(n11453), .IN2(n11454), .IN3(n11455), .IN4(n11456), 
        .QN(WX7125) );
  NAND2X0 U11536 ( .IN1(n11457), .IN2(n10790), .QN(n11456) );
  NAND2X0 U11537 ( .IN1(n11458), .IN2(n10793), .QN(n10790) );
  NAND2X0 U11538 ( .IN1(n11459), .IN2(n11460), .QN(n11458) );
  NAND2X0 U11539 ( .IN1(n16390), .IN2(n9120), .QN(n11460) );
  NAND2X0 U11540 ( .IN1(TM1), .IN2(n8370), .QN(n11459) );
  NAND3X0 U11541 ( .IN1(n11461), .IN2(n11462), .IN3(n11463), .QN(n11457) );
  NAND2X0 U11542 ( .IN1(n9332), .IN2(n10793), .QN(n11463) );
  NAND2X0 U11543 ( .IN1(n11464), .IN2(n11465), .QN(n10793) );
  NAND2X0 U11544 ( .IN1(n7698), .IN2(n11466), .QN(n11465) );
  INVX0 U11545 ( .INP(n11467), .ZN(n11464) );
  NOR2X0 U11546 ( .IN1(n11466), .IN2(n7698), .QN(n11467) );
  NOR2X0 U11547 ( .IN1(n11468), .IN2(n11469), .QN(n11466) );
  NOR2X0 U11548 ( .IN1(WX8611), .IN2(n7699), .QN(n11469) );
  INVX0 U11549 ( .INP(n11470), .ZN(n11468) );
  NAND2X0 U11550 ( .IN1(n7699), .IN2(WX8611), .QN(n11470) );
  NAND2X0 U11551 ( .IN1(n9083), .IN2(n8370), .QN(n11462) );
  NAND2X0 U11552 ( .IN1(n16390), .IN2(n9078), .QN(n11461) );
  NAND2X0 U11553 ( .IN1(n11471), .IN2(n9111), .QN(n11455) );
  NAND2X0 U11554 ( .IN1(n1224), .IN2(n9278), .QN(n11454) );
  NOR2X0 U11555 ( .IN1(n9225), .IN2(n8909), .QN(n1224) );
  NAND2X0 U11556 ( .IN1(n9310), .IN2(CRC_OUT_4_23), .QN(n11453) );
  NAND4X0 U11557 ( .IN1(n11472), .IN2(n11473), .IN3(n11474), .IN4(n11475), 
        .QN(WX7123) );
  NAND2X0 U11558 ( .IN1(n11476), .IN2(n10813), .QN(n11475) );
  NAND2X0 U11559 ( .IN1(n11477), .IN2(n10816), .QN(n10813) );
  NAND2X0 U11560 ( .IN1(n11478), .IN2(n11479), .QN(n11477) );
  NAND2X0 U11561 ( .IN1(n16389), .IN2(n9120), .QN(n11479) );
  NAND2X0 U11562 ( .IN1(TM1), .IN2(n8371), .QN(n11478) );
  NAND3X0 U11563 ( .IN1(n11480), .IN2(n11481), .IN3(n11482), .QN(n11476) );
  NAND2X0 U11564 ( .IN1(n9333), .IN2(n10816), .QN(n11482) );
  NAND2X0 U11565 ( .IN1(n11483), .IN2(n11484), .QN(n10816) );
  NAND2X0 U11566 ( .IN1(n7700), .IN2(n11485), .QN(n11484) );
  INVX0 U11567 ( .INP(n11486), .ZN(n11483) );
  NOR2X0 U11568 ( .IN1(n11485), .IN2(n7700), .QN(n11486) );
  NOR2X0 U11569 ( .IN1(n11487), .IN2(n11488), .QN(n11485) );
  NOR2X0 U11570 ( .IN1(WX8609), .IN2(n7701), .QN(n11488) );
  INVX0 U11571 ( .INP(n11489), .ZN(n11487) );
  NAND2X0 U11572 ( .IN1(n7701), .IN2(WX8609), .QN(n11489) );
  NAND2X0 U11573 ( .IN1(n9082), .IN2(n8371), .QN(n11481) );
  NAND2X0 U11574 ( .IN1(n16389), .IN2(n10069), .QN(n11480) );
  NAND2X0 U11575 ( .IN1(n11490), .IN2(n11491), .QN(n11474) );
  NAND2X0 U11576 ( .IN1(n11492), .IN2(n11493), .QN(n11490) );
  NAND2X0 U11577 ( .IN1(n9092), .IN2(n11494), .QN(n11493) );
  NAND2X0 U11578 ( .IN1(n9092), .IN2(n8429), .QN(n11492) );
  NAND2X0 U11579 ( .IN1(n1223), .IN2(n9278), .QN(n11473) );
  NOR2X0 U11580 ( .IN1(n9225), .IN2(n8910), .QN(n1223) );
  NAND2X0 U11581 ( .IN1(n9310), .IN2(CRC_OUT_4_24), .QN(n11472) );
  NAND4X0 U11582 ( .IN1(n11495), .IN2(n11496), .IN3(n11497), .IN4(n11498), 
        .QN(WX7121) );
  NAND2X0 U11583 ( .IN1(n11499), .IN2(n10836), .QN(n11498) );
  NAND2X0 U11584 ( .IN1(n11500), .IN2(n10839), .QN(n10836) );
  NAND2X0 U11585 ( .IN1(n11501), .IN2(n11502), .QN(n11500) );
  NAND2X0 U11586 ( .IN1(n16388), .IN2(n9120), .QN(n11502) );
  NAND2X0 U11587 ( .IN1(TM1), .IN2(n8372), .QN(n11501) );
  NAND3X0 U11588 ( .IN1(n11503), .IN2(n11504), .IN3(n11505), .QN(n11499) );
  NAND2X0 U11589 ( .IN1(n9333), .IN2(n10839), .QN(n11505) );
  NAND2X0 U11590 ( .IN1(n11506), .IN2(n11507), .QN(n10839) );
  NAND2X0 U11591 ( .IN1(n7702), .IN2(n11508), .QN(n11507) );
  INVX0 U11592 ( .INP(n11509), .ZN(n11506) );
  NOR2X0 U11593 ( .IN1(n11508), .IN2(n7702), .QN(n11509) );
  NOR2X0 U11594 ( .IN1(n11510), .IN2(n11511), .QN(n11508) );
  NOR2X0 U11595 ( .IN1(WX8607), .IN2(n7703), .QN(n11511) );
  INVX0 U11596 ( .INP(n11512), .ZN(n11510) );
  NAND2X0 U11597 ( .IN1(n7703), .IN2(WX8607), .QN(n11512) );
  NAND2X0 U11598 ( .IN1(n10068), .IN2(n8372), .QN(n11504) );
  NAND2X0 U11599 ( .IN1(n16388), .IN2(n9080), .QN(n11503) );
  NAND2X0 U11600 ( .IN1(n11513), .IN2(n9111), .QN(n11497) );
  NAND2X0 U11601 ( .IN1(n1222), .IN2(n9278), .QN(n11496) );
  NOR2X0 U11602 ( .IN1(n9225), .IN2(n8911), .QN(n1222) );
  NAND2X0 U11603 ( .IN1(n9310), .IN2(CRC_OUT_4_25), .QN(n11495) );
  NAND4X0 U11604 ( .IN1(n11514), .IN2(n11515), .IN3(n11516), .IN4(n11517), 
        .QN(WX7119) );
  NAND2X0 U11605 ( .IN1(n11518), .IN2(n11519), .QN(n11517) );
  NAND2X0 U11606 ( .IN1(n11520), .IN2(n11521), .QN(n11518) );
  NAND2X0 U11607 ( .IN1(n9093), .IN2(n11522), .QN(n11521) );
  NAND2X0 U11608 ( .IN1(n9092), .IN2(n8431), .QN(n11520) );
  NAND2X0 U11609 ( .IN1(n10858), .IN2(n2153), .QN(n11516) );
  NOR2X0 U11610 ( .IN1(n11523), .IN2(n11524), .QN(n10858) );
  INVX0 U11611 ( .INP(n11525), .ZN(n11524) );
  NAND2X0 U11612 ( .IN1(n11526), .IN2(n11527), .QN(n11525) );
  NOR2X0 U11613 ( .IN1(n11527), .IN2(n11526), .QN(n11523) );
  NAND2X0 U11614 ( .IN1(n11528), .IN2(n11529), .QN(n11526) );
  NAND2X0 U11615 ( .IN1(n11530), .IN2(WX8541), .QN(n11529) );
  NAND2X0 U11616 ( .IN1(n11531), .IN2(n11532), .QN(n11530) );
  NAND3X0 U11617 ( .IN1(n11531), .IN2(n11532), .IN3(n7705), .QN(n11528) );
  NAND2X0 U11618 ( .IN1(test_so74), .IN2(WX8477), .QN(n11532) );
  NAND2X0 U11619 ( .IN1(n7704), .IN2(n8799), .QN(n11531) );
  NOR2X0 U11620 ( .IN1(n11533), .IN2(n11534), .QN(n11527) );
  INVX0 U11621 ( .INP(n11535), .ZN(n11534) );
  NAND2X0 U11622 ( .IN1(n16387), .IN2(n9120), .QN(n11535) );
  NOR2X0 U11623 ( .IN1(n9118), .IN2(n16387), .QN(n11533) );
  NAND2X0 U11624 ( .IN1(n1221), .IN2(n9278), .QN(n11515) );
  NOR2X0 U11625 ( .IN1(n9225), .IN2(n8912), .QN(n1221) );
  NAND2X0 U11626 ( .IN1(n9311), .IN2(CRC_OUT_4_26), .QN(n11514) );
  NAND4X0 U11627 ( .IN1(n11536), .IN2(n11537), .IN3(n11538), .IN4(n11539), 
        .QN(WX7117) );
  NAND2X0 U11628 ( .IN1(n11540), .IN2(n10878), .QN(n11539) );
  NAND2X0 U11629 ( .IN1(n11541), .IN2(n10881), .QN(n10878) );
  NAND2X0 U11630 ( .IN1(n11542), .IN2(n11543), .QN(n11541) );
  NAND2X0 U11631 ( .IN1(n16386), .IN2(n9120), .QN(n11543) );
  NAND2X0 U11632 ( .IN1(TM1), .IN2(n8374), .QN(n11542) );
  NAND3X0 U11633 ( .IN1(n11544), .IN2(n11545), .IN3(n11546), .QN(n11540) );
  NAND2X0 U11634 ( .IN1(n9333), .IN2(n10881), .QN(n11546) );
  NAND2X0 U11635 ( .IN1(n11547), .IN2(n11548), .QN(n10881) );
  NAND2X0 U11636 ( .IN1(n7706), .IN2(n11549), .QN(n11548) );
  INVX0 U11637 ( .INP(n11550), .ZN(n11547) );
  NOR2X0 U11638 ( .IN1(n11549), .IN2(n7706), .QN(n11550) );
  NOR2X0 U11639 ( .IN1(n11551), .IN2(n11552), .QN(n11549) );
  NOR2X0 U11640 ( .IN1(WX8603), .IN2(n7707), .QN(n11552) );
  INVX0 U11641 ( .INP(n11553), .ZN(n11551) );
  NAND2X0 U11642 ( .IN1(n7707), .IN2(WX8603), .QN(n11553) );
  NAND2X0 U11643 ( .IN1(n9084), .IN2(n8374), .QN(n11545) );
  NAND2X0 U11644 ( .IN1(n16386), .IN2(n9079), .QN(n11544) );
  NAND2X0 U11645 ( .IN1(n11554), .IN2(n11555), .QN(n11538) );
  NAND2X0 U11646 ( .IN1(n11556), .IN2(n11557), .QN(n11554) );
  NAND2X0 U11647 ( .IN1(n9093), .IN2(n11558), .QN(n11557) );
  NAND2X0 U11648 ( .IN1(n8216), .IN2(n9111), .QN(n11556) );
  NAND2X0 U11649 ( .IN1(n1220), .IN2(n9278), .QN(n11537) );
  NOR2X0 U11650 ( .IN1(n9225), .IN2(n8913), .QN(n1220) );
  NAND2X0 U11651 ( .IN1(n9311), .IN2(CRC_OUT_4_27), .QN(n11536) );
  NAND4X0 U11652 ( .IN1(n11559), .IN2(n11560), .IN3(n11561), .IN4(n11562), 
        .QN(WX7115) );
  NAND2X0 U11653 ( .IN1(n11563), .IN2(n11564), .QN(n11562) );
  NAND2X0 U11654 ( .IN1(n11565), .IN2(n11566), .QN(n11563) );
  NAND2X0 U11655 ( .IN1(n9093), .IN2(n11567), .QN(n11566) );
  NAND2X0 U11656 ( .IN1(n9093), .IN2(n8434), .QN(n11565) );
  NAND2X0 U11657 ( .IN1(n10900), .IN2(n2153), .QN(n11561) );
  NOR2X0 U11658 ( .IN1(n11568), .IN2(n11569), .QN(n10900) );
  INVX0 U11659 ( .INP(n11570), .ZN(n11569) );
  NAND2X0 U11660 ( .IN1(n11571), .IN2(n11572), .QN(n11570) );
  NOR2X0 U11661 ( .IN1(n11572), .IN2(n11571), .QN(n11568) );
  NAND2X0 U11662 ( .IN1(n11573), .IN2(n11574), .QN(n11571) );
  NAND2X0 U11663 ( .IN1(n8189), .IN2(n11575), .QN(n11574) );
  INVX0 U11664 ( .INP(n11576), .ZN(n11575) );
  NAND2X0 U11665 ( .IN1(n11576), .IN2(WX8601), .QN(n11573) );
  NAND2X0 U11666 ( .IN1(n11577), .IN2(n11578), .QN(n11576) );
  INVX0 U11667 ( .INP(n11579), .ZN(n11578) );
  NOR2X0 U11668 ( .IN1(n8808), .IN2(n16385), .QN(n11579) );
  NAND2X0 U11669 ( .IN1(n16385), .IN2(n8808), .QN(n11577) );
  NOR2X0 U11670 ( .IN1(n11580), .IN2(n11581), .QN(n11572) );
  INVX0 U11671 ( .INP(n11582), .ZN(n11581) );
  NAND2X0 U11672 ( .IN1(n7708), .IN2(n9120), .QN(n11582) );
  NOR2X0 U11673 ( .IN1(n9117), .IN2(n7708), .QN(n11580) );
  NAND2X0 U11674 ( .IN1(n1219), .IN2(n9278), .QN(n11560) );
  NOR2X0 U11675 ( .IN1(n9225), .IN2(n8914), .QN(n1219) );
  NAND2X0 U11676 ( .IN1(n9311), .IN2(CRC_OUT_4_28), .QN(n11559) );
  NAND4X0 U11677 ( .IN1(n11583), .IN2(n11584), .IN3(n11585), .IN4(n11586), 
        .QN(WX7113) );
  NAND2X0 U11678 ( .IN1(n11587), .IN2(n10920), .QN(n11586) );
  NAND2X0 U11679 ( .IN1(n11588), .IN2(n10923), .QN(n10920) );
  NAND2X0 U11680 ( .IN1(n11589), .IN2(n11590), .QN(n11588) );
  NAND2X0 U11681 ( .IN1(n16384), .IN2(n9120), .QN(n11590) );
  NAND2X0 U11682 ( .IN1(TM1), .IN2(n8376), .QN(n11589) );
  NAND3X0 U11683 ( .IN1(n11591), .IN2(n11592), .IN3(n11593), .QN(n11587) );
  NAND2X0 U11684 ( .IN1(n9333), .IN2(n10923), .QN(n11593) );
  NAND2X0 U11685 ( .IN1(n11594), .IN2(n11595), .QN(n10923) );
  NAND2X0 U11686 ( .IN1(n7709), .IN2(n11596), .QN(n11595) );
  INVX0 U11687 ( .INP(n11597), .ZN(n11594) );
  NOR2X0 U11688 ( .IN1(n11596), .IN2(n7709), .QN(n11597) );
  NOR2X0 U11689 ( .IN1(n11598), .IN2(n11599), .QN(n11596) );
  NOR2X0 U11690 ( .IN1(WX8599), .IN2(n7710), .QN(n11599) );
  INVX0 U11691 ( .INP(n11600), .ZN(n11598) );
  NAND2X0 U11692 ( .IN1(n7710), .IN2(WX8599), .QN(n11600) );
  NAND2X0 U11693 ( .IN1(n9083), .IN2(n8376), .QN(n11592) );
  NAND2X0 U11694 ( .IN1(n16384), .IN2(n9078), .QN(n11591) );
  NAND2X0 U11695 ( .IN1(n11601), .IN2(n11602), .QN(n11585) );
  NAND2X0 U11696 ( .IN1(n11603), .IN2(n11604), .QN(n11601) );
  NAND2X0 U11697 ( .IN1(n9093), .IN2(n11605), .QN(n11604) );
  NAND2X0 U11698 ( .IN1(n9093), .IN2(n8435), .QN(n11603) );
  NAND2X0 U11699 ( .IN1(n1218), .IN2(n9278), .QN(n11584) );
  NOR2X0 U11700 ( .IN1(n9066), .IN2(n9164), .QN(n1218) );
  NAND2X0 U11701 ( .IN1(test_so66), .IN2(n9315), .QN(n11583) );
  NAND4X0 U11702 ( .IN1(n11606), .IN2(n11607), .IN3(n11608), .IN4(n11609), 
        .QN(WX7111) );
  NAND2X0 U11703 ( .IN1(n11610), .IN2(n11611), .QN(n11609) );
  NAND2X0 U11704 ( .IN1(n11612), .IN2(n11613), .QN(n11610) );
  NAND2X0 U11705 ( .IN1(n9093), .IN2(n11614), .QN(n11613) );
  NAND2X0 U11706 ( .IN1(n9093), .IN2(n8436), .QN(n11612) );
  NAND2X0 U11707 ( .IN1(n10942), .IN2(n2153), .QN(n11608) );
  NOR2X0 U11708 ( .IN1(n11615), .IN2(n11616), .QN(n10942) );
  INVX0 U11709 ( .INP(n11617), .ZN(n11616) );
  NAND2X0 U11710 ( .IN1(n11618), .IN2(n11619), .QN(n11617) );
  NOR2X0 U11711 ( .IN1(n11619), .IN2(n11618), .QN(n11615) );
  NAND2X0 U11712 ( .IN1(n11620), .IN2(n11621), .QN(n11618) );
  NAND2X0 U11713 ( .IN1(n8187), .IN2(n11622), .QN(n11621) );
  INVX0 U11714 ( .INP(n11623), .ZN(n11622) );
  NAND2X0 U11715 ( .IN1(n11623), .IN2(WX8597), .QN(n11620) );
  NAND2X0 U11716 ( .IN1(n11624), .IN2(n11625), .QN(n11623) );
  INVX0 U11717 ( .INP(n11626), .ZN(n11625) );
  NOR2X0 U11718 ( .IN1(n8809), .IN2(n16383), .QN(n11626) );
  NAND2X0 U11719 ( .IN1(n16383), .IN2(n8809), .QN(n11624) );
  NOR2X0 U11720 ( .IN1(n11627), .IN2(n11628), .QN(n11619) );
  INVX0 U11721 ( .INP(n11629), .ZN(n11628) );
  NAND2X0 U11722 ( .IN1(n7711), .IN2(n9119), .QN(n11629) );
  NOR2X0 U11723 ( .IN1(n9118), .IN2(n7711), .QN(n11627) );
  NAND2X0 U11724 ( .IN1(n1217), .IN2(n9278), .QN(n11607) );
  NOR2X0 U11725 ( .IN1(n9225), .IN2(n8915), .QN(n1217) );
  NAND2X0 U11726 ( .IN1(n9311), .IN2(CRC_OUT_4_30), .QN(n11606) );
  NAND4X0 U11727 ( .IN1(n11630), .IN2(n11631), .IN3(n11632), .IN4(n11633), 
        .QN(WX7109) );
  NAND2X0 U11728 ( .IN1(n11634), .IN2(n10948), .QN(n11633) );
  NAND2X0 U11729 ( .IN1(n11635), .IN2(n10951), .QN(n10948) );
  NAND2X0 U11730 ( .IN1(n11636), .IN2(n11637), .QN(n11635) );
  NAND2X0 U11731 ( .IN1(n16382), .IN2(n9119), .QN(n11637) );
  NAND2X0 U11732 ( .IN1(TM1), .IN2(n8378), .QN(n11636) );
  NAND3X0 U11733 ( .IN1(n11638), .IN2(n11639), .IN3(n11640), .QN(n11634) );
  NAND2X0 U11734 ( .IN1(n9333), .IN2(n10951), .QN(n11640) );
  NAND2X0 U11735 ( .IN1(n11641), .IN2(n11642), .QN(n10951) );
  NAND2X0 U11736 ( .IN1(n7616), .IN2(n11643), .QN(n11642) );
  INVX0 U11737 ( .INP(n11644), .ZN(n11641) );
  NOR2X0 U11738 ( .IN1(n11643), .IN2(n7616), .QN(n11644) );
  NOR2X0 U11739 ( .IN1(n11645), .IN2(n11646), .QN(n11643) );
  NOR2X0 U11740 ( .IN1(WX8595), .IN2(n7617), .QN(n11646) );
  INVX0 U11741 ( .INP(n11647), .ZN(n11645) );
  NAND2X0 U11742 ( .IN1(n7617), .IN2(WX8595), .QN(n11647) );
  NAND2X0 U11743 ( .IN1(n9082), .IN2(n8378), .QN(n11639) );
  NAND2X0 U11744 ( .IN1(n16382), .IN2(n10069), .QN(n11638) );
  NAND2X0 U11745 ( .IN1(n11648), .IN2(n11649), .QN(n11632) );
  NAND2X0 U11746 ( .IN1(n11650), .IN2(n11651), .QN(n11648) );
  NAND2X0 U11747 ( .IN1(n9093), .IN2(n11652), .QN(n11651) );
  NAND2X0 U11748 ( .IN1(n9093), .IN2(n8437), .QN(n11650) );
  NAND2X0 U11749 ( .IN1(n9310), .IN2(CRC_OUT_4_31), .QN(n11631) );
  NAND2X0 U11750 ( .IN1(n2245), .IN2(WX6950), .QN(n11630) );
  NAND4X0 U11751 ( .IN1(n11653), .IN2(n11654), .IN3(n11655), .IN4(n11656), 
        .QN(WX706) );
  NAND3X0 U11752 ( .IN1(n11657), .IN2(n11658), .IN3(n9322), .QN(n11656) );
  NAND2X0 U11753 ( .IN1(n9094), .IN2(n11659), .QN(n11655) );
  NAND2X0 U11754 ( .IN1(WX544), .IN2(n9278), .QN(n11654) );
  NAND2X0 U11755 ( .IN1(n9311), .IN2(CRC_OUT_9_0), .QN(n11653) );
  NAND4X0 U11756 ( .IN1(n11660), .IN2(n11661), .IN3(n11662), .IN4(n11663), 
        .QN(WX704) );
  NAND2X0 U11757 ( .IN1(n9333), .IN2(n11664), .QN(n11663) );
  NAND2X0 U11758 ( .IN1(n9093), .IN2(n11665), .QN(n11662) );
  NAND2X0 U11759 ( .IN1(WX542), .IN2(n9278), .QN(n11661) );
  NAND2X0 U11760 ( .IN1(test_so9), .IN2(n9315), .QN(n11660) );
  NAND4X0 U11761 ( .IN1(n11666), .IN2(n11667), .IN3(n11668), .IN4(n11669), 
        .QN(WX702) );
  NAND2X0 U11762 ( .IN1(n9333), .IN2(n11670), .QN(n11669) );
  NAND2X0 U11763 ( .IN1(n11671), .IN2(n9110), .QN(n11668) );
  INVX0 U11764 ( .INP(n11672), .ZN(n11671) );
  NAND2X0 U11765 ( .IN1(WX540), .IN2(n9278), .QN(n11667) );
  NAND2X0 U11766 ( .IN1(n9311), .IN2(CRC_OUT_9_2), .QN(n11666) );
  NOR2X0 U11767 ( .IN1(n9226), .IN2(WX6950), .QN(WX7011) );
  NAND4X0 U11768 ( .IN1(n11673), .IN2(n11674), .IN3(n11675), .IN4(n11676), 
        .QN(WX700) );
  NAND2X0 U11769 ( .IN1(n9333), .IN2(n11677), .QN(n11676) );
  NAND2X0 U11770 ( .IN1(n9093), .IN2(n11678), .QN(n11675) );
  NAND2X0 U11771 ( .IN1(WX538), .IN2(n9278), .QN(n11674) );
  NAND2X0 U11772 ( .IN1(n9310), .IN2(CRC_OUT_9_3), .QN(n11673) );
  NAND4X0 U11773 ( .IN1(n11679), .IN2(n11680), .IN3(n11681), .IN4(n11682), 
        .QN(WX698) );
  NAND3X0 U11774 ( .IN1(n11683), .IN2(n11684), .IN3(n9322), .QN(n11682) );
  NAND2X0 U11775 ( .IN1(n9093), .IN2(n11685), .QN(n11681) );
  NAND2X0 U11776 ( .IN1(WX536), .IN2(n9278), .QN(n11680) );
  NAND2X0 U11777 ( .IN1(n9311), .IN2(CRC_OUT_9_4), .QN(n11679) );
  NAND4X0 U11778 ( .IN1(n11686), .IN2(n11687), .IN3(n11688), .IN4(n11689), 
        .QN(WX696) );
  NAND2X0 U11779 ( .IN1(n9333), .IN2(n11690), .QN(n11689) );
  NAND2X0 U11780 ( .IN1(n9094), .IN2(n11691), .QN(n11688) );
  NAND2X0 U11781 ( .IN1(WX534), .IN2(n9278), .QN(n11687) );
  NAND2X0 U11782 ( .IN1(n9312), .IN2(CRC_OUT_9_5), .QN(n11686) );
  NAND4X0 U11783 ( .IN1(n11692), .IN2(n11693), .IN3(n11694), .IN4(n11695), 
        .QN(WX694) );
  NAND2X0 U11784 ( .IN1(n9333), .IN2(n11696), .QN(n11695) );
  NAND2X0 U11785 ( .IN1(n11697), .IN2(n9112), .QN(n11694) );
  INVX0 U11786 ( .INP(n11698), .ZN(n11697) );
  NAND2X0 U11787 ( .IN1(WX532), .IN2(n9278), .QN(n11693) );
  NAND2X0 U11788 ( .IN1(n9311), .IN2(CRC_OUT_9_6), .QN(n11692) );
  NAND4X0 U11789 ( .IN1(n11699), .IN2(n11700), .IN3(n11701), .IN4(n11702), 
        .QN(WX692) );
  NAND2X0 U11790 ( .IN1(n9333), .IN2(n11703), .QN(n11702) );
  NAND2X0 U11791 ( .IN1(n9094), .IN2(n11704), .QN(n11701) );
  NAND2X0 U11792 ( .IN1(WX530), .IN2(n9278), .QN(n11700) );
  NAND2X0 U11793 ( .IN1(n9312), .IN2(CRC_OUT_9_7), .QN(n11699) );
  NAND4X0 U11794 ( .IN1(n11705), .IN2(n11706), .IN3(n11707), .IN4(n11708), 
        .QN(WX690) );
  NAND2X0 U11795 ( .IN1(n9333), .IN2(n11709), .QN(n11708) );
  NAND2X0 U11796 ( .IN1(n9094), .IN2(n11710), .QN(n11707) );
  NAND2X0 U11797 ( .IN1(WX528), .IN2(n9279), .QN(n11706) );
  NAND2X0 U11798 ( .IN1(n9310), .IN2(CRC_OUT_9_8), .QN(n11705) );
  NAND4X0 U11799 ( .IN1(n11711), .IN2(n11712), .IN3(n11713), .IN4(n11714), 
        .QN(WX688) );
  NAND2X0 U11800 ( .IN1(n9333), .IN2(n11715), .QN(n11714) );
  NAND2X0 U11801 ( .IN1(n9094), .IN2(n11716), .QN(n11713) );
  NAND2X0 U11802 ( .IN1(WX526), .IN2(n9279), .QN(n11712) );
  NAND2X0 U11803 ( .IN1(n9312), .IN2(CRC_OUT_9_9), .QN(n11711) );
  NAND4X0 U11804 ( .IN1(n11717), .IN2(n11718), .IN3(n11719), .IN4(n11720), 
        .QN(WX686) );
  NAND3X0 U11805 ( .IN1(n11721), .IN2(n11722), .IN3(n9322), .QN(n11720) );
  NAND2X0 U11806 ( .IN1(n11723), .IN2(n9111), .QN(n11719) );
  INVX0 U11807 ( .INP(n11724), .ZN(n11723) );
  NAND2X0 U11808 ( .IN1(WX524), .IN2(n9279), .QN(n11718) );
  NAND2X0 U11809 ( .IN1(n9312), .IN2(CRC_OUT_9_10), .QN(n11717) );
  NAND4X0 U11810 ( .IN1(n11725), .IN2(n11726), .IN3(n11727), .IN4(n11728), 
        .QN(WX684) );
  NAND2X0 U11811 ( .IN1(n9333), .IN2(n11729), .QN(n11728) );
  NAND2X0 U11812 ( .IN1(n9094), .IN2(n11730), .QN(n11727) );
  NAND2X0 U11813 ( .IN1(WX522), .IN2(n9279), .QN(n11726) );
  NAND2X0 U11814 ( .IN1(n9312), .IN2(CRC_OUT_9_11), .QN(n11725) );
  NAND4X0 U11815 ( .IN1(n11731), .IN2(n11732), .IN3(n11733), .IN4(n11734), 
        .QN(WX682) );
  NAND2X0 U11816 ( .IN1(n9332), .IN2(n11735), .QN(n11734) );
  NAND2X0 U11817 ( .IN1(n9094), .IN2(n11736), .QN(n11733) );
  NAND2X0 U11818 ( .IN1(WX520), .IN2(n9279), .QN(n11732) );
  NAND2X0 U11819 ( .IN1(n9311), .IN2(CRC_OUT_9_12), .QN(n11731) );
  NAND4X0 U11820 ( .IN1(n11737), .IN2(n11738), .IN3(n11739), .IN4(n11740), 
        .QN(WX680) );
  NAND2X0 U11821 ( .IN1(n9333), .IN2(n11741), .QN(n11740) );
  NAND2X0 U11822 ( .IN1(n9094), .IN2(n11742), .QN(n11739) );
  NAND2X0 U11823 ( .IN1(WX518), .IN2(n9279), .QN(n11738) );
  NAND2X0 U11824 ( .IN1(n9309), .IN2(CRC_OUT_9_13), .QN(n11737) );
  NAND4X0 U11825 ( .IN1(n11743), .IN2(n11744), .IN3(n11745), .IN4(n11746), 
        .QN(WX678) );
  NAND3X0 U11826 ( .IN1(n11747), .IN2(n11748), .IN3(n9322), .QN(n11746) );
  NAND2X0 U11827 ( .IN1(n9094), .IN2(n11749), .QN(n11745) );
  NAND2X0 U11828 ( .IN1(WX516), .IN2(n9279), .QN(n11744) );
  NAND2X0 U11829 ( .IN1(n9311), .IN2(CRC_OUT_9_14), .QN(n11743) );
  NAND4X0 U11830 ( .IN1(n11750), .IN2(n11751), .IN3(n11752), .IN4(n11753), 
        .QN(WX676) );
  NAND2X0 U11831 ( .IN1(n9333), .IN2(n11754), .QN(n11753) );
  NAND2X0 U11832 ( .IN1(n9094), .IN2(n11755), .QN(n11752) );
  NAND2X0 U11833 ( .IN1(WX514), .IN2(n9279), .QN(n11751) );
  NAND2X0 U11834 ( .IN1(n9313), .IN2(CRC_OUT_9_15), .QN(n11750) );
  NAND4X0 U11835 ( .IN1(n11756), .IN2(n11757), .IN3(n11758), .IN4(n11759), 
        .QN(WX674) );
  NAND2X0 U11836 ( .IN1(n11760), .IN2(n11761), .QN(n11759) );
  NAND3X0 U11837 ( .IN1(n11762), .IN2(n11763), .IN3(n11764), .QN(n11760) );
  NAND2X0 U11838 ( .IN1(n9333), .IN2(n11765), .QN(n11764) );
  NAND2X0 U11839 ( .IN1(n10068), .IN2(n8653), .QN(n11763) );
  NAND2X0 U11840 ( .IN1(n16321), .IN2(n9080), .QN(n11762) );
  NAND2X0 U11841 ( .IN1(n11766), .IN2(n9110), .QN(n11758) );
  INVX0 U11842 ( .INP(n11767), .ZN(n11766) );
  NAND2X0 U11843 ( .IN1(WX512), .IN2(n9279), .QN(n11757) );
  NAND2X0 U11844 ( .IN1(n9312), .IN2(CRC_OUT_9_16), .QN(n11756) );
  NAND4X0 U11845 ( .IN1(n11768), .IN2(n11769), .IN3(n11770), .IN4(n11771), 
        .QN(WX672) );
  NAND2X0 U11846 ( .IN1(n11772), .IN2(n11773), .QN(n11771) );
  NAND3X0 U11847 ( .IN1(n11774), .IN2(n11775), .IN3(n11776), .QN(n11772) );
  NAND2X0 U11848 ( .IN1(n9334), .IN2(n11777), .QN(n11776) );
  NAND2X0 U11849 ( .IN1(n9084), .IN2(n8654), .QN(n11775) );
  NAND2X0 U11850 ( .IN1(n16320), .IN2(n9079), .QN(n11774) );
  NAND2X0 U11851 ( .IN1(n9094), .IN2(n11778), .QN(n11770) );
  NAND2X0 U11852 ( .IN1(WX510), .IN2(n9279), .QN(n11769) );
  NAND2X0 U11853 ( .IN1(n9313), .IN2(CRC_OUT_9_17), .QN(n11768) );
  NAND4X0 U11854 ( .IN1(n11779), .IN2(n11780), .IN3(n11781), .IN4(n11782), 
        .QN(WX670) );
  NAND2X0 U11855 ( .IN1(n11783), .IN2(n9336), .QN(n11782) );
  NAND2X0 U11856 ( .IN1(n9094), .IN2(n11784), .QN(n11781) );
  NAND2X0 U11857 ( .IN1(WX508), .IN2(n9279), .QN(n11780) );
  NAND2X0 U11858 ( .IN1(n9311), .IN2(CRC_OUT_9_18), .QN(n11779) );
  NAND4X0 U11859 ( .IN1(n11785), .IN2(n11786), .IN3(n11787), .IN4(n11788), 
        .QN(WX668) );
  NAND2X0 U11860 ( .IN1(n11789), .IN2(n11790), .QN(n11788) );
  NAND3X0 U11861 ( .IN1(n11791), .IN2(n11792), .IN3(n11793), .QN(n11789) );
  NAND2X0 U11862 ( .IN1(n9334), .IN2(n11794), .QN(n11793) );
  NAND2X0 U11863 ( .IN1(n9083), .IN2(n8656), .QN(n11792) );
  NAND2X0 U11864 ( .IN1(n16318), .IN2(n9078), .QN(n11791) );
  NAND2X0 U11865 ( .IN1(n9094), .IN2(n11795), .QN(n11787) );
  NAND2X0 U11866 ( .IN1(WX506), .IN2(n9279), .QN(n11786) );
  NAND2X0 U11867 ( .IN1(test_so10), .IN2(n9314), .QN(n11785) );
  NAND4X0 U11868 ( .IN1(n11796), .IN2(n11797), .IN3(n11798), .IN4(n11799), 
        .QN(WX666) );
  NAND2X0 U11869 ( .IN1(n11800), .IN2(n11801), .QN(n11799) );
  NAND3X0 U11870 ( .IN1(n11802), .IN2(n11803), .IN3(n11804), .QN(n11800) );
  NAND2X0 U11871 ( .IN1(n9334), .IN2(n11805), .QN(n11804) );
  NAND2X0 U11872 ( .IN1(n9082), .IN2(n8657), .QN(n11803) );
  NAND2X0 U11873 ( .IN1(n16317), .IN2(n10069), .QN(n11802) );
  NAND2X0 U11874 ( .IN1(n11806), .IN2(n9110), .QN(n11798) );
  INVX0 U11875 ( .INP(n11807), .ZN(n11806) );
  NAND2X0 U11876 ( .IN1(WX504), .IN2(n9279), .QN(n11797) );
  NAND2X0 U11877 ( .IN1(n9313), .IN2(CRC_OUT_9_20), .QN(n11796) );
  NAND4X0 U11878 ( .IN1(n11808), .IN2(n11809), .IN3(n11810), .IN4(n11811), 
        .QN(WX664) );
  NAND2X0 U11879 ( .IN1(n11812), .IN2(n11813), .QN(n11811) );
  NAND3X0 U11880 ( .IN1(n11814), .IN2(n11815), .IN3(n11816), .QN(n11812) );
  NAND2X0 U11881 ( .IN1(n9333), .IN2(n11817), .QN(n11816) );
  NAND2X0 U11882 ( .IN1(n10068), .IN2(n8658), .QN(n11815) );
  NAND2X0 U11883 ( .IN1(n16316), .IN2(n9080), .QN(n11814) );
  NAND2X0 U11884 ( .IN1(n9094), .IN2(n11818), .QN(n11810) );
  NAND2X0 U11885 ( .IN1(WX502), .IN2(n9279), .QN(n11809) );
  NAND2X0 U11886 ( .IN1(n9312), .IN2(CRC_OUT_9_21), .QN(n11808) );
  NAND4X0 U11887 ( .IN1(n11819), .IN2(n11820), .IN3(n11821), .IN4(n11822), 
        .QN(WX662) );
  NAND2X0 U11888 ( .IN1(n11823), .IN2(n11824), .QN(n11822) );
  NAND3X0 U11889 ( .IN1(n11825), .IN2(n11826), .IN3(n11827), .QN(n11823) );
  NAND2X0 U11890 ( .IN1(n9334), .IN2(n11828), .QN(n11827) );
  NAND2X0 U11891 ( .IN1(n9079), .IN2(WX2148), .QN(n11826) );
  NAND2X0 U11892 ( .IN1(n9084), .IN2(n8593), .QN(n11825) );
  NAND2X0 U11893 ( .IN1(n9094), .IN2(n11829), .QN(n11821) );
  NAND2X0 U11894 ( .IN1(WX500), .IN2(n9279), .QN(n11820) );
  NAND2X0 U11895 ( .IN1(n9313), .IN2(CRC_OUT_9_22), .QN(n11819) );
  NAND4X0 U11896 ( .IN1(n11830), .IN2(n11831), .IN3(n11832), .IN4(n11833), 
        .QN(WX660) );
  NAND2X0 U11897 ( .IN1(n11834), .IN2(n11835), .QN(n11833) );
  NAND3X0 U11898 ( .IN1(n11836), .IN2(n11837), .IN3(n11838), .QN(n11834) );
  NAND2X0 U11899 ( .IN1(n9334), .IN2(n11839), .QN(n11838) );
  NAND2X0 U11900 ( .IN1(n9083), .IN2(n8661), .QN(n11837) );
  NAND2X0 U11901 ( .IN1(n16315), .IN2(n9079), .QN(n11836) );
  NAND2X0 U11902 ( .IN1(n9094), .IN2(n11840), .QN(n11832) );
  NAND2X0 U11903 ( .IN1(WX498), .IN2(n9279), .QN(n11831) );
  NAND2X0 U11904 ( .IN1(n9311), .IN2(CRC_OUT_9_23), .QN(n11830) );
  NAND4X0 U11905 ( .IN1(n11841), .IN2(n11842), .IN3(n11843), .IN4(n11844), 
        .QN(WX658) );
  NAND2X0 U11906 ( .IN1(n11845), .IN2(n11846), .QN(n11844) );
  NAND3X0 U11907 ( .IN1(n11847), .IN2(n11848), .IN3(n11849), .QN(n11845) );
  NAND2X0 U11908 ( .IN1(n9334), .IN2(n11850), .QN(n11849) );
  NAND2X0 U11909 ( .IN1(n9082), .IN2(n8662), .QN(n11848) );
  NAND2X0 U11910 ( .IN1(n16314), .IN2(n9078), .QN(n11847) );
  NAND2X0 U11911 ( .IN1(n11851), .IN2(n9111), .QN(n11843) );
  INVX0 U11912 ( .INP(n11852), .ZN(n11851) );
  NAND2X0 U11913 ( .IN1(WX496), .IN2(n9279), .QN(n11842) );
  NAND2X0 U11914 ( .IN1(n9313), .IN2(CRC_OUT_9_24), .QN(n11841) );
  NAND4X0 U11915 ( .IN1(n11853), .IN2(n11854), .IN3(n11855), .IN4(n11856), 
        .QN(WX656) );
  NAND2X0 U11916 ( .IN1(n11857), .IN2(n11858), .QN(n11856) );
  NAND3X0 U11917 ( .IN1(n11859), .IN2(n11860), .IN3(n11861), .QN(n11857) );
  NAND2X0 U11918 ( .IN1(n9334), .IN2(n11862), .QN(n11861) );
  NAND2X0 U11919 ( .IN1(n10068), .IN2(n8663), .QN(n11860) );
  NAND2X0 U11920 ( .IN1(n16313), .IN2(n10069), .QN(n11859) );
  NAND2X0 U11921 ( .IN1(n9094), .IN2(n11863), .QN(n11855) );
  NAND2X0 U11922 ( .IN1(WX494), .IN2(n9280), .QN(n11854) );
  NAND2X0 U11923 ( .IN1(n9312), .IN2(CRC_OUT_9_25), .QN(n11853) );
  NAND4X0 U11924 ( .IN1(n11864), .IN2(n11865), .IN3(n11866), .IN4(n11867), 
        .QN(WX654) );
  NAND2X0 U11925 ( .IN1(n11868), .IN2(n11869), .QN(n11867) );
  NAND3X0 U11926 ( .IN1(n11870), .IN2(n11871), .IN3(n11872), .QN(n11868) );
  NAND2X0 U11927 ( .IN1(n9334), .IN2(n11873), .QN(n11872) );
  NAND2X0 U11928 ( .IN1(n9084), .IN2(n8664), .QN(n11871) );
  NAND2X0 U11929 ( .IN1(n16312), .IN2(n9080), .QN(n11870) );
  NAND2X0 U11930 ( .IN1(n9095), .IN2(n11874), .QN(n11866) );
  NAND2X0 U11931 ( .IN1(WX492), .IN2(n9280), .QN(n11865) );
  NAND2X0 U11932 ( .IN1(n9313), .IN2(CRC_OUT_9_26), .QN(n11864) );
  NAND4X0 U11933 ( .IN1(n11875), .IN2(n11876), .IN3(n11877), .IN4(n11878), 
        .QN(WX652) );
  NAND2X0 U11934 ( .IN1(n11879), .IN2(n11880), .QN(n11878) );
  NAND3X0 U11935 ( .IN1(n11881), .IN2(n11882), .IN3(n11883), .QN(n11879) );
  NAND2X0 U11936 ( .IN1(n9334), .IN2(n11884), .QN(n11883) );
  NAND2X0 U11937 ( .IN1(n9083), .IN2(n8665), .QN(n11882) );
  NAND2X0 U11938 ( .IN1(n16311), .IN2(n9079), .QN(n11881) );
  NAND2X0 U11939 ( .IN1(n9095), .IN2(n11885), .QN(n11877) );
  NAND2X0 U11940 ( .IN1(WX490), .IN2(n9280), .QN(n11876) );
  NAND2X0 U11941 ( .IN1(n9312), .IN2(CRC_OUT_9_27), .QN(n11875) );
  NAND4X0 U11942 ( .IN1(n11886), .IN2(n11887), .IN3(n11888), .IN4(n11889), 
        .QN(WX650) );
  NAND2X0 U11943 ( .IN1(n11890), .IN2(n9336), .QN(n11889) );
  NAND2X0 U11944 ( .IN1(n11891), .IN2(n9110), .QN(n11888) );
  INVX0 U11945 ( .INP(n11892), .ZN(n11891) );
  NAND2X0 U11946 ( .IN1(WX488), .IN2(n9280), .QN(n11887) );
  NAND2X0 U11947 ( .IN1(n9312), .IN2(CRC_OUT_9_28), .QN(n11886) );
  NOR3X0 U11948 ( .IN1(n9143), .IN2(n11893), .IN3(n11894), .QN(WX6498) );
  NOR2X0 U11949 ( .IN1(n8239), .IN2(CRC_OUT_5_30), .QN(n11894) );
  NOR2X0 U11950 ( .IN1(DFF_958_n1), .IN2(WX6009), .QN(n11893) );
  NOR3X0 U11951 ( .IN1(n9143), .IN2(n11895), .IN3(n11896), .QN(WX6496) );
  NOR2X0 U11952 ( .IN1(n8240), .IN2(CRC_OUT_5_29), .QN(n11896) );
  NOR2X0 U11953 ( .IN1(DFF_957_n1), .IN2(WX6011), .QN(n11895) );
  NOR3X0 U11954 ( .IN1(n9142), .IN2(n11897), .IN3(n11898), .QN(WX6494) );
  NOR2X0 U11955 ( .IN1(n8241), .IN2(CRC_OUT_5_28), .QN(n11898) );
  NOR2X0 U11956 ( .IN1(DFF_956_n1), .IN2(WX6013), .QN(n11897) );
  NOR3X0 U11957 ( .IN1(n9142), .IN2(n11899), .IN3(n11900), .QN(WX6492) );
  NOR2X0 U11958 ( .IN1(n8242), .IN2(CRC_OUT_5_27), .QN(n11900) );
  NOR2X0 U11959 ( .IN1(DFF_955_n1), .IN2(WX6015), .QN(n11899) );
  NOR3X0 U11960 ( .IN1(n9142), .IN2(n11901), .IN3(n11902), .QN(WX6490) );
  NOR2X0 U11961 ( .IN1(n8243), .IN2(CRC_OUT_5_26), .QN(n11902) );
  NOR2X0 U11962 ( .IN1(DFF_954_n1), .IN2(WX6017), .QN(n11901) );
  NOR3X0 U11963 ( .IN1(n9142), .IN2(n11903), .IN3(n11904), .QN(WX6488) );
  NOR2X0 U11964 ( .IN1(n8244), .IN2(CRC_OUT_5_25), .QN(n11904) );
  NOR2X0 U11965 ( .IN1(DFF_953_n1), .IN2(WX6019), .QN(n11903) );
  NOR3X0 U11966 ( .IN1(n9142), .IN2(n11905), .IN3(n11906), .QN(WX6486) );
  NOR2X0 U11967 ( .IN1(n8245), .IN2(CRC_OUT_5_24), .QN(n11906) );
  NOR2X0 U11968 ( .IN1(DFF_952_n1), .IN2(WX6021), .QN(n11905) );
  NOR3X0 U11969 ( .IN1(n10681), .IN2(n11907), .IN3(n11908), .QN(WX6484) );
  NOR2X0 U11970 ( .IN1(n8255), .IN2(CRC_OUT_5_23), .QN(n11908) );
  NOR2X0 U11971 ( .IN1(DFF_951_n1), .IN2(WX6023), .QN(n11907) );
  NAND2X0 U11972 ( .IN1(RESET), .IN2(n11909), .QN(n10681) );
  INVX0 U11973 ( .INP(Tj_Trigger), .ZN(n11909) );
  NOR3X0 U11974 ( .IN1(n9142), .IN2(n11910), .IN3(n11911), .QN(WX6482) );
  NOR2X0 U11975 ( .IN1(n8256), .IN2(CRC_OUT_5_22), .QN(n11911) );
  NOR2X0 U11976 ( .IN1(DFF_950_n1), .IN2(WX6025), .QN(n11910) );
  NOR3X0 U11977 ( .IN1(n9142), .IN2(n11912), .IN3(n11913), .QN(WX6480) );
  NOR2X0 U11978 ( .IN1(n8273), .IN2(CRC_OUT_5_21), .QN(n11913) );
  NOR2X0 U11979 ( .IN1(DFF_949_n1), .IN2(WX6027), .QN(n11912) );
  NAND4X0 U11980 ( .IN1(n11914), .IN2(n11915), .IN3(n11916), .IN4(n11917), 
        .QN(WX648) );
  NAND2X0 U11981 ( .IN1(n11918), .IN2(n11919), .QN(n11917) );
  NAND3X0 U11982 ( .IN1(n11920), .IN2(n11921), .IN3(n11922), .QN(n11918) );
  NAND2X0 U11983 ( .IN1(n9334), .IN2(n11923), .QN(n11922) );
  NAND2X0 U11984 ( .IN1(n9082), .IN2(n8667), .QN(n11921) );
  NAND2X0 U11985 ( .IN1(n16309), .IN2(n9078), .QN(n11920) );
  NAND2X0 U11986 ( .IN1(n9095), .IN2(n11924), .QN(n11916) );
  NAND2X0 U11987 ( .IN1(WX486), .IN2(n9280), .QN(n11915) );
  NAND2X0 U11988 ( .IN1(n9313), .IN2(CRC_OUT_9_29), .QN(n11914) );
  NOR3X0 U11989 ( .IN1(n9142), .IN2(n11925), .IN3(n11926), .QN(WX6478) );
  NOR2X0 U11990 ( .IN1(n8274), .IN2(CRC_OUT_5_20), .QN(n11926) );
  NOR2X0 U11991 ( .IN1(DFF_948_n1), .IN2(WX6029), .QN(n11925) );
  NOR3X0 U11992 ( .IN1(n9142), .IN2(n11927), .IN3(n11928), .QN(WX6476) );
  NOR2X0 U11993 ( .IN1(n8291), .IN2(CRC_OUT_5_19), .QN(n11928) );
  NOR2X0 U11994 ( .IN1(DFF_947_n1), .IN2(WX6031), .QN(n11927) );
  NOR3X0 U11995 ( .IN1(n9142), .IN2(n11929), .IN3(n11930), .QN(WX6474) );
  NOR2X0 U11996 ( .IN1(n8292), .IN2(CRC_OUT_5_18), .QN(n11930) );
  NOR2X0 U11997 ( .IN1(DFF_946_n1), .IN2(WX6033), .QN(n11929) );
  NOR2X0 U11998 ( .IN1(n9226), .IN2(n11931), .QN(WX6472) );
  NOR2X0 U11999 ( .IN1(n11932), .IN2(n11933), .QN(n11931) );
  NOR2X0 U12000 ( .IN1(test_so54), .IN2(WX6035), .QN(n11933) );
  NOR2X0 U12001 ( .IN1(n8296), .IN2(n8828), .QN(n11932) );
  NOR3X0 U12002 ( .IN1(n9142), .IN2(n11934), .IN3(n11935), .QN(WX6470) );
  NOR2X0 U12003 ( .IN1(n8297), .IN2(CRC_OUT_5_16), .QN(n11935) );
  NOR2X0 U12004 ( .IN1(DFF_944_n1), .IN2(WX6037), .QN(n11934) );
  NOR3X0 U12005 ( .IN1(n9142), .IN2(n11936), .IN3(n11937), .QN(WX6468) );
  INVX0 U12006 ( .INP(n11938), .ZN(n11937) );
  NAND2X0 U12007 ( .IN1(CRC_OUT_5_15), .IN2(n11939), .QN(n11938) );
  NOR2X0 U12008 ( .IN1(n11939), .IN2(CRC_OUT_5_15), .QN(n11936) );
  NAND2X0 U12009 ( .IN1(n11940), .IN2(n11941), .QN(n11939) );
  NAND2X0 U12010 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .QN(n11941) );
  NAND2X0 U12011 ( .IN1(DFF_959_n1), .IN2(n8827), .QN(n11940) );
  NOR3X0 U12012 ( .IN1(n9141), .IN2(n11942), .IN3(n11943), .QN(WX6466) );
  NOR2X0 U12013 ( .IN1(n8298), .IN2(CRC_OUT_5_14), .QN(n11943) );
  NOR2X0 U12014 ( .IN1(DFF_942_n1), .IN2(WX6041), .QN(n11942) );
  NOR3X0 U12015 ( .IN1(n9141), .IN2(n11944), .IN3(n11945), .QN(WX6464) );
  NOR2X0 U12016 ( .IN1(n8299), .IN2(CRC_OUT_5_13), .QN(n11945) );
  NOR2X0 U12017 ( .IN1(DFF_941_n1), .IN2(WX6043), .QN(n11944) );
  NOR3X0 U12018 ( .IN1(n9141), .IN2(n11946), .IN3(n11947), .QN(WX6462) );
  NOR2X0 U12019 ( .IN1(n8300), .IN2(CRC_OUT_5_12), .QN(n11947) );
  NOR2X0 U12020 ( .IN1(DFF_940_n1), .IN2(WX6045), .QN(n11946) );
  NOR3X0 U12021 ( .IN1(n9141), .IN2(n11948), .IN3(n11949), .QN(WX6460) );
  NOR2X0 U12022 ( .IN1(n8301), .IN2(CRC_OUT_5_11), .QN(n11949) );
  NOR2X0 U12023 ( .IN1(DFF_939_n1), .IN2(WX6047), .QN(n11948) );
  NAND4X0 U12024 ( .IN1(n11950), .IN2(n11951), .IN3(n11952), .IN4(n11953), 
        .QN(WX646) );
  NAND2X0 U12025 ( .IN1(n11954), .IN2(n11955), .QN(n11953) );
  NAND3X0 U12026 ( .IN1(n11956), .IN2(n11957), .IN3(n11958), .QN(n11954) );
  NAND2X0 U12027 ( .IN1(n9334), .IN2(n11959), .QN(n11958) );
  NAND2X0 U12028 ( .IN1(n10068), .IN2(n8668), .QN(n11957) );
  NAND2X0 U12029 ( .IN1(n16308), .IN2(n10069), .QN(n11956) );
  NAND2X0 U12030 ( .IN1(n9095), .IN2(n11960), .QN(n11952) );
  NAND2X0 U12031 ( .IN1(WX484), .IN2(n9280), .QN(n11951) );
  NAND2X0 U12032 ( .IN1(n9314), .IN2(CRC_OUT_9_30), .QN(n11950) );
  NOR2X0 U12033 ( .IN1(n9241), .IN2(n11961), .QN(WX6458) );
  NOR2X0 U12034 ( .IN1(n11962), .IN2(n11963), .QN(n11961) );
  INVX0 U12035 ( .INP(n11964), .ZN(n11963) );
  NAND2X0 U12036 ( .IN1(CRC_OUT_5_10), .IN2(n11965), .QN(n11964) );
  NOR2X0 U12037 ( .IN1(n11965), .IN2(CRC_OUT_5_10), .QN(n11962) );
  NAND2X0 U12038 ( .IN1(n11966), .IN2(n11967), .QN(n11965) );
  NAND2X0 U12039 ( .IN1(n8116), .IN2(CRC_OUT_5_31), .QN(n11967) );
  NAND2X0 U12040 ( .IN1(DFF_959_n1), .IN2(WX6049), .QN(n11966) );
  NOR3X0 U12041 ( .IN1(n9141), .IN2(n11968), .IN3(n11969), .QN(WX6456) );
  NOR2X0 U12042 ( .IN1(n8302), .IN2(CRC_OUT_5_9), .QN(n11969) );
  NOR2X0 U12043 ( .IN1(DFF_937_n1), .IN2(WX6051), .QN(n11968) );
  NOR3X0 U12044 ( .IN1(n9141), .IN2(n11970), .IN3(n11971), .QN(WX6454) );
  NOR2X0 U12045 ( .IN1(n8303), .IN2(CRC_OUT_5_8), .QN(n11971) );
  NOR2X0 U12046 ( .IN1(DFF_936_n1), .IN2(WX6053), .QN(n11970) );
  NOR3X0 U12047 ( .IN1(n9141), .IN2(n11972), .IN3(n11973), .QN(WX6452) );
  NOR2X0 U12048 ( .IN1(n8308), .IN2(CRC_OUT_5_7), .QN(n11973) );
  NOR2X0 U12049 ( .IN1(DFF_935_n1), .IN2(WX6055), .QN(n11972) );
  NOR3X0 U12050 ( .IN1(n9141), .IN2(n11974), .IN3(n11975), .QN(WX6450) );
  NOR2X0 U12051 ( .IN1(n8309), .IN2(CRC_OUT_5_6), .QN(n11975) );
  NOR2X0 U12052 ( .IN1(DFF_934_n1), .IN2(WX6057), .QN(n11974) );
  NOR3X0 U12053 ( .IN1(n9141), .IN2(n11976), .IN3(n11977), .QN(WX6448) );
  NOR2X0 U12054 ( .IN1(n8326), .IN2(CRC_OUT_5_5), .QN(n11977) );
  NOR2X0 U12055 ( .IN1(DFF_933_n1), .IN2(WX6059), .QN(n11976) );
  NOR3X0 U12056 ( .IN1(n9141), .IN2(n11978), .IN3(n11979), .QN(WX6446) );
  NOR2X0 U12057 ( .IN1(n8327), .IN2(CRC_OUT_5_4), .QN(n11979) );
  NOR2X0 U12058 ( .IN1(DFF_932_n1), .IN2(WX6061), .QN(n11978) );
  NOR2X0 U12059 ( .IN1(n9241), .IN2(n11980), .QN(WX6444) );
  NOR2X0 U12060 ( .IN1(n11981), .IN2(n11982), .QN(n11980) );
  INVX0 U12061 ( .INP(n11983), .ZN(n11982) );
  NAND2X0 U12062 ( .IN1(CRC_OUT_5_3), .IN2(n11984), .QN(n11983) );
  NOR2X0 U12063 ( .IN1(n11984), .IN2(CRC_OUT_5_3), .QN(n11981) );
  NAND2X0 U12064 ( .IN1(n11985), .IN2(n11986), .QN(n11984) );
  NAND2X0 U12065 ( .IN1(n8117), .IN2(CRC_OUT_5_31), .QN(n11986) );
  NAND2X0 U12066 ( .IN1(DFF_959_n1), .IN2(WX6063), .QN(n11985) );
  NOR3X0 U12067 ( .IN1(n9141), .IN2(n11987), .IN3(n11988), .QN(WX6442) );
  NOR2X0 U12068 ( .IN1(n8344), .IN2(CRC_OUT_5_2), .QN(n11988) );
  NOR2X0 U12069 ( .IN1(DFF_930_n1), .IN2(WX6065), .QN(n11987) );
  NOR3X0 U12070 ( .IN1(n9140), .IN2(n11989), .IN3(n11990), .QN(WX6440) );
  NOR2X0 U12071 ( .IN1(n8345), .IN2(CRC_OUT_5_1), .QN(n11990) );
  NOR2X0 U12072 ( .IN1(DFF_929_n1), .IN2(WX6067), .QN(n11989) );
  NAND4X0 U12073 ( .IN1(n11991), .IN2(n11992), .IN3(n11993), .IN4(n11994), 
        .QN(WX644) );
  NAND2X0 U12074 ( .IN1(n11995), .IN2(n11996), .QN(n11994) );
  NAND3X0 U12075 ( .IN1(n11997), .IN2(n11998), .IN3(n11999), .QN(n11995) );
  NAND2X0 U12076 ( .IN1(n9334), .IN2(n12000), .QN(n11999) );
  NAND2X0 U12077 ( .IN1(n9084), .IN2(n8669), .QN(n11998) );
  NAND2X0 U12078 ( .IN1(n16307), .IN2(n9080), .QN(n11997) );
  NAND2X0 U12079 ( .IN1(n9095), .IN2(n12001), .QN(n11993) );
  NAND2X0 U12080 ( .IN1(n9313), .IN2(CRC_OUT_9_31), .QN(n11992) );
  NAND2X0 U12081 ( .IN1(n2245), .IN2(WX485), .QN(n11991) );
  NOR2X0 U12082 ( .IN1(n9241), .IN2(n12002), .QN(WX6438) );
  NOR2X0 U12083 ( .IN1(n12003), .IN2(n12004), .QN(n12002) );
  NOR2X0 U12084 ( .IN1(test_so53), .IN2(WX6069), .QN(n12004) );
  INVX0 U12085 ( .INP(n12005), .ZN(n12003) );
  NAND2X0 U12086 ( .IN1(WX6069), .IN2(test_so53), .QN(n12005) );
  NOR3X0 U12087 ( .IN1(n9140), .IN2(n12006), .IN3(n12007), .QN(WX6436) );
  NOR2X0 U12088 ( .IN1(n8130), .IN2(CRC_OUT_5_31), .QN(n12007) );
  NOR2X0 U12089 ( .IN1(DFF_959_n1), .IN2(WX6071), .QN(n12006) );
  NOR2X0 U12090 ( .IN1(n16366), .IN2(n9163), .QN(WX5910) );
  NOR2X0 U12091 ( .IN1(n16365), .IN2(n9162), .QN(WX5908) );
  NOR2X0 U12092 ( .IN1(n16364), .IN2(n9163), .QN(WX5906) );
  NOR2X0 U12093 ( .IN1(n16363), .IN2(n9163), .QN(WX5904) );
  NOR2X0 U12094 ( .IN1(n16362), .IN2(n9163), .QN(WX5902) );
  NOR2X0 U12095 ( .IN1(n16361), .IN2(n9163), .QN(WX5900) );
  NOR2X0 U12096 ( .IN1(n9240), .IN2(n8822), .QN(WX5898) );
  NOR2X0 U12097 ( .IN1(n16360), .IN2(n9163), .QN(WX5896) );
  NOR2X0 U12098 ( .IN1(n16359), .IN2(n9163), .QN(WX5894) );
  NOR2X0 U12099 ( .IN1(n16358), .IN2(n9163), .QN(WX5892) );
  NOR2X0 U12100 ( .IN1(n16357), .IN2(n9163), .QN(WX5890) );
  NOR2X0 U12101 ( .IN1(n16356), .IN2(n9163), .QN(WX5888) );
  NOR2X0 U12102 ( .IN1(n16355), .IN2(n9163), .QN(WX5886) );
  NOR2X0 U12103 ( .IN1(n16354), .IN2(n9163), .QN(WX5884) );
  NOR2X0 U12104 ( .IN1(n16353), .IN2(n9163), .QN(WX5882) );
  NOR2X0 U12105 ( .IN1(n16352), .IN2(n9163), .QN(WX5880) );
  NAND4X0 U12106 ( .IN1(n12008), .IN2(n12009), .IN3(n12010), .IN4(n12011), 
        .QN(WX5878) );
  NAND2X0 U12107 ( .IN1(n9334), .IN2(n11063), .QN(n12011) );
  NAND2X0 U12108 ( .IN1(n12012), .IN2(n12013), .QN(n11063) );
  INVX0 U12109 ( .INP(n12014), .ZN(n12013) );
  NOR2X0 U12110 ( .IN1(n12015), .IN2(n12016), .QN(n12014) );
  NAND2X0 U12111 ( .IN1(n12016), .IN2(n12015), .QN(n12012) );
  NOR2X0 U12112 ( .IN1(n12017), .IN2(n12018), .QN(n12015) );
  NOR2X0 U12113 ( .IN1(WX7364), .IN2(n7946), .QN(n12018) );
  INVX0 U12114 ( .INP(n12019), .ZN(n12017) );
  NAND2X0 U12115 ( .IN1(n7946), .IN2(WX7364), .QN(n12019) );
  NAND2X0 U12116 ( .IN1(n12020), .IN2(n12021), .QN(n12016) );
  NAND2X0 U12117 ( .IN1(n7945), .IN2(WX7236), .QN(n12021) );
  INVX0 U12118 ( .INP(n12022), .ZN(n12020) );
  NOR2X0 U12119 ( .IN1(WX7236), .IN2(n7945), .QN(n12022) );
  NAND2X0 U12120 ( .IN1(n9095), .IN2(n12023), .QN(n12010) );
  NAND2X0 U12121 ( .IN1(n1006), .IN2(n9280), .QN(n12009) );
  NOR2X0 U12122 ( .IN1(n9240), .IN2(n8916), .QN(n1006) );
  NAND2X0 U12123 ( .IN1(test_so53), .IN2(n9315), .QN(n12008) );
  NAND4X0 U12124 ( .IN1(n12024), .IN2(n12025), .IN3(n12026), .IN4(n12027), 
        .QN(WX5876) );
  NAND3X0 U12125 ( .IN1(n12028), .IN2(n12029), .IN3(n9090), .QN(n12027) );
  NAND2X0 U12126 ( .IN1(n9334), .IN2(n11079), .QN(n12026) );
  NAND2X0 U12127 ( .IN1(n12030), .IN2(n12031), .QN(n11079) );
  INVX0 U12128 ( .INP(n12032), .ZN(n12031) );
  NOR2X0 U12129 ( .IN1(n12033), .IN2(n12034), .QN(n12032) );
  NAND2X0 U12130 ( .IN1(n12034), .IN2(n12033), .QN(n12030) );
  NOR2X0 U12131 ( .IN1(n12035), .IN2(n12036), .QN(n12033) );
  NOR2X0 U12132 ( .IN1(WX7362), .IN2(n7948), .QN(n12036) );
  INVX0 U12133 ( .INP(n12037), .ZN(n12035) );
  NAND2X0 U12134 ( .IN1(n7948), .IN2(WX7362), .QN(n12037) );
  NAND2X0 U12135 ( .IN1(n12038), .IN2(n12039), .QN(n12034) );
  NAND2X0 U12136 ( .IN1(n7947), .IN2(WX7234), .QN(n12039) );
  INVX0 U12137 ( .INP(n12040), .ZN(n12038) );
  NOR2X0 U12138 ( .IN1(WX7234), .IN2(n7947), .QN(n12040) );
  NAND2X0 U12139 ( .IN1(n1005), .IN2(n9280), .QN(n12025) );
  NOR2X0 U12140 ( .IN1(n9240), .IN2(n8917), .QN(n1005) );
  NAND2X0 U12141 ( .IN1(n9312), .IN2(CRC_OUT_5_1), .QN(n12024) );
  NAND4X0 U12142 ( .IN1(n12041), .IN2(n12042), .IN3(n12043), .IN4(n12044), 
        .QN(WX5874) );
  NAND2X0 U12143 ( .IN1(n9325), .IN2(n11095), .QN(n12044) );
  NAND2X0 U12144 ( .IN1(n12045), .IN2(n12046), .QN(n11095) );
  INVX0 U12145 ( .INP(n12047), .ZN(n12046) );
  NOR2X0 U12146 ( .IN1(n12048), .IN2(n12049), .QN(n12047) );
  NAND2X0 U12147 ( .IN1(n12049), .IN2(n12048), .QN(n12045) );
  NOR2X0 U12148 ( .IN1(n12050), .IN2(n12051), .QN(n12048) );
  NOR2X0 U12149 ( .IN1(WX7360), .IN2(n7950), .QN(n12051) );
  INVX0 U12150 ( .INP(n12052), .ZN(n12050) );
  NAND2X0 U12151 ( .IN1(n7950), .IN2(WX7360), .QN(n12052) );
  NAND2X0 U12152 ( .IN1(n12053), .IN2(n12054), .QN(n12049) );
  NAND2X0 U12153 ( .IN1(n7949), .IN2(WX7232), .QN(n12054) );
  INVX0 U12154 ( .INP(n12055), .ZN(n12053) );
  NOR2X0 U12155 ( .IN1(WX7232), .IN2(n7949), .QN(n12055) );
  NAND2X0 U12156 ( .IN1(n9095), .IN2(n12056), .QN(n12043) );
  NAND2X0 U12157 ( .IN1(n1004), .IN2(n9280), .QN(n12042) );
  NOR2X0 U12158 ( .IN1(n9240), .IN2(n8918), .QN(n1004) );
  NAND2X0 U12159 ( .IN1(n9314), .IN2(CRC_OUT_5_2), .QN(n12041) );
  NAND4X0 U12160 ( .IN1(n12057), .IN2(n12058), .IN3(n12059), .IN4(n12060), 
        .QN(WX5872) );
  NAND3X0 U12161 ( .IN1(n12061), .IN2(n12062), .IN3(n9091), .QN(n12060) );
  NAND2X0 U12162 ( .IN1(n9323), .IN2(n11111), .QN(n12059) );
  NAND2X0 U12163 ( .IN1(n12063), .IN2(n12064), .QN(n11111) );
  INVX0 U12164 ( .INP(n12065), .ZN(n12064) );
  NOR2X0 U12165 ( .IN1(n12066), .IN2(n12067), .QN(n12065) );
  NAND2X0 U12166 ( .IN1(n12067), .IN2(n12066), .QN(n12063) );
  NOR2X0 U12167 ( .IN1(n12068), .IN2(n12069), .QN(n12066) );
  NOR2X0 U12168 ( .IN1(WX7358), .IN2(n7952), .QN(n12069) );
  INVX0 U12169 ( .INP(n12070), .ZN(n12068) );
  NAND2X0 U12170 ( .IN1(n7952), .IN2(WX7358), .QN(n12070) );
  NAND2X0 U12171 ( .IN1(n12071), .IN2(n12072), .QN(n12067) );
  NAND2X0 U12172 ( .IN1(n7951), .IN2(WX7230), .QN(n12072) );
  INVX0 U12173 ( .INP(n12073), .ZN(n12071) );
  NOR2X0 U12174 ( .IN1(WX7230), .IN2(n7951), .QN(n12073) );
  NAND2X0 U12175 ( .IN1(n1003), .IN2(n9280), .QN(n12058) );
  NOR2X0 U12176 ( .IN1(n9239), .IN2(n8919), .QN(n1003) );
  NAND2X0 U12177 ( .IN1(n9313), .IN2(CRC_OUT_5_3), .QN(n12057) );
  NAND4X0 U12178 ( .IN1(n12074), .IN2(n12075), .IN3(n12076), .IN4(n12077), 
        .QN(WX5870) );
  NAND3X0 U12179 ( .IN1(n11116), .IN2(n11117), .IN3(n9321), .QN(n12077) );
  NAND3X0 U12180 ( .IN1(n12078), .IN2(n12079), .IN3(n12080), .QN(n11117) );
  INVX0 U12181 ( .INP(n12081), .ZN(n12080) );
  NAND2X0 U12182 ( .IN1(n12081), .IN2(n12082), .QN(n11116) );
  NAND2X0 U12183 ( .IN1(n12078), .IN2(n12079), .QN(n12082) );
  NAND2X0 U12184 ( .IN1(n7954), .IN2(WX7228), .QN(n12079) );
  NAND2X0 U12185 ( .IN1(n3635), .IN2(WX7292), .QN(n12078) );
  NOR2X0 U12186 ( .IN1(n12083), .IN2(n12084), .QN(n12081) );
  NOR2X0 U12187 ( .IN1(n8796), .IN2(n7953), .QN(n12084) );
  INVX0 U12188 ( .INP(n12085), .ZN(n12083) );
  NAND2X0 U12189 ( .IN1(n7953), .IN2(n8796), .QN(n12085) );
  NAND2X0 U12190 ( .IN1(n9095), .IN2(n12086), .QN(n12076) );
  NAND2X0 U12191 ( .IN1(n1002), .IN2(n9280), .QN(n12075) );
  NOR2X0 U12192 ( .IN1(n9239), .IN2(n8920), .QN(n1002) );
  NAND2X0 U12193 ( .IN1(n9314), .IN2(CRC_OUT_5_4), .QN(n12074) );
  NAND4X0 U12194 ( .IN1(n12087), .IN2(n12088), .IN3(n12089), .IN4(n12090), 
        .QN(WX5868) );
  NAND3X0 U12195 ( .IN1(n12091), .IN2(n12092), .IN3(n9091), .QN(n12090) );
  NAND2X0 U12196 ( .IN1(n9324), .IN2(n11144), .QN(n12089) );
  NAND2X0 U12197 ( .IN1(n12093), .IN2(n12094), .QN(n11144) );
  INVX0 U12198 ( .INP(n12095), .ZN(n12094) );
  NOR2X0 U12199 ( .IN1(n12096), .IN2(n12097), .QN(n12095) );
  NAND2X0 U12200 ( .IN1(n12097), .IN2(n12096), .QN(n12093) );
  NOR2X0 U12201 ( .IN1(n12098), .IN2(n12099), .QN(n12096) );
  NOR2X0 U12202 ( .IN1(WX7354), .IN2(n7956), .QN(n12099) );
  INVX0 U12203 ( .INP(n12100), .ZN(n12098) );
  NAND2X0 U12204 ( .IN1(n7956), .IN2(WX7354), .QN(n12100) );
  NAND2X0 U12205 ( .IN1(n12101), .IN2(n12102), .QN(n12097) );
  NAND2X0 U12206 ( .IN1(n7955), .IN2(WX7226), .QN(n12102) );
  INVX0 U12207 ( .INP(n12103), .ZN(n12101) );
  NOR2X0 U12208 ( .IN1(WX7226), .IN2(n7955), .QN(n12103) );
  NAND2X0 U12209 ( .IN1(n1001), .IN2(n9280), .QN(n12088) );
  NOR2X0 U12210 ( .IN1(n9239), .IN2(n8921), .QN(n1001) );
  NAND2X0 U12211 ( .IN1(n9313), .IN2(CRC_OUT_5_5), .QN(n12087) );
  NAND4X0 U12212 ( .IN1(n12104), .IN2(n12105), .IN3(n12106), .IN4(n12107), 
        .QN(WX5866) );
  NAND3X0 U12213 ( .IN1(n11149), .IN2(n11150), .IN3(n9321), .QN(n12107) );
  NAND3X0 U12214 ( .IN1(n12108), .IN2(n12109), .IN3(n12110), .QN(n11150) );
  INVX0 U12215 ( .INP(n12111), .ZN(n12110) );
  NAND2X0 U12216 ( .IN1(n12111), .IN2(n12112), .QN(n11149) );
  NAND2X0 U12217 ( .IN1(n12108), .IN2(n12109), .QN(n12112) );
  NAND2X0 U12218 ( .IN1(n8234), .IN2(WX7224), .QN(n12109) );
  NAND2X0 U12219 ( .IN1(n3639), .IN2(WX7352), .QN(n12108) );
  NOR2X0 U12220 ( .IN1(n12113), .IN2(n12114), .QN(n12111) );
  INVX0 U12221 ( .INP(n12115), .ZN(n12114) );
  NAND2X0 U12222 ( .IN1(test_so62), .IN2(WX7160), .QN(n12115) );
  NOR2X0 U12223 ( .IN1(WX7160), .IN2(test_so62), .QN(n12113) );
  NAND2X0 U12224 ( .IN1(n9095), .IN2(n12116), .QN(n12106) );
  NAND2X0 U12225 ( .IN1(n1000), .IN2(n9280), .QN(n12105) );
  NOR2X0 U12226 ( .IN1(n9239), .IN2(n8922), .QN(n1000) );
  NAND2X0 U12227 ( .IN1(n9314), .IN2(CRC_OUT_5_6), .QN(n12104) );
  NAND4X0 U12228 ( .IN1(n12117), .IN2(n12118), .IN3(n12119), .IN4(n12120), 
        .QN(WX5864) );
  NAND2X0 U12229 ( .IN1(n9323), .IN2(n11177), .QN(n12120) );
  NAND2X0 U12230 ( .IN1(n12121), .IN2(n12122), .QN(n11177) );
  INVX0 U12231 ( .INP(n12123), .ZN(n12122) );
  NOR2X0 U12232 ( .IN1(n12124), .IN2(n12125), .QN(n12123) );
  NAND2X0 U12233 ( .IN1(n12125), .IN2(n12124), .QN(n12121) );
  NOR2X0 U12234 ( .IN1(n12126), .IN2(n12127), .QN(n12124) );
  NOR2X0 U12235 ( .IN1(WX7350), .IN2(n7959), .QN(n12127) );
  INVX0 U12236 ( .INP(n12128), .ZN(n12126) );
  NAND2X0 U12237 ( .IN1(n7959), .IN2(WX7350), .QN(n12128) );
  NAND2X0 U12238 ( .IN1(n12129), .IN2(n12130), .QN(n12125) );
  NAND2X0 U12239 ( .IN1(n7958), .IN2(WX7222), .QN(n12130) );
  INVX0 U12240 ( .INP(n12131), .ZN(n12129) );
  NOR2X0 U12241 ( .IN1(WX7222), .IN2(n7958), .QN(n12131) );
  NAND2X0 U12242 ( .IN1(n9095), .IN2(n12132), .QN(n12119) );
  NAND2X0 U12243 ( .IN1(n999), .IN2(n9280), .QN(n12118) );
  NOR2X0 U12244 ( .IN1(n9067), .IN2(n9162), .QN(n999) );
  NAND2X0 U12245 ( .IN1(n9314), .IN2(CRC_OUT_5_7), .QN(n12117) );
  NAND4X0 U12246 ( .IN1(n12133), .IN2(n12134), .IN3(n12135), .IN4(n12136), 
        .QN(WX5862) );
  NAND3X0 U12247 ( .IN1(n11182), .IN2(n11183), .IN3(n9321), .QN(n12136) );
  NAND3X0 U12248 ( .IN1(n12137), .IN2(n12138), .IN3(n12139), .QN(n11183) );
  INVX0 U12249 ( .INP(n12140), .ZN(n12139) );
  NAND2X0 U12250 ( .IN1(n12140), .IN2(n12141), .QN(n11182) );
  NAND2X0 U12251 ( .IN1(n12137), .IN2(n12138), .QN(n12141) );
  NAND2X0 U12252 ( .IN1(n8232), .IN2(WX7284), .QN(n12138) );
  NAND2X0 U12253 ( .IN1(n7961), .IN2(WX7348), .QN(n12137) );
  NOR2X0 U12254 ( .IN1(n12142), .IN2(n12143), .QN(n12140) );
  INVX0 U12255 ( .INP(n12144), .ZN(n12143) );
  NAND2X0 U12256 ( .IN1(test_so60), .IN2(WX7156), .QN(n12144) );
  NOR2X0 U12257 ( .IN1(WX7156), .IN2(test_so60), .QN(n12142) );
  NAND2X0 U12258 ( .IN1(n9095), .IN2(n12145), .QN(n12135) );
  NAND2X0 U12259 ( .IN1(n998), .IN2(n9280), .QN(n12134) );
  NOR2X0 U12260 ( .IN1(n9239), .IN2(n8923), .QN(n998) );
  NAND2X0 U12261 ( .IN1(n9313), .IN2(CRC_OUT_5_8), .QN(n12133) );
  NAND4X0 U12262 ( .IN1(n12146), .IN2(n12147), .IN3(n12148), .IN4(n12149), 
        .QN(WX5860) );
  NAND2X0 U12263 ( .IN1(n9324), .IN2(n11207), .QN(n12149) );
  NAND2X0 U12264 ( .IN1(n12150), .IN2(n12151), .QN(n11207) );
  INVX0 U12265 ( .INP(n12152), .ZN(n12151) );
  NOR2X0 U12266 ( .IN1(n12153), .IN2(n12154), .QN(n12152) );
  NAND2X0 U12267 ( .IN1(n12154), .IN2(n12153), .QN(n12150) );
  NOR2X0 U12268 ( .IN1(n12155), .IN2(n12156), .QN(n12153) );
  NOR2X0 U12269 ( .IN1(WX7346), .IN2(n7963), .QN(n12156) );
  INVX0 U12270 ( .INP(n12157), .ZN(n12155) );
  NAND2X0 U12271 ( .IN1(n7963), .IN2(WX7346), .QN(n12157) );
  NAND2X0 U12272 ( .IN1(n12158), .IN2(n12159), .QN(n12154) );
  NAND2X0 U12273 ( .IN1(n7962), .IN2(WX7218), .QN(n12159) );
  INVX0 U12274 ( .INP(n12160), .ZN(n12158) );
  NOR2X0 U12275 ( .IN1(WX7218), .IN2(n7962), .QN(n12160) );
  NAND2X0 U12276 ( .IN1(n9095), .IN2(n12161), .QN(n12148) );
  NAND2X0 U12277 ( .IN1(n997), .IN2(n9280), .QN(n12147) );
  NOR2X0 U12278 ( .IN1(n9239), .IN2(n8924), .QN(n997) );
  NAND2X0 U12279 ( .IN1(n9314), .IN2(CRC_OUT_5_9), .QN(n12146) );
  NAND4X0 U12280 ( .IN1(n12162), .IN2(n12163), .IN3(n12164), .IN4(n12165), 
        .QN(WX5858) );
  NAND3X0 U12281 ( .IN1(n11212), .IN2(n11213), .IN3(n9321), .QN(n12165) );
  NAND3X0 U12282 ( .IN1(n12166), .IN2(n12167), .IN3(n12168), .QN(n11213) );
  INVX0 U12283 ( .INP(n12169), .ZN(n12168) );
  NAND2X0 U12284 ( .IN1(n12169), .IN2(n12170), .QN(n11212) );
  NAND2X0 U12285 ( .IN1(n12166), .IN2(n12167), .QN(n12170) );
  NAND2X0 U12286 ( .IN1(n8230), .IN2(WX7216), .QN(n12167) );
  NAND2X0 U12287 ( .IN1(n3647), .IN2(WX7344), .QN(n12166) );
  NOR2X0 U12288 ( .IN1(n12171), .IN2(n12172), .QN(n12169) );
  INVX0 U12289 ( .INP(n12173), .ZN(n12172) );
  NAND2X0 U12290 ( .IN1(test_so58), .IN2(WX7280), .QN(n12173) );
  NOR2X0 U12291 ( .IN1(WX7280), .IN2(test_so58), .QN(n12171) );
  NAND2X0 U12292 ( .IN1(n9095), .IN2(n12174), .QN(n12164) );
  NAND2X0 U12293 ( .IN1(n996), .IN2(n9280), .QN(n12163) );
  NOR2X0 U12294 ( .IN1(n9238), .IN2(n8925), .QN(n996) );
  NAND2X0 U12295 ( .IN1(n9313), .IN2(CRC_OUT_5_10), .QN(n12162) );
  NAND4X0 U12296 ( .IN1(n12175), .IN2(n12176), .IN3(n12177), .IN4(n12178), 
        .QN(WX5856) );
  NAND2X0 U12297 ( .IN1(n9323), .IN2(n11237), .QN(n12178) );
  NAND2X0 U12298 ( .IN1(n12179), .IN2(n12180), .QN(n11237) );
  INVX0 U12299 ( .INP(n12181), .ZN(n12180) );
  NOR2X0 U12300 ( .IN1(n12182), .IN2(n12183), .QN(n12181) );
  NAND2X0 U12301 ( .IN1(n12183), .IN2(n12182), .QN(n12179) );
  NOR2X0 U12302 ( .IN1(n12184), .IN2(n12185), .QN(n12182) );
  NOR2X0 U12303 ( .IN1(WX7342), .IN2(n7966), .QN(n12185) );
  INVX0 U12304 ( .INP(n12186), .ZN(n12184) );
  NAND2X0 U12305 ( .IN1(n7966), .IN2(WX7342), .QN(n12186) );
  NAND2X0 U12306 ( .IN1(n12187), .IN2(n12188), .QN(n12183) );
  NAND2X0 U12307 ( .IN1(n7965), .IN2(WX7214), .QN(n12188) );
  INVX0 U12308 ( .INP(n12189), .ZN(n12187) );
  NOR2X0 U12309 ( .IN1(WX7214), .IN2(n7965), .QN(n12189) );
  NAND2X0 U12310 ( .IN1(n9095), .IN2(n12190), .QN(n12177) );
  NAND2X0 U12311 ( .IN1(n995), .IN2(n9281), .QN(n12176) );
  NOR2X0 U12312 ( .IN1(n9237), .IN2(n8926), .QN(n995) );
  NAND2X0 U12313 ( .IN1(n9312), .IN2(CRC_OUT_5_11), .QN(n12175) );
  NAND4X0 U12314 ( .IN1(n12191), .IN2(n12192), .IN3(n12193), .IN4(n12194), 
        .QN(WX5854) );
  NAND2X0 U12315 ( .IN1(n9323), .IN2(n11253), .QN(n12194) );
  NAND2X0 U12316 ( .IN1(n12195), .IN2(n12196), .QN(n11253) );
  INVX0 U12317 ( .INP(n12197), .ZN(n12196) );
  NOR2X0 U12318 ( .IN1(n12198), .IN2(n12199), .QN(n12197) );
  NAND2X0 U12319 ( .IN1(n12199), .IN2(n12198), .QN(n12195) );
  NOR2X0 U12320 ( .IN1(n12200), .IN2(n12201), .QN(n12198) );
  NOR2X0 U12321 ( .IN1(WX7340), .IN2(n7968), .QN(n12201) );
  INVX0 U12322 ( .INP(n12202), .ZN(n12200) );
  NAND2X0 U12323 ( .IN1(n7968), .IN2(WX7340), .QN(n12202) );
  NAND2X0 U12324 ( .IN1(n12203), .IN2(n12204), .QN(n12199) );
  NAND2X0 U12325 ( .IN1(n7967), .IN2(WX7212), .QN(n12204) );
  INVX0 U12326 ( .INP(n12205), .ZN(n12203) );
  NOR2X0 U12327 ( .IN1(WX7212), .IN2(n7967), .QN(n12205) );
  NAND2X0 U12328 ( .IN1(n9095), .IN2(n12206), .QN(n12193) );
  NAND2X0 U12329 ( .IN1(n994), .IN2(n9281), .QN(n12192) );
  NOR2X0 U12330 ( .IN1(n9237), .IN2(n8927), .QN(n994) );
  NAND2X0 U12331 ( .IN1(n9297), .IN2(CRC_OUT_5_12), .QN(n12191) );
  NAND4X0 U12332 ( .IN1(n12207), .IN2(n12208), .IN3(n12209), .IN4(n12210), 
        .QN(WX5852) );
  NAND2X0 U12333 ( .IN1(n9324), .IN2(n11266), .QN(n12210) );
  NAND2X0 U12334 ( .IN1(n12211), .IN2(n12212), .QN(n11266) );
  INVX0 U12335 ( .INP(n12213), .ZN(n12212) );
  NOR2X0 U12336 ( .IN1(n12214), .IN2(n12215), .QN(n12213) );
  NAND2X0 U12337 ( .IN1(n12215), .IN2(n12214), .QN(n12211) );
  NOR2X0 U12338 ( .IN1(n12216), .IN2(n12217), .QN(n12214) );
  NOR2X0 U12339 ( .IN1(WX7338), .IN2(n7970), .QN(n12217) );
  INVX0 U12340 ( .INP(n12218), .ZN(n12216) );
  NAND2X0 U12341 ( .IN1(n7970), .IN2(WX7338), .QN(n12218) );
  NAND2X0 U12342 ( .IN1(n12219), .IN2(n12220), .QN(n12215) );
  NAND2X0 U12343 ( .IN1(n7969), .IN2(WX7210), .QN(n12220) );
  INVX0 U12344 ( .INP(n12221), .ZN(n12219) );
  NOR2X0 U12345 ( .IN1(WX7210), .IN2(n7969), .QN(n12221) );
  NAND2X0 U12346 ( .IN1(n9095), .IN2(n12222), .QN(n12209) );
  NAND2X0 U12347 ( .IN1(n993), .IN2(n9281), .QN(n12208) );
  NOR2X0 U12348 ( .IN1(n9237), .IN2(n8928), .QN(n993) );
  NAND2X0 U12349 ( .IN1(n9292), .IN2(CRC_OUT_5_13), .QN(n12207) );
  NAND4X0 U12350 ( .IN1(n12223), .IN2(n12224), .IN3(n12225), .IN4(n12226), 
        .QN(WX5850) );
  NAND2X0 U12351 ( .IN1(n9323), .IN2(n11282), .QN(n12226) );
  NAND2X0 U12352 ( .IN1(n12227), .IN2(n12228), .QN(n11282) );
  INVX0 U12353 ( .INP(n12229), .ZN(n12228) );
  NOR2X0 U12354 ( .IN1(n12230), .IN2(n12231), .QN(n12229) );
  NAND2X0 U12355 ( .IN1(n12231), .IN2(n12230), .QN(n12227) );
  NOR2X0 U12356 ( .IN1(n12232), .IN2(n12233), .QN(n12230) );
  NOR2X0 U12357 ( .IN1(WX7336), .IN2(n7972), .QN(n12233) );
  INVX0 U12358 ( .INP(n12234), .ZN(n12232) );
  NAND2X0 U12359 ( .IN1(n7972), .IN2(WX7336), .QN(n12234) );
  NAND2X0 U12360 ( .IN1(n12235), .IN2(n12236), .QN(n12231) );
  NAND2X0 U12361 ( .IN1(n7971), .IN2(WX7208), .QN(n12236) );
  INVX0 U12362 ( .INP(n12237), .ZN(n12235) );
  NOR2X0 U12363 ( .IN1(WX7208), .IN2(n7971), .QN(n12237) );
  NAND2X0 U12364 ( .IN1(n9095), .IN2(n12238), .QN(n12225) );
  NAND2X0 U12365 ( .IN1(n992), .IN2(n9281), .QN(n12224) );
  NOR2X0 U12366 ( .IN1(n9237), .IN2(n8929), .QN(n992) );
  NAND2X0 U12367 ( .IN1(n9292), .IN2(CRC_OUT_5_14), .QN(n12223) );
  NAND4X0 U12368 ( .IN1(n12239), .IN2(n12240), .IN3(n12241), .IN4(n12242), 
        .QN(WX5848) );
  NAND2X0 U12369 ( .IN1(n9324), .IN2(n11295), .QN(n12242) );
  NAND2X0 U12370 ( .IN1(n12243), .IN2(n12244), .QN(n11295) );
  INVX0 U12371 ( .INP(n12245), .ZN(n12244) );
  NOR2X0 U12372 ( .IN1(n12246), .IN2(n12247), .QN(n12245) );
  NAND2X0 U12373 ( .IN1(n12247), .IN2(n12246), .QN(n12243) );
  NOR2X0 U12374 ( .IN1(n12248), .IN2(n12249), .QN(n12246) );
  NOR2X0 U12375 ( .IN1(WX7334), .IN2(n7974), .QN(n12249) );
  INVX0 U12376 ( .INP(n12250), .ZN(n12248) );
  NAND2X0 U12377 ( .IN1(n7974), .IN2(WX7334), .QN(n12250) );
  NAND2X0 U12378 ( .IN1(n12251), .IN2(n12252), .QN(n12247) );
  NAND2X0 U12379 ( .IN1(n7973), .IN2(WX7206), .QN(n12252) );
  INVX0 U12380 ( .INP(n12253), .ZN(n12251) );
  NOR2X0 U12381 ( .IN1(WX7206), .IN2(n7973), .QN(n12253) );
  NAND2X0 U12382 ( .IN1(n9095), .IN2(n12254), .QN(n12241) );
  NAND2X0 U12383 ( .IN1(n991), .IN2(n9281), .QN(n12240) );
  NOR2X0 U12384 ( .IN1(n9237), .IN2(n8930), .QN(n991) );
  NAND2X0 U12385 ( .IN1(n9292), .IN2(CRC_OUT_5_15), .QN(n12239) );
  NAND4X0 U12386 ( .IN1(n12255), .IN2(n12256), .IN3(n12257), .IN4(n12258), 
        .QN(WX5846) );
  NAND2X0 U12387 ( .IN1(n12259), .IN2(n11315), .QN(n12258) );
  NAND2X0 U12388 ( .IN1(n12260), .IN2(n11318), .QN(n11315) );
  NAND2X0 U12389 ( .IN1(n12261), .IN2(n12262), .QN(n12260) );
  NAND2X0 U12390 ( .IN1(n16381), .IN2(n9119), .QN(n12262) );
  NAND2X0 U12391 ( .IN1(TM1), .IN2(n8421), .QN(n12261) );
  NAND3X0 U12392 ( .IN1(n12263), .IN2(n12264), .IN3(n12265), .QN(n12259) );
  NAND2X0 U12393 ( .IN1(n9323), .IN2(n11318), .QN(n12265) );
  NAND2X0 U12394 ( .IN1(n12266), .IN2(n12267), .QN(n11318) );
  NAND2X0 U12395 ( .IN1(n7712), .IN2(n12268), .QN(n12267) );
  INVX0 U12396 ( .INP(n12269), .ZN(n12266) );
  NOR2X0 U12397 ( .IN1(n12268), .IN2(n7712), .QN(n12269) );
  NOR2X0 U12398 ( .IN1(n12270), .IN2(n12271), .QN(n12268) );
  NOR2X0 U12399 ( .IN1(WX7332), .IN2(n7713), .QN(n12271) );
  INVX0 U12400 ( .INP(n12272), .ZN(n12270) );
  NAND2X0 U12401 ( .IN1(n7713), .IN2(WX7332), .QN(n12272) );
  NAND2X0 U12402 ( .IN1(n9083), .IN2(n8421), .QN(n12264) );
  NAND2X0 U12403 ( .IN1(n16381), .IN2(n9079), .QN(n12263) );
  NAND2X0 U12404 ( .IN1(n12273), .IN2(n9111), .QN(n12257) );
  NAND2X0 U12405 ( .IN1(n990), .IN2(n9281), .QN(n12256) );
  NOR2X0 U12406 ( .IN1(n9237), .IN2(n8931), .QN(n990) );
  NAND2X0 U12407 ( .IN1(n9292), .IN2(CRC_OUT_5_16), .QN(n12255) );
  NAND4X0 U12408 ( .IN1(n12274), .IN2(n12275), .IN3(n12276), .IN4(n12277), 
        .QN(WX5844) );
  NAND2X0 U12409 ( .IN1(n12278), .IN2(n11338), .QN(n12277) );
  NAND2X0 U12410 ( .IN1(n12279), .IN2(n11341), .QN(n11338) );
  NAND2X0 U12411 ( .IN1(n12280), .IN2(n12281), .QN(n12279) );
  NAND2X0 U12412 ( .IN1(n16380), .IN2(n9119), .QN(n12281) );
  NAND2X0 U12413 ( .IN1(TM1), .IN2(n8422), .QN(n12280) );
  NAND3X0 U12414 ( .IN1(n12282), .IN2(n12283), .IN3(n12284), .QN(n12278) );
  NAND2X0 U12415 ( .IN1(n9324), .IN2(n11341), .QN(n12284) );
  NAND2X0 U12416 ( .IN1(n12285), .IN2(n12286), .QN(n11341) );
  NAND2X0 U12417 ( .IN1(n7714), .IN2(n12287), .QN(n12286) );
  INVX0 U12418 ( .INP(n12288), .ZN(n12285) );
  NOR2X0 U12419 ( .IN1(n12287), .IN2(n7714), .QN(n12288) );
  NOR2X0 U12420 ( .IN1(n12289), .IN2(n12290), .QN(n12287) );
  NOR2X0 U12421 ( .IN1(WX7330), .IN2(n7715), .QN(n12290) );
  INVX0 U12422 ( .INP(n12291), .ZN(n12289) );
  NAND2X0 U12423 ( .IN1(n7715), .IN2(WX7330), .QN(n12291) );
  NAND2X0 U12424 ( .IN1(n9082), .IN2(n8422), .QN(n12283) );
  NAND2X0 U12425 ( .IN1(n16380), .IN2(n9078), .QN(n12282) );
  NAND2X0 U12426 ( .IN1(n12292), .IN2(n12293), .QN(n12276) );
  NAND2X0 U12427 ( .IN1(n12294), .IN2(n12295), .QN(n12292) );
  NAND2X0 U12428 ( .IN1(n9096), .IN2(n12296), .QN(n12295) );
  NAND2X0 U12429 ( .IN1(n9096), .IN2(n8480), .QN(n12294) );
  NAND2X0 U12430 ( .IN1(n989), .IN2(n9281), .QN(n12275) );
  NOR2X0 U12431 ( .IN1(n9237), .IN2(n8932), .QN(n989) );
  NAND2X0 U12432 ( .IN1(test_so54), .IN2(n9315), .QN(n12274) );
  NAND4X0 U12433 ( .IN1(n12297), .IN2(n12298), .IN3(n12299), .IN4(n12300), 
        .QN(WX5842) );
  NAND2X0 U12434 ( .IN1(n12301), .IN2(n11361), .QN(n12300) );
  NAND2X0 U12435 ( .IN1(n12302), .IN2(n11364), .QN(n11361) );
  NAND2X0 U12436 ( .IN1(n12303), .IN2(n12304), .QN(n12302) );
  NAND2X0 U12437 ( .IN1(n16379), .IN2(n9119), .QN(n12304) );
  NAND2X0 U12438 ( .IN1(TM1), .IN2(n8423), .QN(n12303) );
  NAND3X0 U12439 ( .IN1(n12305), .IN2(n12306), .IN3(n12307), .QN(n12301) );
  NAND2X0 U12440 ( .IN1(n9323), .IN2(n11364), .QN(n12307) );
  NAND2X0 U12441 ( .IN1(n12308), .IN2(n12309), .QN(n11364) );
  NAND2X0 U12442 ( .IN1(n7716), .IN2(n12310), .QN(n12309) );
  INVX0 U12443 ( .INP(n12311), .ZN(n12308) );
  NOR2X0 U12444 ( .IN1(n12310), .IN2(n7716), .QN(n12311) );
  NOR2X0 U12445 ( .IN1(n12312), .IN2(n12313), .QN(n12310) );
  NOR2X0 U12446 ( .IN1(WX7328), .IN2(n7717), .QN(n12313) );
  INVX0 U12447 ( .INP(n12314), .ZN(n12312) );
  NAND2X0 U12448 ( .IN1(n7717), .IN2(WX7328), .QN(n12314) );
  NAND2X0 U12449 ( .IN1(n10068), .IN2(n8423), .QN(n12306) );
  NAND2X0 U12450 ( .IN1(n16379), .IN2(n10069), .QN(n12305) );
  NAND2X0 U12451 ( .IN1(n12315), .IN2(n9112), .QN(n12299) );
  NAND2X0 U12452 ( .IN1(n988), .IN2(n9281), .QN(n12298) );
  NOR2X0 U12453 ( .IN1(n9236), .IN2(n8933), .QN(n988) );
  NAND2X0 U12454 ( .IN1(n9292), .IN2(CRC_OUT_5_18), .QN(n12297) );
  NAND4X0 U12455 ( .IN1(n12316), .IN2(n12317), .IN3(n12318), .IN4(n12319), 
        .QN(WX5840) );
  NAND2X0 U12456 ( .IN1(n12320), .IN2(n11384), .QN(n12319) );
  NAND2X0 U12457 ( .IN1(n12321), .IN2(n11387), .QN(n11384) );
  NAND2X0 U12458 ( .IN1(n12322), .IN2(n12323), .QN(n12321) );
  NAND2X0 U12459 ( .IN1(n16378), .IN2(n9119), .QN(n12323) );
  NAND2X0 U12460 ( .IN1(TM1), .IN2(n8424), .QN(n12322) );
  NAND3X0 U12461 ( .IN1(n12324), .IN2(n12325), .IN3(n12326), .QN(n12320) );
  NAND2X0 U12462 ( .IN1(n9323), .IN2(n11387), .QN(n12326) );
  NAND2X0 U12463 ( .IN1(n12327), .IN2(n12328), .QN(n11387) );
  NAND2X0 U12464 ( .IN1(n7718), .IN2(n12329), .QN(n12328) );
  INVX0 U12465 ( .INP(n12330), .ZN(n12327) );
  NOR2X0 U12466 ( .IN1(n12329), .IN2(n7718), .QN(n12330) );
  NOR2X0 U12467 ( .IN1(n12331), .IN2(n12332), .QN(n12329) );
  NOR2X0 U12468 ( .IN1(WX7326), .IN2(n7719), .QN(n12332) );
  INVX0 U12469 ( .INP(n12333), .ZN(n12331) );
  NAND2X0 U12470 ( .IN1(n7719), .IN2(WX7326), .QN(n12333) );
  NAND2X0 U12471 ( .IN1(n9084), .IN2(n8424), .QN(n12325) );
  NAND2X0 U12472 ( .IN1(n16378), .IN2(n9080), .QN(n12324) );
  NAND2X0 U12473 ( .IN1(n12334), .IN2(n12335), .QN(n12318) );
  NAND2X0 U12474 ( .IN1(n12336), .IN2(n12337), .QN(n12334) );
  NAND2X0 U12475 ( .IN1(n9096), .IN2(n12338), .QN(n12337) );
  NAND2X0 U12476 ( .IN1(n9096), .IN2(n8482), .QN(n12336) );
  NAND2X0 U12477 ( .IN1(n987), .IN2(n9281), .QN(n12317) );
  NOR2X0 U12478 ( .IN1(n9236), .IN2(n8934), .QN(n987) );
  NAND2X0 U12479 ( .IN1(n9292), .IN2(CRC_OUT_5_19), .QN(n12316) );
  NAND4X0 U12480 ( .IN1(n12339), .IN2(n12340), .IN3(n12341), .IN4(n12342), 
        .QN(WX5838) );
  NAND2X0 U12481 ( .IN1(n12343), .IN2(n11407), .QN(n12342) );
  NAND2X0 U12482 ( .IN1(n12344), .IN2(n11410), .QN(n11407) );
  NAND2X0 U12483 ( .IN1(n12345), .IN2(n12346), .QN(n12344) );
  NAND2X0 U12484 ( .IN1(n16377), .IN2(n9119), .QN(n12346) );
  NAND2X0 U12485 ( .IN1(TM1), .IN2(n8425), .QN(n12345) );
  NAND3X0 U12486 ( .IN1(n12347), .IN2(n12348), .IN3(n12349), .QN(n12343) );
  NAND2X0 U12487 ( .IN1(n9324), .IN2(n11410), .QN(n12349) );
  NAND2X0 U12488 ( .IN1(n12350), .IN2(n12351), .QN(n11410) );
  NAND2X0 U12489 ( .IN1(n7720), .IN2(n12352), .QN(n12351) );
  INVX0 U12490 ( .INP(n12353), .ZN(n12350) );
  NOR2X0 U12491 ( .IN1(n12352), .IN2(n7720), .QN(n12353) );
  NOR2X0 U12492 ( .IN1(n12354), .IN2(n12355), .QN(n12352) );
  NOR2X0 U12493 ( .IN1(WX7324), .IN2(n7721), .QN(n12355) );
  INVX0 U12494 ( .INP(n12356), .ZN(n12354) );
  NAND2X0 U12495 ( .IN1(n7721), .IN2(WX7324), .QN(n12356) );
  NAND2X0 U12496 ( .IN1(n9083), .IN2(n8425), .QN(n12348) );
  NAND2X0 U12497 ( .IN1(n16377), .IN2(n9079), .QN(n12347) );
  NAND2X0 U12498 ( .IN1(n12357), .IN2(n9112), .QN(n12341) );
  NAND2X0 U12499 ( .IN1(n986), .IN2(n9281), .QN(n12340) );
  NOR2X0 U12500 ( .IN1(n9236), .IN2(n8935), .QN(n986) );
  NAND2X0 U12501 ( .IN1(n9292), .IN2(CRC_OUT_5_20), .QN(n12339) );
  NAND4X0 U12502 ( .IN1(n12358), .IN2(n12359), .IN3(n12360), .IN4(n12361), 
        .QN(WX5836) );
  NAND2X0 U12503 ( .IN1(n12362), .IN2(n12363), .QN(n12361) );
  NAND2X0 U12504 ( .IN1(n12364), .IN2(n12365), .QN(n12362) );
  NAND2X0 U12505 ( .IN1(n9096), .IN2(n12366), .QN(n12365) );
  NAND2X0 U12506 ( .IN1(n9096), .IN2(n8484), .QN(n12364) );
  NAND2X0 U12507 ( .IN1(n11429), .IN2(n9336), .QN(n12360) );
  NOR2X0 U12508 ( .IN1(n12367), .IN2(n12368), .QN(n11429) );
  INVX0 U12509 ( .INP(n12369), .ZN(n12368) );
  NAND2X0 U12510 ( .IN1(n12370), .IN2(n12371), .QN(n12369) );
  NOR2X0 U12511 ( .IN1(n12371), .IN2(n12370), .QN(n12367) );
  NAND2X0 U12512 ( .IN1(n12372), .IN2(n12373), .QN(n12370) );
  NAND2X0 U12513 ( .IN1(n12374), .IN2(WX7258), .QN(n12373) );
  NAND2X0 U12514 ( .IN1(n12375), .IN2(n12376), .QN(n12374) );
  NAND3X0 U12515 ( .IN1(n12375), .IN2(n12376), .IN3(n7723), .QN(n12372) );
  NAND2X0 U12516 ( .IN1(test_so63), .IN2(WX7194), .QN(n12376) );
  NAND2X0 U12517 ( .IN1(n7722), .IN2(n8800), .QN(n12375) );
  NOR2X0 U12518 ( .IN1(n12377), .IN2(n12378), .QN(n12371) );
  INVX0 U12519 ( .INP(n12379), .ZN(n12378) );
  NAND2X0 U12520 ( .IN1(n16376), .IN2(n9119), .QN(n12379) );
  NOR2X0 U12521 ( .IN1(n9117), .IN2(n16376), .QN(n12377) );
  NAND2X0 U12522 ( .IN1(n985), .IN2(n9281), .QN(n12359) );
  NOR2X0 U12523 ( .IN1(n9236), .IN2(n8936), .QN(n985) );
  NAND2X0 U12524 ( .IN1(n9292), .IN2(CRC_OUT_5_21), .QN(n12358) );
  NAND4X0 U12525 ( .IN1(n12380), .IN2(n12381), .IN3(n12382), .IN4(n12383), 
        .QN(WX5834) );
  NAND2X0 U12526 ( .IN1(n12384), .IN2(n11449), .QN(n12383) );
  NAND2X0 U12527 ( .IN1(n12385), .IN2(n11452), .QN(n11449) );
  NAND2X0 U12528 ( .IN1(n12386), .IN2(n12387), .QN(n12385) );
  NAND2X0 U12529 ( .IN1(n16375), .IN2(n9119), .QN(n12387) );
  NAND2X0 U12530 ( .IN1(TM1), .IN2(n8427), .QN(n12386) );
  NAND3X0 U12531 ( .IN1(n12388), .IN2(n12389), .IN3(n12390), .QN(n12384) );
  NAND2X0 U12532 ( .IN1(n9323), .IN2(n11452), .QN(n12390) );
  NAND2X0 U12533 ( .IN1(n12391), .IN2(n12392), .QN(n11452) );
  NAND2X0 U12534 ( .IN1(n7724), .IN2(n12393), .QN(n12392) );
  INVX0 U12535 ( .INP(n12394), .ZN(n12391) );
  NOR2X0 U12536 ( .IN1(n12393), .IN2(n7724), .QN(n12394) );
  NOR2X0 U12537 ( .IN1(n12395), .IN2(n12396), .QN(n12393) );
  NOR2X0 U12538 ( .IN1(WX7320), .IN2(n7725), .QN(n12396) );
  INVX0 U12539 ( .INP(n12397), .ZN(n12395) );
  NAND2X0 U12540 ( .IN1(n7725), .IN2(WX7320), .QN(n12397) );
  NAND2X0 U12541 ( .IN1(n9082), .IN2(n8427), .QN(n12389) );
  NAND2X0 U12542 ( .IN1(n16375), .IN2(n9078), .QN(n12388) );
  NAND2X0 U12543 ( .IN1(n12398), .IN2(n12399), .QN(n12382) );
  NAND2X0 U12544 ( .IN1(n12400), .IN2(n12401), .QN(n12398) );
  NAND2X0 U12545 ( .IN1(n9096), .IN2(n12402), .QN(n12401) );
  NAND2X0 U12546 ( .IN1(n8273), .IN2(n9112), .QN(n12400) );
  NAND2X0 U12547 ( .IN1(n984), .IN2(n9281), .QN(n12381) );
  NOR2X0 U12548 ( .IN1(n9236), .IN2(n8937), .QN(n984) );
  NAND2X0 U12549 ( .IN1(n9292), .IN2(CRC_OUT_5_22), .QN(n12380) );
  NAND4X0 U12550 ( .IN1(n12403), .IN2(n12404), .IN3(n12405), .IN4(n12406), 
        .QN(WX5832) );
  NAND2X0 U12551 ( .IN1(n12407), .IN2(n12408), .QN(n12406) );
  NAND2X0 U12552 ( .IN1(n12409), .IN2(n12410), .QN(n12407) );
  NAND2X0 U12553 ( .IN1(n9096), .IN2(n12411), .QN(n12410) );
  NAND2X0 U12554 ( .IN1(n9096), .IN2(n8487), .QN(n12409) );
  NAND2X0 U12555 ( .IN1(n11471), .IN2(n9336), .QN(n12405) );
  NOR2X0 U12556 ( .IN1(n12412), .IN2(n12413), .QN(n11471) );
  INVX0 U12557 ( .INP(n12414), .ZN(n12413) );
  NAND2X0 U12558 ( .IN1(n12415), .IN2(n12416), .QN(n12414) );
  NOR2X0 U12559 ( .IN1(n12416), .IN2(n12415), .QN(n12412) );
  NAND2X0 U12560 ( .IN1(n12417), .IN2(n12418), .QN(n12415) );
  NAND2X0 U12561 ( .IN1(n8220), .IN2(n12419), .QN(n12418) );
  INVX0 U12562 ( .INP(n12420), .ZN(n12419) );
  NAND2X0 U12563 ( .IN1(n12420), .IN2(WX7318), .QN(n12417) );
  NAND2X0 U12564 ( .IN1(n12421), .IN2(n12422), .QN(n12420) );
  INVX0 U12565 ( .INP(n12423), .ZN(n12422) );
  NOR2X0 U12566 ( .IN1(n8810), .IN2(n16374), .QN(n12423) );
  NAND2X0 U12567 ( .IN1(n16374), .IN2(n8810), .QN(n12421) );
  NOR2X0 U12568 ( .IN1(n12424), .IN2(n12425), .QN(n12416) );
  INVX0 U12569 ( .INP(n12426), .ZN(n12425) );
  NAND2X0 U12570 ( .IN1(n7726), .IN2(n9119), .QN(n12426) );
  NOR2X0 U12571 ( .IN1(n9117), .IN2(n7726), .QN(n12424) );
  NAND2X0 U12572 ( .IN1(n983), .IN2(n9281), .QN(n12404) );
  NOR2X0 U12573 ( .IN1(n9236), .IN2(n8938), .QN(n983) );
  NAND2X0 U12574 ( .IN1(n9292), .IN2(CRC_OUT_5_23), .QN(n12403) );
  NAND4X0 U12575 ( .IN1(n12427), .IN2(n12428), .IN3(n12429), .IN4(n12430), 
        .QN(WX5830) );
  NAND2X0 U12576 ( .IN1(n12431), .IN2(n11491), .QN(n12430) );
  NAND2X0 U12577 ( .IN1(n12432), .IN2(n11494), .QN(n11491) );
  NAND2X0 U12578 ( .IN1(n12433), .IN2(n12434), .QN(n12432) );
  NAND2X0 U12579 ( .IN1(n16373), .IN2(n9119), .QN(n12434) );
  NAND2X0 U12580 ( .IN1(TM1), .IN2(n8429), .QN(n12433) );
  NAND3X0 U12581 ( .IN1(n12435), .IN2(n12436), .IN3(n12437), .QN(n12431) );
  NAND2X0 U12582 ( .IN1(n9323), .IN2(n11494), .QN(n12437) );
  NAND2X0 U12583 ( .IN1(n12438), .IN2(n12439), .QN(n11494) );
  NAND2X0 U12584 ( .IN1(n7727), .IN2(n12440), .QN(n12439) );
  INVX0 U12585 ( .INP(n12441), .ZN(n12438) );
  NOR2X0 U12586 ( .IN1(n12440), .IN2(n7727), .QN(n12441) );
  NOR2X0 U12587 ( .IN1(n12442), .IN2(n12443), .QN(n12440) );
  NOR2X0 U12588 ( .IN1(WX7316), .IN2(n7728), .QN(n12443) );
  INVX0 U12589 ( .INP(n12444), .ZN(n12442) );
  NAND2X0 U12590 ( .IN1(n7728), .IN2(WX7316), .QN(n12444) );
  NAND2X0 U12591 ( .IN1(n10068), .IN2(n8429), .QN(n12436) );
  NAND2X0 U12592 ( .IN1(n16373), .IN2(n10069), .QN(n12435) );
  NAND2X0 U12593 ( .IN1(n12445), .IN2(n12446), .QN(n12429) );
  NAND2X0 U12594 ( .IN1(n12447), .IN2(n12448), .QN(n12445) );
  NAND2X0 U12595 ( .IN1(n9096), .IN2(n12449), .QN(n12448) );
  NAND2X0 U12596 ( .IN1(n9096), .IN2(n8488), .QN(n12447) );
  NAND2X0 U12597 ( .IN1(n982), .IN2(n9281), .QN(n12428) );
  NOR2X0 U12598 ( .IN1(n9068), .IN2(n9162), .QN(n982) );
  NAND2X0 U12599 ( .IN1(n9292), .IN2(CRC_OUT_5_24), .QN(n12427) );
  NAND4X0 U12600 ( .IN1(n12450), .IN2(n12451), .IN3(n12452), .IN4(n12453), 
        .QN(WX5828) );
  NAND2X0 U12601 ( .IN1(n12454), .IN2(n12455), .QN(n12453) );
  NAND2X0 U12602 ( .IN1(n12456), .IN2(n12457), .QN(n12454) );
  NAND2X0 U12603 ( .IN1(n9096), .IN2(n12458), .QN(n12457) );
  NAND2X0 U12604 ( .IN1(n9096), .IN2(n8489), .QN(n12456) );
  NAND2X0 U12605 ( .IN1(n11513), .IN2(n9336), .QN(n12452) );
  NOR2X0 U12606 ( .IN1(n12459), .IN2(n12460), .QN(n11513) );
  INVX0 U12607 ( .INP(n12461), .ZN(n12460) );
  NAND2X0 U12608 ( .IN1(n12462), .IN2(n12463), .QN(n12461) );
  NOR2X0 U12609 ( .IN1(n12463), .IN2(n12462), .QN(n12459) );
  NAND2X0 U12610 ( .IN1(n12464), .IN2(n12465), .QN(n12462) );
  NAND2X0 U12611 ( .IN1(n8218), .IN2(n12466), .QN(n12465) );
  INVX0 U12612 ( .INP(n12467), .ZN(n12466) );
  NAND2X0 U12613 ( .IN1(n12467), .IN2(WX7314), .QN(n12464) );
  NAND2X0 U12614 ( .IN1(n12468), .IN2(n12469), .QN(n12467) );
  INVX0 U12615 ( .INP(n12470), .ZN(n12469) );
  NOR2X0 U12616 ( .IN1(n8811), .IN2(n16372), .QN(n12470) );
  NAND2X0 U12617 ( .IN1(n16372), .IN2(n8811), .QN(n12468) );
  NOR2X0 U12618 ( .IN1(n12471), .IN2(n12472), .QN(n12463) );
  INVX0 U12619 ( .INP(n12473), .ZN(n12472) );
  NAND2X0 U12620 ( .IN1(n7729), .IN2(n9119), .QN(n12473) );
  NOR2X0 U12621 ( .IN1(n9117), .IN2(n7729), .QN(n12471) );
  NAND2X0 U12622 ( .IN1(n981), .IN2(n9281), .QN(n12451) );
  NOR2X0 U12623 ( .IN1(n9236), .IN2(n8939), .QN(n981) );
  NAND2X0 U12624 ( .IN1(n9293), .IN2(CRC_OUT_5_25), .QN(n12450) );
  NAND4X0 U12625 ( .IN1(n12474), .IN2(n12475), .IN3(n12476), .IN4(n12477), 
        .QN(WX5826) );
  NAND2X0 U12626 ( .IN1(n12478), .IN2(n11519), .QN(n12477) );
  NAND2X0 U12627 ( .IN1(n12479), .IN2(n11522), .QN(n11519) );
  NAND2X0 U12628 ( .IN1(n12480), .IN2(n12481), .QN(n12479) );
  NAND2X0 U12629 ( .IN1(n16371), .IN2(n9119), .QN(n12481) );
  NAND2X0 U12630 ( .IN1(TM1), .IN2(n8431), .QN(n12480) );
  NAND3X0 U12631 ( .IN1(n12482), .IN2(n12483), .IN3(n12484), .QN(n12478) );
  NAND2X0 U12632 ( .IN1(n9324), .IN2(n11522), .QN(n12484) );
  NAND2X0 U12633 ( .IN1(n12485), .IN2(n12486), .QN(n11522) );
  NAND2X0 U12634 ( .IN1(n7730), .IN2(n12487), .QN(n12486) );
  INVX0 U12635 ( .INP(n12488), .ZN(n12485) );
  NOR2X0 U12636 ( .IN1(n12487), .IN2(n7730), .QN(n12488) );
  NOR2X0 U12637 ( .IN1(n12489), .IN2(n12490), .QN(n12487) );
  NOR2X0 U12638 ( .IN1(WX7312), .IN2(n7731), .QN(n12490) );
  INVX0 U12639 ( .INP(n12491), .ZN(n12489) );
  NAND2X0 U12640 ( .IN1(n7731), .IN2(WX7312), .QN(n12491) );
  NAND2X0 U12641 ( .IN1(n9084), .IN2(n8431), .QN(n12483) );
  NAND2X0 U12642 ( .IN1(n16371), .IN2(n9080), .QN(n12482) );
  NAND2X0 U12643 ( .IN1(n12492), .IN2(n12493), .QN(n12476) );
  NAND2X0 U12644 ( .IN1(n12494), .IN2(n12495), .QN(n12492) );
  NAND2X0 U12645 ( .IN1(n9109), .IN2(n12496), .QN(n12495) );
  NAND2X0 U12646 ( .IN1(n9106), .IN2(n8490), .QN(n12494) );
  NAND2X0 U12647 ( .IN1(n980), .IN2(n9281), .QN(n12475) );
  NOR2X0 U12648 ( .IN1(n9236), .IN2(n8940), .QN(n980) );
  NAND2X0 U12649 ( .IN1(n9293), .IN2(CRC_OUT_5_26), .QN(n12474) );
  NAND4X0 U12650 ( .IN1(n12497), .IN2(n12498), .IN3(n12499), .IN4(n12500), 
        .QN(WX5824) );
  NAND2X0 U12651 ( .IN1(n12501), .IN2(n11555), .QN(n12500) );
  NAND3X0 U12652 ( .IN1(n12502), .IN2(n12503), .IN3(n11558), .QN(n11555) );
  NAND2X0 U12653 ( .IN1(n8216), .IN2(n9119), .QN(n12503) );
  NAND2X0 U12654 ( .IN1(TM1), .IN2(WX7310), .QN(n12502) );
  NAND3X0 U12655 ( .IN1(n12504), .IN2(n12505), .IN3(n12506), .QN(n12501) );
  NAND2X0 U12656 ( .IN1(n9324), .IN2(n11558), .QN(n12506) );
  NAND2X0 U12657 ( .IN1(n12507), .IN2(n12508), .QN(n11558) );
  NAND2X0 U12658 ( .IN1(n12509), .IN2(WX7246), .QN(n12508) );
  NAND2X0 U12659 ( .IN1(n12510), .IN2(n12511), .QN(n12509) );
  NAND3X0 U12660 ( .IN1(n12510), .IN2(n12511), .IN3(n7733), .QN(n12507) );
  NAND2X0 U12661 ( .IN1(test_so57), .IN2(WX7182), .QN(n12511) );
  NAND2X0 U12662 ( .IN1(n7732), .IN2(n8821), .QN(n12510) );
  NAND2X0 U12663 ( .IN1(n9078), .IN2(WX7310), .QN(n12505) );
  NAND2X0 U12664 ( .IN1(n9083), .IN2(n8216), .QN(n12504) );
  NAND2X0 U12665 ( .IN1(n12512), .IN2(n12513), .QN(n12499) );
  NAND2X0 U12666 ( .IN1(n12514), .IN2(n12515), .QN(n12512) );
  NAND2X0 U12667 ( .IN1(n9106), .IN2(n12516), .QN(n12515) );
  NAND2X0 U12668 ( .IN1(n9106), .IN2(n8491), .QN(n12514) );
  NAND2X0 U12669 ( .IN1(n979), .IN2(n9281), .QN(n12498) );
  NOR2X0 U12670 ( .IN1(n9236), .IN2(n8941), .QN(n979) );
  NAND2X0 U12671 ( .IN1(n9293), .IN2(CRC_OUT_5_27), .QN(n12497) );
  NAND4X0 U12672 ( .IN1(n12517), .IN2(n12518), .IN3(n12519), .IN4(n12520), 
        .QN(WX5822) );
  NAND2X0 U12673 ( .IN1(n12521), .IN2(n11564), .QN(n12520) );
  NAND2X0 U12674 ( .IN1(n12522), .IN2(n11567), .QN(n11564) );
  NAND2X0 U12675 ( .IN1(n12523), .IN2(n12524), .QN(n12522) );
  NAND2X0 U12676 ( .IN1(n16370), .IN2(n9119), .QN(n12524) );
  NAND2X0 U12677 ( .IN1(TM1), .IN2(n8434), .QN(n12523) );
  NAND3X0 U12678 ( .IN1(n12525), .IN2(n12526), .IN3(n12527), .QN(n12521) );
  NAND2X0 U12679 ( .IN1(n9324), .IN2(n11567), .QN(n12527) );
  NAND2X0 U12680 ( .IN1(n12528), .IN2(n12529), .QN(n11567) );
  NAND2X0 U12681 ( .IN1(n7734), .IN2(n12530), .QN(n12529) );
  INVX0 U12682 ( .INP(n12531), .ZN(n12528) );
  NOR2X0 U12683 ( .IN1(n12530), .IN2(n7734), .QN(n12531) );
  NOR2X0 U12684 ( .IN1(n12532), .IN2(n12533), .QN(n12530) );
  NOR2X0 U12685 ( .IN1(WX7308), .IN2(n7735), .QN(n12533) );
  INVX0 U12686 ( .INP(n12534), .ZN(n12532) );
  NAND2X0 U12687 ( .IN1(n7735), .IN2(WX7308), .QN(n12534) );
  NAND2X0 U12688 ( .IN1(n9082), .IN2(n8434), .QN(n12526) );
  NAND2X0 U12689 ( .IN1(n16370), .IN2(n9079), .QN(n12525) );
  NAND2X0 U12690 ( .IN1(n12535), .IN2(n12536), .QN(n12519) );
  NAND2X0 U12691 ( .IN1(n12537), .IN2(n12538), .QN(n12535) );
  NAND2X0 U12692 ( .IN1(n9106), .IN2(n12539), .QN(n12538) );
  NAND2X0 U12693 ( .IN1(n9106), .IN2(n8492), .QN(n12537) );
  NAND2X0 U12694 ( .IN1(n978), .IN2(n9282), .QN(n12518) );
  NOR2X0 U12695 ( .IN1(n9236), .IN2(n8942), .QN(n978) );
  NAND2X0 U12696 ( .IN1(n9293), .IN2(CRC_OUT_5_28), .QN(n12517) );
  NAND4X0 U12697 ( .IN1(n12540), .IN2(n12541), .IN3(n12542), .IN4(n12543), 
        .QN(WX5820) );
  NAND2X0 U12698 ( .IN1(n12544), .IN2(n11602), .QN(n12543) );
  NAND2X0 U12699 ( .IN1(n12545), .IN2(n11605), .QN(n11602) );
  NAND2X0 U12700 ( .IN1(n12546), .IN2(n12547), .QN(n12545) );
  NAND2X0 U12701 ( .IN1(n16369), .IN2(n9119), .QN(n12547) );
  NAND2X0 U12702 ( .IN1(TM1), .IN2(n8435), .QN(n12546) );
  NAND3X0 U12703 ( .IN1(n12548), .IN2(n12549), .IN3(n12550), .QN(n12544) );
  NAND2X0 U12704 ( .IN1(n9324), .IN2(n11605), .QN(n12550) );
  NAND2X0 U12705 ( .IN1(n12551), .IN2(n12552), .QN(n11605) );
  NAND2X0 U12706 ( .IN1(n7736), .IN2(n12553), .QN(n12552) );
  INVX0 U12707 ( .INP(n12554), .ZN(n12551) );
  NOR2X0 U12708 ( .IN1(n12553), .IN2(n7736), .QN(n12554) );
  NOR2X0 U12709 ( .IN1(n12555), .IN2(n12556), .QN(n12553) );
  NOR2X0 U12710 ( .IN1(WX7306), .IN2(n7737), .QN(n12556) );
  INVX0 U12711 ( .INP(n12557), .ZN(n12555) );
  NAND2X0 U12712 ( .IN1(n7737), .IN2(WX7306), .QN(n12557) );
  NAND2X0 U12713 ( .IN1(n10068), .IN2(n8435), .QN(n12549) );
  NAND2X0 U12714 ( .IN1(n16369), .IN2(n9078), .QN(n12548) );
  NAND2X0 U12715 ( .IN1(n12558), .IN2(n12559), .QN(n12542) );
  NAND2X0 U12716 ( .IN1(n12560), .IN2(n12561), .QN(n12558) );
  NAND2X0 U12717 ( .IN1(n9106), .IN2(n12562), .QN(n12561) );
  NAND2X0 U12718 ( .IN1(n9107), .IN2(n8493), .QN(n12560) );
  NAND2X0 U12719 ( .IN1(n977), .IN2(n9282), .QN(n12541) );
  NOR2X0 U12720 ( .IN1(n9236), .IN2(n8943), .QN(n977) );
  NAND2X0 U12721 ( .IN1(n9293), .IN2(CRC_OUT_5_29), .QN(n12540) );
  NAND4X0 U12722 ( .IN1(n12563), .IN2(n12564), .IN3(n12565), .IN4(n12566), 
        .QN(WX5818) );
  NAND2X0 U12723 ( .IN1(n12567), .IN2(n11611), .QN(n12566) );
  NAND2X0 U12724 ( .IN1(n12568), .IN2(n11614), .QN(n11611) );
  NAND2X0 U12725 ( .IN1(n12569), .IN2(n12570), .QN(n12568) );
  NAND2X0 U12726 ( .IN1(n16368), .IN2(n9118), .QN(n12570) );
  NAND2X0 U12727 ( .IN1(TM1), .IN2(n8436), .QN(n12569) );
  NAND3X0 U12728 ( .IN1(n12571), .IN2(n12572), .IN3(n12573), .QN(n12567) );
  NAND2X0 U12729 ( .IN1(n9324), .IN2(n11614), .QN(n12573) );
  NAND2X0 U12730 ( .IN1(n12574), .IN2(n12575), .QN(n11614) );
  NAND2X0 U12731 ( .IN1(n7738), .IN2(n12576), .QN(n12575) );
  INVX0 U12732 ( .INP(n12577), .ZN(n12574) );
  NOR2X0 U12733 ( .IN1(n12576), .IN2(n7738), .QN(n12577) );
  NOR2X0 U12734 ( .IN1(n12578), .IN2(n12579), .QN(n12576) );
  NOR2X0 U12735 ( .IN1(WX7304), .IN2(n7739), .QN(n12579) );
  INVX0 U12736 ( .INP(n12580), .ZN(n12578) );
  NAND2X0 U12737 ( .IN1(n7739), .IN2(WX7304), .QN(n12580) );
  NAND2X0 U12738 ( .IN1(n9084), .IN2(n8436), .QN(n12572) );
  NAND2X0 U12739 ( .IN1(n16368), .IN2(n10069), .QN(n12571) );
  NAND2X0 U12740 ( .IN1(n12581), .IN2(n12582), .QN(n12565) );
  NAND2X0 U12741 ( .IN1(n12583), .IN2(n12584), .QN(n12581) );
  NAND2X0 U12742 ( .IN1(n9107), .IN2(n12585), .QN(n12584) );
  NAND2X0 U12743 ( .IN1(n9107), .IN2(n8494), .QN(n12583) );
  NAND2X0 U12744 ( .IN1(n976), .IN2(n9282), .QN(n12564) );
  NOR2X0 U12745 ( .IN1(n9236), .IN2(n8944), .QN(n976) );
  NAND2X0 U12746 ( .IN1(n9293), .IN2(CRC_OUT_5_30), .QN(n12563) );
  NAND4X0 U12747 ( .IN1(n12586), .IN2(n12587), .IN3(n12588), .IN4(n12589), 
        .QN(WX5816) );
  NAND2X0 U12748 ( .IN1(n12590), .IN2(n11649), .QN(n12589) );
  NAND2X0 U12749 ( .IN1(n12591), .IN2(n11652), .QN(n11649) );
  NAND2X0 U12750 ( .IN1(n12592), .IN2(n12593), .QN(n12591) );
  NAND2X0 U12751 ( .IN1(n16367), .IN2(n9118), .QN(n12593) );
  NAND2X0 U12752 ( .IN1(TM1), .IN2(n8437), .QN(n12592) );
  NAND3X0 U12753 ( .IN1(n12594), .IN2(n12595), .IN3(n12596), .QN(n12590) );
  NAND2X0 U12754 ( .IN1(n9324), .IN2(n11652), .QN(n12596) );
  NAND2X0 U12755 ( .IN1(n12597), .IN2(n12598), .QN(n11652) );
  NAND2X0 U12756 ( .IN1(n7618), .IN2(n12599), .QN(n12598) );
  INVX0 U12757 ( .INP(n12600), .ZN(n12597) );
  NOR2X0 U12758 ( .IN1(n12599), .IN2(n7618), .QN(n12600) );
  NOR2X0 U12759 ( .IN1(n12601), .IN2(n12602), .QN(n12599) );
  NOR2X0 U12760 ( .IN1(WX7302), .IN2(n7619), .QN(n12602) );
  INVX0 U12761 ( .INP(n12603), .ZN(n12601) );
  NAND2X0 U12762 ( .IN1(n7619), .IN2(WX7302), .QN(n12603) );
  NAND2X0 U12763 ( .IN1(n9083), .IN2(n8437), .QN(n12595) );
  NAND2X0 U12764 ( .IN1(n16367), .IN2(n9080), .QN(n12594) );
  NAND2X0 U12765 ( .IN1(n12604), .IN2(n12605), .QN(n12588) );
  NAND2X0 U12766 ( .IN1(n12606), .IN2(n12607), .QN(n12604) );
  NAND2X0 U12767 ( .IN1(n9107), .IN2(n12608), .QN(n12607) );
  NAND2X0 U12768 ( .IN1(n9107), .IN2(n8495), .QN(n12606) );
  NAND2X0 U12769 ( .IN1(n9293), .IN2(CRC_OUT_5_31), .QN(n12587) );
  NAND2X0 U12770 ( .IN1(n2245), .IN2(WX5657), .QN(n12586) );
  NOR2X0 U12771 ( .IN1(n9236), .IN2(WX5657), .QN(WX5718) );
  NOR2X0 U12772 ( .IN1(n9235), .IN2(WX485), .QN(WX546) );
  NOR3X0 U12773 ( .IN1(n9140), .IN2(n12609), .IN3(n12610), .QN(WX5205) );
  NOR2X0 U12774 ( .IN1(n8355), .IN2(CRC_OUT_6_30), .QN(n12610) );
  NOR2X0 U12775 ( .IN1(DFF_766_n1), .IN2(WX4716), .QN(n12609) );
  NOR3X0 U12776 ( .IN1(n9140), .IN2(n12611), .IN3(n12612), .QN(WX5203) );
  NOR2X0 U12777 ( .IN1(n8356), .IN2(CRC_OUT_6_29), .QN(n12612) );
  NOR2X0 U12778 ( .IN1(DFF_765_n1), .IN2(WX4718), .QN(n12611) );
  NOR3X0 U12779 ( .IN1(n9140), .IN2(n12613), .IN3(n12614), .QN(WX5201) );
  NOR2X0 U12780 ( .IN1(n8357), .IN2(CRC_OUT_6_28), .QN(n12614) );
  NOR2X0 U12781 ( .IN1(DFF_764_n1), .IN2(WX4720), .QN(n12613) );
  NOR2X0 U12782 ( .IN1(n9235), .IN2(n12615), .QN(WX5199) );
  NOR2X0 U12783 ( .IN1(n12616), .IN2(n12617), .QN(n12615) );
  NOR2X0 U12784 ( .IN1(test_so40), .IN2(CRC_OUT_6_27), .QN(n12617) );
  NOR2X0 U12785 ( .IN1(DFF_763_n1), .IN2(n8801), .QN(n12616) );
  NOR3X0 U12786 ( .IN1(n9140), .IN2(n12618), .IN3(n12619), .QN(WX5197) );
  NOR2X0 U12787 ( .IN1(n8358), .IN2(CRC_OUT_6_26), .QN(n12619) );
  NOR2X0 U12788 ( .IN1(DFF_762_n1), .IN2(WX4724), .QN(n12618) );
  NOR3X0 U12789 ( .IN1(n9140), .IN2(n12620), .IN3(n12621), .QN(WX5195) );
  NOR2X0 U12790 ( .IN1(n8359), .IN2(CRC_OUT_6_25), .QN(n12621) );
  NOR2X0 U12791 ( .IN1(DFF_761_n1), .IN2(WX4726), .QN(n12620) );
  NOR3X0 U12792 ( .IN1(n9140), .IN2(n12622), .IN3(n12623), .QN(WX5193) );
  NOR2X0 U12793 ( .IN1(n8360), .IN2(CRC_OUT_6_24), .QN(n12623) );
  NOR2X0 U12794 ( .IN1(DFF_760_n1), .IN2(WX4728), .QN(n12622) );
  NOR3X0 U12795 ( .IN1(n9140), .IN2(n12624), .IN3(n12625), .QN(WX5191) );
  NOR2X0 U12796 ( .IN1(n8361), .IN2(CRC_OUT_6_23), .QN(n12625) );
  NOR2X0 U12797 ( .IN1(DFF_759_n1), .IN2(WX4730), .QN(n12624) );
  NOR2X0 U12798 ( .IN1(n9235), .IN2(n12626), .QN(WX5189) );
  NOR2X0 U12799 ( .IN1(n12627), .IN2(n12628), .QN(n12626) );
  NOR2X0 U12800 ( .IN1(test_so43), .IN2(WX4732), .QN(n12628) );
  INVX0 U12801 ( .INP(n12629), .ZN(n12627) );
  NAND2X0 U12802 ( .IN1(WX4732), .IN2(test_so43), .QN(n12629) );
  NOR3X0 U12803 ( .IN1(n9140), .IN2(n12630), .IN3(n12631), .QN(WX5187) );
  NOR2X0 U12804 ( .IN1(n8379), .IN2(CRC_OUT_6_21), .QN(n12631) );
  NOR2X0 U12805 ( .IN1(DFF_757_n1), .IN2(WX4734), .QN(n12630) );
  NOR3X0 U12806 ( .IN1(n9140), .IN2(n12632), .IN3(n12633), .QN(WX5185) );
  NOR2X0 U12807 ( .IN1(n8380), .IN2(CRC_OUT_6_20), .QN(n12633) );
  NOR2X0 U12808 ( .IN1(DFF_756_n1), .IN2(WX4736), .QN(n12632) );
  NOR3X0 U12809 ( .IN1(n9140), .IN2(n12634), .IN3(n12635), .QN(WX5183) );
  NOR2X0 U12810 ( .IN1(n8397), .IN2(CRC_OUT_6_19), .QN(n12635) );
  NOR2X0 U12811 ( .IN1(DFF_755_n1), .IN2(WX4738), .QN(n12634) );
  NOR3X0 U12812 ( .IN1(n9139), .IN2(n12636), .IN3(n12637), .QN(WX5181) );
  NOR2X0 U12813 ( .IN1(n8398), .IN2(CRC_OUT_6_18), .QN(n12637) );
  NOR2X0 U12814 ( .IN1(DFF_754_n1), .IN2(WX4740), .QN(n12636) );
  NOR3X0 U12815 ( .IN1(n9139), .IN2(n12638), .IN3(n12639), .QN(WX5179) );
  NOR2X0 U12816 ( .IN1(n8412), .IN2(CRC_OUT_6_17), .QN(n12639) );
  NOR2X0 U12817 ( .IN1(DFF_753_n1), .IN2(WX4742), .QN(n12638) );
  NOR3X0 U12818 ( .IN1(n9139), .IN2(n12640), .IN3(n12641), .QN(WX5177) );
  NOR2X0 U12819 ( .IN1(n8413), .IN2(CRC_OUT_6_16), .QN(n12641) );
  NOR2X0 U12820 ( .IN1(DFF_752_n1), .IN2(WX4744), .QN(n12640) );
  NOR2X0 U12821 ( .IN1(n9234), .IN2(n12642), .QN(WX5175) );
  NOR2X0 U12822 ( .IN1(n12643), .IN2(n12644), .QN(n12642) );
  INVX0 U12823 ( .INP(n12645), .ZN(n12644) );
  NAND2X0 U12824 ( .IN1(CRC_OUT_6_15), .IN2(n12646), .QN(n12645) );
  NOR2X0 U12825 ( .IN1(n12646), .IN2(CRC_OUT_6_15), .QN(n12643) );
  NAND2X0 U12826 ( .IN1(n12647), .IN2(n12648), .QN(n12646) );
  NAND2X0 U12827 ( .IN1(n8118), .IN2(CRC_OUT_6_31), .QN(n12648) );
  NAND2X0 U12828 ( .IN1(DFF_767_n1), .IN2(WX4746), .QN(n12647) );
  NOR3X0 U12829 ( .IN1(n9139), .IN2(n12649), .IN3(n12650), .QN(WX5173) );
  NOR2X0 U12830 ( .IN1(n8414), .IN2(CRC_OUT_6_14), .QN(n12650) );
  NOR2X0 U12831 ( .IN1(DFF_750_n1), .IN2(WX4748), .QN(n12649) );
  NOR3X0 U12832 ( .IN1(n9139), .IN2(n12651), .IN3(n12652), .QN(WX5171) );
  NOR2X0 U12833 ( .IN1(n8415), .IN2(CRC_OUT_6_13), .QN(n12652) );
  NOR2X0 U12834 ( .IN1(DFF_749_n1), .IN2(WX4750), .QN(n12651) );
  NOR3X0 U12835 ( .IN1(n9139), .IN2(n12653), .IN3(n12654), .QN(WX5169) );
  NOR2X0 U12836 ( .IN1(n8416), .IN2(CRC_OUT_6_12), .QN(n12654) );
  NOR2X0 U12837 ( .IN1(DFF_748_n1), .IN2(WX4752), .QN(n12653) );
  NOR3X0 U12838 ( .IN1(n9139), .IN2(n12655), .IN3(n12656), .QN(WX5167) );
  NOR2X0 U12839 ( .IN1(n8417), .IN2(CRC_OUT_6_11), .QN(n12656) );
  NOR2X0 U12840 ( .IN1(DFF_747_n1), .IN2(WX4754), .QN(n12655) );
  NOR3X0 U12841 ( .IN1(n9139), .IN2(n12657), .IN3(n12658), .QN(WX5165) );
  INVX0 U12842 ( .INP(n12659), .ZN(n12658) );
  NAND2X0 U12843 ( .IN1(CRC_OUT_6_10), .IN2(n12660), .QN(n12659) );
  NOR2X0 U12844 ( .IN1(n12660), .IN2(CRC_OUT_6_10), .QN(n12657) );
  NAND2X0 U12845 ( .IN1(n12661), .IN2(n12662), .QN(n12660) );
  NAND2X0 U12846 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .QN(n12662) );
  NAND2X0 U12847 ( .IN1(DFF_767_n1), .IN2(n8797), .QN(n12661) );
  NOR3X0 U12848 ( .IN1(n9139), .IN2(n12663), .IN3(n12664), .QN(WX5163) );
  NOR2X0 U12849 ( .IN1(n8418), .IN2(CRC_OUT_6_9), .QN(n12664) );
  NOR2X0 U12850 ( .IN1(DFF_745_n1), .IN2(WX4758), .QN(n12663) );
  NOR3X0 U12851 ( .IN1(n9139), .IN2(n12665), .IN3(n12666), .QN(WX5161) );
  NOR2X0 U12852 ( .IN1(n8419), .IN2(CRC_OUT_6_8), .QN(n12666) );
  NOR2X0 U12853 ( .IN1(DFF_744_n1), .IN2(WX4760), .QN(n12665) );
  NOR3X0 U12854 ( .IN1(n9139), .IN2(n12667), .IN3(n12668), .QN(WX5159) );
  NOR2X0 U12855 ( .IN1(n8420), .IN2(CRC_OUT_6_7), .QN(n12668) );
  NOR2X0 U12856 ( .IN1(DFF_743_n1), .IN2(WX4762), .QN(n12667) );
  NOR3X0 U12857 ( .IN1(n9139), .IN2(n12669), .IN3(n12670), .QN(WX5157) );
  NOR2X0 U12858 ( .IN1(n8432), .IN2(CRC_OUT_6_6), .QN(n12670) );
  NOR2X0 U12859 ( .IN1(DFF_742_n1), .IN2(WX4764), .QN(n12669) );
  NOR2X0 U12860 ( .IN1(n9232), .IN2(n12671), .QN(WX5155) );
  NOR2X0 U12861 ( .IN1(n12672), .IN2(n12673), .QN(n12671) );
  NOR2X0 U12862 ( .IN1(test_so42), .IN2(WX4766), .QN(n12673) );
  INVX0 U12863 ( .INP(n12674), .ZN(n12672) );
  NAND2X0 U12864 ( .IN1(WX4766), .IN2(test_so42), .QN(n12674) );
  NOR3X0 U12865 ( .IN1(n9138), .IN2(n12675), .IN3(n12676), .QN(WX5153) );
  NOR2X0 U12866 ( .IN1(n8450), .IN2(CRC_OUT_6_4), .QN(n12676) );
  NOR2X0 U12867 ( .IN1(DFF_740_n1), .IN2(WX4768), .QN(n12675) );
  NOR2X0 U12868 ( .IN1(n9232), .IN2(n12677), .QN(WX5151) );
  NOR2X0 U12869 ( .IN1(n12678), .IN2(n12679), .QN(n12677) );
  INVX0 U12870 ( .INP(n12680), .ZN(n12679) );
  NAND2X0 U12871 ( .IN1(CRC_OUT_6_3), .IN2(n12681), .QN(n12680) );
  NOR2X0 U12872 ( .IN1(n12681), .IN2(CRC_OUT_6_3), .QN(n12678) );
  NAND2X0 U12873 ( .IN1(n12682), .IN2(n12683), .QN(n12681) );
  NAND2X0 U12874 ( .IN1(n8119), .IN2(CRC_OUT_6_31), .QN(n12683) );
  NAND2X0 U12875 ( .IN1(DFF_767_n1), .IN2(WX4770), .QN(n12682) );
  NOR3X0 U12876 ( .IN1(n9138), .IN2(n12684), .IN3(n12685), .QN(WX5149) );
  NOR2X0 U12877 ( .IN1(n8451), .IN2(CRC_OUT_6_2), .QN(n12685) );
  NOR2X0 U12878 ( .IN1(DFF_738_n1), .IN2(WX4772), .QN(n12684) );
  NOR3X0 U12879 ( .IN1(n9138), .IN2(n12686), .IN3(n12687), .QN(WX5147) );
  NOR2X0 U12880 ( .IN1(n8468), .IN2(CRC_OUT_6_1), .QN(n12687) );
  NOR2X0 U12881 ( .IN1(DFF_737_n1), .IN2(WX4774), .QN(n12686) );
  NOR3X0 U12882 ( .IN1(n9138), .IN2(n12688), .IN3(n12689), .QN(WX5145) );
  NOR2X0 U12883 ( .IN1(n8469), .IN2(CRC_OUT_6_0), .QN(n12689) );
  NOR2X0 U12884 ( .IN1(DFF_736_n1), .IN2(WX4776), .QN(n12688) );
  NOR3X0 U12885 ( .IN1(n9138), .IN2(n12690), .IN3(n12691), .QN(WX5143) );
  NOR2X0 U12886 ( .IN1(n8131), .IN2(CRC_OUT_6_31), .QN(n12691) );
  NOR2X0 U12887 ( .IN1(DFF_767_n1), .IN2(WX4778), .QN(n12690) );
  NOR2X0 U12888 ( .IN1(n16351), .IN2(n9162), .QN(WX4617) );
  NOR2X0 U12889 ( .IN1(n9237), .IN2(n8823), .QN(WX4615) );
  NOR2X0 U12890 ( .IN1(n16350), .IN2(n9162), .QN(WX4613) );
  NOR2X0 U12891 ( .IN1(n16349), .IN2(n9162), .QN(WX4611) );
  NOR2X0 U12892 ( .IN1(n16348), .IN2(n9162), .QN(WX4609) );
  NOR2X0 U12893 ( .IN1(n16347), .IN2(n9162), .QN(WX4607) );
  NOR2X0 U12894 ( .IN1(n16346), .IN2(n9161), .QN(WX4605) );
  NOR2X0 U12895 ( .IN1(n16345), .IN2(n9161), .QN(WX4603) );
  NOR2X0 U12896 ( .IN1(n16344), .IN2(n9161), .QN(WX4601) );
  NOR2X0 U12897 ( .IN1(n16343), .IN2(n9161), .QN(WX4599) );
  NOR2X0 U12898 ( .IN1(n16342), .IN2(n9161), .QN(WX4597) );
  NOR2X0 U12899 ( .IN1(n16341), .IN2(n9161), .QN(WX4595) );
  NOR2X0 U12900 ( .IN1(n16340), .IN2(n9161), .QN(WX4593) );
  NOR2X0 U12901 ( .IN1(n16339), .IN2(n9161), .QN(WX4591) );
  NOR2X0 U12902 ( .IN1(n16338), .IN2(n9161), .QN(WX4589) );
  NOR2X0 U12903 ( .IN1(n16337), .IN2(n9161), .QN(WX4587) );
  NAND4X0 U12904 ( .IN1(n12692), .IN2(n12693), .IN3(n12694), .IN4(n12695), 
        .QN(WX4585) );
  NAND3X0 U12905 ( .IN1(n12696), .IN2(n12697), .IN3(n9090), .QN(n12695) );
  NAND2X0 U12906 ( .IN1(n9324), .IN2(n12023), .QN(n12694) );
  NAND2X0 U12907 ( .IN1(n12698), .IN2(n12699), .QN(n12023) );
  INVX0 U12908 ( .INP(n12700), .ZN(n12699) );
  NOR2X0 U12909 ( .IN1(n12701), .IN2(n12702), .QN(n12700) );
  NAND2X0 U12910 ( .IN1(n12702), .IN2(n12701), .QN(n12698) );
  NOR2X0 U12911 ( .IN1(n12703), .IN2(n12704), .QN(n12701) );
  NOR2X0 U12912 ( .IN1(WX6071), .IN2(n7976), .QN(n12704) );
  INVX0 U12913 ( .INP(n12705), .ZN(n12703) );
  NAND2X0 U12914 ( .IN1(n7976), .IN2(WX6071), .QN(n12705) );
  NAND2X0 U12915 ( .IN1(n12706), .IN2(n12707), .QN(n12702) );
  NAND2X0 U12916 ( .IN1(n7975), .IN2(WX5943), .QN(n12707) );
  INVX0 U12917 ( .INP(n12708), .ZN(n12706) );
  NOR2X0 U12918 ( .IN1(WX5943), .IN2(n7975), .QN(n12708) );
  NAND2X0 U12919 ( .IN1(n765), .IN2(n9282), .QN(n12693) );
  NOR2X0 U12920 ( .IN1(n9232), .IN2(n8945), .QN(n765) );
  NAND2X0 U12921 ( .IN1(n9293), .IN2(CRC_OUT_6_0), .QN(n12692) );
  NAND4X0 U12922 ( .IN1(n12709), .IN2(n12710), .IN3(n12711), .IN4(n12712), 
        .QN(WX4583) );
  NAND3X0 U12923 ( .IN1(n12028), .IN2(n12029), .IN3(n9322), .QN(n12712) );
  NAND3X0 U12924 ( .IN1(n12713), .IN2(n12714), .IN3(n12715), .QN(n12029) );
  INVX0 U12925 ( .INP(n12716), .ZN(n12715) );
  NAND2X0 U12926 ( .IN1(n12716), .IN2(n12717), .QN(n12028) );
  NAND2X0 U12927 ( .IN1(n12713), .IN2(n12714), .QN(n12717) );
  NAND2X0 U12928 ( .IN1(n8354), .IN2(WX5941), .QN(n12714) );
  NAND2X0 U12929 ( .IN1(n3661), .IN2(WX6069), .QN(n12713) );
  NOR2X0 U12930 ( .IN1(n12718), .IN2(n12719), .QN(n12716) );
  INVX0 U12931 ( .INP(n12720), .ZN(n12719) );
  NAND2X0 U12932 ( .IN1(test_so51), .IN2(WX5877), .QN(n12720) );
  NOR2X0 U12933 ( .IN1(WX5877), .IN2(test_so51), .QN(n12718) );
  NAND2X0 U12934 ( .IN1(n9107), .IN2(n12721), .QN(n12711) );
  NAND2X0 U12935 ( .IN1(n764), .IN2(n9282), .QN(n12710) );
  NOR2X0 U12936 ( .IN1(n9232), .IN2(n8946), .QN(n764) );
  NAND2X0 U12937 ( .IN1(n9293), .IN2(CRC_OUT_6_1), .QN(n12709) );
  NAND4X0 U12938 ( .IN1(n12722), .IN2(n12723), .IN3(n12724), .IN4(n12725), 
        .QN(WX4581) );
  NAND2X0 U12939 ( .IN1(n9324), .IN2(n12056), .QN(n12725) );
  NAND2X0 U12940 ( .IN1(n12726), .IN2(n12727), .QN(n12056) );
  INVX0 U12941 ( .INP(n12728), .ZN(n12727) );
  NOR2X0 U12942 ( .IN1(n12729), .IN2(n12730), .QN(n12728) );
  NAND2X0 U12943 ( .IN1(n12730), .IN2(n12729), .QN(n12726) );
  NOR2X0 U12944 ( .IN1(n12731), .IN2(n12732), .QN(n12729) );
  NOR2X0 U12945 ( .IN1(WX6067), .IN2(n7979), .QN(n12732) );
  INVX0 U12946 ( .INP(n12733), .ZN(n12731) );
  NAND2X0 U12947 ( .IN1(n7979), .IN2(WX6067), .QN(n12733) );
  NAND2X0 U12948 ( .IN1(n12734), .IN2(n12735), .QN(n12730) );
  NAND2X0 U12949 ( .IN1(n7978), .IN2(WX5939), .QN(n12735) );
  INVX0 U12950 ( .INP(n12736), .ZN(n12734) );
  NOR2X0 U12951 ( .IN1(WX5939), .IN2(n7978), .QN(n12736) );
  NAND2X0 U12952 ( .IN1(n9107), .IN2(n12737), .QN(n12724) );
  NAND2X0 U12953 ( .IN1(n763), .IN2(n9282), .QN(n12723) );
  NOR2X0 U12954 ( .IN1(n9069), .IN2(n9161), .QN(n763) );
  NAND2X0 U12955 ( .IN1(n9293), .IN2(CRC_OUT_6_2), .QN(n12722) );
  NAND4X0 U12956 ( .IN1(n12738), .IN2(n12739), .IN3(n12740), .IN4(n12741), 
        .QN(WX4579) );
  NAND3X0 U12957 ( .IN1(n12061), .IN2(n12062), .IN3(n9321), .QN(n12741) );
  NAND3X0 U12958 ( .IN1(n12742), .IN2(n12743), .IN3(n12744), .QN(n12062) );
  INVX0 U12959 ( .INP(n12745), .ZN(n12744) );
  NAND2X0 U12960 ( .IN1(n12745), .IN2(n12746), .QN(n12061) );
  NAND2X0 U12961 ( .IN1(n12742), .IN2(n12743), .QN(n12746) );
  NAND2X0 U12962 ( .IN1(n8344), .IN2(WX6001), .QN(n12743) );
  NAND2X0 U12963 ( .IN1(n7981), .IN2(WX6065), .QN(n12742) );
  NOR2X0 U12964 ( .IN1(n12747), .IN2(n12748), .QN(n12745) );
  INVX0 U12965 ( .INP(n12749), .ZN(n12748) );
  NAND2X0 U12966 ( .IN1(test_so49), .IN2(WX5873), .QN(n12749) );
  NOR2X0 U12967 ( .IN1(WX5873), .IN2(test_so49), .QN(n12747) );
  NAND2X0 U12968 ( .IN1(n9107), .IN2(n12750), .QN(n12740) );
  NAND2X0 U12969 ( .IN1(n762), .IN2(n9282), .QN(n12739) );
  NOR2X0 U12970 ( .IN1(n9232), .IN2(n8947), .QN(n762) );
  NAND2X0 U12971 ( .IN1(n9293), .IN2(CRC_OUT_6_3), .QN(n12738) );
  NAND4X0 U12972 ( .IN1(n12751), .IN2(n12752), .IN3(n12753), .IN4(n12754), 
        .QN(WX4577) );
  NAND2X0 U12973 ( .IN1(n9324), .IN2(n12086), .QN(n12754) );
  NAND2X0 U12974 ( .IN1(n12755), .IN2(n12756), .QN(n12086) );
  INVX0 U12975 ( .INP(n12757), .ZN(n12756) );
  NOR2X0 U12976 ( .IN1(n12758), .IN2(n12759), .QN(n12757) );
  NAND2X0 U12977 ( .IN1(n12759), .IN2(n12758), .QN(n12755) );
  NOR2X0 U12978 ( .IN1(n12760), .IN2(n12761), .QN(n12758) );
  NOR2X0 U12979 ( .IN1(WX6063), .IN2(n7983), .QN(n12761) );
  INVX0 U12980 ( .INP(n12762), .ZN(n12760) );
  NAND2X0 U12981 ( .IN1(n7983), .IN2(WX6063), .QN(n12762) );
  NAND2X0 U12982 ( .IN1(n12763), .IN2(n12764), .QN(n12759) );
  NAND2X0 U12983 ( .IN1(n7982), .IN2(WX5935), .QN(n12764) );
  INVX0 U12984 ( .INP(n12765), .ZN(n12763) );
  NOR2X0 U12985 ( .IN1(WX5935), .IN2(n7982), .QN(n12765) );
  NAND2X0 U12986 ( .IN1(n9107), .IN2(n12766), .QN(n12753) );
  NAND2X0 U12987 ( .IN1(n761), .IN2(n9282), .QN(n12752) );
  NOR2X0 U12988 ( .IN1(n9232), .IN2(n8948), .QN(n761) );
  NAND2X0 U12989 ( .IN1(n9293), .IN2(CRC_OUT_6_4), .QN(n12751) );
  NAND4X0 U12990 ( .IN1(n12767), .IN2(n12768), .IN3(n12769), .IN4(n12770), 
        .QN(WX4575) );
  NAND3X0 U12991 ( .IN1(n12091), .IN2(n12092), .IN3(n9322), .QN(n12770) );
  NAND3X0 U12992 ( .IN1(n12771), .IN2(n12772), .IN3(n12773), .QN(n12092) );
  INVX0 U12993 ( .INP(n12774), .ZN(n12773) );
  NAND2X0 U12994 ( .IN1(n12774), .IN2(n12775), .QN(n12091) );
  NAND2X0 U12995 ( .IN1(n12771), .IN2(n12772), .QN(n12775) );
  NAND2X0 U12996 ( .IN1(n8327), .IN2(WX5933), .QN(n12772) );
  NAND2X0 U12997 ( .IN1(n3669), .IN2(WX6061), .QN(n12771) );
  NOR2X0 U12998 ( .IN1(n12776), .IN2(n12777), .QN(n12774) );
  INVX0 U12999 ( .INP(n12778), .ZN(n12777) );
  NAND2X0 U13000 ( .IN1(test_so47), .IN2(WX5997), .QN(n12778) );
  NOR2X0 U13001 ( .IN1(WX5997), .IN2(test_so47), .QN(n12776) );
  NAND2X0 U13002 ( .IN1(n9107), .IN2(n12779), .QN(n12769) );
  NAND2X0 U13003 ( .IN1(n760), .IN2(n9282), .QN(n12768) );
  NOR2X0 U13004 ( .IN1(n9232), .IN2(n8949), .QN(n760) );
  NAND2X0 U13005 ( .IN1(test_so42), .IN2(n9315), .QN(n12767) );
  NAND4X0 U13006 ( .IN1(n12780), .IN2(n12781), .IN3(n12782), .IN4(n12783), 
        .QN(WX4573) );
  NAND2X0 U13007 ( .IN1(n9325), .IN2(n12116), .QN(n12783) );
  NAND2X0 U13008 ( .IN1(n12784), .IN2(n12785), .QN(n12116) );
  INVX0 U13009 ( .INP(n12786), .ZN(n12785) );
  NOR2X0 U13010 ( .IN1(n12787), .IN2(n12788), .QN(n12786) );
  NAND2X0 U13011 ( .IN1(n12788), .IN2(n12787), .QN(n12784) );
  NOR2X0 U13012 ( .IN1(n12789), .IN2(n12790), .QN(n12787) );
  NOR2X0 U13013 ( .IN1(WX6059), .IN2(n7986), .QN(n12790) );
  INVX0 U13014 ( .INP(n12791), .ZN(n12789) );
  NAND2X0 U13015 ( .IN1(n7986), .IN2(WX6059), .QN(n12791) );
  NAND2X0 U13016 ( .IN1(n12792), .IN2(n12793), .QN(n12788) );
  NAND2X0 U13017 ( .IN1(n7985), .IN2(WX5931), .QN(n12793) );
  INVX0 U13018 ( .INP(n12794), .ZN(n12792) );
  NOR2X0 U13019 ( .IN1(WX5931), .IN2(n7985), .QN(n12794) );
  NAND2X0 U13020 ( .IN1(n9107), .IN2(n12795), .QN(n12782) );
  NAND2X0 U13021 ( .IN1(n759), .IN2(n9282), .QN(n12781) );
  NOR2X0 U13022 ( .IN1(n9232), .IN2(n8950), .QN(n759) );
  NAND2X0 U13023 ( .IN1(n9294), .IN2(CRC_OUT_6_6), .QN(n12780) );
  NAND4X0 U13024 ( .IN1(n12796), .IN2(n12797), .IN3(n12798), .IN4(n12799), 
        .QN(WX4571) );
  NAND2X0 U13025 ( .IN1(n9324), .IN2(n12132), .QN(n12799) );
  NAND2X0 U13026 ( .IN1(n12800), .IN2(n12801), .QN(n12132) );
  INVX0 U13027 ( .INP(n12802), .ZN(n12801) );
  NOR2X0 U13028 ( .IN1(n12803), .IN2(n12804), .QN(n12802) );
  NAND2X0 U13029 ( .IN1(n12804), .IN2(n12803), .QN(n12800) );
  NOR2X0 U13030 ( .IN1(n12805), .IN2(n12806), .QN(n12803) );
  NOR2X0 U13031 ( .IN1(WX6057), .IN2(n7988), .QN(n12806) );
  INVX0 U13032 ( .INP(n12807), .ZN(n12805) );
  NAND2X0 U13033 ( .IN1(n7988), .IN2(WX6057), .QN(n12807) );
  NAND2X0 U13034 ( .IN1(n12808), .IN2(n12809), .QN(n12804) );
  NAND2X0 U13035 ( .IN1(n7987), .IN2(WX5929), .QN(n12809) );
  INVX0 U13036 ( .INP(n12810), .ZN(n12808) );
  NOR2X0 U13037 ( .IN1(WX5929), .IN2(n7987), .QN(n12810) );
  NAND2X0 U13038 ( .IN1(n9107), .IN2(n12811), .QN(n12798) );
  NAND2X0 U13039 ( .IN1(n758), .IN2(n9282), .QN(n12797) );
  NOR2X0 U13040 ( .IN1(n9232), .IN2(n8951), .QN(n758) );
  NAND2X0 U13041 ( .IN1(n9294), .IN2(CRC_OUT_6_7), .QN(n12796) );
  NAND4X0 U13042 ( .IN1(n12812), .IN2(n12813), .IN3(n12814), .IN4(n12815), 
        .QN(WX4569) );
  NAND2X0 U13043 ( .IN1(n9324), .IN2(n12145), .QN(n12815) );
  NAND2X0 U13044 ( .IN1(n12816), .IN2(n12817), .QN(n12145) );
  INVX0 U13045 ( .INP(n12818), .ZN(n12817) );
  NOR2X0 U13046 ( .IN1(n12819), .IN2(n12820), .QN(n12818) );
  NAND2X0 U13047 ( .IN1(n12820), .IN2(n12819), .QN(n12816) );
  NOR2X0 U13048 ( .IN1(n12821), .IN2(n12822), .QN(n12819) );
  NOR2X0 U13049 ( .IN1(WX6055), .IN2(n7990), .QN(n12822) );
  INVX0 U13050 ( .INP(n12823), .ZN(n12821) );
  NAND2X0 U13051 ( .IN1(n7990), .IN2(WX6055), .QN(n12823) );
  NAND2X0 U13052 ( .IN1(n12824), .IN2(n12825), .QN(n12820) );
  NAND2X0 U13053 ( .IN1(n7989), .IN2(WX5927), .QN(n12825) );
  INVX0 U13054 ( .INP(n12826), .ZN(n12824) );
  NOR2X0 U13055 ( .IN1(WX5927), .IN2(n7989), .QN(n12826) );
  NAND2X0 U13056 ( .IN1(n9107), .IN2(n12827), .QN(n12814) );
  NAND2X0 U13057 ( .IN1(n757), .IN2(n9282), .QN(n12813) );
  NOR2X0 U13058 ( .IN1(n9233), .IN2(n8952), .QN(n757) );
  NAND2X0 U13059 ( .IN1(n9294), .IN2(CRC_OUT_6_8), .QN(n12812) );
  NAND4X0 U13060 ( .IN1(n12828), .IN2(n12829), .IN3(n12830), .IN4(n12831), 
        .QN(WX4567) );
  NAND2X0 U13061 ( .IN1(n9324), .IN2(n12161), .QN(n12831) );
  NAND2X0 U13062 ( .IN1(n12832), .IN2(n12833), .QN(n12161) );
  INVX0 U13063 ( .INP(n12834), .ZN(n12833) );
  NOR2X0 U13064 ( .IN1(n12835), .IN2(n12836), .QN(n12834) );
  NAND2X0 U13065 ( .IN1(n12836), .IN2(n12835), .QN(n12832) );
  NOR2X0 U13066 ( .IN1(n12837), .IN2(n12838), .QN(n12835) );
  NOR2X0 U13067 ( .IN1(WX6053), .IN2(n7992), .QN(n12838) );
  INVX0 U13068 ( .INP(n12839), .ZN(n12837) );
  NAND2X0 U13069 ( .IN1(n7992), .IN2(WX6053), .QN(n12839) );
  NAND2X0 U13070 ( .IN1(n12840), .IN2(n12841), .QN(n12836) );
  NAND2X0 U13071 ( .IN1(n7991), .IN2(WX5925), .QN(n12841) );
  INVX0 U13072 ( .INP(n12842), .ZN(n12840) );
  NOR2X0 U13073 ( .IN1(WX5925), .IN2(n7991), .QN(n12842) );
  NAND2X0 U13074 ( .IN1(n9107), .IN2(n12843), .QN(n12830) );
  NAND2X0 U13075 ( .IN1(n756), .IN2(n9282), .QN(n12829) );
  NOR2X0 U13076 ( .IN1(n9233), .IN2(n8953), .QN(n756) );
  NAND2X0 U13077 ( .IN1(n9294), .IN2(CRC_OUT_6_9), .QN(n12828) );
  NAND4X0 U13078 ( .IN1(n12844), .IN2(n12845), .IN3(n12846), .IN4(n12847), 
        .QN(WX4565) );
  NAND2X0 U13079 ( .IN1(n9325), .IN2(n12174), .QN(n12847) );
  NAND2X0 U13080 ( .IN1(n12848), .IN2(n12849), .QN(n12174) );
  INVX0 U13081 ( .INP(n12850), .ZN(n12849) );
  NOR2X0 U13082 ( .IN1(n12851), .IN2(n12852), .QN(n12850) );
  NAND2X0 U13083 ( .IN1(n12852), .IN2(n12851), .QN(n12848) );
  NOR2X0 U13084 ( .IN1(n12853), .IN2(n12854), .QN(n12851) );
  NOR2X0 U13085 ( .IN1(WX6051), .IN2(n7994), .QN(n12854) );
  INVX0 U13086 ( .INP(n12855), .ZN(n12853) );
  NAND2X0 U13087 ( .IN1(n7994), .IN2(WX6051), .QN(n12855) );
  NAND2X0 U13088 ( .IN1(n12856), .IN2(n12857), .QN(n12852) );
  NAND2X0 U13089 ( .IN1(n7993), .IN2(WX5923), .QN(n12857) );
  INVX0 U13090 ( .INP(n12858), .ZN(n12856) );
  NOR2X0 U13091 ( .IN1(WX5923), .IN2(n7993), .QN(n12858) );
  NAND2X0 U13092 ( .IN1(n9107), .IN2(n12859), .QN(n12846) );
  NAND2X0 U13093 ( .IN1(n755), .IN2(n9282), .QN(n12845) );
  NOR2X0 U13094 ( .IN1(n9233), .IN2(n8954), .QN(n755) );
  NAND2X0 U13095 ( .IN1(n9294), .IN2(CRC_OUT_6_10), .QN(n12844) );
  NAND4X0 U13096 ( .IN1(n12860), .IN2(n12861), .IN3(n12862), .IN4(n12863), 
        .QN(WX4563) );
  NAND3X0 U13097 ( .IN1(n12864), .IN2(n12865), .IN3(n9091), .QN(n12863) );
  NAND2X0 U13098 ( .IN1(n9325), .IN2(n12190), .QN(n12862) );
  NAND2X0 U13099 ( .IN1(n12866), .IN2(n12867), .QN(n12190) );
  INVX0 U13100 ( .INP(n12868), .ZN(n12867) );
  NOR2X0 U13101 ( .IN1(n12869), .IN2(n12870), .QN(n12868) );
  NAND2X0 U13102 ( .IN1(n12870), .IN2(n12869), .QN(n12866) );
  NOR2X0 U13103 ( .IN1(n12871), .IN2(n12872), .QN(n12869) );
  NOR2X0 U13104 ( .IN1(WX6049), .IN2(n7996), .QN(n12872) );
  INVX0 U13105 ( .INP(n12873), .ZN(n12871) );
  NAND2X0 U13106 ( .IN1(n7996), .IN2(WX6049), .QN(n12873) );
  NAND2X0 U13107 ( .IN1(n12874), .IN2(n12875), .QN(n12870) );
  NAND2X0 U13108 ( .IN1(n7995), .IN2(WX5921), .QN(n12875) );
  INVX0 U13109 ( .INP(n12876), .ZN(n12874) );
  NOR2X0 U13110 ( .IN1(WX5921), .IN2(n7995), .QN(n12876) );
  NAND2X0 U13111 ( .IN1(n754), .IN2(n9282), .QN(n12861) );
  NOR2X0 U13112 ( .IN1(n9233), .IN2(n8955), .QN(n754) );
  NAND2X0 U13113 ( .IN1(n9294), .IN2(CRC_OUT_6_11), .QN(n12860) );
  NAND4X0 U13114 ( .IN1(n12877), .IN2(n12878), .IN3(n12879), .IN4(n12880), 
        .QN(WX4561) );
  NAND2X0 U13115 ( .IN1(n9325), .IN2(n12206), .QN(n12880) );
  NAND2X0 U13116 ( .IN1(n12881), .IN2(n12882), .QN(n12206) );
  INVX0 U13117 ( .INP(n12883), .ZN(n12882) );
  NOR2X0 U13118 ( .IN1(n12884), .IN2(n12885), .QN(n12883) );
  NAND2X0 U13119 ( .IN1(n12885), .IN2(n12884), .QN(n12881) );
  NOR2X0 U13120 ( .IN1(n12886), .IN2(n12887), .QN(n12884) );
  NOR2X0 U13121 ( .IN1(WX6047), .IN2(n7998), .QN(n12887) );
  INVX0 U13122 ( .INP(n12888), .ZN(n12886) );
  NAND2X0 U13123 ( .IN1(n7998), .IN2(WX6047), .QN(n12888) );
  NAND2X0 U13124 ( .IN1(n12889), .IN2(n12890), .QN(n12885) );
  NAND2X0 U13125 ( .IN1(n7997), .IN2(WX5919), .QN(n12890) );
  INVX0 U13126 ( .INP(n12891), .ZN(n12889) );
  NOR2X0 U13127 ( .IN1(WX5919), .IN2(n7997), .QN(n12891) );
  NAND2X0 U13128 ( .IN1(n9107), .IN2(n12892), .QN(n12879) );
  NAND2X0 U13129 ( .IN1(n753), .IN2(n9282), .QN(n12878) );
  NOR2X0 U13130 ( .IN1(n9233), .IN2(n8956), .QN(n753) );
  NAND2X0 U13131 ( .IN1(n9294), .IN2(CRC_OUT_6_12), .QN(n12877) );
  NAND4X0 U13132 ( .IN1(n12893), .IN2(n12894), .IN3(n12895), .IN4(n12896), 
        .QN(WX4559) );
  NAND3X0 U13133 ( .IN1(n12897), .IN2(n12898), .IN3(n9091), .QN(n12896) );
  NAND2X0 U13134 ( .IN1(n9325), .IN2(n12222), .QN(n12895) );
  NAND2X0 U13135 ( .IN1(n12899), .IN2(n12900), .QN(n12222) );
  INVX0 U13136 ( .INP(n12901), .ZN(n12900) );
  NOR2X0 U13137 ( .IN1(n12902), .IN2(n12903), .QN(n12901) );
  NAND2X0 U13138 ( .IN1(n12903), .IN2(n12902), .QN(n12899) );
  NOR2X0 U13139 ( .IN1(n12904), .IN2(n12905), .QN(n12902) );
  NOR2X0 U13140 ( .IN1(WX6045), .IN2(n8000), .QN(n12905) );
  INVX0 U13141 ( .INP(n12906), .ZN(n12904) );
  NAND2X0 U13142 ( .IN1(n8000), .IN2(WX6045), .QN(n12906) );
  NAND2X0 U13143 ( .IN1(n12907), .IN2(n12908), .QN(n12903) );
  NAND2X0 U13144 ( .IN1(n7999), .IN2(WX5917), .QN(n12908) );
  INVX0 U13145 ( .INP(n12909), .ZN(n12907) );
  NOR2X0 U13146 ( .IN1(WX5917), .IN2(n7999), .QN(n12909) );
  NAND2X0 U13147 ( .IN1(n752), .IN2(n9282), .QN(n12894) );
  NOR2X0 U13148 ( .IN1(n9233), .IN2(n8957), .QN(n752) );
  NAND2X0 U13149 ( .IN1(n9294), .IN2(CRC_OUT_6_13), .QN(n12893) );
  NAND4X0 U13150 ( .IN1(n12910), .IN2(n12911), .IN3(n12912), .IN4(n12913), 
        .QN(WX4557) );
  NAND2X0 U13151 ( .IN1(n9325), .IN2(n12238), .QN(n12913) );
  NAND2X0 U13152 ( .IN1(n12914), .IN2(n12915), .QN(n12238) );
  INVX0 U13153 ( .INP(n12916), .ZN(n12915) );
  NOR2X0 U13154 ( .IN1(n12917), .IN2(n12918), .QN(n12916) );
  NAND2X0 U13155 ( .IN1(n12918), .IN2(n12917), .QN(n12914) );
  NOR2X0 U13156 ( .IN1(n12919), .IN2(n12920), .QN(n12917) );
  NOR2X0 U13157 ( .IN1(WX6043), .IN2(n8002), .QN(n12920) );
  INVX0 U13158 ( .INP(n12921), .ZN(n12919) );
  NAND2X0 U13159 ( .IN1(n8002), .IN2(WX6043), .QN(n12921) );
  NAND2X0 U13160 ( .IN1(n12922), .IN2(n12923), .QN(n12918) );
  NAND2X0 U13161 ( .IN1(n8001), .IN2(WX5915), .QN(n12923) );
  INVX0 U13162 ( .INP(n12924), .ZN(n12922) );
  NOR2X0 U13163 ( .IN1(WX5915), .IN2(n8001), .QN(n12924) );
  NAND2X0 U13164 ( .IN1(n9107), .IN2(n12925), .QN(n12912) );
  NAND2X0 U13165 ( .IN1(n751), .IN2(n9283), .QN(n12911) );
  NOR2X0 U13166 ( .IN1(n9233), .IN2(n8958), .QN(n751) );
  NAND2X0 U13167 ( .IN1(n9294), .IN2(CRC_OUT_6_14), .QN(n12910) );
  NAND4X0 U13168 ( .IN1(n12926), .IN2(n12927), .IN3(n12928), .IN4(n12929), 
        .QN(WX4555) );
  NAND3X0 U13169 ( .IN1(n12930), .IN2(n12931), .IN3(n9091), .QN(n12929) );
  NAND2X0 U13170 ( .IN1(n9325), .IN2(n12254), .QN(n12928) );
  NAND2X0 U13171 ( .IN1(n12932), .IN2(n12933), .QN(n12254) );
  INVX0 U13172 ( .INP(n12934), .ZN(n12933) );
  NOR2X0 U13173 ( .IN1(n12935), .IN2(n12936), .QN(n12934) );
  NAND2X0 U13174 ( .IN1(n12936), .IN2(n12935), .QN(n12932) );
  NOR2X0 U13175 ( .IN1(n12937), .IN2(n12938), .QN(n12935) );
  NOR2X0 U13176 ( .IN1(WX6041), .IN2(n8004), .QN(n12938) );
  INVX0 U13177 ( .INP(n12939), .ZN(n12937) );
  NAND2X0 U13178 ( .IN1(n8004), .IN2(WX6041), .QN(n12939) );
  NAND2X0 U13179 ( .IN1(n12940), .IN2(n12941), .QN(n12936) );
  NAND2X0 U13180 ( .IN1(n8003), .IN2(WX5913), .QN(n12941) );
  INVX0 U13181 ( .INP(n12942), .ZN(n12940) );
  NOR2X0 U13182 ( .IN1(WX5913), .IN2(n8003), .QN(n12942) );
  NAND2X0 U13183 ( .IN1(n750), .IN2(n9283), .QN(n12927) );
  NOR2X0 U13184 ( .IN1(n9233), .IN2(n8959), .QN(n750) );
  NAND2X0 U13185 ( .IN1(n9294), .IN2(CRC_OUT_6_15), .QN(n12926) );
  NAND4X0 U13186 ( .IN1(n12943), .IN2(n12944), .IN3(n12945), .IN4(n12946), 
        .QN(WX4553) );
  NAND2X0 U13187 ( .IN1(n12947), .IN2(n12948), .QN(n12946) );
  NAND2X0 U13188 ( .IN1(n12949), .IN2(n12950), .QN(n12947) );
  NAND2X0 U13189 ( .IN1(n9107), .IN2(n12951), .QN(n12950) );
  NAND2X0 U13190 ( .IN1(n9108), .IN2(n8537), .QN(n12949) );
  NAND2X0 U13191 ( .IN1(n12273), .IN2(n2153), .QN(n12945) );
  NOR2X0 U13192 ( .IN1(n12952), .IN2(n12953), .QN(n12273) );
  INVX0 U13193 ( .INP(n12954), .ZN(n12953) );
  NAND2X0 U13194 ( .IN1(n12955), .IN2(n12956), .QN(n12954) );
  NOR2X0 U13195 ( .IN1(n12956), .IN2(n12955), .QN(n12952) );
  NAND2X0 U13196 ( .IN1(n12957), .IN2(n12958), .QN(n12955) );
  NAND2X0 U13197 ( .IN1(n12959), .IN2(WX5975), .QN(n12958) );
  NAND2X0 U13198 ( .IN1(n12960), .IN2(n12961), .QN(n12959) );
  NAND3X0 U13199 ( .IN1(n12960), .IN2(n12961), .IN3(n7741), .QN(n12957) );
  NAND2X0 U13200 ( .IN1(test_so52), .IN2(WX5911), .QN(n12961) );
  NAND2X0 U13201 ( .IN1(n7740), .IN2(n8827), .QN(n12960) );
  NOR2X0 U13202 ( .IN1(n12962), .IN2(n12963), .QN(n12956) );
  INVX0 U13203 ( .INP(n12964), .ZN(n12963) );
  NAND2X0 U13204 ( .IN1(n16366), .IN2(n9118), .QN(n12964) );
  NOR2X0 U13205 ( .IN1(n9117), .IN2(n16366), .QN(n12962) );
  NAND2X0 U13206 ( .IN1(n749), .IN2(n9283), .QN(n12944) );
  NOR2X0 U13207 ( .IN1(n9233), .IN2(n8960), .QN(n749) );
  NAND2X0 U13208 ( .IN1(n9294), .IN2(CRC_OUT_6_16), .QN(n12943) );
  NAND4X0 U13209 ( .IN1(n12965), .IN2(n12966), .IN3(n12967), .IN4(n12968), 
        .QN(WX4551) );
  NAND2X0 U13210 ( .IN1(n12969), .IN2(n12293), .QN(n12968) );
  NAND2X0 U13211 ( .IN1(n12970), .IN2(n12296), .QN(n12293) );
  NAND2X0 U13212 ( .IN1(n12971), .IN2(n12972), .QN(n12970) );
  NAND2X0 U13213 ( .IN1(n16365), .IN2(n9118), .QN(n12972) );
  NAND2X0 U13214 ( .IN1(TM1), .IN2(n8480), .QN(n12971) );
  NAND3X0 U13215 ( .IN1(n12973), .IN2(n12974), .IN3(n12975), .QN(n12969) );
  NAND2X0 U13216 ( .IN1(n9325), .IN2(n12296), .QN(n12975) );
  NAND2X0 U13217 ( .IN1(n12976), .IN2(n12977), .QN(n12296) );
  NAND2X0 U13218 ( .IN1(n7742), .IN2(n12978), .QN(n12977) );
  INVX0 U13219 ( .INP(n12979), .ZN(n12976) );
  NOR2X0 U13220 ( .IN1(n12978), .IN2(n7742), .QN(n12979) );
  NOR2X0 U13221 ( .IN1(n12980), .IN2(n12981), .QN(n12978) );
  NOR2X0 U13222 ( .IN1(WX6037), .IN2(n7743), .QN(n12981) );
  INVX0 U13223 ( .INP(n12982), .ZN(n12980) );
  NAND2X0 U13224 ( .IN1(n7743), .IN2(WX6037), .QN(n12982) );
  NAND2X0 U13225 ( .IN1(n9082), .IN2(n8480), .QN(n12974) );
  NAND2X0 U13226 ( .IN1(n16365), .IN2(n9079), .QN(n12973) );
  NAND2X0 U13227 ( .IN1(n12983), .IN2(n12984), .QN(n12967) );
  NAND2X0 U13228 ( .IN1(n12985), .IN2(n12986), .QN(n12983) );
  NAND2X0 U13229 ( .IN1(n9108), .IN2(n12987), .QN(n12986) );
  NAND2X0 U13230 ( .IN1(n8413), .IN2(n9111), .QN(n12985) );
  NAND2X0 U13231 ( .IN1(n748), .IN2(n9283), .QN(n12966) );
  NOR2X0 U13232 ( .IN1(n9233), .IN2(n8961), .QN(n748) );
  NAND2X0 U13233 ( .IN1(n9294), .IN2(CRC_OUT_6_17), .QN(n12965) );
  NAND4X0 U13234 ( .IN1(n12988), .IN2(n12989), .IN3(n12990), .IN4(n12991), 
        .QN(WX4549) );
  NAND2X0 U13235 ( .IN1(n12992), .IN2(n12993), .QN(n12991) );
  NAND2X0 U13236 ( .IN1(n12994), .IN2(n12995), .QN(n12992) );
  NAND2X0 U13237 ( .IN1(n9108), .IN2(n12996), .QN(n12995) );
  NAND2X0 U13238 ( .IN1(n9108), .IN2(n8540), .QN(n12994) );
  NAND2X0 U13239 ( .IN1(n12315), .IN2(n2153), .QN(n12990) );
  NOR2X0 U13240 ( .IN1(n12997), .IN2(n12998), .QN(n12315) );
  INVX0 U13241 ( .INP(n12999), .ZN(n12998) );
  NAND2X0 U13242 ( .IN1(n13000), .IN2(n13001), .QN(n12999) );
  NOR2X0 U13243 ( .IN1(n13001), .IN2(n13000), .QN(n12997) );
  NAND2X0 U13244 ( .IN1(n13002), .IN2(n13003), .QN(n13000) );
  NAND2X0 U13245 ( .IN1(n8296), .IN2(n13004), .QN(n13003) );
  INVX0 U13246 ( .INP(n13005), .ZN(n13004) );
  NAND2X0 U13247 ( .IN1(n13005), .IN2(WX6035), .QN(n13002) );
  NAND2X0 U13248 ( .IN1(n13006), .IN2(n13007), .QN(n13005) );
  INVX0 U13249 ( .INP(n13008), .ZN(n13007) );
  NOR2X0 U13250 ( .IN1(n8812), .IN2(n16364), .QN(n13008) );
  NAND2X0 U13251 ( .IN1(n16364), .IN2(n8812), .QN(n13006) );
  NOR2X0 U13252 ( .IN1(n13009), .IN2(n13010), .QN(n13001) );
  INVX0 U13253 ( .INP(n13011), .ZN(n13010) );
  NAND2X0 U13254 ( .IN1(n7744), .IN2(n9118), .QN(n13011) );
  NOR2X0 U13255 ( .IN1(n9116), .IN2(n7744), .QN(n13009) );
  NAND2X0 U13256 ( .IN1(n747), .IN2(n9283), .QN(n12989) );
  NOR2X0 U13257 ( .IN1(n9233), .IN2(n8962), .QN(n747) );
  NAND2X0 U13258 ( .IN1(n9295), .IN2(CRC_OUT_6_18), .QN(n12988) );
  NAND4X0 U13259 ( .IN1(n13012), .IN2(n13013), .IN3(n13014), .IN4(n13015), 
        .QN(WX4547) );
  NAND2X0 U13260 ( .IN1(n13016), .IN2(n12335), .QN(n13015) );
  NAND2X0 U13261 ( .IN1(n13017), .IN2(n12338), .QN(n12335) );
  NAND2X0 U13262 ( .IN1(n13018), .IN2(n13019), .QN(n13017) );
  NAND2X0 U13263 ( .IN1(n16363), .IN2(n9119), .QN(n13019) );
  NAND2X0 U13264 ( .IN1(TM1), .IN2(n8482), .QN(n13018) );
  NAND3X0 U13265 ( .IN1(n13020), .IN2(n13021), .IN3(n13022), .QN(n13016) );
  NAND2X0 U13266 ( .IN1(n9325), .IN2(n12338), .QN(n13022) );
  NAND2X0 U13267 ( .IN1(n13023), .IN2(n13024), .QN(n12338) );
  NAND2X0 U13268 ( .IN1(n7745), .IN2(n13025), .QN(n13024) );
  INVX0 U13269 ( .INP(n13026), .ZN(n13023) );
  NOR2X0 U13270 ( .IN1(n13025), .IN2(n7745), .QN(n13026) );
  NOR2X0 U13271 ( .IN1(n13027), .IN2(n13028), .QN(n13025) );
  NOR2X0 U13272 ( .IN1(WX6033), .IN2(n7746), .QN(n13028) );
  INVX0 U13273 ( .INP(n13029), .ZN(n13027) );
  NAND2X0 U13274 ( .IN1(n7746), .IN2(WX6033), .QN(n13029) );
  NAND2X0 U13275 ( .IN1(n10068), .IN2(n8482), .QN(n13021) );
  NAND2X0 U13276 ( .IN1(n16363), .IN2(n9078), .QN(n13020) );
  NAND2X0 U13277 ( .IN1(n13030), .IN2(n13031), .QN(n13014) );
  NAND2X0 U13278 ( .IN1(n13032), .IN2(n13033), .QN(n13030) );
  NAND2X0 U13279 ( .IN1(n9108), .IN2(n13034), .QN(n13033) );
  NAND2X0 U13280 ( .IN1(n9108), .IN2(n8541), .QN(n13032) );
  NAND2X0 U13281 ( .IN1(n746), .IN2(n9283), .QN(n13013) );
  NOR2X0 U13282 ( .IN1(n9070), .IN2(n9161), .QN(n746) );
  NAND2X0 U13283 ( .IN1(n9295), .IN2(CRC_OUT_6_19), .QN(n13012) );
  NAND4X0 U13284 ( .IN1(n13035), .IN2(n13036), .IN3(n13037), .IN4(n13038), 
        .QN(WX4545) );
  NAND2X0 U13285 ( .IN1(n13039), .IN2(n13040), .QN(n13038) );
  NAND2X0 U13286 ( .IN1(n13041), .IN2(n13042), .QN(n13039) );
  NAND2X0 U13287 ( .IN1(n9108), .IN2(n13043), .QN(n13042) );
  NAND2X0 U13288 ( .IN1(n9108), .IN2(n8542), .QN(n13041) );
  NAND2X0 U13289 ( .IN1(n12357), .IN2(n2153), .QN(n13037) );
  NOR2X0 U13290 ( .IN1(n13044), .IN2(n13045), .QN(n12357) );
  INVX0 U13291 ( .INP(n13046), .ZN(n13045) );
  NAND2X0 U13292 ( .IN1(n13047), .IN2(n13048), .QN(n13046) );
  NOR2X0 U13293 ( .IN1(n13048), .IN2(n13047), .QN(n13044) );
  NAND2X0 U13294 ( .IN1(n13049), .IN2(n13050), .QN(n13047) );
  NAND2X0 U13295 ( .IN1(n8291), .IN2(n13051), .QN(n13050) );
  INVX0 U13296 ( .INP(n13052), .ZN(n13051) );
  NAND2X0 U13297 ( .IN1(n13052), .IN2(WX6031), .QN(n13049) );
  NAND2X0 U13298 ( .IN1(n13053), .IN2(n13054), .QN(n13052) );
  INVX0 U13299 ( .INP(n13055), .ZN(n13054) );
  NOR2X0 U13300 ( .IN1(n8813), .IN2(n16362), .QN(n13055) );
  NAND2X0 U13301 ( .IN1(n16362), .IN2(n8813), .QN(n13053) );
  NOR2X0 U13302 ( .IN1(n13056), .IN2(n13057), .QN(n13048) );
  INVX0 U13303 ( .INP(n13058), .ZN(n13057) );
  NAND2X0 U13304 ( .IN1(n7747), .IN2(n9118), .QN(n13058) );
  NOR2X0 U13305 ( .IN1(n9117), .IN2(n7747), .QN(n13056) );
  NAND2X0 U13306 ( .IN1(n745), .IN2(n9283), .QN(n13036) );
  NOR2X0 U13307 ( .IN1(n9233), .IN2(n8963), .QN(n745) );
  NAND2X0 U13308 ( .IN1(n9295), .IN2(CRC_OUT_6_20), .QN(n13035) );
  NAND4X0 U13309 ( .IN1(n13059), .IN2(n13060), .IN3(n13061), .IN4(n13062), 
        .QN(WX4543) );
  NAND2X0 U13310 ( .IN1(n13063), .IN2(n12363), .QN(n13062) );
  NAND2X0 U13311 ( .IN1(n13064), .IN2(n12366), .QN(n12363) );
  NAND2X0 U13312 ( .IN1(n13065), .IN2(n13066), .QN(n13064) );
  NAND2X0 U13313 ( .IN1(n16361), .IN2(n9118), .QN(n13066) );
  NAND2X0 U13314 ( .IN1(TM1), .IN2(n8484), .QN(n13065) );
  NAND3X0 U13315 ( .IN1(n13067), .IN2(n13068), .IN3(n13069), .QN(n13063) );
  NAND2X0 U13316 ( .IN1(n9325), .IN2(n12366), .QN(n13069) );
  NAND2X0 U13317 ( .IN1(n13070), .IN2(n13071), .QN(n12366) );
  NAND2X0 U13318 ( .IN1(n7748), .IN2(n13072), .QN(n13071) );
  INVX0 U13319 ( .INP(n13073), .ZN(n13070) );
  NOR2X0 U13320 ( .IN1(n13072), .IN2(n7748), .QN(n13073) );
  NOR2X0 U13321 ( .IN1(n13074), .IN2(n13075), .QN(n13072) );
  NOR2X0 U13322 ( .IN1(WX6029), .IN2(n7749), .QN(n13075) );
  INVX0 U13323 ( .INP(n13076), .ZN(n13074) );
  NAND2X0 U13324 ( .IN1(n7749), .IN2(WX6029), .QN(n13076) );
  NAND2X0 U13325 ( .IN1(n9084), .IN2(n8484), .QN(n13068) );
  NAND2X0 U13326 ( .IN1(n16361), .IN2(n10069), .QN(n13067) );
  NAND2X0 U13327 ( .IN1(n13077), .IN2(n13078), .QN(n13061) );
  NAND2X0 U13328 ( .IN1(n13079), .IN2(n13080), .QN(n13077) );
  NAND2X0 U13329 ( .IN1(n9108), .IN2(n13081), .QN(n13080) );
  NAND2X0 U13330 ( .IN1(n9108), .IN2(n8543), .QN(n13079) );
  NAND2X0 U13331 ( .IN1(n744), .IN2(n9283), .QN(n13060) );
  NOR2X0 U13332 ( .IN1(n9233), .IN2(n8964), .QN(n744) );
  NAND2X0 U13333 ( .IN1(n9295), .IN2(CRC_OUT_6_21), .QN(n13059) );
  NAND4X0 U13334 ( .IN1(n13082), .IN2(n13083), .IN3(n13084), .IN4(n13085), 
        .QN(WX4541) );
  NAND2X0 U13335 ( .IN1(n13086), .IN2(n12399), .QN(n13085) );
  NAND3X0 U13336 ( .IN1(n13087), .IN2(n13088), .IN3(n12402), .QN(n12399) );
  NAND2X0 U13337 ( .IN1(n8273), .IN2(n9119), .QN(n13088) );
  NAND2X0 U13338 ( .IN1(TM1), .IN2(WX6027), .QN(n13087) );
  NAND3X0 U13339 ( .IN1(n13089), .IN2(n13090), .IN3(n13091), .QN(n13086) );
  NAND2X0 U13340 ( .IN1(n9325), .IN2(n12402), .QN(n13091) );
  NAND2X0 U13341 ( .IN1(n13092), .IN2(n13093), .QN(n12402) );
  NAND2X0 U13342 ( .IN1(n13094), .IN2(WX5963), .QN(n13093) );
  NAND2X0 U13343 ( .IN1(n13095), .IN2(n13096), .QN(n13094) );
  NAND3X0 U13344 ( .IN1(n13095), .IN2(n13096), .IN3(n7751), .QN(n13092) );
  NAND2X0 U13345 ( .IN1(test_so46), .IN2(WX5899), .QN(n13096) );
  NAND2X0 U13346 ( .IN1(n7750), .IN2(n8822), .QN(n13095) );
  NAND2X0 U13347 ( .IN1(n10069), .IN2(WX6027), .QN(n13090) );
  NAND2X0 U13348 ( .IN1(n9083), .IN2(n8273), .QN(n13089) );
  NAND2X0 U13349 ( .IN1(n13097), .IN2(n13098), .QN(n13084) );
  NAND2X0 U13350 ( .IN1(n13099), .IN2(n13100), .QN(n13097) );
  NAND2X0 U13351 ( .IN1(n9108), .IN2(n13101), .QN(n13100) );
  NAND2X0 U13352 ( .IN1(n9108), .IN2(n8544), .QN(n13099) );
  NAND2X0 U13353 ( .IN1(n743), .IN2(n9283), .QN(n13083) );
  NOR2X0 U13354 ( .IN1(n9233), .IN2(n8965), .QN(n743) );
  NAND2X0 U13355 ( .IN1(test_so43), .IN2(n9314), .QN(n13082) );
  NAND4X0 U13356 ( .IN1(n13102), .IN2(n13103), .IN3(n13104), .IN4(n13105), 
        .QN(WX4539) );
  NAND2X0 U13357 ( .IN1(n13106), .IN2(n12408), .QN(n13105) );
  NAND2X0 U13358 ( .IN1(n13107), .IN2(n12411), .QN(n12408) );
  NAND2X0 U13359 ( .IN1(n13108), .IN2(n13109), .QN(n13107) );
  NAND2X0 U13360 ( .IN1(n16360), .IN2(n9118), .QN(n13109) );
  NAND2X0 U13361 ( .IN1(TM1), .IN2(n8487), .QN(n13108) );
  NAND3X0 U13362 ( .IN1(n13110), .IN2(n13111), .IN3(n13112), .QN(n13106) );
  NAND2X0 U13363 ( .IN1(n9325), .IN2(n12411), .QN(n13112) );
  NAND2X0 U13364 ( .IN1(n13113), .IN2(n13114), .QN(n12411) );
  NAND2X0 U13365 ( .IN1(n7752), .IN2(n13115), .QN(n13114) );
  INVX0 U13366 ( .INP(n13116), .ZN(n13113) );
  NOR2X0 U13367 ( .IN1(n13115), .IN2(n7752), .QN(n13116) );
  NOR2X0 U13368 ( .IN1(n13117), .IN2(n13118), .QN(n13115) );
  NOR2X0 U13369 ( .IN1(WX6025), .IN2(n7753), .QN(n13118) );
  INVX0 U13370 ( .INP(n13119), .ZN(n13117) );
  NAND2X0 U13371 ( .IN1(n7753), .IN2(WX6025), .QN(n13119) );
  NAND2X0 U13372 ( .IN1(n9082), .IN2(n8487), .QN(n13111) );
  NAND2X0 U13373 ( .IN1(n16360), .IN2(n9080), .QN(n13110) );
  NAND2X0 U13374 ( .IN1(n13120), .IN2(n13121), .QN(n13104) );
  NAND2X0 U13375 ( .IN1(n13122), .IN2(n13123), .QN(n13120) );
  NAND2X0 U13376 ( .IN1(n9108), .IN2(n13124), .QN(n13123) );
  NAND2X0 U13377 ( .IN1(n9108), .IN2(n8545), .QN(n13122) );
  NAND2X0 U13378 ( .IN1(n742), .IN2(n9283), .QN(n13103) );
  NOR2X0 U13379 ( .IN1(n9233), .IN2(n8966), .QN(n742) );
  NAND2X0 U13380 ( .IN1(n9295), .IN2(CRC_OUT_6_23), .QN(n13102) );
  NAND4X0 U13381 ( .IN1(n13125), .IN2(n13126), .IN3(n13127), .IN4(n13128), 
        .QN(WX4537) );
  NAND2X0 U13382 ( .IN1(n13129), .IN2(n12446), .QN(n13128) );
  NAND2X0 U13383 ( .IN1(n13130), .IN2(n12449), .QN(n12446) );
  NAND2X0 U13384 ( .IN1(n13131), .IN2(n13132), .QN(n13130) );
  NAND2X0 U13385 ( .IN1(n16359), .IN2(n9118), .QN(n13132) );
  NAND2X0 U13386 ( .IN1(TM1), .IN2(n8488), .QN(n13131) );
  NAND3X0 U13387 ( .IN1(n13133), .IN2(n13134), .IN3(n13135), .QN(n13129) );
  NAND2X0 U13388 ( .IN1(n9325), .IN2(n12449), .QN(n13135) );
  NAND2X0 U13389 ( .IN1(n13136), .IN2(n13137), .QN(n12449) );
  NAND2X0 U13390 ( .IN1(n7754), .IN2(n13138), .QN(n13137) );
  INVX0 U13391 ( .INP(n13139), .ZN(n13136) );
  NOR2X0 U13392 ( .IN1(n13138), .IN2(n7754), .QN(n13139) );
  NOR2X0 U13393 ( .IN1(n13140), .IN2(n13141), .QN(n13138) );
  NOR2X0 U13394 ( .IN1(WX6023), .IN2(n7755), .QN(n13141) );
  INVX0 U13395 ( .INP(n13142), .ZN(n13140) );
  NAND2X0 U13396 ( .IN1(n7755), .IN2(WX6023), .QN(n13142) );
  NAND2X0 U13397 ( .IN1(n10068), .IN2(n8488), .QN(n13134) );
  NAND2X0 U13398 ( .IN1(n16359), .IN2(n9079), .QN(n13133) );
  NAND2X0 U13399 ( .IN1(n13143), .IN2(n13144), .QN(n13127) );
  NAND2X0 U13400 ( .IN1(n13145), .IN2(n13146), .QN(n13143) );
  NAND2X0 U13401 ( .IN1(n9108), .IN2(n13147), .QN(n13146) );
  NAND2X0 U13402 ( .IN1(n9108), .IN2(n8546), .QN(n13145) );
  NAND2X0 U13403 ( .IN1(n741), .IN2(n9283), .QN(n13126) );
  NOR2X0 U13404 ( .IN1(n9233), .IN2(n8967), .QN(n741) );
  NAND2X0 U13405 ( .IN1(n9295), .IN2(CRC_OUT_6_24), .QN(n13125) );
  NAND4X0 U13406 ( .IN1(n13148), .IN2(n13149), .IN3(n13150), .IN4(n13151), 
        .QN(WX4535) );
  NAND2X0 U13407 ( .IN1(n13152), .IN2(n12455), .QN(n13151) );
  NAND2X0 U13408 ( .IN1(n13153), .IN2(n12458), .QN(n12455) );
  NAND2X0 U13409 ( .IN1(n13154), .IN2(n13155), .QN(n13153) );
  NAND2X0 U13410 ( .IN1(n16358), .IN2(n9118), .QN(n13155) );
  NAND2X0 U13411 ( .IN1(TM1), .IN2(n8489), .QN(n13154) );
  NAND3X0 U13412 ( .IN1(n13156), .IN2(n13157), .IN3(n13158), .QN(n13152) );
  NAND2X0 U13413 ( .IN1(n9325), .IN2(n12458), .QN(n13158) );
  NAND2X0 U13414 ( .IN1(n13159), .IN2(n13160), .QN(n12458) );
  NAND2X0 U13415 ( .IN1(n7756), .IN2(n13161), .QN(n13160) );
  INVX0 U13416 ( .INP(n13162), .ZN(n13159) );
  NOR2X0 U13417 ( .IN1(n13161), .IN2(n7756), .QN(n13162) );
  NOR2X0 U13418 ( .IN1(n13163), .IN2(n13164), .QN(n13161) );
  NOR2X0 U13419 ( .IN1(WX6021), .IN2(n7757), .QN(n13164) );
  INVX0 U13420 ( .INP(n13165), .ZN(n13163) );
  NAND2X0 U13421 ( .IN1(n7757), .IN2(WX6021), .QN(n13165) );
  NAND2X0 U13422 ( .IN1(n9084), .IN2(n8489), .QN(n13157) );
  NAND2X0 U13423 ( .IN1(n16358), .IN2(n9078), .QN(n13156) );
  NAND2X0 U13424 ( .IN1(n13166), .IN2(n13167), .QN(n13150) );
  NAND2X0 U13425 ( .IN1(n13168), .IN2(n13169), .QN(n13166) );
  NAND2X0 U13426 ( .IN1(n9108), .IN2(n13170), .QN(n13169) );
  NAND2X0 U13427 ( .IN1(n9108), .IN2(n8547), .QN(n13168) );
  NAND2X0 U13428 ( .IN1(n740), .IN2(n9283), .QN(n13149) );
  NOR2X0 U13429 ( .IN1(n9234), .IN2(n8968), .QN(n740) );
  NAND2X0 U13430 ( .IN1(n9295), .IN2(CRC_OUT_6_25), .QN(n13148) );
  NAND4X0 U13431 ( .IN1(n13171), .IN2(n13172), .IN3(n13173), .IN4(n13174), 
        .QN(WX4533) );
  NAND2X0 U13432 ( .IN1(n13175), .IN2(n12493), .QN(n13174) );
  NAND2X0 U13433 ( .IN1(n13176), .IN2(n12496), .QN(n12493) );
  NAND2X0 U13434 ( .IN1(n13177), .IN2(n13178), .QN(n13176) );
  NAND2X0 U13435 ( .IN1(n16357), .IN2(n9118), .QN(n13178) );
  NAND2X0 U13436 ( .IN1(TM1), .IN2(n8490), .QN(n13177) );
  NAND3X0 U13437 ( .IN1(n13179), .IN2(n13180), .IN3(n13181), .QN(n13175) );
  NAND2X0 U13438 ( .IN1(n9325), .IN2(n12496), .QN(n13181) );
  NAND2X0 U13439 ( .IN1(n13182), .IN2(n13183), .QN(n12496) );
  NAND2X0 U13440 ( .IN1(n7758), .IN2(n13184), .QN(n13183) );
  INVX0 U13441 ( .INP(n13185), .ZN(n13182) );
  NOR2X0 U13442 ( .IN1(n13184), .IN2(n7758), .QN(n13185) );
  NOR2X0 U13443 ( .IN1(n13186), .IN2(n13187), .QN(n13184) );
  NOR2X0 U13444 ( .IN1(WX6019), .IN2(n7759), .QN(n13187) );
  INVX0 U13445 ( .INP(n13188), .ZN(n13186) );
  NAND2X0 U13446 ( .IN1(n7759), .IN2(WX6019), .QN(n13188) );
  NAND2X0 U13447 ( .IN1(n9083), .IN2(n8490), .QN(n13180) );
  NAND2X0 U13448 ( .IN1(n16357), .IN2(n10069), .QN(n13179) );
  NAND2X0 U13449 ( .IN1(n13189), .IN2(n13190), .QN(n13173) );
  NAND2X0 U13450 ( .IN1(n13191), .IN2(n13192), .QN(n13189) );
  NAND2X0 U13451 ( .IN1(n9109), .IN2(n13193), .QN(n13192) );
  NAND2X0 U13452 ( .IN1(n9109), .IN2(n8548), .QN(n13191) );
  NAND2X0 U13453 ( .IN1(n739), .IN2(n9283), .QN(n13172) );
  NOR2X0 U13454 ( .IN1(n9234), .IN2(n8969), .QN(n739) );
  NAND2X0 U13455 ( .IN1(n9295), .IN2(CRC_OUT_6_26), .QN(n13171) );
  NAND4X0 U13456 ( .IN1(n13194), .IN2(n13195), .IN3(n13196), .IN4(n13197), 
        .QN(WX4531) );
  NAND2X0 U13457 ( .IN1(n13198), .IN2(n12513), .QN(n13197) );
  NAND2X0 U13458 ( .IN1(n13199), .IN2(n12516), .QN(n12513) );
  NAND2X0 U13459 ( .IN1(n13200), .IN2(n13201), .QN(n13199) );
  NAND2X0 U13460 ( .IN1(n16356), .IN2(n9119), .QN(n13201) );
  NAND2X0 U13461 ( .IN1(TM1), .IN2(n8491), .QN(n13200) );
  NAND3X0 U13462 ( .IN1(n13202), .IN2(n13203), .IN3(n13204), .QN(n13198) );
  NAND2X0 U13463 ( .IN1(n9325), .IN2(n12516), .QN(n13204) );
  NAND2X0 U13464 ( .IN1(n13205), .IN2(n13206), .QN(n12516) );
  NAND2X0 U13465 ( .IN1(n7760), .IN2(n13207), .QN(n13206) );
  INVX0 U13466 ( .INP(n13208), .ZN(n13205) );
  NOR2X0 U13467 ( .IN1(n13207), .IN2(n7760), .QN(n13208) );
  NOR2X0 U13468 ( .IN1(n13209), .IN2(n13210), .QN(n13207) );
  NOR2X0 U13469 ( .IN1(WX6017), .IN2(n7761), .QN(n13210) );
  INVX0 U13470 ( .INP(n13211), .ZN(n13209) );
  NAND2X0 U13471 ( .IN1(n7761), .IN2(WX6017), .QN(n13211) );
  NAND2X0 U13472 ( .IN1(n9082), .IN2(n8491), .QN(n13203) );
  NAND2X0 U13473 ( .IN1(n16356), .IN2(n9080), .QN(n13202) );
  NAND2X0 U13474 ( .IN1(n13212), .IN2(n13213), .QN(n13196) );
  NAND2X0 U13475 ( .IN1(n13214), .IN2(n13215), .QN(n13212) );
  NAND2X0 U13476 ( .IN1(n9109), .IN2(n13216), .QN(n13215) );
  NAND2X0 U13477 ( .IN1(n9109), .IN2(n8549), .QN(n13214) );
  NAND2X0 U13478 ( .IN1(n738), .IN2(n9283), .QN(n13195) );
  NOR2X0 U13479 ( .IN1(n9234), .IN2(n8970), .QN(n738) );
  NAND2X0 U13480 ( .IN1(n9295), .IN2(CRC_OUT_6_27), .QN(n13194) );
  NAND4X0 U13481 ( .IN1(n13217), .IN2(n13218), .IN3(n13219), .IN4(n13220), 
        .QN(WX4529) );
  NAND2X0 U13482 ( .IN1(n13221), .IN2(n12536), .QN(n13220) );
  NAND2X0 U13483 ( .IN1(n13222), .IN2(n12539), .QN(n12536) );
  NAND2X0 U13484 ( .IN1(n13223), .IN2(n13224), .QN(n13222) );
  NAND2X0 U13485 ( .IN1(n16355), .IN2(n9118), .QN(n13224) );
  NAND2X0 U13486 ( .IN1(TM1), .IN2(n8492), .QN(n13223) );
  NAND3X0 U13487 ( .IN1(n13225), .IN2(n13226), .IN3(n13227), .QN(n13221) );
  NAND2X0 U13488 ( .IN1(n9325), .IN2(n12539), .QN(n13227) );
  NAND2X0 U13489 ( .IN1(n13228), .IN2(n13229), .QN(n12539) );
  NAND2X0 U13490 ( .IN1(n7762), .IN2(n13230), .QN(n13229) );
  INVX0 U13491 ( .INP(n13231), .ZN(n13228) );
  NOR2X0 U13492 ( .IN1(n13230), .IN2(n7762), .QN(n13231) );
  NOR2X0 U13493 ( .IN1(n13232), .IN2(n13233), .QN(n13230) );
  NOR2X0 U13494 ( .IN1(WX6015), .IN2(n7763), .QN(n13233) );
  INVX0 U13495 ( .INP(n13234), .ZN(n13232) );
  NAND2X0 U13496 ( .IN1(n7763), .IN2(WX6015), .QN(n13234) );
  NAND2X0 U13497 ( .IN1(n10068), .IN2(n8492), .QN(n13226) );
  NAND2X0 U13498 ( .IN1(n16355), .IN2(n9079), .QN(n13225) );
  NAND2X0 U13499 ( .IN1(n13235), .IN2(n9111), .QN(n13219) );
  NAND2X0 U13500 ( .IN1(n737), .IN2(n9283), .QN(n13218) );
  NOR2X0 U13501 ( .IN1(n9234), .IN2(n8971), .QN(n737) );
  NAND2X0 U13502 ( .IN1(n9295), .IN2(CRC_OUT_6_28), .QN(n13217) );
  NAND4X0 U13503 ( .IN1(n13236), .IN2(n13237), .IN3(n13238), .IN4(n13239), 
        .QN(WX4527) );
  NAND2X0 U13504 ( .IN1(n13240), .IN2(n12559), .QN(n13239) );
  NAND2X0 U13505 ( .IN1(n13241), .IN2(n12562), .QN(n12559) );
  NAND2X0 U13506 ( .IN1(n13242), .IN2(n13243), .QN(n13241) );
  NAND2X0 U13507 ( .IN1(n16354), .IN2(n9118), .QN(n13243) );
  NAND2X0 U13508 ( .IN1(TM1), .IN2(n8493), .QN(n13242) );
  NAND3X0 U13509 ( .IN1(n13244), .IN2(n13245), .IN3(n13246), .QN(n13240) );
  NAND2X0 U13510 ( .IN1(n9326), .IN2(n12562), .QN(n13246) );
  NAND2X0 U13511 ( .IN1(n13247), .IN2(n13248), .QN(n12562) );
  NAND2X0 U13512 ( .IN1(n7764), .IN2(n13249), .QN(n13248) );
  INVX0 U13513 ( .INP(n13250), .ZN(n13247) );
  NOR2X0 U13514 ( .IN1(n13249), .IN2(n7764), .QN(n13250) );
  NOR2X0 U13515 ( .IN1(n13251), .IN2(n13252), .QN(n13249) );
  NOR2X0 U13516 ( .IN1(WX6013), .IN2(n7765), .QN(n13252) );
  INVX0 U13517 ( .INP(n13253), .ZN(n13251) );
  NAND2X0 U13518 ( .IN1(n7765), .IN2(WX6013), .QN(n13253) );
  NAND2X0 U13519 ( .IN1(n9084), .IN2(n8493), .QN(n13245) );
  NAND2X0 U13520 ( .IN1(n16354), .IN2(n9078), .QN(n13244) );
  NAND2X0 U13521 ( .IN1(n13254), .IN2(n13255), .QN(n13238) );
  NAND2X0 U13522 ( .IN1(n13256), .IN2(n13257), .QN(n13254) );
  NAND2X0 U13523 ( .IN1(n9109), .IN2(n13258), .QN(n13257) );
  NAND2X0 U13524 ( .IN1(n9109), .IN2(n8551), .QN(n13256) );
  NAND2X0 U13525 ( .IN1(n736), .IN2(n9283), .QN(n13237) );
  NOR2X0 U13526 ( .IN1(n9234), .IN2(n8972), .QN(n736) );
  NAND2X0 U13527 ( .IN1(n9295), .IN2(CRC_OUT_6_29), .QN(n13236) );
  NAND4X0 U13528 ( .IN1(n13259), .IN2(n13260), .IN3(n13261), .IN4(n13262), 
        .QN(WX4525) );
  NAND2X0 U13529 ( .IN1(n13263), .IN2(n12582), .QN(n13262) );
  NAND2X0 U13530 ( .IN1(n13264), .IN2(n12585), .QN(n12582) );
  NAND2X0 U13531 ( .IN1(n13265), .IN2(n13266), .QN(n13264) );
  NAND2X0 U13532 ( .IN1(n16353), .IN2(n9119), .QN(n13266) );
  NAND2X0 U13533 ( .IN1(TM1), .IN2(n8494), .QN(n13265) );
  NAND3X0 U13534 ( .IN1(n13267), .IN2(n13268), .IN3(n13269), .QN(n13263) );
  NAND2X0 U13535 ( .IN1(n9326), .IN2(n12585), .QN(n13269) );
  NAND2X0 U13536 ( .IN1(n13270), .IN2(n13271), .QN(n12585) );
  NAND2X0 U13537 ( .IN1(n7766), .IN2(n13272), .QN(n13271) );
  INVX0 U13538 ( .INP(n13273), .ZN(n13270) );
  NOR2X0 U13539 ( .IN1(n13272), .IN2(n7766), .QN(n13273) );
  NOR2X0 U13540 ( .IN1(n13274), .IN2(n13275), .QN(n13272) );
  NOR2X0 U13541 ( .IN1(WX6011), .IN2(n7767), .QN(n13275) );
  INVX0 U13542 ( .INP(n13276), .ZN(n13274) );
  NAND2X0 U13543 ( .IN1(n7767), .IN2(WX6011), .QN(n13276) );
  NAND2X0 U13544 ( .IN1(n9083), .IN2(n8494), .QN(n13268) );
  NAND2X0 U13545 ( .IN1(n16353), .IN2(n10069), .QN(n13267) );
  NAND2X0 U13546 ( .IN1(n13277), .IN2(n9110), .QN(n13261) );
  NAND2X0 U13547 ( .IN1(n735), .IN2(n9283), .QN(n13260) );
  NOR2X0 U13548 ( .IN1(n9234), .IN2(n8973), .QN(n735) );
  NAND2X0 U13549 ( .IN1(n9295), .IN2(CRC_OUT_6_30), .QN(n13259) );
  NAND4X0 U13550 ( .IN1(n13278), .IN2(n13279), .IN3(n13280), .IN4(n13281), 
        .QN(WX4523) );
  NAND2X0 U13551 ( .IN1(n13282), .IN2(n12605), .QN(n13281) );
  NAND2X0 U13552 ( .IN1(n13283), .IN2(n12608), .QN(n12605) );
  NAND2X0 U13553 ( .IN1(n13284), .IN2(n13285), .QN(n13283) );
  NAND2X0 U13554 ( .IN1(n16352), .IN2(n9119), .QN(n13285) );
  NAND2X0 U13555 ( .IN1(TM1), .IN2(n8495), .QN(n13284) );
  NAND3X0 U13556 ( .IN1(n13286), .IN2(n13287), .IN3(n13288), .QN(n13282) );
  NAND2X0 U13557 ( .IN1(n9326), .IN2(n12608), .QN(n13288) );
  NAND2X0 U13558 ( .IN1(n13289), .IN2(n13290), .QN(n12608) );
  NAND2X0 U13559 ( .IN1(n7620), .IN2(n13291), .QN(n13290) );
  INVX0 U13560 ( .INP(n13292), .ZN(n13289) );
  NOR2X0 U13561 ( .IN1(n13291), .IN2(n7620), .QN(n13292) );
  NOR2X0 U13562 ( .IN1(n13293), .IN2(n13294), .QN(n13291) );
  NOR2X0 U13563 ( .IN1(WX6009), .IN2(n7621), .QN(n13294) );
  INVX0 U13564 ( .INP(n13295), .ZN(n13293) );
  NAND2X0 U13565 ( .IN1(n7621), .IN2(WX6009), .QN(n13295) );
  NAND2X0 U13566 ( .IN1(n9082), .IN2(n8495), .QN(n13287) );
  NAND2X0 U13567 ( .IN1(n16352), .IN2(n9080), .QN(n13286) );
  NAND2X0 U13568 ( .IN1(n13296), .IN2(n13297), .QN(n13280) );
  NAND2X0 U13569 ( .IN1(n13298), .IN2(n13299), .QN(n13296) );
  NAND2X0 U13570 ( .IN1(n9109), .IN2(n13300), .QN(n13299) );
  NAND2X0 U13571 ( .IN1(n9109), .IN2(n8553), .QN(n13298) );
  NAND2X0 U13572 ( .IN1(n9296), .IN2(CRC_OUT_6_31), .QN(n13279) );
  NAND2X0 U13573 ( .IN1(n2245), .IN2(WX4364), .QN(n13278) );
  NOR2X0 U13574 ( .IN1(n9234), .IN2(WX4364), .QN(WX4425) );
  NOR3X0 U13575 ( .IN1(n9138), .IN2(n13301), .IN3(n13302), .QN(WX3912) );
  NOR2X0 U13576 ( .IN1(n8471), .IN2(CRC_OUT_7_30), .QN(n13302) );
  NOR2X0 U13577 ( .IN1(DFF_574_n1), .IN2(WX3423), .QN(n13301) );
  NOR3X0 U13578 ( .IN1(n9138), .IN2(n13303), .IN3(n13304), .QN(WX3910) );
  NOR2X0 U13579 ( .IN1(n8472), .IN2(CRC_OUT_7_29), .QN(n13304) );
  NOR2X0 U13580 ( .IN1(DFF_573_n1), .IN2(WX3425), .QN(n13303) );
  NOR3X0 U13581 ( .IN1(n9138), .IN2(n13305), .IN3(n13306), .QN(WX3908) );
  NOR2X0 U13582 ( .IN1(n8473), .IN2(CRC_OUT_7_28), .QN(n13306) );
  NOR2X0 U13583 ( .IN1(DFF_572_n1), .IN2(WX3427), .QN(n13305) );
  NOR2X0 U13584 ( .IN1(n9234), .IN2(n13307), .QN(WX3906) );
  NOR2X0 U13585 ( .IN1(n13308), .IN2(n13309), .QN(n13307) );
  NOR2X0 U13586 ( .IN1(test_so32), .IN2(WX3429), .QN(n13309) );
  INVX0 U13587 ( .INP(n13310), .ZN(n13308) );
  NAND2X0 U13588 ( .IN1(WX3429), .IN2(test_so32), .QN(n13310) );
  NOR3X0 U13589 ( .IN1(n9138), .IN2(n13311), .IN3(n13312), .QN(WX3904) );
  NOR2X0 U13590 ( .IN1(n8475), .IN2(CRC_OUT_7_26), .QN(n13312) );
  NOR2X0 U13591 ( .IN1(DFF_570_n1), .IN2(WX3431), .QN(n13311) );
  NOR3X0 U13592 ( .IN1(n9138), .IN2(n13313), .IN3(n13314), .QN(WX3902) );
  NOR2X0 U13593 ( .IN1(n8476), .IN2(CRC_OUT_7_25), .QN(n13314) );
  NOR2X0 U13594 ( .IN1(DFF_569_n1), .IN2(WX3433), .QN(n13313) );
  NOR3X0 U13595 ( .IN1(n9138), .IN2(n13315), .IN3(n13316), .QN(WX3900) );
  NOR2X0 U13596 ( .IN1(n8477), .IN2(CRC_OUT_7_24), .QN(n13316) );
  NOR2X0 U13597 ( .IN1(DFF_568_n1), .IN2(WX3435), .QN(n13315) );
  NOR3X0 U13598 ( .IN1(n9138), .IN2(n13317), .IN3(n13318), .QN(WX3898) );
  NOR2X0 U13599 ( .IN1(n8478), .IN2(CRC_OUT_7_23), .QN(n13318) );
  NOR2X0 U13600 ( .IN1(DFF_567_n1), .IN2(WX3437), .QN(n13317) );
  NOR2X0 U13601 ( .IN1(n9234), .IN2(n13319), .QN(WX3896) );
  NOR2X0 U13602 ( .IN1(n13320), .IN2(n13321), .QN(n13319) );
  NOR2X0 U13603 ( .IN1(test_so29), .IN2(CRC_OUT_7_22), .QN(n13321) );
  NOR2X0 U13604 ( .IN1(DFF_566_n1), .IN2(n8802), .QN(n13320) );
  NOR3X0 U13605 ( .IN1(n9137), .IN2(n13322), .IN3(n13323), .QN(WX3894) );
  NOR2X0 U13606 ( .IN1(n8485), .IN2(CRC_OUT_7_21), .QN(n13323) );
  NOR2X0 U13607 ( .IN1(DFF_565_n1), .IN2(WX3441), .QN(n13322) );
  NOR3X0 U13608 ( .IN1(n9137), .IN2(n13324), .IN3(n13325), .QN(WX3892) );
  NOR2X0 U13609 ( .IN1(n8486), .IN2(CRC_OUT_7_20), .QN(n13325) );
  NOR2X0 U13610 ( .IN1(DFF_564_n1), .IN2(WX3443), .QN(n13324) );
  NOR3X0 U13611 ( .IN1(n9137), .IN2(n13326), .IN3(n13327), .QN(WX3890) );
  NOR2X0 U13612 ( .IN1(n8503), .IN2(CRC_OUT_7_19), .QN(n13327) );
  NOR2X0 U13613 ( .IN1(DFF_563_n1), .IN2(WX3445), .QN(n13326) );
  NOR3X0 U13614 ( .IN1(n9137), .IN2(n13328), .IN3(n13329), .QN(WX3888) );
  NOR2X0 U13615 ( .IN1(n8504), .IN2(CRC_OUT_7_18), .QN(n13329) );
  NOR2X0 U13616 ( .IN1(DFF_562_n1), .IN2(WX3447), .QN(n13328) );
  NOR3X0 U13617 ( .IN1(n9137), .IN2(n13330), .IN3(n13331), .QN(WX3886) );
  NOR2X0 U13618 ( .IN1(n8521), .IN2(CRC_OUT_7_17), .QN(n13331) );
  NOR2X0 U13619 ( .IN1(DFF_561_n1), .IN2(WX3449), .QN(n13330) );
  NOR3X0 U13620 ( .IN1(n9137), .IN2(n13332), .IN3(n13333), .QN(WX3884) );
  NOR2X0 U13621 ( .IN1(n8522), .IN2(CRC_OUT_7_16), .QN(n13333) );
  NOR2X0 U13622 ( .IN1(DFF_560_n1), .IN2(WX3451), .QN(n13332) );
  NOR2X0 U13623 ( .IN1(n9235), .IN2(n13334), .QN(WX3882) );
  NOR2X0 U13624 ( .IN1(n13335), .IN2(n13336), .QN(n13334) );
  INVX0 U13625 ( .INP(n13337), .ZN(n13336) );
  NAND2X0 U13626 ( .IN1(CRC_OUT_7_15), .IN2(n13338), .QN(n13337) );
  NOR2X0 U13627 ( .IN1(n13338), .IN2(CRC_OUT_7_15), .QN(n13335) );
  NAND2X0 U13628 ( .IN1(n13339), .IN2(n13340), .QN(n13338) );
  NAND2X0 U13629 ( .IN1(n8120), .IN2(CRC_OUT_7_31), .QN(n13340) );
  NAND2X0 U13630 ( .IN1(DFF_575_n1), .IN2(WX3453), .QN(n13339) );
  NOR3X0 U13631 ( .IN1(n9137), .IN2(n13341), .IN3(n13342), .QN(WX3880) );
  NOR2X0 U13632 ( .IN1(n8529), .IN2(CRC_OUT_7_14), .QN(n13342) );
  NOR2X0 U13633 ( .IN1(DFF_558_n1), .IN2(WX3455), .QN(n13341) );
  NOR3X0 U13634 ( .IN1(n9137), .IN2(n13343), .IN3(n13344), .QN(WX3878) );
  NOR2X0 U13635 ( .IN1(n8530), .IN2(CRC_OUT_7_13), .QN(n13344) );
  NOR2X0 U13636 ( .IN1(DFF_557_n1), .IN2(WX3457), .QN(n13343) );
  NOR3X0 U13637 ( .IN1(n9137), .IN2(n13345), .IN3(n13346), .QN(WX3876) );
  NOR2X0 U13638 ( .IN1(n8531), .IN2(CRC_OUT_7_12), .QN(n13346) );
  NOR2X0 U13639 ( .IN1(DFF_556_n1), .IN2(WX3459), .QN(n13345) );
  NOR3X0 U13640 ( .IN1(n9137), .IN2(n13347), .IN3(n13348), .QN(WX3874) );
  NOR2X0 U13641 ( .IN1(n8532), .IN2(CRC_OUT_7_11), .QN(n13348) );
  NOR2X0 U13642 ( .IN1(DFF_555_n1), .IN2(WX3461), .QN(n13347) );
  NOR3X0 U13643 ( .IN1(n9137), .IN2(n13349), .IN3(n13350), .QN(WX3872) );
  NOR2X0 U13644 ( .IN1(DFF_575_n1), .IN2(n13351), .QN(n13350) );
  INVX0 U13645 ( .INP(n13352), .ZN(n13349) );
  NAND2X0 U13646 ( .IN1(n13351), .IN2(DFF_575_n1), .QN(n13352) );
  NOR2X0 U13647 ( .IN1(n13353), .IN2(n13354), .QN(n13351) );
  INVX0 U13648 ( .INP(n13355), .ZN(n13354) );
  NAND2X0 U13649 ( .IN1(test_so31), .IN2(WX3463), .QN(n13355) );
  NOR2X0 U13650 ( .IN1(WX3463), .IN2(test_so31), .QN(n13353) );
  NOR3X0 U13651 ( .IN1(n9137), .IN2(n13356), .IN3(n13357), .QN(WX3870) );
  NOR2X0 U13652 ( .IN1(n8533), .IN2(CRC_OUT_7_9), .QN(n13357) );
  NOR2X0 U13653 ( .IN1(DFF_553_n1), .IN2(WX3465), .QN(n13356) );
  NOR3X0 U13654 ( .IN1(n9136), .IN2(n13358), .IN3(n13359), .QN(WX3868) );
  NOR2X0 U13655 ( .IN1(n8534), .IN2(CRC_OUT_7_8), .QN(n13359) );
  NOR2X0 U13656 ( .IN1(DFF_552_n1), .IN2(WX3467), .QN(n13358) );
  NOR3X0 U13657 ( .IN1(n9136), .IN2(n13360), .IN3(n13361), .QN(WX3866) );
  NOR2X0 U13658 ( .IN1(n8535), .IN2(CRC_OUT_7_7), .QN(n13361) );
  NOR2X0 U13659 ( .IN1(DFF_551_n1), .IN2(WX3469), .QN(n13360) );
  NOR3X0 U13660 ( .IN1(n9136), .IN2(n13362), .IN3(n13363), .QN(WX3864) );
  NOR2X0 U13661 ( .IN1(n8536), .IN2(CRC_OUT_7_6), .QN(n13363) );
  NOR2X0 U13662 ( .IN1(DFF_550_n1), .IN2(WX3471), .QN(n13362) );
  NOR2X0 U13663 ( .IN1(n9235), .IN2(n13364), .QN(WX3862) );
  NOR2X0 U13664 ( .IN1(n13365), .IN2(n13366), .QN(n13364) );
  NOR2X0 U13665 ( .IN1(test_so30), .IN2(CRC_OUT_7_5), .QN(n13366) );
  NOR2X0 U13666 ( .IN1(DFF_549_n1), .IN2(n8792), .QN(n13365) );
  NOR3X0 U13667 ( .IN1(n9136), .IN2(n13367), .IN3(n13368), .QN(WX3860) );
  NOR2X0 U13668 ( .IN1(n8538), .IN2(CRC_OUT_7_4), .QN(n13368) );
  NOR2X0 U13669 ( .IN1(DFF_548_n1), .IN2(WX3475), .QN(n13367) );
  NOR2X0 U13670 ( .IN1(n9236), .IN2(n13369), .QN(WX3858) );
  NOR2X0 U13671 ( .IN1(n13370), .IN2(n13371), .QN(n13369) );
  INVX0 U13672 ( .INP(n13372), .ZN(n13371) );
  NAND2X0 U13673 ( .IN1(CRC_OUT_7_3), .IN2(n13373), .QN(n13372) );
  NOR2X0 U13674 ( .IN1(n13373), .IN2(CRC_OUT_7_3), .QN(n13370) );
  NAND2X0 U13675 ( .IN1(n13374), .IN2(n13375), .QN(n13373) );
  NAND2X0 U13676 ( .IN1(n8122), .IN2(CRC_OUT_7_31), .QN(n13375) );
  NAND2X0 U13677 ( .IN1(DFF_575_n1), .IN2(WX3477), .QN(n13374) );
  NOR3X0 U13678 ( .IN1(n9136), .IN2(n13376), .IN3(n13377), .QN(WX3856) );
  NOR2X0 U13679 ( .IN1(n8539), .IN2(CRC_OUT_7_2), .QN(n13377) );
  NOR2X0 U13680 ( .IN1(DFF_546_n1), .IN2(WX3479), .QN(n13376) );
  NOR3X0 U13681 ( .IN1(n9136), .IN2(n13378), .IN3(n13379), .QN(WX3854) );
  NOR2X0 U13682 ( .IN1(n8556), .IN2(CRC_OUT_7_1), .QN(n13379) );
  NOR2X0 U13683 ( .IN1(DFF_545_n1), .IN2(WX3481), .QN(n13378) );
  NOR3X0 U13684 ( .IN1(n9136), .IN2(n13380), .IN3(n13381), .QN(WX3852) );
  NOR2X0 U13685 ( .IN1(n8557), .IN2(CRC_OUT_7_0), .QN(n13381) );
  NOR2X0 U13686 ( .IN1(DFF_544_n1), .IN2(WX3483), .QN(n13380) );
  NOR3X0 U13687 ( .IN1(n9136), .IN2(n13382), .IN3(n13383), .QN(WX3850) );
  NOR2X0 U13688 ( .IN1(n8132), .IN2(CRC_OUT_7_31), .QN(n13383) );
  NOR2X0 U13689 ( .IN1(DFF_575_n1), .IN2(WX3485), .QN(n13382) );
  NOR2X0 U13690 ( .IN1(n9236), .IN2(n8824), .QN(WX3324) );
  NOR2X0 U13691 ( .IN1(n16336), .IN2(n9160), .QN(WX3322) );
  NOR2X0 U13692 ( .IN1(n16335), .IN2(n9160), .QN(WX3320) );
  NOR2X0 U13693 ( .IN1(n16334), .IN2(n9160), .QN(WX3318) );
  NOR2X0 U13694 ( .IN1(n16333), .IN2(n9160), .QN(WX3316) );
  NOR2X0 U13695 ( .IN1(n16332), .IN2(n9160), .QN(WX3314) );
  NOR2X0 U13696 ( .IN1(n16331), .IN2(n9160), .QN(WX3312) );
  NOR2X0 U13697 ( .IN1(n16330), .IN2(n9160), .QN(WX3310) );
  NOR2X0 U13698 ( .IN1(n16329), .IN2(n9160), .QN(WX3308) );
  NOR2X0 U13699 ( .IN1(n16328), .IN2(n9159), .QN(WX3306) );
  NOR2X0 U13700 ( .IN1(n16327), .IN2(n9159), .QN(WX3304) );
  NOR2X0 U13701 ( .IN1(n16326), .IN2(n9159), .QN(WX3302) );
  NOR2X0 U13702 ( .IN1(n16325), .IN2(n9159), .QN(WX3300) );
  NOR2X0 U13703 ( .IN1(n16324), .IN2(n9159), .QN(WX3298) );
  NOR2X0 U13704 ( .IN1(n16323), .IN2(n9159), .QN(WX3296) );
  NOR2X0 U13705 ( .IN1(n16322), .IN2(n9159), .QN(WX3294) );
  NAND4X0 U13706 ( .IN1(n13384), .IN2(n13385), .IN3(n13386), .IN4(n13387), 
        .QN(WX3292) );
  NAND3X0 U13707 ( .IN1(n12696), .IN2(n12697), .IN3(n9321), .QN(n13387) );
  NAND3X0 U13708 ( .IN1(n13388), .IN2(n13389), .IN3(n13390), .QN(n12697) );
  INVX0 U13709 ( .INP(n13391), .ZN(n13390) );
  NAND2X0 U13710 ( .IN1(n13391), .IN2(n13392), .QN(n12696) );
  NAND2X0 U13711 ( .IN1(n13388), .IN2(n13389), .QN(n13392) );
  NAND2X0 U13712 ( .IN1(n8131), .IN2(WX4650), .QN(n13389) );
  NAND2X0 U13713 ( .IN1(n3691), .IN2(WX4778), .QN(n13388) );
  NOR2X0 U13714 ( .IN1(n13393), .IN2(n13394), .QN(n13391) );
  INVX0 U13715 ( .INP(n13395), .ZN(n13394) );
  NAND2X0 U13716 ( .IN1(test_so36), .IN2(WX4714), .QN(n13395) );
  NOR2X0 U13717 ( .IN1(WX4714), .IN2(test_so36), .QN(n13393) );
  NAND2X0 U13718 ( .IN1(n9109), .IN2(n13396), .QN(n13386) );
  NAND2X0 U13719 ( .IN1(n524), .IN2(n9284), .QN(n13385) );
  NOR2X0 U13720 ( .IN1(n9237), .IN2(n8974), .QN(n524) );
  NAND2X0 U13721 ( .IN1(n9296), .IN2(CRC_OUT_7_0), .QN(n13384) );
  NAND4X0 U13722 ( .IN1(n13397), .IN2(n13398), .IN3(n13399), .IN4(n13400), 
        .QN(WX3290) );
  NAND2X0 U13723 ( .IN1(n9326), .IN2(n12721), .QN(n13400) );
  NAND2X0 U13724 ( .IN1(n13401), .IN2(n13402), .QN(n12721) );
  INVX0 U13725 ( .INP(n13403), .ZN(n13402) );
  NOR2X0 U13726 ( .IN1(n13404), .IN2(n13405), .QN(n13403) );
  NAND2X0 U13727 ( .IN1(n13405), .IN2(n13404), .QN(n13401) );
  NOR2X0 U13728 ( .IN1(n13406), .IN2(n13407), .QN(n13404) );
  NOR2X0 U13729 ( .IN1(WX4776), .IN2(n8007), .QN(n13407) );
  INVX0 U13730 ( .INP(n13408), .ZN(n13406) );
  NAND2X0 U13731 ( .IN1(n8007), .IN2(WX4776), .QN(n13408) );
  NAND2X0 U13732 ( .IN1(n13409), .IN2(n13410), .QN(n13405) );
  NAND2X0 U13733 ( .IN1(n8006), .IN2(WX4648), .QN(n13410) );
  INVX0 U13734 ( .INP(n13411), .ZN(n13409) );
  NOR2X0 U13735 ( .IN1(WX4648), .IN2(n8006), .QN(n13411) );
  NAND2X0 U13736 ( .IN1(n9109), .IN2(n13412), .QN(n13399) );
  NAND2X0 U13737 ( .IN1(n523), .IN2(n9284), .QN(n13398) );
  NOR2X0 U13738 ( .IN1(n9237), .IN2(n8975), .QN(n523) );
  NAND2X0 U13739 ( .IN1(n9296), .IN2(CRC_OUT_7_1), .QN(n13397) );
  NAND4X0 U13740 ( .IN1(n13413), .IN2(n13414), .IN3(n13415), .IN4(n13416), 
        .QN(WX3288) );
  NAND2X0 U13741 ( .IN1(n9326), .IN2(n12737), .QN(n13416) );
  NAND2X0 U13742 ( .IN1(n13417), .IN2(n13418), .QN(n12737) );
  INVX0 U13743 ( .INP(n13419), .ZN(n13418) );
  NOR2X0 U13744 ( .IN1(n13420), .IN2(n13421), .QN(n13419) );
  NAND2X0 U13745 ( .IN1(n13421), .IN2(n13420), .QN(n13417) );
  NOR2X0 U13746 ( .IN1(n13422), .IN2(n13423), .QN(n13420) );
  NOR2X0 U13747 ( .IN1(WX4774), .IN2(n8009), .QN(n13423) );
  INVX0 U13748 ( .INP(n13424), .ZN(n13422) );
  NAND2X0 U13749 ( .IN1(n8009), .IN2(WX4774), .QN(n13424) );
  NAND2X0 U13750 ( .IN1(n13425), .IN2(n13426), .QN(n13421) );
  NAND2X0 U13751 ( .IN1(n8008), .IN2(WX4646), .QN(n13426) );
  INVX0 U13752 ( .INP(n13427), .ZN(n13425) );
  NOR2X0 U13753 ( .IN1(WX4646), .IN2(n8008), .QN(n13427) );
  NAND2X0 U13754 ( .IN1(n9110), .IN2(n13428), .QN(n13415) );
  NAND2X0 U13755 ( .IN1(n522), .IN2(n9284), .QN(n13414) );
  NOR2X0 U13756 ( .IN1(n9071), .IN2(n9159), .QN(n522) );
  NAND2X0 U13757 ( .IN1(n9296), .IN2(CRC_OUT_7_2), .QN(n13413) );
  NAND4X0 U13758 ( .IN1(n13429), .IN2(n13430), .IN3(n13431), .IN4(n13432), 
        .QN(WX3286) );
  NAND2X0 U13759 ( .IN1(n9326), .IN2(n12750), .QN(n13432) );
  NAND2X0 U13760 ( .IN1(n13433), .IN2(n13434), .QN(n12750) );
  INVX0 U13761 ( .INP(n13435), .ZN(n13434) );
  NOR2X0 U13762 ( .IN1(n13436), .IN2(n13437), .QN(n13435) );
  NAND2X0 U13763 ( .IN1(n13437), .IN2(n13436), .QN(n13433) );
  NOR2X0 U13764 ( .IN1(n13438), .IN2(n13439), .QN(n13436) );
  NOR2X0 U13765 ( .IN1(WX4772), .IN2(n8011), .QN(n13439) );
  INVX0 U13766 ( .INP(n13440), .ZN(n13438) );
  NAND2X0 U13767 ( .IN1(n8011), .IN2(WX4772), .QN(n13440) );
  NAND2X0 U13768 ( .IN1(n13441), .IN2(n13442), .QN(n13437) );
  NAND2X0 U13769 ( .IN1(n8010), .IN2(WX4644), .QN(n13442) );
  INVX0 U13770 ( .INP(n13443), .ZN(n13441) );
  NOR2X0 U13771 ( .IN1(WX4644), .IN2(n8010), .QN(n13443) );
  NAND2X0 U13772 ( .IN1(n9109), .IN2(n13444), .QN(n13431) );
  NAND2X0 U13773 ( .IN1(n521), .IN2(n9284), .QN(n13430) );
  NOR2X0 U13774 ( .IN1(n9237), .IN2(n8976), .QN(n521) );
  NAND2X0 U13775 ( .IN1(n9296), .IN2(CRC_OUT_7_3), .QN(n13429) );
  NAND4X0 U13776 ( .IN1(n13445), .IN2(n13446), .IN3(n13447), .IN4(n13448), 
        .QN(WX3284) );
  NAND2X0 U13777 ( .IN1(n9326), .IN2(n12766), .QN(n13448) );
  NAND2X0 U13778 ( .IN1(n13449), .IN2(n13450), .QN(n12766) );
  INVX0 U13779 ( .INP(n13451), .ZN(n13450) );
  NOR2X0 U13780 ( .IN1(n13452), .IN2(n13453), .QN(n13451) );
  NAND2X0 U13781 ( .IN1(n13453), .IN2(n13452), .QN(n13449) );
  NOR2X0 U13782 ( .IN1(n13454), .IN2(n13455), .QN(n13452) );
  NOR2X0 U13783 ( .IN1(WX4770), .IN2(n8013), .QN(n13455) );
  INVX0 U13784 ( .INP(n13456), .ZN(n13454) );
  NAND2X0 U13785 ( .IN1(n8013), .IN2(WX4770), .QN(n13456) );
  NAND2X0 U13786 ( .IN1(n13457), .IN2(n13458), .QN(n13453) );
  NAND2X0 U13787 ( .IN1(n8012), .IN2(WX4642), .QN(n13458) );
  INVX0 U13788 ( .INP(n13459), .ZN(n13457) );
  NOR2X0 U13789 ( .IN1(WX4642), .IN2(n8012), .QN(n13459) );
  NAND2X0 U13790 ( .IN1(n9110), .IN2(n13460), .QN(n13447) );
  NAND2X0 U13791 ( .IN1(n520), .IN2(n9284), .QN(n13446) );
  NOR2X0 U13792 ( .IN1(n9237), .IN2(n8977), .QN(n520) );
  NAND2X0 U13793 ( .IN1(n9296), .IN2(CRC_OUT_7_4), .QN(n13445) );
  NAND4X0 U13794 ( .IN1(n13461), .IN2(n13462), .IN3(n13463), .IN4(n13464), 
        .QN(WX3282) );
  NAND2X0 U13795 ( .IN1(n9326), .IN2(n12779), .QN(n13464) );
  NAND2X0 U13796 ( .IN1(n13465), .IN2(n13466), .QN(n12779) );
  INVX0 U13797 ( .INP(n13467), .ZN(n13466) );
  NOR2X0 U13798 ( .IN1(n13468), .IN2(n13469), .QN(n13467) );
  NAND2X0 U13799 ( .IN1(n13469), .IN2(n13468), .QN(n13465) );
  NOR2X0 U13800 ( .IN1(n13470), .IN2(n13471), .QN(n13468) );
  NOR2X0 U13801 ( .IN1(WX4768), .IN2(n8015), .QN(n13471) );
  INVX0 U13802 ( .INP(n13472), .ZN(n13470) );
  NAND2X0 U13803 ( .IN1(n8015), .IN2(WX4768), .QN(n13472) );
  NAND2X0 U13804 ( .IN1(n13473), .IN2(n13474), .QN(n13469) );
  NAND2X0 U13805 ( .IN1(n8014), .IN2(WX4640), .QN(n13474) );
  INVX0 U13806 ( .INP(n13475), .ZN(n13473) );
  NOR2X0 U13807 ( .IN1(WX4640), .IN2(n8014), .QN(n13475) );
  NAND2X0 U13808 ( .IN1(n9109), .IN2(n13476), .QN(n13463) );
  NAND2X0 U13809 ( .IN1(n519), .IN2(n9284), .QN(n13462) );
  NOR2X0 U13810 ( .IN1(n9237), .IN2(n8978), .QN(n519) );
  NAND2X0 U13811 ( .IN1(n9296), .IN2(CRC_OUT_7_5), .QN(n13461) );
  NAND4X0 U13812 ( .IN1(n13477), .IN2(n13478), .IN3(n13479), .IN4(n13480), 
        .QN(WX3280) );
  NAND3X0 U13813 ( .IN1(n13481), .IN2(n13482), .IN3(n9091), .QN(n13480) );
  NAND2X0 U13814 ( .IN1(n9326), .IN2(n12795), .QN(n13479) );
  NAND2X0 U13815 ( .IN1(n13483), .IN2(n13484), .QN(n12795) );
  INVX0 U13816 ( .INP(n13485), .ZN(n13484) );
  NOR2X0 U13817 ( .IN1(n13486), .IN2(n13487), .QN(n13485) );
  NAND2X0 U13818 ( .IN1(n13487), .IN2(n13486), .QN(n13483) );
  NOR2X0 U13819 ( .IN1(n13488), .IN2(n13489), .QN(n13486) );
  NOR2X0 U13820 ( .IN1(WX4766), .IN2(n8017), .QN(n13489) );
  INVX0 U13821 ( .INP(n13490), .ZN(n13488) );
  NAND2X0 U13822 ( .IN1(n8017), .IN2(WX4766), .QN(n13490) );
  NAND2X0 U13823 ( .IN1(n13491), .IN2(n13492), .QN(n13487) );
  NAND2X0 U13824 ( .IN1(n8016), .IN2(WX4638), .QN(n13492) );
  INVX0 U13825 ( .INP(n13493), .ZN(n13491) );
  NOR2X0 U13826 ( .IN1(WX4638), .IN2(n8016), .QN(n13493) );
  NAND2X0 U13827 ( .IN1(n518), .IN2(n9284), .QN(n13478) );
  NOR2X0 U13828 ( .IN1(n9237), .IN2(n8979), .QN(n518) );
  NAND2X0 U13829 ( .IN1(n9296), .IN2(CRC_OUT_7_6), .QN(n13477) );
  NAND4X0 U13830 ( .IN1(n13494), .IN2(n13495), .IN3(n13496), .IN4(n13497), 
        .QN(WX3278) );
  NAND2X0 U13831 ( .IN1(n9326), .IN2(n12811), .QN(n13497) );
  NAND2X0 U13832 ( .IN1(n13498), .IN2(n13499), .QN(n12811) );
  INVX0 U13833 ( .INP(n13500), .ZN(n13499) );
  NOR2X0 U13834 ( .IN1(n13501), .IN2(n13502), .QN(n13500) );
  NAND2X0 U13835 ( .IN1(n13502), .IN2(n13501), .QN(n13498) );
  NOR2X0 U13836 ( .IN1(n13503), .IN2(n13504), .QN(n13501) );
  NOR2X0 U13837 ( .IN1(WX4764), .IN2(n8019), .QN(n13504) );
  INVX0 U13838 ( .INP(n13505), .ZN(n13503) );
  NAND2X0 U13839 ( .IN1(n8019), .IN2(WX4764), .QN(n13505) );
  NAND2X0 U13840 ( .IN1(n13506), .IN2(n13507), .QN(n13502) );
  NAND2X0 U13841 ( .IN1(n8018), .IN2(WX4636), .QN(n13507) );
  INVX0 U13842 ( .INP(n13508), .ZN(n13506) );
  NOR2X0 U13843 ( .IN1(WX4636), .IN2(n8018), .QN(n13508) );
  NAND2X0 U13844 ( .IN1(n9109), .IN2(n13509), .QN(n13496) );
  NAND2X0 U13845 ( .IN1(n517), .IN2(n9284), .QN(n13495) );
  NOR2X0 U13846 ( .IN1(n9237), .IN2(n8980), .QN(n517) );
  NAND2X0 U13847 ( .IN1(n9296), .IN2(CRC_OUT_7_7), .QN(n13494) );
  NAND4X0 U13848 ( .IN1(n13510), .IN2(n13511), .IN3(n13512), .IN4(n13513), 
        .QN(WX3276) );
  NAND3X0 U13849 ( .IN1(n13514), .IN2(n13515), .IN3(n9090), .QN(n13513) );
  NAND2X0 U13850 ( .IN1(n9326), .IN2(n12827), .QN(n13512) );
  NAND2X0 U13851 ( .IN1(n13516), .IN2(n13517), .QN(n12827) );
  INVX0 U13852 ( .INP(n13518), .ZN(n13517) );
  NOR2X0 U13853 ( .IN1(n13519), .IN2(n13520), .QN(n13518) );
  NAND2X0 U13854 ( .IN1(n13520), .IN2(n13519), .QN(n13516) );
  NOR2X0 U13855 ( .IN1(n13521), .IN2(n13522), .QN(n13519) );
  NOR2X0 U13856 ( .IN1(WX4762), .IN2(n8021), .QN(n13522) );
  INVX0 U13857 ( .INP(n13523), .ZN(n13521) );
  NAND2X0 U13858 ( .IN1(n8021), .IN2(WX4762), .QN(n13523) );
  NAND2X0 U13859 ( .IN1(n13524), .IN2(n13525), .QN(n13520) );
  NAND2X0 U13860 ( .IN1(n8020), .IN2(WX4634), .QN(n13525) );
  INVX0 U13861 ( .INP(n13526), .ZN(n13524) );
  NOR2X0 U13862 ( .IN1(WX4634), .IN2(n8020), .QN(n13526) );
  NAND2X0 U13863 ( .IN1(n516), .IN2(n9284), .QN(n13511) );
  NOR2X0 U13864 ( .IN1(n9237), .IN2(n8981), .QN(n516) );
  NAND2X0 U13865 ( .IN1(n9296), .IN2(CRC_OUT_7_8), .QN(n13510) );
  NAND4X0 U13866 ( .IN1(n13527), .IN2(n13528), .IN3(n13529), .IN4(n13530), 
        .QN(WX3274) );
  NAND2X0 U13867 ( .IN1(n9326), .IN2(n12843), .QN(n13530) );
  NAND2X0 U13868 ( .IN1(n13531), .IN2(n13532), .QN(n12843) );
  INVX0 U13869 ( .INP(n13533), .ZN(n13532) );
  NOR2X0 U13870 ( .IN1(n13534), .IN2(n13535), .QN(n13533) );
  NAND2X0 U13871 ( .IN1(n13535), .IN2(n13534), .QN(n13531) );
  NOR2X0 U13872 ( .IN1(n13536), .IN2(n13537), .QN(n13534) );
  NOR2X0 U13873 ( .IN1(WX4760), .IN2(n8023), .QN(n13537) );
  INVX0 U13874 ( .INP(n13538), .ZN(n13536) );
  NAND2X0 U13875 ( .IN1(n8023), .IN2(WX4760), .QN(n13538) );
  NAND2X0 U13876 ( .IN1(n13539), .IN2(n13540), .QN(n13535) );
  NAND2X0 U13877 ( .IN1(n8022), .IN2(WX4632), .QN(n13540) );
  INVX0 U13878 ( .INP(n13541), .ZN(n13539) );
  NOR2X0 U13879 ( .IN1(WX4632), .IN2(n8022), .QN(n13541) );
  NAND2X0 U13880 ( .IN1(n9110), .IN2(n13542), .QN(n13529) );
  NAND2X0 U13881 ( .IN1(n515), .IN2(n9284), .QN(n13528) );
  NOR2X0 U13882 ( .IN1(n9238), .IN2(n8982), .QN(n515) );
  NAND2X0 U13883 ( .IN1(n9296), .IN2(CRC_OUT_7_9), .QN(n13527) );
  NAND4X0 U13884 ( .IN1(n13543), .IN2(n13544), .IN3(n13545), .IN4(n13546), 
        .QN(WX3272) );
  NAND2X0 U13885 ( .IN1(n9326), .IN2(n12859), .QN(n13546) );
  NAND2X0 U13886 ( .IN1(n13547), .IN2(n13548), .QN(n12859) );
  INVX0 U13887 ( .INP(n13549), .ZN(n13548) );
  NOR2X0 U13888 ( .IN1(n13550), .IN2(n13551), .QN(n13549) );
  NAND2X0 U13889 ( .IN1(n13551), .IN2(n13550), .QN(n13547) );
  NOR2X0 U13890 ( .IN1(n13552), .IN2(n13553), .QN(n13550) );
  NOR2X0 U13891 ( .IN1(WX4758), .IN2(n8025), .QN(n13553) );
  INVX0 U13892 ( .INP(n13554), .ZN(n13552) );
  NAND2X0 U13893 ( .IN1(n8025), .IN2(WX4758), .QN(n13554) );
  NAND2X0 U13894 ( .IN1(n13555), .IN2(n13556), .QN(n13551) );
  NAND2X0 U13895 ( .IN1(n8024), .IN2(WX4630), .QN(n13556) );
  INVX0 U13896 ( .INP(n13557), .ZN(n13555) );
  NOR2X0 U13897 ( .IN1(WX4630), .IN2(n8024), .QN(n13557) );
  NAND2X0 U13898 ( .IN1(n9109), .IN2(n13558), .QN(n13545) );
  NAND2X0 U13899 ( .IN1(n514), .IN2(n9284), .QN(n13544) );
  NOR2X0 U13900 ( .IN1(n9238), .IN2(n8983), .QN(n514) );
  NAND2X0 U13901 ( .IN1(test_so31), .IN2(n9315), .QN(n13543) );
  NAND4X0 U13902 ( .IN1(n13559), .IN2(n13560), .IN3(n13561), .IN4(n13562), 
        .QN(WX3270) );
  NAND3X0 U13903 ( .IN1(n12864), .IN2(n12865), .IN3(n9323), .QN(n13562) );
  NAND3X0 U13904 ( .IN1(n13563), .IN2(n13564), .IN3(n13565), .QN(n12865) );
  INVX0 U13905 ( .INP(n13566), .ZN(n13565) );
  NAND2X0 U13906 ( .IN1(n13566), .IN2(n13567), .QN(n12864) );
  NAND2X0 U13907 ( .IN1(n13563), .IN2(n13564), .QN(n13567) );
  NAND2X0 U13908 ( .IN1(n8027), .IN2(WX4628), .QN(n13564) );
  NAND2X0 U13909 ( .IN1(n3713), .IN2(WX4692), .QN(n13563) );
  NOR2X0 U13910 ( .IN1(n13568), .IN2(n13569), .QN(n13566) );
  NOR2X0 U13911 ( .IN1(n8797), .IN2(n8026), .QN(n13569) );
  INVX0 U13912 ( .INP(n13570), .ZN(n13568) );
  NAND2X0 U13913 ( .IN1(n8026), .IN2(n8797), .QN(n13570) );
  NAND2X0 U13914 ( .IN1(n9110), .IN2(n13571), .QN(n13561) );
  NAND2X0 U13915 ( .IN1(n513), .IN2(n9284), .QN(n13560) );
  NOR2X0 U13916 ( .IN1(n9238), .IN2(n8984), .QN(n513) );
  NAND2X0 U13917 ( .IN1(n9296), .IN2(CRC_OUT_7_11), .QN(n13559) );
  NAND4X0 U13918 ( .IN1(n13572), .IN2(n13573), .IN3(n13574), .IN4(n13575), 
        .QN(WX3268) );
  NAND3X0 U13919 ( .IN1(n13576), .IN2(n13577), .IN3(n9090), .QN(n13575) );
  NAND2X0 U13920 ( .IN1(n9326), .IN2(n12892), .QN(n13574) );
  NAND2X0 U13921 ( .IN1(n13578), .IN2(n13579), .QN(n12892) );
  INVX0 U13922 ( .INP(n13580), .ZN(n13579) );
  NOR2X0 U13923 ( .IN1(n13581), .IN2(n13582), .QN(n13580) );
  NAND2X0 U13924 ( .IN1(n13582), .IN2(n13581), .QN(n13578) );
  NOR2X0 U13925 ( .IN1(n13583), .IN2(n13584), .QN(n13581) );
  NOR2X0 U13926 ( .IN1(WX4754), .IN2(n8029), .QN(n13584) );
  INVX0 U13927 ( .INP(n13585), .ZN(n13583) );
  NAND2X0 U13928 ( .IN1(n8029), .IN2(WX4754), .QN(n13585) );
  NAND2X0 U13929 ( .IN1(n13586), .IN2(n13587), .QN(n13582) );
  NAND2X0 U13930 ( .IN1(n8028), .IN2(WX4626), .QN(n13587) );
  INVX0 U13931 ( .INP(n13588), .ZN(n13586) );
  NOR2X0 U13932 ( .IN1(WX4626), .IN2(n8028), .QN(n13588) );
  NAND2X0 U13933 ( .IN1(n512), .IN2(n9284), .QN(n13573) );
  NOR2X0 U13934 ( .IN1(n9238), .IN2(n8985), .QN(n512) );
  NAND2X0 U13935 ( .IN1(n9297), .IN2(CRC_OUT_7_12), .QN(n13572) );
  NAND4X0 U13936 ( .IN1(n13589), .IN2(n13590), .IN3(n13591), .IN4(n13592), 
        .QN(WX3266) );
  NAND3X0 U13937 ( .IN1(n12897), .IN2(n12898), .IN3(n9323), .QN(n13592) );
  NAND3X0 U13938 ( .IN1(n13593), .IN2(n13594), .IN3(n13595), .QN(n12898) );
  INVX0 U13939 ( .INP(n13596), .ZN(n13595) );
  NAND2X0 U13940 ( .IN1(n13596), .IN2(n13597), .QN(n12897) );
  NAND2X0 U13941 ( .IN1(n13593), .IN2(n13594), .QN(n13597) );
  NAND2X0 U13942 ( .IN1(n8416), .IN2(WX4624), .QN(n13594) );
  NAND2X0 U13943 ( .IN1(n3717), .IN2(WX4752), .QN(n13593) );
  NOR2X0 U13944 ( .IN1(n13598), .IN2(n13599), .QN(n13596) );
  INVX0 U13945 ( .INP(n13600), .ZN(n13599) );
  NAND2X0 U13946 ( .IN1(test_so39), .IN2(WX4560), .QN(n13600) );
  NOR2X0 U13947 ( .IN1(WX4560), .IN2(test_so39), .QN(n13598) );
  NAND2X0 U13948 ( .IN1(n9109), .IN2(n13601), .QN(n13591) );
  NAND2X0 U13949 ( .IN1(n511), .IN2(n9284), .QN(n13590) );
  NOR2X0 U13950 ( .IN1(n9238), .IN2(n8986), .QN(n511) );
  NAND2X0 U13951 ( .IN1(n9297), .IN2(CRC_OUT_7_13), .QN(n13589) );
  NAND4X0 U13952 ( .IN1(n13602), .IN2(n13603), .IN3(n13604), .IN4(n13605), 
        .QN(WX3264) );
  NAND2X0 U13953 ( .IN1(n9326), .IN2(n12925), .QN(n13605) );
  NAND2X0 U13954 ( .IN1(n13606), .IN2(n13607), .QN(n12925) );
  INVX0 U13955 ( .INP(n13608), .ZN(n13607) );
  NOR2X0 U13956 ( .IN1(n13609), .IN2(n13610), .QN(n13608) );
  NAND2X0 U13957 ( .IN1(n13610), .IN2(n13609), .QN(n13606) );
  NOR2X0 U13958 ( .IN1(n13611), .IN2(n13612), .QN(n13609) );
  NOR2X0 U13959 ( .IN1(WX4750), .IN2(n8032), .QN(n13612) );
  INVX0 U13960 ( .INP(n13613), .ZN(n13611) );
  NAND2X0 U13961 ( .IN1(n8032), .IN2(WX4750), .QN(n13613) );
  NAND2X0 U13962 ( .IN1(n13614), .IN2(n13615), .QN(n13610) );
  NAND2X0 U13963 ( .IN1(n8031), .IN2(WX4622), .QN(n13615) );
  INVX0 U13964 ( .INP(n13616), .ZN(n13614) );
  NOR2X0 U13965 ( .IN1(WX4622), .IN2(n8031), .QN(n13616) );
  NAND2X0 U13966 ( .IN1(n9110), .IN2(n13617), .QN(n13604) );
  NAND2X0 U13967 ( .IN1(n510), .IN2(n9284), .QN(n13603) );
  NOR2X0 U13968 ( .IN1(n9238), .IN2(n8987), .QN(n510) );
  NAND2X0 U13969 ( .IN1(n9297), .IN2(CRC_OUT_7_14), .QN(n13602) );
  NAND4X0 U13970 ( .IN1(n13618), .IN2(n13619), .IN3(n13620), .IN4(n13621), 
        .QN(WX3262) );
  NAND3X0 U13971 ( .IN1(n12930), .IN2(n12931), .IN3(n9322), .QN(n13621) );
  NAND3X0 U13972 ( .IN1(n13622), .IN2(n13623), .IN3(n13624), .QN(n12931) );
  INVX0 U13973 ( .INP(n13625), .ZN(n13624) );
  NAND2X0 U13974 ( .IN1(n13625), .IN2(n13626), .QN(n12930) );
  NAND2X0 U13975 ( .IN1(n13622), .IN2(n13623), .QN(n13626) );
  NAND2X0 U13976 ( .IN1(n8414), .IN2(WX4684), .QN(n13623) );
  NAND2X0 U13977 ( .IN1(n8034), .IN2(WX4748), .QN(n13622) );
  NOR2X0 U13978 ( .IN1(n13627), .IN2(n13628), .QN(n13625) );
  INVX0 U13979 ( .INP(n13629), .ZN(n13628) );
  NAND2X0 U13980 ( .IN1(test_so37), .IN2(WX4556), .QN(n13629) );
  NOR2X0 U13981 ( .IN1(WX4556), .IN2(test_so37), .QN(n13627) );
  NAND2X0 U13982 ( .IN1(n9110), .IN2(n13630), .QN(n13620) );
  NAND2X0 U13983 ( .IN1(n506), .IN2(n9284), .QN(n13619) );
  NOR2X0 U13984 ( .IN1(n9238), .IN2(n8988), .QN(n506) );
  NAND2X0 U13985 ( .IN1(n9297), .IN2(CRC_OUT_7_15), .QN(n13618) );
  NAND4X0 U13986 ( .IN1(n13631), .IN2(n13632), .IN3(n13633), .IN4(n13634), 
        .QN(WX3260) );
  NAND2X0 U13987 ( .IN1(n13635), .IN2(n12948), .QN(n13634) );
  NAND2X0 U13988 ( .IN1(n13636), .IN2(n12951), .QN(n12948) );
  NAND2X0 U13989 ( .IN1(n13637), .IN2(n13638), .QN(n13636) );
  NAND2X0 U13990 ( .IN1(n16351), .IN2(n9119), .QN(n13638) );
  NAND2X0 U13991 ( .IN1(TM1), .IN2(n8537), .QN(n13637) );
  NAND3X0 U13992 ( .IN1(n13639), .IN2(n13640), .IN3(n13641), .QN(n13635) );
  NAND2X0 U13993 ( .IN1(n9326), .IN2(n12951), .QN(n13641) );
  NAND2X0 U13994 ( .IN1(n13642), .IN2(n13643), .QN(n12951) );
  NAND2X0 U13995 ( .IN1(n7768), .IN2(n13644), .QN(n13643) );
  INVX0 U13996 ( .INP(n13645), .ZN(n13642) );
  NOR2X0 U13997 ( .IN1(n13644), .IN2(n7768), .QN(n13645) );
  NOR2X0 U13998 ( .IN1(n13646), .IN2(n13647), .QN(n13644) );
  NOR2X0 U13999 ( .IN1(WX4746), .IN2(n7769), .QN(n13647) );
  INVX0 U14000 ( .INP(n13648), .ZN(n13646) );
  NAND2X0 U14001 ( .IN1(n7769), .IN2(WX4746), .QN(n13648) );
  NAND2X0 U14002 ( .IN1(n10068), .IN2(n8537), .QN(n13640) );
  NAND2X0 U14003 ( .IN1(n16351), .IN2(n9079), .QN(n13639) );
  NAND2X0 U14004 ( .IN1(n13649), .IN2(n13650), .QN(n13633) );
  NAND2X0 U14005 ( .IN1(n13651), .IN2(n13652), .QN(n13649) );
  NAND2X0 U14006 ( .IN1(n9110), .IN2(n13653), .QN(n13652) );
  NAND2X0 U14007 ( .IN1(n8120), .IN2(n9111), .QN(n13651) );
  NAND2X0 U14008 ( .IN1(n505), .IN2(n9284), .QN(n13632) );
  NOR2X0 U14009 ( .IN1(n9238), .IN2(n8989), .QN(n505) );
  NAND2X0 U14010 ( .IN1(n9297), .IN2(CRC_OUT_7_16), .QN(n13631) );
  NAND4X0 U14011 ( .IN1(n13654), .IN2(n13655), .IN3(n13656), .IN4(n13657), 
        .QN(WX3258) );
  NAND2X0 U14012 ( .IN1(n13658), .IN2(n12984), .QN(n13657) );
  NAND3X0 U14013 ( .IN1(n13659), .IN2(n13660), .IN3(n12987), .QN(n12984) );
  NAND2X0 U14014 ( .IN1(n8413), .IN2(n9119), .QN(n13660) );
  NAND2X0 U14015 ( .IN1(TM1), .IN2(WX4744), .QN(n13659) );
  NAND3X0 U14016 ( .IN1(n13661), .IN2(n13662), .IN3(n13663), .QN(n13658) );
  NAND2X0 U14017 ( .IN1(n9326), .IN2(n12987), .QN(n13663) );
  NAND2X0 U14018 ( .IN1(n13664), .IN2(n13665), .QN(n12987) );
  NAND2X0 U14019 ( .IN1(n13666), .IN2(WX4680), .QN(n13665) );
  NAND2X0 U14020 ( .IN1(n13667), .IN2(n13668), .QN(n13666) );
  NAND3X0 U14021 ( .IN1(n13667), .IN2(n13668), .IN3(n7771), .QN(n13664) );
  NAND2X0 U14022 ( .IN1(test_so35), .IN2(WX4616), .QN(n13668) );
  NAND2X0 U14023 ( .IN1(n7770), .IN2(n8823), .QN(n13667) );
  NAND2X0 U14024 ( .IN1(n9080), .IN2(WX4744), .QN(n13662) );
  NAND2X0 U14025 ( .IN1(n9084), .IN2(n8413), .QN(n13661) );
  NAND2X0 U14026 ( .IN1(n13669), .IN2(n13670), .QN(n13656) );
  NAND2X0 U14027 ( .IN1(n13671), .IN2(n13672), .QN(n13669) );
  NAND2X0 U14028 ( .IN1(n9110), .IN2(n13673), .QN(n13672) );
  NAND2X0 U14029 ( .IN1(n9110), .IN2(n8597), .QN(n13671) );
  NAND2X0 U14030 ( .IN1(n504), .IN2(n9285), .QN(n13655) );
  NOR2X0 U14031 ( .IN1(n9238), .IN2(n8990), .QN(n504) );
  NAND2X0 U14032 ( .IN1(n9297), .IN2(CRC_OUT_7_17), .QN(n13654) );
  NAND4X0 U14033 ( .IN1(n13674), .IN2(n13675), .IN3(n13676), .IN4(n13677), 
        .QN(WX3256) );
  NAND2X0 U14034 ( .IN1(n13678), .IN2(n12993), .QN(n13677) );
  NAND2X0 U14035 ( .IN1(n13679), .IN2(n12996), .QN(n12993) );
  NAND2X0 U14036 ( .IN1(n13680), .IN2(n13681), .QN(n13679) );
  NAND2X0 U14037 ( .IN1(n16350), .IN2(n9121), .QN(n13681) );
  NAND2X0 U14038 ( .IN1(TM1), .IN2(n8540), .QN(n13680) );
  NAND3X0 U14039 ( .IN1(n13682), .IN2(n13683), .IN3(n13684), .QN(n13678) );
  NAND2X0 U14040 ( .IN1(n9326), .IN2(n12996), .QN(n13684) );
  NAND2X0 U14041 ( .IN1(n13685), .IN2(n13686), .QN(n12996) );
  NAND2X0 U14042 ( .IN1(n7772), .IN2(n13687), .QN(n13686) );
  INVX0 U14043 ( .INP(n13688), .ZN(n13685) );
  NOR2X0 U14044 ( .IN1(n13687), .IN2(n7772), .QN(n13688) );
  NOR2X0 U14045 ( .IN1(n13689), .IN2(n13690), .QN(n13687) );
  NOR2X0 U14046 ( .IN1(WX4742), .IN2(n7773), .QN(n13690) );
  INVX0 U14047 ( .INP(n13691), .ZN(n13689) );
  NAND2X0 U14048 ( .IN1(n7773), .IN2(WX4742), .QN(n13691) );
  NAND2X0 U14049 ( .IN1(n9083), .IN2(n8540), .QN(n13683) );
  NAND2X0 U14050 ( .IN1(n16350), .IN2(n9078), .QN(n13682) );
  NAND2X0 U14051 ( .IN1(n13692), .IN2(n13693), .QN(n13676) );
  NAND2X0 U14052 ( .IN1(n13694), .IN2(n13695), .QN(n13692) );
  NAND2X0 U14053 ( .IN1(n9109), .IN2(n13696), .QN(n13695) );
  NAND2X0 U14054 ( .IN1(n9110), .IN2(n8598), .QN(n13694) );
  NAND2X0 U14055 ( .IN1(n503), .IN2(n9285), .QN(n13675) );
  NOR2X0 U14056 ( .IN1(n9238), .IN2(n8991), .QN(n503) );
  NAND2X0 U14057 ( .IN1(n9297), .IN2(CRC_OUT_7_18), .QN(n13674) );
  NAND4X0 U14058 ( .IN1(n13697), .IN2(n13698), .IN3(n13699), .IN4(n13700), 
        .QN(WX3254) );
  NAND2X0 U14059 ( .IN1(n13701), .IN2(n13031), .QN(n13700) );
  NAND2X0 U14060 ( .IN1(n13702), .IN2(n13034), .QN(n13031) );
  NAND2X0 U14061 ( .IN1(n13703), .IN2(n13704), .QN(n13702) );
  NAND2X0 U14062 ( .IN1(n16349), .IN2(n9121), .QN(n13704) );
  NAND2X0 U14063 ( .IN1(TM1), .IN2(n8541), .QN(n13703) );
  NAND3X0 U14064 ( .IN1(n13705), .IN2(n13706), .IN3(n13707), .QN(n13701) );
  NAND2X0 U14065 ( .IN1(n9327), .IN2(n13034), .QN(n13707) );
  NAND2X0 U14066 ( .IN1(n13708), .IN2(n13709), .QN(n13034) );
  NAND2X0 U14067 ( .IN1(n7774), .IN2(n13710), .QN(n13709) );
  INVX0 U14068 ( .INP(n13711), .ZN(n13708) );
  NOR2X0 U14069 ( .IN1(n13710), .IN2(n7774), .QN(n13711) );
  NOR2X0 U14070 ( .IN1(n13712), .IN2(n13713), .QN(n13710) );
  NOR2X0 U14071 ( .IN1(WX4740), .IN2(n7775), .QN(n13713) );
  INVX0 U14072 ( .INP(n13714), .ZN(n13712) );
  NAND2X0 U14073 ( .IN1(n7775), .IN2(WX4740), .QN(n13714) );
  NAND2X0 U14074 ( .IN1(n9082), .IN2(n8541), .QN(n13706) );
  NAND2X0 U14075 ( .IN1(n16349), .IN2(n10069), .QN(n13705) );
  NAND2X0 U14076 ( .IN1(n13715), .IN2(n13716), .QN(n13699) );
  NAND2X0 U14077 ( .IN1(n13717), .IN2(n13718), .QN(n13715) );
  NAND2X0 U14078 ( .IN1(n9110), .IN2(n13719), .QN(n13718) );
  NAND2X0 U14079 ( .IN1(n9110), .IN2(n8599), .QN(n13717) );
  NAND2X0 U14080 ( .IN1(n502), .IN2(n9285), .QN(n13698) );
  NOR2X0 U14081 ( .IN1(n9238), .IN2(n8992), .QN(n502) );
  NAND2X0 U14082 ( .IN1(n9297), .IN2(CRC_OUT_7_19), .QN(n13697) );
  NAND4X0 U14083 ( .IN1(n13720), .IN2(n13721), .IN3(n13722), .IN4(n13723), 
        .QN(WX3252) );
  NAND2X0 U14084 ( .IN1(n13724), .IN2(n13040), .QN(n13723) );
  NAND2X0 U14085 ( .IN1(n13725), .IN2(n13043), .QN(n13040) );
  NAND2X0 U14086 ( .IN1(n13726), .IN2(n13727), .QN(n13725) );
  NAND2X0 U14087 ( .IN1(n16348), .IN2(n9121), .QN(n13727) );
  NAND2X0 U14088 ( .IN1(TM1), .IN2(n8542), .QN(n13726) );
  NAND3X0 U14089 ( .IN1(n13728), .IN2(n13729), .IN3(n13730), .QN(n13724) );
  NAND2X0 U14090 ( .IN1(n9327), .IN2(n13043), .QN(n13730) );
  NAND2X0 U14091 ( .IN1(n13731), .IN2(n13732), .QN(n13043) );
  NAND2X0 U14092 ( .IN1(n7776), .IN2(n13733), .QN(n13732) );
  INVX0 U14093 ( .INP(n13734), .ZN(n13731) );
  NOR2X0 U14094 ( .IN1(n13733), .IN2(n7776), .QN(n13734) );
  NOR2X0 U14095 ( .IN1(n13735), .IN2(n13736), .QN(n13733) );
  NOR2X0 U14096 ( .IN1(WX4738), .IN2(n7777), .QN(n13736) );
  INVX0 U14097 ( .INP(n13737), .ZN(n13735) );
  NAND2X0 U14098 ( .IN1(n7777), .IN2(WX4738), .QN(n13737) );
  NAND2X0 U14099 ( .IN1(n10068), .IN2(n8542), .QN(n13729) );
  NAND2X0 U14100 ( .IN1(n16348), .IN2(n9080), .QN(n13728) );
  NAND2X0 U14101 ( .IN1(n13738), .IN2(n13739), .QN(n13722) );
  NAND2X0 U14102 ( .IN1(n13740), .IN2(n13741), .QN(n13738) );
  NAND2X0 U14103 ( .IN1(n9109), .IN2(n13742), .QN(n13741) );
  NAND2X0 U14104 ( .IN1(n9106), .IN2(n8600), .QN(n13740) );
  NAND2X0 U14105 ( .IN1(n501), .IN2(n9285), .QN(n13721) );
  NOR2X0 U14106 ( .IN1(n9072), .IN2(n9159), .QN(n501) );
  NAND2X0 U14107 ( .IN1(n9297), .IN2(CRC_OUT_7_20), .QN(n13720) );
  NAND4X0 U14108 ( .IN1(n13743), .IN2(n13744), .IN3(n13745), .IN4(n13746), 
        .QN(WX3250) );
  NAND2X0 U14109 ( .IN1(n13747), .IN2(n13078), .QN(n13746) );
  NAND2X0 U14110 ( .IN1(n13748), .IN2(n13081), .QN(n13078) );
  NAND2X0 U14111 ( .IN1(n13749), .IN2(n13750), .QN(n13748) );
  NAND2X0 U14112 ( .IN1(n16347), .IN2(n9121), .QN(n13750) );
  NAND2X0 U14113 ( .IN1(TM1), .IN2(n8543), .QN(n13749) );
  NAND3X0 U14114 ( .IN1(n13751), .IN2(n13752), .IN3(n13753), .QN(n13747) );
  NAND2X0 U14115 ( .IN1(n9327), .IN2(n13081), .QN(n13753) );
  NAND2X0 U14116 ( .IN1(n13754), .IN2(n13755), .QN(n13081) );
  NAND2X0 U14117 ( .IN1(n7778), .IN2(n13756), .QN(n13755) );
  INVX0 U14118 ( .INP(n13757), .ZN(n13754) );
  NOR2X0 U14119 ( .IN1(n13756), .IN2(n7778), .QN(n13757) );
  NOR2X0 U14120 ( .IN1(n13758), .IN2(n13759), .QN(n13756) );
  NOR2X0 U14121 ( .IN1(WX4736), .IN2(n7779), .QN(n13759) );
  INVX0 U14122 ( .INP(n13760), .ZN(n13758) );
  NAND2X0 U14123 ( .IN1(n7779), .IN2(WX4736), .QN(n13760) );
  NAND2X0 U14124 ( .IN1(n9084), .IN2(n8543), .QN(n13752) );
  NAND2X0 U14125 ( .IN1(n16347), .IN2(n9079), .QN(n13751) );
  NAND2X0 U14126 ( .IN1(n13761), .IN2(n13762), .QN(n13745) );
  NAND2X0 U14127 ( .IN1(n13763), .IN2(n13764), .QN(n13761) );
  NAND2X0 U14128 ( .IN1(n9106), .IN2(n13765), .QN(n13764) );
  NAND2X0 U14129 ( .IN1(n9106), .IN2(n8601), .QN(n13763) );
  NAND2X0 U14130 ( .IN1(n500), .IN2(n9285), .QN(n13744) );
  NOR2X0 U14131 ( .IN1(n9238), .IN2(n8993), .QN(n500) );
  NAND2X0 U14132 ( .IN1(n9297), .IN2(CRC_OUT_7_21), .QN(n13743) );
  NAND4X0 U14133 ( .IN1(n13766), .IN2(n13767), .IN3(n13768), .IN4(n13769), 
        .QN(WX3248) );
  NAND2X0 U14134 ( .IN1(n13770), .IN2(n13098), .QN(n13769) );
  NAND2X0 U14135 ( .IN1(n13771), .IN2(n13101), .QN(n13098) );
  NAND2X0 U14136 ( .IN1(n13772), .IN2(n13773), .QN(n13771) );
  NAND2X0 U14137 ( .IN1(n16346), .IN2(n9121), .QN(n13773) );
  NAND2X0 U14138 ( .IN1(TM1), .IN2(n8544), .QN(n13772) );
  NAND3X0 U14139 ( .IN1(n13774), .IN2(n13775), .IN3(n13776), .QN(n13770) );
  NAND2X0 U14140 ( .IN1(n9327), .IN2(n13101), .QN(n13776) );
  NAND2X0 U14141 ( .IN1(n13777), .IN2(n13778), .QN(n13101) );
  NAND2X0 U14142 ( .IN1(n7780), .IN2(n13779), .QN(n13778) );
  INVX0 U14143 ( .INP(n13780), .ZN(n13777) );
  NOR2X0 U14144 ( .IN1(n13779), .IN2(n7780), .QN(n13780) );
  NOR2X0 U14145 ( .IN1(n13781), .IN2(n13782), .QN(n13779) );
  NOR2X0 U14146 ( .IN1(WX4734), .IN2(n7781), .QN(n13782) );
  INVX0 U14147 ( .INP(n13783), .ZN(n13781) );
  NAND2X0 U14148 ( .IN1(n7781), .IN2(WX4734), .QN(n13783) );
  NAND2X0 U14149 ( .IN1(n9083), .IN2(n8544), .QN(n13775) );
  NAND2X0 U14150 ( .IN1(n16346), .IN2(n9078), .QN(n13774) );
  NAND2X0 U14151 ( .IN1(n13784), .IN2(n13785), .QN(n13768) );
  NAND2X0 U14152 ( .IN1(n13786), .IN2(n13787), .QN(n13784) );
  NAND2X0 U14153 ( .IN1(n9106), .IN2(n13788), .QN(n13787) );
  NAND2X0 U14154 ( .IN1(n9106), .IN2(n8602), .QN(n13786) );
  NAND2X0 U14155 ( .IN1(n499), .IN2(n9285), .QN(n13767) );
  NOR2X0 U14156 ( .IN1(n9238), .IN2(n8994), .QN(n499) );
  NAND2X0 U14157 ( .IN1(n9297), .IN2(CRC_OUT_7_22), .QN(n13766) );
  NAND4X0 U14158 ( .IN1(n13789), .IN2(n13790), .IN3(n13791), .IN4(n13792), 
        .QN(WX3246) );
  NAND2X0 U14159 ( .IN1(n13793), .IN2(n13121), .QN(n13792) );
  NAND2X0 U14160 ( .IN1(n13794), .IN2(n13124), .QN(n13121) );
  NAND2X0 U14161 ( .IN1(n13795), .IN2(n13796), .QN(n13794) );
  NAND2X0 U14162 ( .IN1(n16345), .IN2(n9121), .QN(n13796) );
  NAND2X0 U14163 ( .IN1(TM1), .IN2(n8545), .QN(n13795) );
  NAND3X0 U14164 ( .IN1(n13797), .IN2(n13798), .IN3(n13799), .QN(n13793) );
  NAND2X0 U14165 ( .IN1(n9329), .IN2(n13124), .QN(n13799) );
  NAND2X0 U14166 ( .IN1(n13800), .IN2(n13801), .QN(n13124) );
  NAND2X0 U14167 ( .IN1(n7782), .IN2(n13802), .QN(n13801) );
  INVX0 U14168 ( .INP(n13803), .ZN(n13800) );
  NOR2X0 U14169 ( .IN1(n13802), .IN2(n7782), .QN(n13803) );
  NOR2X0 U14170 ( .IN1(n13804), .IN2(n13805), .QN(n13802) );
  NOR2X0 U14171 ( .IN1(WX4732), .IN2(n7783), .QN(n13805) );
  INVX0 U14172 ( .INP(n13806), .ZN(n13804) );
  NAND2X0 U14173 ( .IN1(n7783), .IN2(WX4732), .QN(n13806) );
  NAND2X0 U14174 ( .IN1(n9082), .IN2(n8545), .QN(n13798) );
  NAND2X0 U14175 ( .IN1(n16345), .IN2(n10069), .QN(n13797) );
  NAND2X0 U14176 ( .IN1(n13807), .IN2(n9112), .QN(n13791) );
  NAND2X0 U14177 ( .IN1(n498), .IN2(n9285), .QN(n13790) );
  NOR2X0 U14178 ( .IN1(n9238), .IN2(n8995), .QN(n498) );
  NAND2X0 U14179 ( .IN1(n9303), .IN2(CRC_OUT_7_23), .QN(n13789) );
  NAND4X0 U14180 ( .IN1(n13808), .IN2(n13809), .IN3(n13810), .IN4(n13811), 
        .QN(WX3244) );
  NAND2X0 U14181 ( .IN1(n13812), .IN2(n13144), .QN(n13811) );
  NAND2X0 U14182 ( .IN1(n13813), .IN2(n13147), .QN(n13144) );
  NAND2X0 U14183 ( .IN1(n13814), .IN2(n13815), .QN(n13813) );
  NAND2X0 U14184 ( .IN1(n16344), .IN2(n9121), .QN(n13815) );
  NAND2X0 U14185 ( .IN1(TM1), .IN2(n8546), .QN(n13814) );
  NAND3X0 U14186 ( .IN1(n13816), .IN2(n13817), .IN3(n13818), .QN(n13812) );
  NAND2X0 U14187 ( .IN1(n9327), .IN2(n13147), .QN(n13818) );
  NAND2X0 U14188 ( .IN1(n13819), .IN2(n13820), .QN(n13147) );
  NAND2X0 U14189 ( .IN1(n7784), .IN2(n13821), .QN(n13820) );
  INVX0 U14190 ( .INP(n13822), .ZN(n13819) );
  NOR2X0 U14191 ( .IN1(n13821), .IN2(n7784), .QN(n13822) );
  NOR2X0 U14192 ( .IN1(n13823), .IN2(n13824), .QN(n13821) );
  NOR2X0 U14193 ( .IN1(WX4730), .IN2(n7785), .QN(n13824) );
  INVX0 U14194 ( .INP(n13825), .ZN(n13823) );
  NAND2X0 U14195 ( .IN1(n7785), .IN2(WX4730), .QN(n13825) );
  NAND2X0 U14196 ( .IN1(n10068), .IN2(n8546), .QN(n13817) );
  NAND2X0 U14197 ( .IN1(n16344), .IN2(n9080), .QN(n13816) );
  NAND2X0 U14198 ( .IN1(n13826), .IN2(n13827), .QN(n13810) );
  NAND2X0 U14199 ( .IN1(n13828), .IN2(n13829), .QN(n13826) );
  NAND2X0 U14200 ( .IN1(n9106), .IN2(n13830), .QN(n13829) );
  NAND2X0 U14201 ( .IN1(n9106), .IN2(n8604), .QN(n13828) );
  NAND2X0 U14202 ( .IN1(n497), .IN2(n9285), .QN(n13809) );
  NOR2X0 U14203 ( .IN1(n9238), .IN2(n8996), .QN(n497) );
  NAND2X0 U14204 ( .IN1(n9298), .IN2(CRC_OUT_7_24), .QN(n13808) );
  NAND4X0 U14205 ( .IN1(n13831), .IN2(n13832), .IN3(n13833), .IN4(n13834), 
        .QN(WX3242) );
  NAND2X0 U14206 ( .IN1(n13835), .IN2(n13167), .QN(n13834) );
  NAND2X0 U14207 ( .IN1(n13836), .IN2(n13170), .QN(n13167) );
  NAND2X0 U14208 ( .IN1(n13837), .IN2(n13838), .QN(n13836) );
  NAND2X0 U14209 ( .IN1(n16343), .IN2(n9121), .QN(n13838) );
  NAND2X0 U14210 ( .IN1(TM1), .IN2(n8547), .QN(n13837) );
  NAND3X0 U14211 ( .IN1(n13839), .IN2(n13840), .IN3(n13841), .QN(n13835) );
  NAND2X0 U14212 ( .IN1(n9327), .IN2(n13170), .QN(n13841) );
  NAND2X0 U14213 ( .IN1(n13842), .IN2(n13843), .QN(n13170) );
  NAND2X0 U14214 ( .IN1(n7786), .IN2(n13844), .QN(n13843) );
  INVX0 U14215 ( .INP(n13845), .ZN(n13842) );
  NOR2X0 U14216 ( .IN1(n13844), .IN2(n7786), .QN(n13845) );
  NOR2X0 U14217 ( .IN1(n13846), .IN2(n13847), .QN(n13844) );
  NOR2X0 U14218 ( .IN1(WX4728), .IN2(n7787), .QN(n13847) );
  INVX0 U14219 ( .INP(n13848), .ZN(n13846) );
  NAND2X0 U14220 ( .IN1(n7787), .IN2(WX4728), .QN(n13848) );
  NAND2X0 U14221 ( .IN1(n9084), .IN2(n8547), .QN(n13840) );
  NAND2X0 U14222 ( .IN1(n16343), .IN2(n9079), .QN(n13839) );
  NAND2X0 U14223 ( .IN1(n13849), .IN2(n13850), .QN(n13833) );
  NAND2X0 U14224 ( .IN1(n13851), .IN2(n13852), .QN(n13849) );
  NAND2X0 U14225 ( .IN1(n9106), .IN2(n13853), .QN(n13852) );
  NAND2X0 U14226 ( .IN1(n9106), .IN2(n8605), .QN(n13851) );
  NAND2X0 U14227 ( .IN1(n496), .IN2(n9285), .QN(n13832) );
  NOR2X0 U14228 ( .IN1(n9239), .IN2(n8997), .QN(n496) );
  NAND2X0 U14229 ( .IN1(n9298), .IN2(CRC_OUT_7_25), .QN(n13831) );
  NAND4X0 U14230 ( .IN1(n13854), .IN2(n13855), .IN3(n13856), .IN4(n13857), 
        .QN(WX3240) );
  NAND2X0 U14231 ( .IN1(n13858), .IN2(n13190), .QN(n13857) );
  NAND2X0 U14232 ( .IN1(n13859), .IN2(n13193), .QN(n13190) );
  NAND2X0 U14233 ( .IN1(n13860), .IN2(n13861), .QN(n13859) );
  NAND2X0 U14234 ( .IN1(n16342), .IN2(n9121), .QN(n13861) );
  NAND2X0 U14235 ( .IN1(TM1), .IN2(n8548), .QN(n13860) );
  NAND3X0 U14236 ( .IN1(n13862), .IN2(n13863), .IN3(n13864), .QN(n13858) );
  NAND2X0 U14237 ( .IN1(n9327), .IN2(n13193), .QN(n13864) );
  NAND2X0 U14238 ( .IN1(n13865), .IN2(n13866), .QN(n13193) );
  NAND2X0 U14239 ( .IN1(n7788), .IN2(n13867), .QN(n13866) );
  INVX0 U14240 ( .INP(n13868), .ZN(n13865) );
  NOR2X0 U14241 ( .IN1(n13867), .IN2(n7788), .QN(n13868) );
  NOR2X0 U14242 ( .IN1(n13869), .IN2(n13870), .QN(n13867) );
  NOR2X0 U14243 ( .IN1(WX4726), .IN2(n7789), .QN(n13870) );
  INVX0 U14244 ( .INP(n13871), .ZN(n13869) );
  NAND2X0 U14245 ( .IN1(n7789), .IN2(WX4726), .QN(n13871) );
  NAND2X0 U14246 ( .IN1(n9083), .IN2(n8548), .QN(n13863) );
  NAND2X0 U14247 ( .IN1(n16342), .IN2(n9078), .QN(n13862) );
  NAND2X0 U14248 ( .IN1(n13872), .IN2(n9112), .QN(n13856) );
  NAND2X0 U14249 ( .IN1(n495), .IN2(n9285), .QN(n13855) );
  NOR2X0 U14250 ( .IN1(n9239), .IN2(n8998), .QN(n495) );
  NAND2X0 U14251 ( .IN1(n9298), .IN2(CRC_OUT_7_26), .QN(n13854) );
  NAND4X0 U14252 ( .IN1(n13873), .IN2(n13874), .IN3(n13875), .IN4(n13876), 
        .QN(WX3238) );
  NAND2X0 U14253 ( .IN1(n13877), .IN2(n13213), .QN(n13876) );
  NAND2X0 U14254 ( .IN1(n13878), .IN2(n13216), .QN(n13213) );
  NAND2X0 U14255 ( .IN1(n13879), .IN2(n13880), .QN(n13878) );
  NAND2X0 U14256 ( .IN1(n16341), .IN2(n9121), .QN(n13880) );
  NAND2X0 U14257 ( .IN1(TM1), .IN2(n8549), .QN(n13879) );
  NAND3X0 U14258 ( .IN1(n13881), .IN2(n13882), .IN3(n13883), .QN(n13877) );
  NAND2X0 U14259 ( .IN1(n9327), .IN2(n13216), .QN(n13883) );
  NAND2X0 U14260 ( .IN1(n13884), .IN2(n13885), .QN(n13216) );
  NAND2X0 U14261 ( .IN1(n7790), .IN2(n13886), .QN(n13885) );
  INVX0 U14262 ( .INP(n13887), .ZN(n13884) );
  NOR2X0 U14263 ( .IN1(n13886), .IN2(n7790), .QN(n13887) );
  NOR2X0 U14264 ( .IN1(n13888), .IN2(n13889), .QN(n13886) );
  NOR2X0 U14265 ( .IN1(WX4724), .IN2(n7791), .QN(n13889) );
  INVX0 U14266 ( .INP(n13890), .ZN(n13888) );
  NAND2X0 U14267 ( .IN1(n7791), .IN2(WX4724), .QN(n13890) );
  NAND2X0 U14268 ( .IN1(n9082), .IN2(n8549), .QN(n13882) );
  NAND2X0 U14269 ( .IN1(n16341), .IN2(n10069), .QN(n13881) );
  NAND2X0 U14270 ( .IN1(n13891), .IN2(n13892), .QN(n13875) );
  NAND2X0 U14271 ( .IN1(n13893), .IN2(n13894), .QN(n13891) );
  NAND2X0 U14272 ( .IN1(n9106), .IN2(n13895), .QN(n13894) );
  NAND2X0 U14273 ( .IN1(n9106), .IN2(n8607), .QN(n13893) );
  NAND2X0 U14274 ( .IN1(n494), .IN2(n9285), .QN(n13874) );
  NOR2X0 U14275 ( .IN1(n9239), .IN2(n8999), .QN(n494) );
  NAND2X0 U14276 ( .IN1(test_so32), .IN2(n9314), .QN(n13873) );
  NAND4X0 U14277 ( .IN1(n13896), .IN2(n13897), .IN3(n13898), .IN4(n13899), 
        .QN(WX3236) );
  NAND2X0 U14278 ( .IN1(n13900), .IN2(n13901), .QN(n13899) );
  NAND2X0 U14279 ( .IN1(n13902), .IN2(n13903), .QN(n13900) );
  NAND2X0 U14280 ( .IN1(n9105), .IN2(n13904), .QN(n13903) );
  NAND2X0 U14281 ( .IN1(n9105), .IN2(n8608), .QN(n13902) );
  NAND2X0 U14282 ( .IN1(n13235), .IN2(n9336), .QN(n13898) );
  NOR2X0 U14283 ( .IN1(n13905), .IN2(n13906), .QN(n13235) );
  INVX0 U14284 ( .INP(n13907), .ZN(n13906) );
  NAND2X0 U14285 ( .IN1(n13908), .IN2(n13909), .QN(n13907) );
  NOR2X0 U14286 ( .IN1(n13909), .IN2(n13908), .QN(n13905) );
  NAND2X0 U14287 ( .IN1(n13910), .IN2(n13911), .QN(n13908) );
  NAND2X0 U14288 ( .IN1(n13912), .IN2(WX4658), .QN(n13911) );
  NAND2X0 U14289 ( .IN1(n13913), .IN2(n13914), .QN(n13912) );
  NAND3X0 U14290 ( .IN1(n13913), .IN2(n13914), .IN3(n7793), .QN(n13910) );
  NAND2X0 U14291 ( .IN1(test_so40), .IN2(WX4594), .QN(n13914) );
  NAND2X0 U14292 ( .IN1(n7792), .IN2(n8801), .QN(n13913) );
  NOR2X0 U14293 ( .IN1(n13915), .IN2(n13916), .QN(n13909) );
  INVX0 U14294 ( .INP(n13917), .ZN(n13916) );
  NAND2X0 U14295 ( .IN1(n16340), .IN2(n9121), .QN(n13917) );
  NOR2X0 U14296 ( .IN1(n9117), .IN2(n16340), .QN(n13915) );
  NAND2X0 U14297 ( .IN1(n493), .IN2(n9285), .QN(n13897) );
  NOR2X0 U14298 ( .IN1(n9239), .IN2(n9000), .QN(n493) );
  NAND2X0 U14299 ( .IN1(n9298), .IN2(CRC_OUT_7_28), .QN(n13896) );
  NAND4X0 U14300 ( .IN1(n13918), .IN2(n13919), .IN3(n13920), .IN4(n13921), 
        .QN(WX3234) );
  NAND2X0 U14301 ( .IN1(n13922), .IN2(n13255), .QN(n13921) );
  NAND2X0 U14302 ( .IN1(n13923), .IN2(n13258), .QN(n13255) );
  NAND2X0 U14303 ( .IN1(n13924), .IN2(n13925), .QN(n13923) );
  NAND2X0 U14304 ( .IN1(n16339), .IN2(n9121), .QN(n13925) );
  NAND2X0 U14305 ( .IN1(TM1), .IN2(n8551), .QN(n13924) );
  NAND3X0 U14306 ( .IN1(n13926), .IN2(n13927), .IN3(n13928), .QN(n13922) );
  NAND2X0 U14307 ( .IN1(n9327), .IN2(n13258), .QN(n13928) );
  NAND2X0 U14308 ( .IN1(n13929), .IN2(n13930), .QN(n13258) );
  NAND2X0 U14309 ( .IN1(n7794), .IN2(n13931), .QN(n13930) );
  INVX0 U14310 ( .INP(n13932), .ZN(n13929) );
  NOR2X0 U14311 ( .IN1(n13931), .IN2(n7794), .QN(n13932) );
  NOR2X0 U14312 ( .IN1(n13933), .IN2(n13934), .QN(n13931) );
  NOR2X0 U14313 ( .IN1(WX4720), .IN2(n7795), .QN(n13934) );
  INVX0 U14314 ( .INP(n13935), .ZN(n13933) );
  NAND2X0 U14315 ( .IN1(n7795), .IN2(WX4720), .QN(n13935) );
  NAND2X0 U14316 ( .IN1(n10068), .IN2(n8551), .QN(n13927) );
  NAND2X0 U14317 ( .IN1(n16339), .IN2(n9080), .QN(n13926) );
  NAND2X0 U14318 ( .IN1(n13936), .IN2(n13937), .QN(n13920) );
  NAND2X0 U14319 ( .IN1(n13938), .IN2(n13939), .QN(n13936) );
  NAND2X0 U14320 ( .IN1(n9105), .IN2(n13940), .QN(n13939) );
  NAND2X0 U14321 ( .IN1(n9105), .IN2(n8609), .QN(n13938) );
  NAND2X0 U14322 ( .IN1(n492), .IN2(n9285), .QN(n13919) );
  NOR2X0 U14323 ( .IN1(n9239), .IN2(n9001), .QN(n492) );
  NAND2X0 U14324 ( .IN1(n9298), .IN2(CRC_OUT_7_29), .QN(n13918) );
  NAND4X0 U14325 ( .IN1(n13941), .IN2(n13942), .IN3(n13943), .IN4(n13944), 
        .QN(WX3232) );
  NAND2X0 U14326 ( .IN1(n13277), .IN2(n9336), .QN(n13944) );
  NOR2X0 U14327 ( .IN1(n13945), .IN2(n13946), .QN(n13277) );
  INVX0 U14328 ( .INP(n13947), .ZN(n13946) );
  NAND2X0 U14329 ( .IN1(n13948), .IN2(n13949), .QN(n13947) );
  NOR2X0 U14330 ( .IN1(n13949), .IN2(n13948), .QN(n13945) );
  NAND2X0 U14331 ( .IN1(n13950), .IN2(n13951), .QN(n13948) );
  NAND2X0 U14332 ( .IN1(n8356), .IN2(n13952), .QN(n13951) );
  INVX0 U14333 ( .INP(n13953), .ZN(n13952) );
  NAND2X0 U14334 ( .IN1(n13953), .IN2(WX4718), .QN(n13950) );
  NAND2X0 U14335 ( .IN1(n13954), .IN2(n13955), .QN(n13953) );
  INVX0 U14336 ( .INP(n13956), .ZN(n13955) );
  NOR2X0 U14337 ( .IN1(n8814), .IN2(n16338), .QN(n13956) );
  NAND2X0 U14338 ( .IN1(n16338), .IN2(n8814), .QN(n13954) );
  NOR2X0 U14339 ( .IN1(n13957), .IN2(n13958), .QN(n13949) );
  INVX0 U14340 ( .INP(n13959), .ZN(n13958) );
  NAND2X0 U14341 ( .IN1(n7796), .IN2(n9121), .QN(n13959) );
  NOR2X0 U14342 ( .IN1(n9117), .IN2(n7796), .QN(n13957) );
  NAND2X0 U14343 ( .IN1(n13960), .IN2(n9111), .QN(n13943) );
  NAND2X0 U14344 ( .IN1(n491), .IN2(n9285), .QN(n13942) );
  NOR2X0 U14345 ( .IN1(n9239), .IN2(n9002), .QN(n491) );
  NAND2X0 U14346 ( .IN1(n9298), .IN2(CRC_OUT_7_30), .QN(n13941) );
  NAND4X0 U14347 ( .IN1(n13961), .IN2(n13962), .IN3(n13963), .IN4(n13964), 
        .QN(WX3230) );
  NAND2X0 U14348 ( .IN1(n13965), .IN2(n13297), .QN(n13964) );
  NAND2X0 U14349 ( .IN1(n13966), .IN2(n13300), .QN(n13297) );
  NAND2X0 U14350 ( .IN1(n13967), .IN2(n13968), .QN(n13966) );
  NAND2X0 U14351 ( .IN1(n16337), .IN2(n9121), .QN(n13968) );
  NAND2X0 U14352 ( .IN1(TM1), .IN2(n8553), .QN(n13967) );
  NAND3X0 U14353 ( .IN1(n13969), .IN2(n13970), .IN3(n13971), .QN(n13965) );
  NAND2X0 U14354 ( .IN1(n9327), .IN2(n13300), .QN(n13971) );
  NAND2X0 U14355 ( .IN1(n13972), .IN2(n13973), .QN(n13300) );
  NAND2X0 U14356 ( .IN1(n7622), .IN2(n13974), .QN(n13973) );
  INVX0 U14357 ( .INP(n13975), .ZN(n13972) );
  NOR2X0 U14358 ( .IN1(n13974), .IN2(n7622), .QN(n13975) );
  NOR2X0 U14359 ( .IN1(n13976), .IN2(n13977), .QN(n13974) );
  NOR2X0 U14360 ( .IN1(WX4716), .IN2(n7623), .QN(n13977) );
  INVX0 U14361 ( .INP(n13978), .ZN(n13976) );
  NAND2X0 U14362 ( .IN1(n7623), .IN2(WX4716), .QN(n13978) );
  NAND2X0 U14363 ( .IN1(n9084), .IN2(n8553), .QN(n13970) );
  NAND2X0 U14364 ( .IN1(n16337), .IN2(n9079), .QN(n13969) );
  NAND2X0 U14365 ( .IN1(n13979), .IN2(n13980), .QN(n13963) );
  NAND2X0 U14366 ( .IN1(n13981), .IN2(n13982), .QN(n13979) );
  NAND2X0 U14367 ( .IN1(n9105), .IN2(n13983), .QN(n13982) );
  NAND2X0 U14368 ( .IN1(n9105), .IN2(n8611), .QN(n13981) );
  NAND2X0 U14369 ( .IN1(n9298), .IN2(CRC_OUT_7_31), .QN(n13962) );
  NAND2X0 U14370 ( .IN1(n2245), .IN2(WX3071), .QN(n13961) );
  NOR2X0 U14371 ( .IN1(n9239), .IN2(WX3071), .QN(WX3132) );
  NOR3X0 U14372 ( .IN1(n9136), .IN2(n13984), .IN3(n13985), .QN(WX2619) );
  NOR2X0 U14373 ( .IN1(n8574), .IN2(CRC_OUT_8_30), .QN(n13985) );
  NOR2X0 U14374 ( .IN1(DFF_382_n1), .IN2(WX2130), .QN(n13984) );
  NOR3X0 U14375 ( .IN1(n9136), .IN2(n13986), .IN3(n13987), .QN(WX2617) );
  NOR2X0 U14376 ( .IN1(n8575), .IN2(CRC_OUT_8_29), .QN(n13987) );
  NOR2X0 U14377 ( .IN1(DFF_381_n1), .IN2(WX2132), .QN(n13986) );
  NOR3X0 U14378 ( .IN1(n9136), .IN2(n13988), .IN3(n13989), .QN(WX2615) );
  NOR2X0 U14379 ( .IN1(n8587), .IN2(CRC_OUT_8_28), .QN(n13989) );
  NOR2X0 U14380 ( .IN1(DFF_380_n1), .IN2(WX2134), .QN(n13988) );
  NOR2X0 U14381 ( .IN1(n9239), .IN2(n13990), .QN(WX2613) );
  NOR2X0 U14382 ( .IN1(n13991), .IN2(n13992), .QN(n13990) );
  NOR2X0 U14383 ( .IN1(test_so18), .IN2(CRC_OUT_8_27), .QN(n13992) );
  NOR2X0 U14384 ( .IN1(DFF_379_n1), .IN2(n8803), .QN(n13991) );
  NOR3X0 U14385 ( .IN1(n9141), .IN2(n13993), .IN3(n13994), .QN(WX2611) );
  NOR2X0 U14386 ( .IN1(n8588), .IN2(CRC_OUT_8_26), .QN(n13994) );
  NOR2X0 U14387 ( .IN1(DFF_378_n1), .IN2(WX2138), .QN(n13993) );
  NOR2X0 U14388 ( .IN1(n9239), .IN2(n13995), .QN(WX2609) );
  NOR2X0 U14389 ( .IN1(n13996), .IN2(n13997), .QN(n13995) );
  NOR2X0 U14390 ( .IN1(test_so21), .IN2(WX2140), .QN(n13997) );
  INVX0 U14391 ( .INP(n13998), .ZN(n13996) );
  NAND2X0 U14392 ( .IN1(WX2140), .IN2(test_so21), .QN(n13998) );
  NOR3X0 U14393 ( .IN1(n9155), .IN2(n13999), .IN3(n14000), .QN(WX2607) );
  NOR2X0 U14394 ( .IN1(n8590), .IN2(CRC_OUT_8_24), .QN(n14000) );
  NOR2X0 U14395 ( .IN1(DFF_376_n1), .IN2(WX2142), .QN(n13999) );
  NOR3X0 U14396 ( .IN1(n9155), .IN2(n14001), .IN3(n14002), .QN(WX2605) );
  NOR2X0 U14397 ( .IN1(n8591), .IN2(CRC_OUT_8_23), .QN(n14002) );
  NOR2X0 U14398 ( .IN1(DFF_375_n1), .IN2(WX2144), .QN(n14001) );
  NOR3X0 U14399 ( .IN1(n9155), .IN2(n14003), .IN3(n14004), .QN(WX2603) );
  NOR2X0 U14400 ( .IN1(n8592), .IN2(CRC_OUT_8_22), .QN(n14004) );
  NOR2X0 U14401 ( .IN1(DFF_374_n1), .IN2(WX2146), .QN(n14003) );
  NOR3X0 U14402 ( .IN1(n9155), .IN2(n14005), .IN3(n14006), .QN(WX2601) );
  NOR2X0 U14403 ( .IN1(n8593), .IN2(CRC_OUT_8_21), .QN(n14006) );
  NOR2X0 U14404 ( .IN1(DFF_373_n1), .IN2(WX2148), .QN(n14005) );
  NOR3X0 U14405 ( .IN1(n9155), .IN2(n14007), .IN3(n14008), .QN(WX2599) );
  NOR2X0 U14406 ( .IN1(n8594), .IN2(CRC_OUT_8_20), .QN(n14008) );
  NOR2X0 U14407 ( .IN1(DFF_372_n1), .IN2(WX2150), .QN(n14007) );
  NOR3X0 U14408 ( .IN1(n9155), .IN2(n14009), .IN3(n14010), .QN(WX2597) );
  NOR2X0 U14409 ( .IN1(n8595), .IN2(CRC_OUT_8_19), .QN(n14010) );
  NOR2X0 U14410 ( .IN1(DFF_371_n1), .IN2(WX2152), .QN(n14009) );
  NOR3X0 U14411 ( .IN1(n9155), .IN2(n14011), .IN3(n14012), .QN(WX2595) );
  NOR2X0 U14412 ( .IN1(n8596), .IN2(CRC_OUT_8_18), .QN(n14012) );
  NOR2X0 U14413 ( .IN1(DFF_370_n1), .IN2(WX2154), .QN(n14011) );
  NOR3X0 U14414 ( .IN1(n9155), .IN2(n14013), .IN3(n14014), .QN(WX2593) );
  NOR2X0 U14415 ( .IN1(n8614), .IN2(CRC_OUT_8_17), .QN(n14014) );
  NOR2X0 U14416 ( .IN1(DFF_369_n1), .IN2(WX2156), .QN(n14013) );
  NOR3X0 U14417 ( .IN1(n9155), .IN2(n14015), .IN3(n14016), .QN(WX2591) );
  NOR2X0 U14418 ( .IN1(n8615), .IN2(CRC_OUT_8_16), .QN(n14016) );
  NOR2X0 U14419 ( .IN1(DFF_368_n1), .IN2(WX2158), .QN(n14015) );
  NOR2X0 U14420 ( .IN1(n9240), .IN2(n14017), .QN(WX2589) );
  NOR2X0 U14421 ( .IN1(n14018), .IN2(n14019), .QN(n14017) );
  INVX0 U14422 ( .INP(n14020), .ZN(n14019) );
  NAND2X0 U14423 ( .IN1(CRC_OUT_8_15), .IN2(n14021), .QN(n14020) );
  NOR2X0 U14424 ( .IN1(n14021), .IN2(CRC_OUT_8_15), .QN(n14018) );
  NAND2X0 U14425 ( .IN1(n14022), .IN2(n14023), .QN(n14021) );
  NAND2X0 U14426 ( .IN1(n8123), .IN2(CRC_OUT_8_31), .QN(n14023) );
  NAND2X0 U14427 ( .IN1(DFF_383_n1), .IN2(WX2160), .QN(n14022) );
  NOR3X0 U14428 ( .IN1(n9154), .IN2(n14024), .IN3(n14025), .QN(WX2587) );
  NOR2X0 U14429 ( .IN1(n8633), .IN2(CRC_OUT_8_14), .QN(n14025) );
  NOR2X0 U14430 ( .IN1(DFF_366_n1), .IN2(WX2162), .QN(n14024) );
  NOR3X0 U14431 ( .IN1(n9154), .IN2(n14026), .IN3(n14027), .QN(WX2585) );
  NOR2X0 U14432 ( .IN1(n8634), .IN2(CRC_OUT_8_13), .QN(n14027) );
  NOR2X0 U14433 ( .IN1(DFF_365_n1), .IN2(WX2164), .QN(n14026) );
  NOR3X0 U14434 ( .IN1(n9154), .IN2(n14028), .IN3(n14029), .QN(WX2583) );
  NOR2X0 U14435 ( .IN1(n8645), .IN2(CRC_OUT_8_12), .QN(n14029) );
  NOR2X0 U14436 ( .IN1(DFF_364_n1), .IN2(WX2166), .QN(n14028) );
  NOR3X0 U14437 ( .IN1(n9154), .IN2(n14030), .IN3(n14031), .QN(WX2581) );
  NOR2X0 U14438 ( .IN1(n8646), .IN2(CRC_OUT_8_11), .QN(n14031) );
  NOR2X0 U14439 ( .IN1(DFF_363_n1), .IN2(WX2168), .QN(n14030) );
  NOR2X0 U14440 ( .IN1(n9240), .IN2(n14032), .QN(WX2579) );
  NOR2X0 U14441 ( .IN1(n14033), .IN2(n14034), .QN(n14032) );
  INVX0 U14442 ( .INP(n14035), .ZN(n14034) );
  NAND2X0 U14443 ( .IN1(CRC_OUT_8_10), .IN2(n14036), .QN(n14035) );
  NOR2X0 U14444 ( .IN1(n14036), .IN2(CRC_OUT_8_10), .QN(n14033) );
  NAND2X0 U14445 ( .IN1(n14037), .IN2(n14038), .QN(n14036) );
  NAND2X0 U14446 ( .IN1(n8124), .IN2(CRC_OUT_8_31), .QN(n14038) );
  NAND2X0 U14447 ( .IN1(DFF_383_n1), .IN2(WX2170), .QN(n14037) );
  NOR2X0 U14448 ( .IN1(n9240), .IN2(n14039), .QN(WX2577) );
  NOR2X0 U14449 ( .IN1(n14040), .IN2(n14041), .QN(n14039) );
  NOR2X0 U14450 ( .IN1(test_so19), .IN2(CRC_OUT_8_9), .QN(n14041) );
  NOR2X0 U14451 ( .IN1(DFF_361_n1), .IN2(n8793), .QN(n14040) );
  NOR3X0 U14452 ( .IN1(n9155), .IN2(n14042), .IN3(n14043), .QN(WX2575) );
  NOR2X0 U14453 ( .IN1(n8647), .IN2(CRC_OUT_8_8), .QN(n14043) );
  NOR2X0 U14454 ( .IN1(DFF_360_n1), .IN2(WX2174), .QN(n14042) );
  NOR2X0 U14455 ( .IN1(n9240), .IN2(n14044), .QN(WX2573) );
  NOR2X0 U14456 ( .IN1(n14045), .IN2(n14046), .QN(n14044) );
  NOR2X0 U14457 ( .IN1(test_so20), .IN2(WX2176), .QN(n14046) );
  INVX0 U14458 ( .INP(n14047), .ZN(n14045) );
  NAND2X0 U14459 ( .IN1(WX2176), .IN2(test_so20), .QN(n14047) );
  NOR3X0 U14460 ( .IN1(n9154), .IN2(n14048), .IN3(n14049), .QN(WX2571) );
  NOR2X0 U14461 ( .IN1(n8649), .IN2(CRC_OUT_8_6), .QN(n14049) );
  NOR2X0 U14462 ( .IN1(DFF_358_n1), .IN2(WX2178), .QN(n14048) );
  NOR3X0 U14463 ( .IN1(n9153), .IN2(n14050), .IN3(n14051), .QN(WX2569) );
  NOR2X0 U14464 ( .IN1(n8650), .IN2(CRC_OUT_8_5), .QN(n14051) );
  NOR2X0 U14465 ( .IN1(DFF_357_n1), .IN2(WX2180), .QN(n14050) );
  NOR3X0 U14466 ( .IN1(n9155), .IN2(n14052), .IN3(n14053), .QN(WX2567) );
  NOR2X0 U14467 ( .IN1(n8651), .IN2(CRC_OUT_8_4), .QN(n14053) );
  NOR2X0 U14468 ( .IN1(DFF_356_n1), .IN2(WX2182), .QN(n14052) );
  NOR2X0 U14469 ( .IN1(n9241), .IN2(n14054), .QN(WX2565) );
  NOR2X0 U14470 ( .IN1(n14055), .IN2(n14056), .QN(n14054) );
  INVX0 U14471 ( .INP(n14057), .ZN(n14056) );
  NAND2X0 U14472 ( .IN1(CRC_OUT_8_3), .IN2(n14058), .QN(n14057) );
  NOR2X0 U14473 ( .IN1(n14058), .IN2(CRC_OUT_8_3), .QN(n14055) );
  NAND2X0 U14474 ( .IN1(n14059), .IN2(n14060), .QN(n14058) );
  NAND2X0 U14475 ( .IN1(n8125), .IN2(CRC_OUT_8_31), .QN(n14060) );
  NAND2X0 U14476 ( .IN1(DFF_383_n1), .IN2(WX2184), .QN(n14059) );
  NOR3X0 U14477 ( .IN1(n9154), .IN2(n14061), .IN3(n14062), .QN(WX2563) );
  NOR2X0 U14478 ( .IN1(n8652), .IN2(CRC_OUT_8_2), .QN(n14062) );
  NOR2X0 U14479 ( .IN1(DFF_354_n1), .IN2(WX2186), .QN(n14061) );
  NOR3X0 U14480 ( .IN1(n9154), .IN2(n14063), .IN3(n14064), .QN(WX2561) );
  NOR2X0 U14481 ( .IN1(n8659), .IN2(CRC_OUT_8_1), .QN(n14064) );
  NOR2X0 U14482 ( .IN1(DFF_353_n1), .IN2(WX2188), .QN(n14063) );
  NOR3X0 U14483 ( .IN1(n9153), .IN2(n14065), .IN3(n14066), .QN(WX2559) );
  NOR2X0 U14484 ( .IN1(n8660), .IN2(CRC_OUT_8_0), .QN(n14066) );
  NOR2X0 U14485 ( .IN1(DFF_352_n1), .IN2(WX2190), .QN(n14065) );
  NOR3X0 U14486 ( .IN1(n9154), .IN2(n14067), .IN3(n14068), .QN(WX2557) );
  NOR2X0 U14487 ( .IN1(n8133), .IN2(CRC_OUT_8_31), .QN(n14068) );
  NOR2X0 U14488 ( .IN1(DFF_383_n1), .IN2(WX2192), .QN(n14067) );
  NOR2X0 U14489 ( .IN1(n16321), .IN2(n9160), .QN(WX2031) );
  NOR2X0 U14490 ( .IN1(n16320), .IN2(n9160), .QN(WX2029) );
  NOR2X0 U14491 ( .IN1(n16319), .IN2(n9160), .QN(WX2027) );
  NOR2X0 U14492 ( .IN1(n16318), .IN2(n9160), .QN(WX2025) );
  NOR2X0 U14493 ( .IN1(n16317), .IN2(n9160), .QN(WX2023) );
  NOR2X0 U14494 ( .IN1(n16316), .IN2(n9160), .QN(WX2021) );
  NOR2X0 U14495 ( .IN1(n9241), .IN2(n8825), .QN(WX2019) );
  NOR2X0 U14496 ( .IN1(n16315), .IN2(n9160), .QN(WX2017) );
  NOR2X0 U14497 ( .IN1(n16314), .IN2(n9161), .QN(WX2015) );
  NOR2X0 U14498 ( .IN1(n16313), .IN2(n9161), .QN(WX2013) );
  NOR2X0 U14499 ( .IN1(n16312), .IN2(n9161), .QN(WX2011) );
  NOR2X0 U14500 ( .IN1(n16311), .IN2(n9162), .QN(WX2009) );
  NOR2X0 U14501 ( .IN1(n16310), .IN2(n9162), .QN(WX2007) );
  NOR2X0 U14502 ( .IN1(n16309), .IN2(n9162), .QN(WX2005) );
  NOR2X0 U14503 ( .IN1(n16308), .IN2(n9162), .QN(WX2003) );
  NOR2X0 U14504 ( .IN1(n16307), .IN2(n9162), .QN(WX2001) );
  NAND4X0 U14505 ( .IN1(n14069), .IN2(n14070), .IN3(n14071), .IN4(n14072), 
        .QN(WX1999) );
  NAND3X0 U14506 ( .IN1(n11657), .IN2(n11658), .IN3(n9090), .QN(n14072) );
  NAND3X0 U14507 ( .IN1(n14073), .IN2(n14074), .IN3(n14075), .QN(n11658) );
  INVX0 U14508 ( .INP(n14076), .ZN(n14075) );
  NAND2X0 U14509 ( .IN1(n14076), .IN2(n14077), .QN(n11657) );
  NAND2X0 U14510 ( .IN1(n14073), .IN2(n14074), .QN(n14077) );
  NAND2X0 U14511 ( .IN1(n8133), .IN2(WX2128), .QN(n14074) );
  NAND2X0 U14512 ( .IN1(n8067), .IN2(WX2192), .QN(n14073) );
  NOR2X0 U14513 ( .IN1(n14078), .IN2(n14079), .QN(n14076) );
  INVX0 U14514 ( .INP(n14080), .ZN(n14079) );
  NAND2X0 U14515 ( .IN1(test_so16), .IN2(WX2000), .QN(n14080) );
  NOR2X0 U14516 ( .IN1(WX2000), .IN2(test_so16), .QN(n14078) );
  NAND2X0 U14517 ( .IN1(n9327), .IN2(n13396), .QN(n14071) );
  NAND2X0 U14518 ( .IN1(n14081), .IN2(n14082), .QN(n13396) );
  INVX0 U14519 ( .INP(n14083), .ZN(n14082) );
  NOR2X0 U14520 ( .IN1(n14084), .IN2(n14085), .QN(n14083) );
  NAND2X0 U14521 ( .IN1(n14085), .IN2(n14084), .QN(n14081) );
  NOR2X0 U14522 ( .IN1(n14086), .IN2(n14087), .QN(n14084) );
  NOR2X0 U14523 ( .IN1(WX3485), .IN2(n8036), .QN(n14087) );
  INVX0 U14524 ( .INP(n14088), .ZN(n14086) );
  NAND2X0 U14525 ( .IN1(n8036), .IN2(WX3485), .QN(n14088) );
  NAND2X0 U14526 ( .IN1(n14089), .IN2(n14090), .QN(n14085) );
  NAND2X0 U14527 ( .IN1(n8035), .IN2(WX3357), .QN(n14090) );
  INVX0 U14528 ( .INP(n14091), .ZN(n14089) );
  NOR2X0 U14529 ( .IN1(WX3357), .IN2(n8035), .QN(n14091) );
  NAND2X0 U14530 ( .IN1(n280), .IN2(n9285), .QN(n14070) );
  NOR2X0 U14531 ( .IN1(n9241), .IN2(n9003), .QN(n280) );
  NAND2X0 U14532 ( .IN1(n9298), .IN2(CRC_OUT_8_0), .QN(n14069) );
  NAND4X0 U14533 ( .IN1(n14092), .IN2(n14093), .IN3(n14094), .IN4(n14095), 
        .QN(WX1997) );
  NAND2X0 U14534 ( .IN1(n9327), .IN2(n13412), .QN(n14095) );
  NAND2X0 U14535 ( .IN1(n14096), .IN2(n14097), .QN(n13412) );
  INVX0 U14536 ( .INP(n14098), .ZN(n14097) );
  NOR2X0 U14537 ( .IN1(n14099), .IN2(n14100), .QN(n14098) );
  NAND2X0 U14538 ( .IN1(n14100), .IN2(n14099), .QN(n14096) );
  NOR2X0 U14539 ( .IN1(n14101), .IN2(n14102), .QN(n14099) );
  NOR2X0 U14540 ( .IN1(WX3483), .IN2(n8038), .QN(n14102) );
  INVX0 U14541 ( .INP(n14103), .ZN(n14101) );
  NAND2X0 U14542 ( .IN1(n8038), .IN2(WX3483), .QN(n14103) );
  NAND2X0 U14543 ( .IN1(n14104), .IN2(n14105), .QN(n14100) );
  NAND2X0 U14544 ( .IN1(n8037), .IN2(WX3355), .QN(n14105) );
  INVX0 U14545 ( .INP(n14106), .ZN(n14104) );
  NOR2X0 U14546 ( .IN1(WX3355), .IN2(n8037), .QN(n14106) );
  NAND2X0 U14547 ( .IN1(n9105), .IN2(n11664), .QN(n14094) );
  NAND2X0 U14548 ( .IN1(n14107), .IN2(n14108), .QN(n11664) );
  INVX0 U14549 ( .INP(n14109), .ZN(n14108) );
  NOR2X0 U14550 ( .IN1(n14110), .IN2(n14111), .QN(n14109) );
  NAND2X0 U14551 ( .IN1(n14111), .IN2(n14110), .QN(n14107) );
  NOR2X0 U14552 ( .IN1(n14112), .IN2(n14113), .QN(n14110) );
  NOR2X0 U14553 ( .IN1(WX2190), .IN2(n8069), .QN(n14113) );
  INVX0 U14554 ( .INP(n14114), .ZN(n14112) );
  NAND2X0 U14555 ( .IN1(n8069), .IN2(WX2190), .QN(n14114) );
  NAND2X0 U14556 ( .IN1(n14115), .IN2(n14116), .QN(n14111) );
  NAND2X0 U14557 ( .IN1(n8068), .IN2(WX2062), .QN(n14116) );
  INVX0 U14558 ( .INP(n14117), .ZN(n14115) );
  NOR2X0 U14559 ( .IN1(WX2062), .IN2(n8068), .QN(n14117) );
  NAND2X0 U14560 ( .IN1(n279), .IN2(n9285), .QN(n14093) );
  NOR2X0 U14561 ( .IN1(n9241), .IN2(n9004), .QN(n279) );
  NAND2X0 U14562 ( .IN1(n9298), .IN2(CRC_OUT_8_1), .QN(n14092) );
  NAND4X0 U14563 ( .IN1(n14118), .IN2(n14119), .IN3(n14120), .IN4(n14121), 
        .QN(WX1995) );
  NAND2X0 U14564 ( .IN1(n9327), .IN2(n13428), .QN(n14121) );
  NAND2X0 U14565 ( .IN1(n14122), .IN2(n14123), .QN(n13428) );
  INVX0 U14566 ( .INP(n14124), .ZN(n14123) );
  NOR2X0 U14567 ( .IN1(n14125), .IN2(n14126), .QN(n14124) );
  NAND2X0 U14568 ( .IN1(n14126), .IN2(n14125), .QN(n14122) );
  NOR2X0 U14569 ( .IN1(n14127), .IN2(n14128), .QN(n14125) );
  NOR2X0 U14570 ( .IN1(WX3481), .IN2(n8040), .QN(n14128) );
  INVX0 U14571 ( .INP(n14129), .ZN(n14127) );
  NAND2X0 U14572 ( .IN1(n8040), .IN2(WX3481), .QN(n14129) );
  NAND2X0 U14573 ( .IN1(n14130), .IN2(n14131), .QN(n14126) );
  NAND2X0 U14574 ( .IN1(n8039), .IN2(WX3353), .QN(n14131) );
  INVX0 U14575 ( .INP(n14132), .ZN(n14130) );
  NOR2X0 U14576 ( .IN1(WX3353), .IN2(n8039), .QN(n14132) );
  NAND2X0 U14577 ( .IN1(n9105), .IN2(n11670), .QN(n14120) );
  NAND2X0 U14578 ( .IN1(n14133), .IN2(n14134), .QN(n11670) );
  INVX0 U14579 ( .INP(n14135), .ZN(n14134) );
  NOR2X0 U14580 ( .IN1(n14136), .IN2(n14137), .QN(n14135) );
  NAND2X0 U14581 ( .IN1(n14137), .IN2(n14136), .QN(n14133) );
  NOR2X0 U14582 ( .IN1(n14138), .IN2(n14139), .QN(n14136) );
  NOR2X0 U14583 ( .IN1(WX2188), .IN2(n8071), .QN(n14139) );
  INVX0 U14584 ( .INP(n14140), .ZN(n14138) );
  NAND2X0 U14585 ( .IN1(n8071), .IN2(WX2188), .QN(n14140) );
  NAND2X0 U14586 ( .IN1(n14141), .IN2(n14142), .QN(n14137) );
  NAND2X0 U14587 ( .IN1(n8070), .IN2(WX2060), .QN(n14142) );
  INVX0 U14588 ( .INP(n14143), .ZN(n14141) );
  NOR2X0 U14589 ( .IN1(WX2060), .IN2(n8070), .QN(n14143) );
  NAND2X0 U14590 ( .IN1(n278), .IN2(n9285), .QN(n14119) );
  NOR2X0 U14591 ( .IN1(n9241), .IN2(n9005), .QN(n278) );
  NAND2X0 U14592 ( .IN1(n9298), .IN2(CRC_OUT_8_2), .QN(n14118) );
  NAND4X0 U14593 ( .IN1(n14144), .IN2(n14145), .IN3(n14146), .IN4(n14147), 
        .QN(WX1993) );
  NAND2X0 U14594 ( .IN1(n9327), .IN2(n13444), .QN(n14147) );
  NAND2X0 U14595 ( .IN1(n14148), .IN2(n14149), .QN(n13444) );
  INVX0 U14596 ( .INP(n14150), .ZN(n14149) );
  NOR2X0 U14597 ( .IN1(n14151), .IN2(n14152), .QN(n14150) );
  NAND2X0 U14598 ( .IN1(n14152), .IN2(n14151), .QN(n14148) );
  NOR2X0 U14599 ( .IN1(n14153), .IN2(n14154), .QN(n14151) );
  NOR2X0 U14600 ( .IN1(WX3479), .IN2(n8042), .QN(n14154) );
  INVX0 U14601 ( .INP(n14155), .ZN(n14153) );
  NAND2X0 U14602 ( .IN1(n8042), .IN2(WX3479), .QN(n14155) );
  NAND2X0 U14603 ( .IN1(n14156), .IN2(n14157), .QN(n14152) );
  NAND2X0 U14604 ( .IN1(n8041), .IN2(WX3351), .QN(n14157) );
  INVX0 U14605 ( .INP(n14158), .ZN(n14156) );
  NOR2X0 U14606 ( .IN1(WX3351), .IN2(n8041), .QN(n14158) );
  NAND2X0 U14607 ( .IN1(n9105), .IN2(n11677), .QN(n14146) );
  NAND2X0 U14608 ( .IN1(n14159), .IN2(n14160), .QN(n11677) );
  INVX0 U14609 ( .INP(n14161), .ZN(n14160) );
  NOR2X0 U14610 ( .IN1(n14162), .IN2(n14163), .QN(n14161) );
  NAND2X0 U14611 ( .IN1(n14163), .IN2(n14162), .QN(n14159) );
  NOR2X0 U14612 ( .IN1(n14164), .IN2(n14165), .QN(n14162) );
  NOR2X0 U14613 ( .IN1(WX2186), .IN2(n8073), .QN(n14165) );
  INVX0 U14614 ( .INP(n14166), .ZN(n14164) );
  NAND2X0 U14615 ( .IN1(n8073), .IN2(WX2186), .QN(n14166) );
  NAND2X0 U14616 ( .IN1(n14167), .IN2(n14168), .QN(n14163) );
  NAND2X0 U14617 ( .IN1(n8072), .IN2(WX2058), .QN(n14168) );
  INVX0 U14618 ( .INP(n14169), .ZN(n14167) );
  NOR2X0 U14619 ( .IN1(WX2058), .IN2(n8072), .QN(n14169) );
  NAND2X0 U14620 ( .IN1(n277), .IN2(n9286), .QN(n14145) );
  NOR2X0 U14621 ( .IN1(n9241), .IN2(n9006), .QN(n277) );
  NAND2X0 U14622 ( .IN1(n9298), .IN2(CRC_OUT_8_3), .QN(n14144) );
  NAND4X0 U14623 ( .IN1(n14170), .IN2(n14171), .IN3(n14172), .IN4(n14173), 
        .QN(WX1991) );
  NAND3X0 U14624 ( .IN1(n11683), .IN2(n11684), .IN3(n9091), .QN(n14173) );
  NAND3X0 U14625 ( .IN1(n14174), .IN2(n14175), .IN3(n14176), .QN(n11684) );
  INVX0 U14626 ( .INP(n14177), .ZN(n14176) );
  NAND2X0 U14627 ( .IN1(n14177), .IN2(n14178), .QN(n11683) );
  NAND2X0 U14628 ( .IN1(n14174), .IN2(n14175), .QN(n14178) );
  NAND2X0 U14629 ( .IN1(n8125), .IN2(WX2056), .QN(n14175) );
  NAND2X0 U14630 ( .IN1(n3763), .IN2(WX2184), .QN(n14174) );
  NOR2X0 U14631 ( .IN1(n14179), .IN2(n14180), .QN(n14177) );
  INVX0 U14632 ( .INP(n14181), .ZN(n14180) );
  NAND2X0 U14633 ( .IN1(test_so14), .IN2(WX2120), .QN(n14181) );
  NOR2X0 U14634 ( .IN1(WX2120), .IN2(test_so14), .QN(n14179) );
  NAND2X0 U14635 ( .IN1(n9327), .IN2(n13460), .QN(n14172) );
  NAND2X0 U14636 ( .IN1(n14182), .IN2(n14183), .QN(n13460) );
  INVX0 U14637 ( .INP(n14184), .ZN(n14183) );
  NOR2X0 U14638 ( .IN1(n14185), .IN2(n14186), .QN(n14184) );
  NAND2X0 U14639 ( .IN1(n14186), .IN2(n14185), .QN(n14182) );
  NOR2X0 U14640 ( .IN1(n14187), .IN2(n14188), .QN(n14185) );
  NOR2X0 U14641 ( .IN1(WX3477), .IN2(n8044), .QN(n14188) );
  INVX0 U14642 ( .INP(n14189), .ZN(n14187) );
  NAND2X0 U14643 ( .IN1(n8044), .IN2(WX3477), .QN(n14189) );
  NAND2X0 U14644 ( .IN1(n14190), .IN2(n14191), .QN(n14186) );
  NAND2X0 U14645 ( .IN1(n8043), .IN2(WX3349), .QN(n14191) );
  INVX0 U14646 ( .INP(n14192), .ZN(n14190) );
  NOR2X0 U14647 ( .IN1(WX3349), .IN2(n8043), .QN(n14192) );
  NAND2X0 U14648 ( .IN1(n276), .IN2(n9286), .QN(n14171) );
  NOR2X0 U14649 ( .IN1(n9241), .IN2(n9007), .QN(n276) );
  NAND2X0 U14650 ( .IN1(n9298), .IN2(CRC_OUT_8_4), .QN(n14170) );
  NAND4X0 U14651 ( .IN1(n14193), .IN2(n14194), .IN3(n14195), .IN4(n14196), 
        .QN(WX1989) );
  NAND2X0 U14652 ( .IN1(n9327), .IN2(n13476), .QN(n14196) );
  NAND2X0 U14653 ( .IN1(n14197), .IN2(n14198), .QN(n13476) );
  INVX0 U14654 ( .INP(n14199), .ZN(n14198) );
  NOR2X0 U14655 ( .IN1(n14200), .IN2(n14201), .QN(n14199) );
  NAND2X0 U14656 ( .IN1(n14201), .IN2(n14200), .QN(n14197) );
  NOR2X0 U14657 ( .IN1(n14202), .IN2(n14203), .QN(n14200) );
  NOR2X0 U14658 ( .IN1(WX3475), .IN2(n8046), .QN(n14203) );
  INVX0 U14659 ( .INP(n14204), .ZN(n14202) );
  NAND2X0 U14660 ( .IN1(n8046), .IN2(WX3475), .QN(n14204) );
  NAND2X0 U14661 ( .IN1(n14205), .IN2(n14206), .QN(n14201) );
  NAND2X0 U14662 ( .IN1(n8045), .IN2(WX3347), .QN(n14206) );
  INVX0 U14663 ( .INP(n14207), .ZN(n14205) );
  NOR2X0 U14664 ( .IN1(WX3347), .IN2(n8045), .QN(n14207) );
  NAND2X0 U14665 ( .IN1(n9105), .IN2(n11690), .QN(n14195) );
  NAND2X0 U14666 ( .IN1(n14208), .IN2(n14209), .QN(n11690) );
  INVX0 U14667 ( .INP(n14210), .ZN(n14209) );
  NOR2X0 U14668 ( .IN1(n14211), .IN2(n14212), .QN(n14210) );
  NAND2X0 U14669 ( .IN1(n14212), .IN2(n14211), .QN(n14208) );
  NOR2X0 U14670 ( .IN1(n14213), .IN2(n14214), .QN(n14211) );
  NOR2X0 U14671 ( .IN1(WX2182), .IN2(n8076), .QN(n14214) );
  INVX0 U14672 ( .INP(n14215), .ZN(n14213) );
  NAND2X0 U14673 ( .IN1(n8076), .IN2(WX2182), .QN(n14215) );
  NAND2X0 U14674 ( .IN1(n14216), .IN2(n14217), .QN(n14212) );
  NAND2X0 U14675 ( .IN1(n8075), .IN2(WX2054), .QN(n14217) );
  INVX0 U14676 ( .INP(n14218), .ZN(n14216) );
  NOR2X0 U14677 ( .IN1(WX2054), .IN2(n8075), .QN(n14218) );
  NAND2X0 U14678 ( .IN1(n275), .IN2(n9286), .QN(n14194) );
  NOR2X0 U14679 ( .IN1(n9241), .IN2(n9008), .QN(n275) );
  NAND2X0 U14680 ( .IN1(n9299), .IN2(CRC_OUT_8_5), .QN(n14193) );
  NAND4X0 U14681 ( .IN1(n14219), .IN2(n14220), .IN3(n14221), .IN4(n14222), 
        .QN(WX1987) );
  NAND3X0 U14682 ( .IN1(n13481), .IN2(n13482), .IN3(n9322), .QN(n14222) );
  NAND3X0 U14683 ( .IN1(n14223), .IN2(n14224), .IN3(n14225), .QN(n13482) );
  INVX0 U14684 ( .INP(n14226), .ZN(n14225) );
  NAND2X0 U14685 ( .IN1(n14226), .IN2(n14227), .QN(n13481) );
  NAND2X0 U14686 ( .IN1(n14223), .IN2(n14224), .QN(n14227) );
  NAND2X0 U14687 ( .IN1(n8048), .IN2(WX3345), .QN(n14224) );
  NAND2X0 U14688 ( .IN1(n3735), .IN2(WX3409), .QN(n14223) );
  NOR2X0 U14689 ( .IN1(n14228), .IN2(n14229), .QN(n14226) );
  NOR2X0 U14690 ( .IN1(n8792), .IN2(n8047), .QN(n14229) );
  INVX0 U14691 ( .INP(n14230), .ZN(n14228) );
  NAND2X0 U14692 ( .IN1(n8047), .IN2(n8792), .QN(n14230) );
  NAND2X0 U14693 ( .IN1(n9105), .IN2(n11696), .QN(n14221) );
  NAND2X0 U14694 ( .IN1(n14231), .IN2(n14232), .QN(n11696) );
  INVX0 U14695 ( .INP(n14233), .ZN(n14232) );
  NOR2X0 U14696 ( .IN1(n14234), .IN2(n14235), .QN(n14233) );
  NAND2X0 U14697 ( .IN1(n14235), .IN2(n14234), .QN(n14231) );
  NOR2X0 U14698 ( .IN1(n14236), .IN2(n14237), .QN(n14234) );
  NOR2X0 U14699 ( .IN1(WX2180), .IN2(n8078), .QN(n14237) );
  INVX0 U14700 ( .INP(n14238), .ZN(n14236) );
  NAND2X0 U14701 ( .IN1(n8078), .IN2(WX2180), .QN(n14238) );
  NAND2X0 U14702 ( .IN1(n14239), .IN2(n14240), .QN(n14235) );
  NAND2X0 U14703 ( .IN1(n8077), .IN2(WX2052), .QN(n14240) );
  INVX0 U14704 ( .INP(n14241), .ZN(n14239) );
  NOR2X0 U14705 ( .IN1(WX2052), .IN2(n8077), .QN(n14241) );
  NAND2X0 U14706 ( .IN1(n274), .IN2(n9286), .QN(n14220) );
  NOR2X0 U14707 ( .IN1(n9242), .IN2(n9009), .QN(n274) );
  NAND2X0 U14708 ( .IN1(n9299), .IN2(CRC_OUT_8_6), .QN(n14219) );
  NAND4X0 U14709 ( .IN1(n14242), .IN2(n14243), .IN3(n14244), .IN4(n14245), 
        .QN(WX1985) );
  NAND2X0 U14710 ( .IN1(n9327), .IN2(n13509), .QN(n14245) );
  NAND2X0 U14711 ( .IN1(n14246), .IN2(n14247), .QN(n13509) );
  INVX0 U14712 ( .INP(n14248), .ZN(n14247) );
  NOR2X0 U14713 ( .IN1(n14249), .IN2(n14250), .QN(n14248) );
  NAND2X0 U14714 ( .IN1(n14250), .IN2(n14249), .QN(n14246) );
  NOR2X0 U14715 ( .IN1(n14251), .IN2(n14252), .QN(n14249) );
  NOR2X0 U14716 ( .IN1(WX3471), .IN2(n8050), .QN(n14252) );
  INVX0 U14717 ( .INP(n14253), .ZN(n14251) );
  NAND2X0 U14718 ( .IN1(n8050), .IN2(WX3471), .QN(n14253) );
  NAND2X0 U14719 ( .IN1(n14254), .IN2(n14255), .QN(n14250) );
  NAND2X0 U14720 ( .IN1(n8049), .IN2(WX3343), .QN(n14255) );
  INVX0 U14721 ( .INP(n14256), .ZN(n14254) );
  NOR2X0 U14722 ( .IN1(WX3343), .IN2(n8049), .QN(n14256) );
  NAND2X0 U14723 ( .IN1(n9105), .IN2(n11703), .QN(n14244) );
  NAND2X0 U14724 ( .IN1(n14257), .IN2(n14258), .QN(n11703) );
  INVX0 U14725 ( .INP(n14259), .ZN(n14258) );
  NOR2X0 U14726 ( .IN1(n14260), .IN2(n14261), .QN(n14259) );
  NAND2X0 U14727 ( .IN1(n14261), .IN2(n14260), .QN(n14257) );
  NOR2X0 U14728 ( .IN1(n14262), .IN2(n14263), .QN(n14260) );
  NOR2X0 U14729 ( .IN1(WX2178), .IN2(n8080), .QN(n14263) );
  INVX0 U14730 ( .INP(n14264), .ZN(n14262) );
  NAND2X0 U14731 ( .IN1(n8080), .IN2(WX2178), .QN(n14264) );
  NAND2X0 U14732 ( .IN1(n14265), .IN2(n14266), .QN(n14261) );
  NAND2X0 U14733 ( .IN1(n8079), .IN2(WX2050), .QN(n14266) );
  INVX0 U14734 ( .INP(n14267), .ZN(n14265) );
  NOR2X0 U14735 ( .IN1(WX2050), .IN2(n8079), .QN(n14267) );
  NAND2X0 U14736 ( .IN1(n273), .IN2(n9286), .QN(n14243) );
  NOR2X0 U14737 ( .IN1(n9242), .IN2(n9010), .QN(n273) );
  NAND2X0 U14738 ( .IN1(test_so20), .IN2(n9315), .QN(n14242) );
  NAND4X0 U14739 ( .IN1(n14268), .IN2(n14269), .IN3(n14270), .IN4(n14271), 
        .QN(WX1983) );
  NAND3X0 U14740 ( .IN1(n13514), .IN2(n13515), .IN3(n9322), .QN(n14271) );
  NAND3X0 U14741 ( .IN1(n14272), .IN2(n14273), .IN3(n14274), .QN(n13515) );
  INVX0 U14742 ( .INP(n14275), .ZN(n14274) );
  NAND2X0 U14743 ( .IN1(n14275), .IN2(n14276), .QN(n13514) );
  NAND2X0 U14744 ( .IN1(n14272), .IN2(n14273), .QN(n14276) );
  NAND2X0 U14745 ( .IN1(n8535), .IN2(WX3341), .QN(n14273) );
  NAND2X0 U14746 ( .IN1(n3739), .IN2(WX3469), .QN(n14272) );
  NOR2X0 U14747 ( .IN1(n14277), .IN2(n14278), .QN(n14275) );
  INVX0 U14748 ( .INP(n14279), .ZN(n14278) );
  NAND2X0 U14749 ( .IN1(test_so28), .IN2(WX3277), .QN(n14279) );
  NOR2X0 U14750 ( .IN1(WX3277), .IN2(test_so28), .QN(n14277) );
  NAND2X0 U14751 ( .IN1(n9105), .IN2(n11709), .QN(n14270) );
  NAND2X0 U14752 ( .IN1(n14280), .IN2(n14281), .QN(n11709) );
  INVX0 U14753 ( .INP(n14282), .ZN(n14281) );
  NOR2X0 U14754 ( .IN1(n14283), .IN2(n14284), .QN(n14282) );
  NAND2X0 U14755 ( .IN1(n14284), .IN2(n14283), .QN(n14280) );
  NOR2X0 U14756 ( .IN1(n14285), .IN2(n14286), .QN(n14283) );
  NOR2X0 U14757 ( .IN1(WX2176), .IN2(n8082), .QN(n14286) );
  INVX0 U14758 ( .INP(n14287), .ZN(n14285) );
  NAND2X0 U14759 ( .IN1(n8082), .IN2(WX2176), .QN(n14287) );
  NAND2X0 U14760 ( .IN1(n14288), .IN2(n14289), .QN(n14284) );
  NAND2X0 U14761 ( .IN1(n8081), .IN2(WX2048), .QN(n14289) );
  INVX0 U14762 ( .INP(n14290), .ZN(n14288) );
  NOR2X0 U14763 ( .IN1(WX2048), .IN2(n8081), .QN(n14290) );
  NAND2X0 U14764 ( .IN1(n272), .IN2(n9286), .QN(n14269) );
  NOR2X0 U14765 ( .IN1(n9073), .IN2(n9162), .QN(n272) );
  NAND2X0 U14766 ( .IN1(n9299), .IN2(CRC_OUT_8_8), .QN(n14268) );
  NAND4X0 U14767 ( .IN1(n14291), .IN2(n14292), .IN3(n14293), .IN4(n14294), 
        .QN(WX1981) );
  NAND2X0 U14768 ( .IN1(n9327), .IN2(n13542), .QN(n14294) );
  NAND2X0 U14769 ( .IN1(n14295), .IN2(n14296), .QN(n13542) );
  INVX0 U14770 ( .INP(n14297), .ZN(n14296) );
  NOR2X0 U14771 ( .IN1(n14298), .IN2(n14299), .QN(n14297) );
  NAND2X0 U14772 ( .IN1(n14299), .IN2(n14298), .QN(n14295) );
  NOR2X0 U14773 ( .IN1(n14300), .IN2(n14301), .QN(n14298) );
  NOR2X0 U14774 ( .IN1(WX3467), .IN2(n8053), .QN(n14301) );
  INVX0 U14775 ( .INP(n14302), .ZN(n14300) );
  NAND2X0 U14776 ( .IN1(n8053), .IN2(WX3467), .QN(n14302) );
  NAND2X0 U14777 ( .IN1(n14303), .IN2(n14304), .QN(n14299) );
  NAND2X0 U14778 ( .IN1(n8052), .IN2(WX3339), .QN(n14304) );
  INVX0 U14779 ( .INP(n14305), .ZN(n14303) );
  NOR2X0 U14780 ( .IN1(WX3339), .IN2(n8052), .QN(n14305) );
  NAND2X0 U14781 ( .IN1(n9105), .IN2(n11715), .QN(n14293) );
  NAND2X0 U14782 ( .IN1(n14306), .IN2(n14307), .QN(n11715) );
  INVX0 U14783 ( .INP(n14308), .ZN(n14307) );
  NOR2X0 U14784 ( .IN1(n14309), .IN2(n14310), .QN(n14308) );
  NAND2X0 U14785 ( .IN1(n14310), .IN2(n14309), .QN(n14306) );
  NOR2X0 U14786 ( .IN1(n14311), .IN2(n14312), .QN(n14309) );
  NOR2X0 U14787 ( .IN1(WX2174), .IN2(n8084), .QN(n14312) );
  INVX0 U14788 ( .INP(n14313), .ZN(n14311) );
  NAND2X0 U14789 ( .IN1(n8084), .IN2(WX2174), .QN(n14313) );
  NAND2X0 U14790 ( .IN1(n14314), .IN2(n14315), .QN(n14310) );
  NAND2X0 U14791 ( .IN1(n8083), .IN2(WX2046), .QN(n14315) );
  INVX0 U14792 ( .INP(n14316), .ZN(n14314) );
  NOR2X0 U14793 ( .IN1(WX2046), .IN2(n8083), .QN(n14316) );
  NAND2X0 U14794 ( .IN1(n271), .IN2(n9286), .QN(n14292) );
  NOR2X0 U14795 ( .IN1(n9242), .IN2(n9011), .QN(n271) );
  NAND2X0 U14796 ( .IN1(n9299), .IN2(CRC_OUT_8_9), .QN(n14291) );
  NAND4X0 U14797 ( .IN1(n14317), .IN2(n14318), .IN3(n14319), .IN4(n14320), 
        .QN(WX1979) );
  NAND3X0 U14798 ( .IN1(n11721), .IN2(n11722), .IN3(n9091), .QN(n14320) );
  NAND3X0 U14799 ( .IN1(n14321), .IN2(n14322), .IN3(n14323), .QN(n11722) );
  INVX0 U14800 ( .INP(n14324), .ZN(n14323) );
  NAND2X0 U14801 ( .IN1(n14324), .IN2(n14325), .QN(n11721) );
  NAND2X0 U14802 ( .IN1(n14321), .IN2(n14322), .QN(n14325) );
  NAND2X0 U14803 ( .IN1(n8086), .IN2(WX2044), .QN(n14322) );
  NAND2X0 U14804 ( .IN1(n3775), .IN2(WX2108), .QN(n14321) );
  NOR2X0 U14805 ( .IN1(n14326), .IN2(n14327), .QN(n14324) );
  NOR2X0 U14806 ( .IN1(n8793), .IN2(n8085), .QN(n14327) );
  INVX0 U14807 ( .INP(n14328), .ZN(n14326) );
  NAND2X0 U14808 ( .IN1(n8085), .IN2(n8793), .QN(n14328) );
  NAND2X0 U14809 ( .IN1(n9328), .IN2(n13558), .QN(n14319) );
  NAND2X0 U14810 ( .IN1(n14329), .IN2(n14330), .QN(n13558) );
  INVX0 U14811 ( .INP(n14331), .ZN(n14330) );
  NOR2X0 U14812 ( .IN1(n14332), .IN2(n14333), .QN(n14331) );
  NAND2X0 U14813 ( .IN1(n14333), .IN2(n14332), .QN(n14329) );
  NOR2X0 U14814 ( .IN1(n14334), .IN2(n14335), .QN(n14332) );
  NOR2X0 U14815 ( .IN1(WX3465), .IN2(n8055), .QN(n14335) );
  INVX0 U14816 ( .INP(n14336), .ZN(n14334) );
  NAND2X0 U14817 ( .IN1(n8055), .IN2(WX3465), .QN(n14336) );
  NAND2X0 U14818 ( .IN1(n14337), .IN2(n14338), .QN(n14333) );
  NAND2X0 U14819 ( .IN1(n8054), .IN2(WX3337), .QN(n14338) );
  INVX0 U14820 ( .INP(n14339), .ZN(n14337) );
  NOR2X0 U14821 ( .IN1(WX3337), .IN2(n8054), .QN(n14339) );
  NAND2X0 U14822 ( .IN1(n270), .IN2(n9286), .QN(n14318) );
  NOR2X0 U14823 ( .IN1(n9242), .IN2(n9012), .QN(n270) );
  NAND2X0 U14824 ( .IN1(n9299), .IN2(CRC_OUT_8_10), .QN(n14317) );
  NAND4X0 U14825 ( .IN1(n14340), .IN2(n14341), .IN3(n14342), .IN4(n14343), 
        .QN(WX1977) );
  NAND2X0 U14826 ( .IN1(n9328), .IN2(n13571), .QN(n14343) );
  NAND2X0 U14827 ( .IN1(n14344), .IN2(n14345), .QN(n13571) );
  INVX0 U14828 ( .INP(n14346), .ZN(n14345) );
  NOR2X0 U14829 ( .IN1(n14347), .IN2(n14348), .QN(n14346) );
  NAND2X0 U14830 ( .IN1(n14348), .IN2(n14347), .QN(n14344) );
  NOR2X0 U14831 ( .IN1(n14349), .IN2(n14350), .QN(n14347) );
  NOR2X0 U14832 ( .IN1(WX3463), .IN2(n8057), .QN(n14350) );
  INVX0 U14833 ( .INP(n14351), .ZN(n14349) );
  NAND2X0 U14834 ( .IN1(n8057), .IN2(WX3463), .QN(n14351) );
  NAND2X0 U14835 ( .IN1(n14352), .IN2(n14353), .QN(n14348) );
  NAND2X0 U14836 ( .IN1(n8056), .IN2(WX3335), .QN(n14353) );
  INVX0 U14837 ( .INP(n14354), .ZN(n14352) );
  NOR2X0 U14838 ( .IN1(WX3335), .IN2(n8056), .QN(n14354) );
  NAND2X0 U14839 ( .IN1(n9105), .IN2(n11729), .QN(n14342) );
  NAND2X0 U14840 ( .IN1(n14355), .IN2(n14356), .QN(n11729) );
  INVX0 U14841 ( .INP(n14357), .ZN(n14356) );
  NOR2X0 U14842 ( .IN1(n14358), .IN2(n14359), .QN(n14357) );
  NAND2X0 U14843 ( .IN1(n14359), .IN2(n14358), .QN(n14355) );
  NOR2X0 U14844 ( .IN1(n14360), .IN2(n14361), .QN(n14358) );
  NOR2X0 U14845 ( .IN1(WX2170), .IN2(n8088), .QN(n14361) );
  INVX0 U14846 ( .INP(n14362), .ZN(n14360) );
  NAND2X0 U14847 ( .IN1(n8088), .IN2(WX2170), .QN(n14362) );
  NAND2X0 U14848 ( .IN1(n14363), .IN2(n14364), .QN(n14359) );
  NAND2X0 U14849 ( .IN1(n8087), .IN2(WX2042), .QN(n14364) );
  INVX0 U14850 ( .INP(n14365), .ZN(n14363) );
  NOR2X0 U14851 ( .IN1(WX2042), .IN2(n8087), .QN(n14365) );
  NAND2X0 U14852 ( .IN1(n269), .IN2(n9286), .QN(n14341) );
  NOR2X0 U14853 ( .IN1(n9242), .IN2(n9013), .QN(n269) );
  NAND2X0 U14854 ( .IN1(n9299), .IN2(CRC_OUT_8_11), .QN(n14340) );
  NAND4X0 U14855 ( .IN1(n14366), .IN2(n14367), .IN3(n14368), .IN4(n14369), 
        .QN(WX1975) );
  NAND3X0 U14856 ( .IN1(n13576), .IN2(n13577), .IN3(n9321), .QN(n14369) );
  NAND3X0 U14857 ( .IN1(n14370), .IN2(n14371), .IN3(n14372), .QN(n13577) );
  INVX0 U14858 ( .INP(n14373), .ZN(n14372) );
  NAND2X0 U14859 ( .IN1(n14373), .IN2(n14374), .QN(n13576) );
  NAND2X0 U14860 ( .IN1(n14370), .IN2(n14371), .QN(n14374) );
  NAND2X0 U14861 ( .IN1(n8532), .IN2(WX3397), .QN(n14371) );
  NAND2X0 U14862 ( .IN1(n8059), .IN2(WX3461), .QN(n14370) );
  NOR2X0 U14863 ( .IN1(n14375), .IN2(n14376), .QN(n14373) );
  INVX0 U14864 ( .INP(n14377), .ZN(n14376) );
  NAND2X0 U14865 ( .IN1(test_so26), .IN2(WX3269), .QN(n14377) );
  NOR2X0 U14866 ( .IN1(WX3269), .IN2(test_so26), .QN(n14375) );
  NAND2X0 U14867 ( .IN1(n9105), .IN2(n11735), .QN(n14368) );
  NAND2X0 U14868 ( .IN1(n14378), .IN2(n14379), .QN(n11735) );
  INVX0 U14869 ( .INP(n14380), .ZN(n14379) );
  NOR2X0 U14870 ( .IN1(n14381), .IN2(n14382), .QN(n14380) );
  NAND2X0 U14871 ( .IN1(n14382), .IN2(n14381), .QN(n14378) );
  NOR2X0 U14872 ( .IN1(n14383), .IN2(n14384), .QN(n14381) );
  NOR2X0 U14873 ( .IN1(WX2168), .IN2(n8090), .QN(n14384) );
  INVX0 U14874 ( .INP(n14385), .ZN(n14383) );
  NAND2X0 U14875 ( .IN1(n8090), .IN2(WX2168), .QN(n14385) );
  NAND2X0 U14876 ( .IN1(n14386), .IN2(n14387), .QN(n14382) );
  NAND2X0 U14877 ( .IN1(n8089), .IN2(WX2040), .QN(n14387) );
  INVX0 U14878 ( .INP(n14388), .ZN(n14386) );
  NOR2X0 U14879 ( .IN1(WX2040), .IN2(n8089), .QN(n14388) );
  NAND2X0 U14880 ( .IN1(n268), .IN2(n9286), .QN(n14367) );
  NOR2X0 U14881 ( .IN1(n9242), .IN2(n9014), .QN(n268) );
  NAND2X0 U14882 ( .IN1(n9299), .IN2(CRC_OUT_8_12), .QN(n14366) );
  NAND4X0 U14883 ( .IN1(n14389), .IN2(n14390), .IN3(n14391), .IN4(n14392), 
        .QN(WX1973) );
  NAND2X0 U14884 ( .IN1(n9328), .IN2(n13601), .QN(n14392) );
  NAND2X0 U14885 ( .IN1(n14393), .IN2(n14394), .QN(n13601) );
  INVX0 U14886 ( .INP(n14395), .ZN(n14394) );
  NOR2X0 U14887 ( .IN1(n14396), .IN2(n14397), .QN(n14395) );
  NAND2X0 U14888 ( .IN1(n14397), .IN2(n14396), .QN(n14393) );
  NOR2X0 U14889 ( .IN1(n14398), .IN2(n14399), .QN(n14396) );
  NOR2X0 U14890 ( .IN1(WX3459), .IN2(n8061), .QN(n14399) );
  INVX0 U14891 ( .INP(n14400), .ZN(n14398) );
  NAND2X0 U14892 ( .IN1(n8061), .IN2(WX3459), .QN(n14400) );
  NAND2X0 U14893 ( .IN1(n14401), .IN2(n14402), .QN(n14397) );
  NAND2X0 U14894 ( .IN1(n8060), .IN2(WX3331), .QN(n14402) );
  INVX0 U14895 ( .INP(n14403), .ZN(n14401) );
  NOR2X0 U14896 ( .IN1(WX3331), .IN2(n8060), .QN(n14403) );
  NAND2X0 U14897 ( .IN1(n9105), .IN2(n11741), .QN(n14391) );
  NAND2X0 U14898 ( .IN1(n14404), .IN2(n14405), .QN(n11741) );
  INVX0 U14899 ( .INP(n14406), .ZN(n14405) );
  NOR2X0 U14900 ( .IN1(n14407), .IN2(n14408), .QN(n14406) );
  NAND2X0 U14901 ( .IN1(n14408), .IN2(n14407), .QN(n14404) );
  NOR2X0 U14902 ( .IN1(n14409), .IN2(n14410), .QN(n14407) );
  NOR2X0 U14903 ( .IN1(WX2166), .IN2(n8092), .QN(n14410) );
  INVX0 U14904 ( .INP(n14411), .ZN(n14409) );
  NAND2X0 U14905 ( .IN1(n8092), .IN2(WX2166), .QN(n14411) );
  NAND2X0 U14906 ( .IN1(n14412), .IN2(n14413), .QN(n14408) );
  NAND2X0 U14907 ( .IN1(n8091), .IN2(WX2038), .QN(n14413) );
  INVX0 U14908 ( .INP(n14414), .ZN(n14412) );
  NOR2X0 U14909 ( .IN1(WX2038), .IN2(n8091), .QN(n14414) );
  NAND2X0 U14910 ( .IN1(n267), .IN2(n9286), .QN(n14390) );
  NOR2X0 U14911 ( .IN1(n9242), .IN2(n9015), .QN(n267) );
  NAND2X0 U14912 ( .IN1(n9299), .IN2(CRC_OUT_8_13), .QN(n14389) );
  NAND4X0 U14913 ( .IN1(n14415), .IN2(n14416), .IN3(n14417), .IN4(n14418), 
        .QN(WX1971) );
  NAND3X0 U14914 ( .IN1(n11747), .IN2(n11748), .IN3(n9091), .QN(n14418) );
  NAND3X0 U14915 ( .IN1(n14419), .IN2(n14420), .IN3(n14421), .QN(n11748) );
  INVX0 U14916 ( .INP(n14422), .ZN(n14421) );
  NAND2X0 U14917 ( .IN1(n14422), .IN2(n14423), .QN(n11747) );
  NAND2X0 U14918 ( .IN1(n14419), .IN2(n14420), .QN(n14423) );
  NAND2X0 U14919 ( .IN1(n8634), .IN2(WX2036), .QN(n14420) );
  NAND2X0 U14920 ( .IN1(n3783), .IN2(WX2164), .QN(n14419) );
  NOR2X0 U14921 ( .IN1(n14424), .IN2(n14425), .QN(n14422) );
  INVX0 U14922 ( .INP(n14426), .ZN(n14425) );
  NAND2X0 U14923 ( .IN1(test_so17), .IN2(WX1972), .QN(n14426) );
  NOR2X0 U14924 ( .IN1(WX1972), .IN2(test_so17), .QN(n14424) );
  NAND2X0 U14925 ( .IN1(n9328), .IN2(n13617), .QN(n14417) );
  NAND2X0 U14926 ( .IN1(n14427), .IN2(n14428), .QN(n13617) );
  INVX0 U14927 ( .INP(n14429), .ZN(n14428) );
  NOR2X0 U14928 ( .IN1(n14430), .IN2(n14431), .QN(n14429) );
  NAND2X0 U14929 ( .IN1(n14431), .IN2(n14430), .QN(n14427) );
  NOR2X0 U14930 ( .IN1(n14432), .IN2(n14433), .QN(n14430) );
  NOR2X0 U14931 ( .IN1(WX3457), .IN2(n8063), .QN(n14433) );
  INVX0 U14932 ( .INP(n14434), .ZN(n14432) );
  NAND2X0 U14933 ( .IN1(n8063), .IN2(WX3457), .QN(n14434) );
  NAND2X0 U14934 ( .IN1(n14435), .IN2(n14436), .QN(n14431) );
  NAND2X0 U14935 ( .IN1(n8062), .IN2(WX3329), .QN(n14436) );
  INVX0 U14936 ( .INP(n14437), .ZN(n14435) );
  NOR2X0 U14937 ( .IN1(WX3329), .IN2(n8062), .QN(n14437) );
  NAND2X0 U14938 ( .IN1(n266), .IN2(n9286), .QN(n14416) );
  NOR2X0 U14939 ( .IN1(n9242), .IN2(n9016), .QN(n266) );
  NAND2X0 U14940 ( .IN1(n9299), .IN2(CRC_OUT_8_14), .QN(n14415) );
  NAND4X0 U14941 ( .IN1(n14438), .IN2(n14439), .IN3(n14440), .IN4(n14441), 
        .QN(WX1969) );
  NAND2X0 U14942 ( .IN1(n9328), .IN2(n13630), .QN(n14441) );
  NAND2X0 U14943 ( .IN1(n14442), .IN2(n14443), .QN(n13630) );
  INVX0 U14944 ( .INP(n14444), .ZN(n14443) );
  NOR2X0 U14945 ( .IN1(n14445), .IN2(n14446), .QN(n14444) );
  NAND2X0 U14946 ( .IN1(n14446), .IN2(n14445), .QN(n14442) );
  NOR2X0 U14947 ( .IN1(n14447), .IN2(n14448), .QN(n14445) );
  NOR2X0 U14948 ( .IN1(WX3455), .IN2(n8065), .QN(n14448) );
  INVX0 U14949 ( .INP(n14449), .ZN(n14447) );
  NAND2X0 U14950 ( .IN1(n8065), .IN2(WX3455), .QN(n14449) );
  NAND2X0 U14951 ( .IN1(n14450), .IN2(n14451), .QN(n14446) );
  NAND2X0 U14952 ( .IN1(n8064), .IN2(WX3327), .QN(n14451) );
  INVX0 U14953 ( .INP(n14452), .ZN(n14450) );
  NOR2X0 U14954 ( .IN1(WX3327), .IN2(n8064), .QN(n14452) );
  NAND2X0 U14955 ( .IN1(n9105), .IN2(n11754), .QN(n14440) );
  NAND2X0 U14956 ( .IN1(n14453), .IN2(n14454), .QN(n11754) );
  INVX0 U14957 ( .INP(n14455), .ZN(n14454) );
  NOR2X0 U14958 ( .IN1(n14456), .IN2(n14457), .QN(n14455) );
  NAND2X0 U14959 ( .IN1(n14457), .IN2(n14456), .QN(n14453) );
  NOR2X0 U14960 ( .IN1(n14458), .IN2(n14459), .QN(n14456) );
  NOR2X0 U14961 ( .IN1(WX2162), .IN2(n8095), .QN(n14459) );
  INVX0 U14962 ( .INP(n14460), .ZN(n14458) );
  NAND2X0 U14963 ( .IN1(n8095), .IN2(WX2162), .QN(n14460) );
  NAND2X0 U14964 ( .IN1(n14461), .IN2(n14462), .QN(n14457) );
  NAND2X0 U14965 ( .IN1(n8094), .IN2(WX2034), .QN(n14462) );
  INVX0 U14966 ( .INP(n14463), .ZN(n14461) );
  NOR2X0 U14967 ( .IN1(WX2034), .IN2(n8094), .QN(n14463) );
  NAND2X0 U14968 ( .IN1(n265), .IN2(n9286), .QN(n14439) );
  NOR2X0 U14969 ( .IN1(n9227), .IN2(n9017), .QN(n265) );
  NAND2X0 U14970 ( .IN1(n9299), .IN2(CRC_OUT_8_15), .QN(n14438) );
  NAND4X0 U14971 ( .IN1(n14464), .IN2(n14465), .IN3(n14466), .IN4(n14467), 
        .QN(WX1967) );
  NAND2X0 U14972 ( .IN1(n14468), .IN2(n13650), .QN(n14467) );
  NAND3X0 U14973 ( .IN1(n14469), .IN2(n14470), .IN3(n13653), .QN(n13650) );
  NAND2X0 U14974 ( .IN1(n8120), .IN2(n9121), .QN(n14470) );
  NAND2X0 U14975 ( .IN1(TM1), .IN2(WX3453), .QN(n14469) );
  NAND3X0 U14976 ( .IN1(n14471), .IN2(n14472), .IN3(n14473), .QN(n14468) );
  NAND2X0 U14977 ( .IN1(n9328), .IN2(n13653), .QN(n14473) );
  NAND2X0 U14978 ( .IN1(n14474), .IN2(n14475), .QN(n13653) );
  NAND2X0 U14979 ( .IN1(n14476), .IN2(WX3389), .QN(n14475) );
  NAND2X0 U14980 ( .IN1(n14477), .IN2(n14478), .QN(n14476) );
  NAND3X0 U14981 ( .IN1(n14477), .IN2(n14478), .IN3(n7798), .QN(n14474) );
  NAND2X0 U14982 ( .IN1(test_so24), .IN2(WX3325), .QN(n14478) );
  NAND2X0 U14983 ( .IN1(n7797), .IN2(n8824), .QN(n14477) );
  NAND2X0 U14984 ( .IN1(n9079), .IN2(WX3453), .QN(n14472) );
  NAND2X0 U14985 ( .IN1(n9083), .IN2(n8120), .QN(n14471) );
  NAND2X0 U14986 ( .IN1(n14479), .IN2(n11761), .QN(n14466) );
  NAND2X0 U14987 ( .IN1(n14480), .IN2(n11765), .QN(n11761) );
  NAND2X0 U14988 ( .IN1(n14481), .IN2(n14482), .QN(n14480) );
  NAND2X0 U14989 ( .IN1(n16321), .IN2(n9121), .QN(n14482) );
  NAND2X0 U14990 ( .IN1(TM1), .IN2(n8653), .QN(n14481) );
  NAND2X0 U14991 ( .IN1(n14483), .IN2(n14484), .QN(n14479) );
  NAND2X0 U14992 ( .IN1(n9104), .IN2(n11765), .QN(n14484) );
  NAND2X0 U14993 ( .IN1(n14485), .IN2(n14486), .QN(n11765) );
  NAND2X0 U14994 ( .IN1(n7825), .IN2(n14487), .QN(n14486) );
  INVX0 U14995 ( .INP(n14488), .ZN(n14485) );
  NOR2X0 U14996 ( .IN1(n14487), .IN2(n7825), .QN(n14488) );
  NOR2X0 U14997 ( .IN1(n14489), .IN2(n14490), .QN(n14487) );
  NOR2X0 U14998 ( .IN1(WX2160), .IN2(n7826), .QN(n14490) );
  INVX0 U14999 ( .INP(n14491), .ZN(n14489) );
  NAND2X0 U15000 ( .IN1(n7826), .IN2(WX2160), .QN(n14491) );
  NAND2X0 U15001 ( .IN1(n9104), .IN2(n8653), .QN(n14483) );
  NAND2X0 U15002 ( .IN1(n264), .IN2(n9286), .QN(n14465) );
  NOR2X0 U15003 ( .IN1(n9227), .IN2(n9018), .QN(n264) );
  NAND2X0 U15004 ( .IN1(n9299), .IN2(CRC_OUT_8_16), .QN(n14464) );
  NAND4X0 U15005 ( .IN1(n14492), .IN2(n14493), .IN3(n14494), .IN4(n14495), 
        .QN(WX1965) );
  NAND2X0 U15006 ( .IN1(n14496), .IN2(n13670), .QN(n14495) );
  NAND2X0 U15007 ( .IN1(n14497), .IN2(n13673), .QN(n13670) );
  NAND2X0 U15008 ( .IN1(n14498), .IN2(n14499), .QN(n14497) );
  NAND2X0 U15009 ( .IN1(n16336), .IN2(n9122), .QN(n14499) );
  NAND2X0 U15010 ( .IN1(TM1), .IN2(n8597), .QN(n14498) );
  NAND3X0 U15011 ( .IN1(n14500), .IN2(n14501), .IN3(n14502), .QN(n14496) );
  NAND2X0 U15012 ( .IN1(n9328), .IN2(n13673), .QN(n14502) );
  NAND2X0 U15013 ( .IN1(n14503), .IN2(n14504), .QN(n13673) );
  NAND2X0 U15014 ( .IN1(n7799), .IN2(n14505), .QN(n14504) );
  INVX0 U15015 ( .INP(n14506), .ZN(n14503) );
  NOR2X0 U15016 ( .IN1(n14505), .IN2(n7799), .QN(n14506) );
  NOR2X0 U15017 ( .IN1(n14507), .IN2(n14508), .QN(n14505) );
  NOR2X0 U15018 ( .IN1(WX3451), .IN2(n7800), .QN(n14508) );
  INVX0 U15019 ( .INP(n14509), .ZN(n14507) );
  NAND2X0 U15020 ( .IN1(n7800), .IN2(WX3451), .QN(n14509) );
  NAND2X0 U15021 ( .IN1(n9082), .IN2(n8597), .QN(n14501) );
  NAND2X0 U15022 ( .IN1(n16336), .IN2(n9078), .QN(n14500) );
  NAND2X0 U15023 ( .IN1(n14510), .IN2(n11773), .QN(n14494) );
  NAND2X0 U15024 ( .IN1(n14511), .IN2(n11777), .QN(n11773) );
  NAND2X0 U15025 ( .IN1(n14512), .IN2(n14513), .QN(n14511) );
  NAND2X0 U15026 ( .IN1(n16320), .IN2(n9122), .QN(n14513) );
  NAND2X0 U15027 ( .IN1(TM1), .IN2(n8654), .QN(n14512) );
  NAND2X0 U15028 ( .IN1(n14514), .IN2(n14515), .QN(n14510) );
  NAND2X0 U15029 ( .IN1(n9104), .IN2(n11777), .QN(n14515) );
  NAND2X0 U15030 ( .IN1(n14516), .IN2(n14517), .QN(n11777) );
  NAND2X0 U15031 ( .IN1(n7827), .IN2(n14518), .QN(n14517) );
  INVX0 U15032 ( .INP(n14519), .ZN(n14516) );
  NOR2X0 U15033 ( .IN1(n14518), .IN2(n7827), .QN(n14519) );
  NOR2X0 U15034 ( .IN1(n14520), .IN2(n14521), .QN(n14518) );
  NOR2X0 U15035 ( .IN1(WX2158), .IN2(n7828), .QN(n14521) );
  INVX0 U15036 ( .INP(n14522), .ZN(n14520) );
  NAND2X0 U15037 ( .IN1(n7828), .IN2(WX2158), .QN(n14522) );
  NAND2X0 U15038 ( .IN1(n9104), .IN2(n8654), .QN(n14514) );
  NAND2X0 U15039 ( .IN1(n263), .IN2(n9286), .QN(n14493) );
  NOR2X0 U15040 ( .IN1(n9227), .IN2(n9019), .QN(n263) );
  NAND2X0 U15041 ( .IN1(n9299), .IN2(CRC_OUT_8_17), .QN(n14492) );
  NAND4X0 U15042 ( .IN1(n14523), .IN2(n14524), .IN3(n14525), .IN4(n14526), 
        .QN(WX1963) );
  NAND2X0 U15043 ( .IN1(n14527), .IN2(n13693), .QN(n14526) );
  NAND2X0 U15044 ( .IN1(n14528), .IN2(n13696), .QN(n13693) );
  NAND2X0 U15045 ( .IN1(n14529), .IN2(n14530), .QN(n14528) );
  NAND2X0 U15046 ( .IN1(n16335), .IN2(n9122), .QN(n14530) );
  NAND2X0 U15047 ( .IN1(TM1), .IN2(n8598), .QN(n14529) );
  NAND3X0 U15048 ( .IN1(n14531), .IN2(n14532), .IN3(n14533), .QN(n14527) );
  NAND2X0 U15049 ( .IN1(n9328), .IN2(n13696), .QN(n14533) );
  NAND2X0 U15050 ( .IN1(n14534), .IN2(n14535), .QN(n13696) );
  NAND2X0 U15051 ( .IN1(n7801), .IN2(n14536), .QN(n14535) );
  INVX0 U15052 ( .INP(n14537), .ZN(n14534) );
  NOR2X0 U15053 ( .IN1(n14536), .IN2(n7801), .QN(n14537) );
  NOR2X0 U15054 ( .IN1(n14538), .IN2(n14539), .QN(n14536) );
  NOR2X0 U15055 ( .IN1(WX3449), .IN2(n7802), .QN(n14539) );
  INVX0 U15056 ( .INP(n14540), .ZN(n14538) );
  NAND2X0 U15057 ( .IN1(n7802), .IN2(WX3449), .QN(n14540) );
  NAND2X0 U15058 ( .IN1(n10068), .IN2(n8598), .QN(n14532) );
  NAND2X0 U15059 ( .IN1(n16335), .IN2(n10069), .QN(n14531) );
  NAND2X0 U15060 ( .IN1(n11783), .IN2(n9111), .QN(n14525) );
  NOR2X0 U15061 ( .IN1(n14541), .IN2(n14542), .QN(n11783) );
  INVX0 U15062 ( .INP(n14543), .ZN(n14542) );
  NAND2X0 U15063 ( .IN1(n14544), .IN2(n14545), .QN(n14543) );
  NOR2X0 U15064 ( .IN1(n14545), .IN2(n14544), .QN(n14541) );
  NAND2X0 U15065 ( .IN1(n14546), .IN2(n14547), .QN(n14544) );
  NAND2X0 U15066 ( .IN1(n8614), .IN2(n14548), .QN(n14547) );
  INVX0 U15067 ( .INP(n14549), .ZN(n14548) );
  NAND2X0 U15068 ( .IN1(n14549), .IN2(WX2156), .QN(n14546) );
  NAND2X0 U15069 ( .IN1(n14550), .IN2(n14551), .QN(n14549) );
  INVX0 U15070 ( .INP(n14552), .ZN(n14551) );
  NOR2X0 U15071 ( .IN1(n8815), .IN2(n16319), .QN(n14552) );
  NAND2X0 U15072 ( .IN1(n16319), .IN2(n8815), .QN(n14550) );
  NOR2X0 U15073 ( .IN1(n14553), .IN2(n14554), .QN(n14545) );
  INVX0 U15074 ( .INP(n14555), .ZN(n14554) );
  NAND2X0 U15075 ( .IN1(n7829), .IN2(n9122), .QN(n14555) );
  NOR2X0 U15076 ( .IN1(n9117), .IN2(n7829), .QN(n14553) );
  NAND2X0 U15077 ( .IN1(n262), .IN2(n9286), .QN(n14524) );
  NOR2X0 U15078 ( .IN1(n9227), .IN2(n9020), .QN(n262) );
  NAND2X0 U15079 ( .IN1(n9300), .IN2(CRC_OUT_8_18), .QN(n14523) );
  NAND4X0 U15080 ( .IN1(n14556), .IN2(n14557), .IN3(n14558), .IN4(n14559), 
        .QN(WX1961) );
  NAND2X0 U15081 ( .IN1(n14560), .IN2(n13716), .QN(n14559) );
  NAND2X0 U15082 ( .IN1(n14561), .IN2(n13719), .QN(n13716) );
  NAND2X0 U15083 ( .IN1(n14562), .IN2(n14563), .QN(n14561) );
  NAND2X0 U15084 ( .IN1(n16334), .IN2(n9122), .QN(n14563) );
  NAND2X0 U15085 ( .IN1(TM1), .IN2(n8599), .QN(n14562) );
  NAND3X0 U15086 ( .IN1(n14564), .IN2(n14565), .IN3(n14566), .QN(n14560) );
  NAND2X0 U15087 ( .IN1(n9328), .IN2(n13719), .QN(n14566) );
  NAND2X0 U15088 ( .IN1(n14567), .IN2(n14568), .QN(n13719) );
  NAND2X0 U15089 ( .IN1(n7803), .IN2(n14569), .QN(n14568) );
  INVX0 U15090 ( .INP(n14570), .ZN(n14567) );
  NOR2X0 U15091 ( .IN1(n14569), .IN2(n7803), .QN(n14570) );
  NOR2X0 U15092 ( .IN1(n14571), .IN2(n14572), .QN(n14569) );
  NOR2X0 U15093 ( .IN1(WX3447), .IN2(n7804), .QN(n14572) );
  INVX0 U15094 ( .INP(n14573), .ZN(n14571) );
  NAND2X0 U15095 ( .IN1(n7804), .IN2(WX3447), .QN(n14573) );
  NAND2X0 U15096 ( .IN1(n9084), .IN2(n8599), .QN(n14565) );
  NAND2X0 U15097 ( .IN1(n16334), .IN2(n9080), .QN(n14564) );
  NAND2X0 U15098 ( .IN1(n14574), .IN2(n11790), .QN(n14558) );
  NAND2X0 U15099 ( .IN1(n14575), .IN2(n11794), .QN(n11790) );
  NAND2X0 U15100 ( .IN1(n14576), .IN2(n14577), .QN(n14575) );
  NAND2X0 U15101 ( .IN1(n16318), .IN2(n9122), .QN(n14577) );
  NAND2X0 U15102 ( .IN1(TM1), .IN2(n8656), .QN(n14576) );
  NAND2X0 U15103 ( .IN1(n14578), .IN2(n14579), .QN(n14574) );
  NAND2X0 U15104 ( .IN1(n9104), .IN2(n11794), .QN(n14579) );
  NAND2X0 U15105 ( .IN1(n14580), .IN2(n14581), .QN(n11794) );
  NAND2X0 U15106 ( .IN1(n7830), .IN2(n14582), .QN(n14581) );
  INVX0 U15107 ( .INP(n14583), .ZN(n14580) );
  NOR2X0 U15108 ( .IN1(n14582), .IN2(n7830), .QN(n14583) );
  NOR2X0 U15109 ( .IN1(n14584), .IN2(n14585), .QN(n14582) );
  NOR2X0 U15110 ( .IN1(WX2154), .IN2(n7831), .QN(n14585) );
  INVX0 U15111 ( .INP(n14586), .ZN(n14584) );
  NAND2X0 U15112 ( .IN1(n7831), .IN2(WX2154), .QN(n14586) );
  NAND2X0 U15113 ( .IN1(n9104), .IN2(n8656), .QN(n14578) );
  NAND2X0 U15114 ( .IN1(n261), .IN2(n9286), .QN(n14557) );
  NOR2X0 U15115 ( .IN1(n9227), .IN2(n9021), .QN(n261) );
  NAND2X0 U15116 ( .IN1(n9300), .IN2(CRC_OUT_8_19), .QN(n14556) );
  NAND4X0 U15117 ( .IN1(n14587), .IN2(n14588), .IN3(n14589), .IN4(n14590), 
        .QN(WX1959) );
  NAND2X0 U15118 ( .IN1(n14591), .IN2(n13739), .QN(n14590) );
  NAND2X0 U15119 ( .IN1(n14592), .IN2(n13742), .QN(n13739) );
  NAND2X0 U15120 ( .IN1(n14593), .IN2(n14594), .QN(n14592) );
  NAND2X0 U15121 ( .IN1(n16333), .IN2(n9122), .QN(n14594) );
  NAND2X0 U15122 ( .IN1(TM1), .IN2(n8600), .QN(n14593) );
  NAND3X0 U15123 ( .IN1(n14595), .IN2(n14596), .IN3(n14597), .QN(n14591) );
  NAND2X0 U15124 ( .IN1(n9328), .IN2(n13742), .QN(n14597) );
  NAND2X0 U15125 ( .IN1(n14598), .IN2(n14599), .QN(n13742) );
  NAND2X0 U15126 ( .IN1(n7805), .IN2(n14600), .QN(n14599) );
  INVX0 U15127 ( .INP(n14601), .ZN(n14598) );
  NOR2X0 U15128 ( .IN1(n14600), .IN2(n7805), .QN(n14601) );
  NOR2X0 U15129 ( .IN1(n14602), .IN2(n14603), .QN(n14600) );
  NOR2X0 U15130 ( .IN1(WX3445), .IN2(n7806), .QN(n14603) );
  INVX0 U15131 ( .INP(n14604), .ZN(n14602) );
  NAND2X0 U15132 ( .IN1(n7806), .IN2(WX3445), .QN(n14604) );
  NAND2X0 U15133 ( .IN1(n9083), .IN2(n8600), .QN(n14596) );
  NAND2X0 U15134 ( .IN1(n16333), .IN2(n9079), .QN(n14595) );
  NAND2X0 U15135 ( .IN1(n14605), .IN2(n11801), .QN(n14589) );
  NAND2X0 U15136 ( .IN1(n14606), .IN2(n11805), .QN(n11801) );
  NAND2X0 U15137 ( .IN1(n14607), .IN2(n14608), .QN(n14606) );
  NAND2X0 U15138 ( .IN1(n16317), .IN2(n9122), .QN(n14608) );
  NAND2X0 U15139 ( .IN1(TM1), .IN2(n8657), .QN(n14607) );
  NAND2X0 U15140 ( .IN1(n14609), .IN2(n14610), .QN(n14605) );
  NAND2X0 U15141 ( .IN1(n9104), .IN2(n11805), .QN(n14610) );
  NAND2X0 U15142 ( .IN1(n14611), .IN2(n14612), .QN(n11805) );
  NAND2X0 U15143 ( .IN1(n7832), .IN2(n14613), .QN(n14612) );
  INVX0 U15144 ( .INP(n14614), .ZN(n14611) );
  NOR2X0 U15145 ( .IN1(n14613), .IN2(n7832), .QN(n14614) );
  NOR2X0 U15146 ( .IN1(n14615), .IN2(n14616), .QN(n14613) );
  NOR2X0 U15147 ( .IN1(WX2152), .IN2(n7833), .QN(n14616) );
  INVX0 U15148 ( .INP(n14617), .ZN(n14615) );
  NAND2X0 U15149 ( .IN1(n7833), .IN2(WX2152), .QN(n14617) );
  NAND2X0 U15150 ( .IN1(n9104), .IN2(n8657), .QN(n14609) );
  NAND2X0 U15151 ( .IN1(n260), .IN2(n9287), .QN(n14588) );
  NOR2X0 U15152 ( .IN1(n9227), .IN2(n9022), .QN(n260) );
  NAND2X0 U15153 ( .IN1(n9300), .IN2(CRC_OUT_8_20), .QN(n14587) );
  NAND4X0 U15154 ( .IN1(n14618), .IN2(n14619), .IN3(n14620), .IN4(n14621), 
        .QN(WX1957) );
  NAND2X0 U15155 ( .IN1(n14622), .IN2(n13762), .QN(n14621) );
  NAND2X0 U15156 ( .IN1(n14623), .IN2(n13765), .QN(n13762) );
  NAND2X0 U15157 ( .IN1(n14624), .IN2(n14625), .QN(n14623) );
  NAND2X0 U15158 ( .IN1(n16332), .IN2(n9122), .QN(n14625) );
  NAND2X0 U15159 ( .IN1(TM1), .IN2(n8601), .QN(n14624) );
  NAND3X0 U15160 ( .IN1(n14626), .IN2(n14627), .IN3(n14628), .QN(n14622) );
  NAND2X0 U15161 ( .IN1(n9328), .IN2(n13765), .QN(n14628) );
  NAND2X0 U15162 ( .IN1(n14629), .IN2(n14630), .QN(n13765) );
  NAND2X0 U15163 ( .IN1(n7807), .IN2(n14631), .QN(n14630) );
  INVX0 U15164 ( .INP(n14632), .ZN(n14629) );
  NOR2X0 U15165 ( .IN1(n14631), .IN2(n7807), .QN(n14632) );
  NOR2X0 U15166 ( .IN1(n14633), .IN2(n14634), .QN(n14631) );
  NOR2X0 U15167 ( .IN1(WX3443), .IN2(n7808), .QN(n14634) );
  INVX0 U15168 ( .INP(n14635), .ZN(n14633) );
  NAND2X0 U15169 ( .IN1(n7808), .IN2(WX3443), .QN(n14635) );
  NAND2X0 U15170 ( .IN1(n9082), .IN2(n8601), .QN(n14627) );
  NAND2X0 U15171 ( .IN1(n16332), .IN2(n9078), .QN(n14626) );
  NAND2X0 U15172 ( .IN1(n14636), .IN2(n11813), .QN(n14620) );
  NAND2X0 U15173 ( .IN1(n14637), .IN2(n11817), .QN(n11813) );
  NAND2X0 U15174 ( .IN1(n14638), .IN2(n14639), .QN(n14637) );
  NAND2X0 U15175 ( .IN1(n16316), .IN2(n9122), .QN(n14639) );
  NAND2X0 U15176 ( .IN1(TM1), .IN2(n8658), .QN(n14638) );
  NAND2X0 U15177 ( .IN1(n14640), .IN2(n14641), .QN(n14636) );
  NAND2X0 U15178 ( .IN1(n9104), .IN2(n11817), .QN(n14641) );
  NAND2X0 U15179 ( .IN1(n14642), .IN2(n14643), .QN(n11817) );
  NAND2X0 U15180 ( .IN1(n7834), .IN2(n14644), .QN(n14643) );
  INVX0 U15181 ( .INP(n14645), .ZN(n14642) );
  NOR2X0 U15182 ( .IN1(n14644), .IN2(n7834), .QN(n14645) );
  NOR2X0 U15183 ( .IN1(n14646), .IN2(n14647), .QN(n14644) );
  NOR2X0 U15184 ( .IN1(WX2150), .IN2(n7835), .QN(n14647) );
  INVX0 U15185 ( .INP(n14648), .ZN(n14646) );
  NAND2X0 U15186 ( .IN1(n7835), .IN2(WX2150), .QN(n14648) );
  NAND2X0 U15187 ( .IN1(n9104), .IN2(n8658), .QN(n14640) );
  NAND2X0 U15188 ( .IN1(n259), .IN2(n9287), .QN(n14619) );
  NOR2X0 U15189 ( .IN1(n9227), .IN2(n9023), .QN(n259) );
  NAND2X0 U15190 ( .IN1(n9300), .IN2(CRC_OUT_8_21), .QN(n14618) );
  NAND4X0 U15191 ( .IN1(n14649), .IN2(n14650), .IN3(n14651), .IN4(n14652), 
        .QN(WX1955) );
  NAND2X0 U15192 ( .IN1(n14653), .IN2(n13785), .QN(n14652) );
  NAND2X0 U15193 ( .IN1(n14654), .IN2(n13788), .QN(n13785) );
  NAND2X0 U15194 ( .IN1(n14655), .IN2(n14656), .QN(n14654) );
  NAND2X0 U15195 ( .IN1(n16331), .IN2(n9122), .QN(n14656) );
  NAND2X0 U15196 ( .IN1(TM1), .IN2(n8602), .QN(n14655) );
  NAND3X0 U15197 ( .IN1(n14657), .IN2(n14658), .IN3(n14659), .QN(n14653) );
  NAND2X0 U15198 ( .IN1(n9328), .IN2(n13788), .QN(n14659) );
  NAND2X0 U15199 ( .IN1(n14660), .IN2(n14661), .QN(n13788) );
  NAND2X0 U15200 ( .IN1(n7809), .IN2(n14662), .QN(n14661) );
  INVX0 U15201 ( .INP(n14663), .ZN(n14660) );
  NOR2X0 U15202 ( .IN1(n14662), .IN2(n7809), .QN(n14663) );
  NOR2X0 U15203 ( .IN1(n14664), .IN2(n14665), .QN(n14662) );
  NOR2X0 U15204 ( .IN1(WX3441), .IN2(n7810), .QN(n14665) );
  INVX0 U15205 ( .INP(n14666), .ZN(n14664) );
  NAND2X0 U15206 ( .IN1(n7810), .IN2(WX3441), .QN(n14666) );
  NAND2X0 U15207 ( .IN1(n10068), .IN2(n8602), .QN(n14658) );
  NAND2X0 U15208 ( .IN1(n16331), .IN2(n10069), .QN(n14657) );
  NAND2X0 U15209 ( .IN1(n14667), .IN2(n11824), .QN(n14651) );
  NAND3X0 U15210 ( .IN1(n14668), .IN2(n14669), .IN3(n11828), .QN(n11824) );
  NAND2X0 U15211 ( .IN1(n8593), .IN2(n9122), .QN(n14669) );
  NAND2X0 U15212 ( .IN1(TM1), .IN2(WX2148), .QN(n14668) );
  NAND2X0 U15213 ( .IN1(n14670), .IN2(n14671), .QN(n14667) );
  NAND2X0 U15214 ( .IN1(n9104), .IN2(n11828), .QN(n14671) );
  NAND2X0 U15215 ( .IN1(n14672), .IN2(n14673), .QN(n11828) );
  NAND2X0 U15216 ( .IN1(n14674), .IN2(WX2084), .QN(n14673) );
  NAND2X0 U15217 ( .IN1(n14675), .IN2(n14676), .QN(n14674) );
  NAND3X0 U15218 ( .IN1(n14675), .IN2(n14676), .IN3(n7837), .QN(n14672) );
  NAND2X0 U15219 ( .IN1(test_so13), .IN2(WX2020), .QN(n14676) );
  NAND2X0 U15220 ( .IN1(n7836), .IN2(n8825), .QN(n14675) );
  NAND2X0 U15221 ( .IN1(n8593), .IN2(n9110), .QN(n14670) );
  NAND2X0 U15222 ( .IN1(n258), .IN2(n9287), .QN(n14650) );
  NOR2X0 U15223 ( .IN1(n9227), .IN2(n9024), .QN(n258) );
  NAND2X0 U15224 ( .IN1(n9300), .IN2(CRC_OUT_8_22), .QN(n14649) );
  NAND4X0 U15225 ( .IN1(n14677), .IN2(n14678), .IN3(n14679), .IN4(n14680), 
        .QN(WX1953) );
  NAND2X0 U15226 ( .IN1(n14681), .IN2(n11835), .QN(n14680) );
  NAND2X0 U15227 ( .IN1(n14682), .IN2(n11839), .QN(n11835) );
  NAND2X0 U15228 ( .IN1(n14683), .IN2(n14684), .QN(n14682) );
  NAND2X0 U15229 ( .IN1(n16315), .IN2(n9122), .QN(n14684) );
  NAND2X0 U15230 ( .IN1(TM1), .IN2(n8661), .QN(n14683) );
  NAND2X0 U15231 ( .IN1(n14685), .IN2(n14686), .QN(n14681) );
  NAND2X0 U15232 ( .IN1(n9104), .IN2(n11839), .QN(n14686) );
  NAND2X0 U15233 ( .IN1(n14687), .IN2(n14688), .QN(n11839) );
  NAND2X0 U15234 ( .IN1(n7838), .IN2(n14689), .QN(n14688) );
  INVX0 U15235 ( .INP(n14690), .ZN(n14687) );
  NOR2X0 U15236 ( .IN1(n14689), .IN2(n7838), .QN(n14690) );
  NOR2X0 U15237 ( .IN1(n14691), .IN2(n14692), .QN(n14689) );
  NOR2X0 U15238 ( .IN1(WX2146), .IN2(n7839), .QN(n14692) );
  INVX0 U15239 ( .INP(n14693), .ZN(n14691) );
  NAND2X0 U15240 ( .IN1(n7839), .IN2(WX2146), .QN(n14693) );
  NAND2X0 U15241 ( .IN1(n9104), .IN2(n8661), .QN(n14685) );
  NAND2X0 U15242 ( .IN1(n13807), .IN2(n9336), .QN(n14679) );
  NOR2X0 U15243 ( .IN1(n14694), .IN2(n14695), .QN(n13807) );
  INVX0 U15244 ( .INP(n14696), .ZN(n14695) );
  NAND2X0 U15245 ( .IN1(n14697), .IN2(n14698), .QN(n14696) );
  NOR2X0 U15246 ( .IN1(n14698), .IN2(n14697), .QN(n14694) );
  NAND2X0 U15247 ( .IN1(n14699), .IN2(n14700), .QN(n14697) );
  NAND2X0 U15248 ( .IN1(n14701), .IN2(WX3375), .QN(n14700) );
  NAND2X0 U15249 ( .IN1(n14702), .IN2(n14703), .QN(n14701) );
  NAND3X0 U15250 ( .IN1(n14702), .IN2(n14703), .IN3(n7812), .QN(n14699) );
  NAND2X0 U15251 ( .IN1(test_so29), .IN2(WX3311), .QN(n14703) );
  NAND2X0 U15252 ( .IN1(n7811), .IN2(n8802), .QN(n14702) );
  NOR2X0 U15253 ( .IN1(n14704), .IN2(n14705), .QN(n14698) );
  INVX0 U15254 ( .INP(n14706), .ZN(n14705) );
  NAND2X0 U15255 ( .IN1(n16330), .IN2(n9122), .QN(n14706) );
  NOR2X0 U15256 ( .IN1(n9118), .IN2(n16330), .QN(n14704) );
  NAND2X0 U15257 ( .IN1(n257), .IN2(n9287), .QN(n14678) );
  NOR2X0 U15258 ( .IN1(n9226), .IN2(n9025), .QN(n257) );
  NAND2X0 U15259 ( .IN1(n9300), .IN2(CRC_OUT_8_23), .QN(n14677) );
  NAND4X0 U15260 ( .IN1(n14707), .IN2(n14708), .IN3(n14709), .IN4(n14710), 
        .QN(WX1951) );
  NAND2X0 U15261 ( .IN1(n14711), .IN2(n13827), .QN(n14710) );
  NAND2X0 U15262 ( .IN1(n14712), .IN2(n13830), .QN(n13827) );
  NAND2X0 U15263 ( .IN1(n14713), .IN2(n14714), .QN(n14712) );
  NAND2X0 U15264 ( .IN1(n16329), .IN2(n9122), .QN(n14714) );
  NAND2X0 U15265 ( .IN1(TM1), .IN2(n8604), .QN(n14713) );
  NAND3X0 U15266 ( .IN1(n14715), .IN2(n14716), .IN3(n14717), .QN(n14711) );
  NAND2X0 U15267 ( .IN1(n9328), .IN2(n13830), .QN(n14717) );
  NAND2X0 U15268 ( .IN1(n14718), .IN2(n14719), .QN(n13830) );
  NAND2X0 U15269 ( .IN1(n7813), .IN2(n14720), .QN(n14719) );
  INVX0 U15270 ( .INP(n14721), .ZN(n14718) );
  NOR2X0 U15271 ( .IN1(n14720), .IN2(n7813), .QN(n14721) );
  NOR2X0 U15272 ( .IN1(n14722), .IN2(n14723), .QN(n14720) );
  NOR2X0 U15273 ( .IN1(WX3437), .IN2(n7814), .QN(n14723) );
  INVX0 U15274 ( .INP(n14724), .ZN(n14722) );
  NAND2X0 U15275 ( .IN1(n7814), .IN2(WX3437), .QN(n14724) );
  NAND2X0 U15276 ( .IN1(n9084), .IN2(n8604), .QN(n14716) );
  NAND2X0 U15277 ( .IN1(n16329), .IN2(n9080), .QN(n14715) );
  NAND2X0 U15278 ( .IN1(n14725), .IN2(n11846), .QN(n14709) );
  NAND2X0 U15279 ( .IN1(n14726), .IN2(n11850), .QN(n11846) );
  NAND2X0 U15280 ( .IN1(n14727), .IN2(n14728), .QN(n14726) );
  NAND2X0 U15281 ( .IN1(n16314), .IN2(n9122), .QN(n14728) );
  NAND2X0 U15282 ( .IN1(TM1), .IN2(n8662), .QN(n14727) );
  NAND2X0 U15283 ( .IN1(n14729), .IN2(n14730), .QN(n14725) );
  NAND2X0 U15284 ( .IN1(n9104), .IN2(n11850), .QN(n14730) );
  NAND2X0 U15285 ( .IN1(n14731), .IN2(n14732), .QN(n11850) );
  NAND2X0 U15286 ( .IN1(n7840), .IN2(n14733), .QN(n14732) );
  INVX0 U15287 ( .INP(n14734), .ZN(n14731) );
  NOR2X0 U15288 ( .IN1(n14733), .IN2(n7840), .QN(n14734) );
  NOR2X0 U15289 ( .IN1(n14735), .IN2(n14736), .QN(n14733) );
  NOR2X0 U15290 ( .IN1(WX2144), .IN2(n7841), .QN(n14736) );
  INVX0 U15291 ( .INP(n14737), .ZN(n14735) );
  NAND2X0 U15292 ( .IN1(n7841), .IN2(WX2144), .QN(n14737) );
  NAND2X0 U15293 ( .IN1(n9104), .IN2(n8662), .QN(n14729) );
  NAND2X0 U15294 ( .IN1(n256), .IN2(n9287), .QN(n14708) );
  NOR2X0 U15295 ( .IN1(n9226), .IN2(n9026), .QN(n256) );
  NAND2X0 U15296 ( .IN1(n9300), .IN2(CRC_OUT_8_24), .QN(n14707) );
  NAND4X0 U15297 ( .IN1(n14738), .IN2(n14739), .IN3(n14740), .IN4(n14741), 
        .QN(WX1949) );
  NAND2X0 U15298 ( .IN1(n14742), .IN2(n13850), .QN(n14741) );
  NAND2X0 U15299 ( .IN1(n14743), .IN2(n13853), .QN(n13850) );
  NAND2X0 U15300 ( .IN1(n14744), .IN2(n14745), .QN(n14743) );
  NAND2X0 U15301 ( .IN1(n16328), .IN2(n9122), .QN(n14745) );
  NAND2X0 U15302 ( .IN1(TM1), .IN2(n8605), .QN(n14744) );
  NAND3X0 U15303 ( .IN1(n14746), .IN2(n14747), .IN3(n14748), .QN(n14742) );
  NAND2X0 U15304 ( .IN1(n9328), .IN2(n13853), .QN(n14748) );
  NAND2X0 U15305 ( .IN1(n14749), .IN2(n14750), .QN(n13853) );
  NAND2X0 U15306 ( .IN1(n7815), .IN2(n14751), .QN(n14750) );
  INVX0 U15307 ( .INP(n14752), .ZN(n14749) );
  NOR2X0 U15308 ( .IN1(n14751), .IN2(n7815), .QN(n14752) );
  NOR2X0 U15309 ( .IN1(n14753), .IN2(n14754), .QN(n14751) );
  NOR2X0 U15310 ( .IN1(WX3435), .IN2(n7816), .QN(n14754) );
  INVX0 U15311 ( .INP(n14755), .ZN(n14753) );
  NAND2X0 U15312 ( .IN1(n7816), .IN2(WX3435), .QN(n14755) );
  NAND2X0 U15313 ( .IN1(n9083), .IN2(n8605), .QN(n14747) );
  NAND2X0 U15314 ( .IN1(n16328), .IN2(n9079), .QN(n14746) );
  NAND2X0 U15315 ( .IN1(n14756), .IN2(n11858), .QN(n14740) );
  NAND2X0 U15316 ( .IN1(n14757), .IN2(n11862), .QN(n11858) );
  NAND2X0 U15317 ( .IN1(n14758), .IN2(n14759), .QN(n14757) );
  NAND2X0 U15318 ( .IN1(n16313), .IN2(n9122), .QN(n14759) );
  NAND2X0 U15319 ( .IN1(TM1), .IN2(n8663), .QN(n14758) );
  NAND2X0 U15320 ( .IN1(n14760), .IN2(n14761), .QN(n14756) );
  NAND2X0 U15321 ( .IN1(n9104), .IN2(n11862), .QN(n14761) );
  NAND2X0 U15322 ( .IN1(n14762), .IN2(n14763), .QN(n11862) );
  NAND2X0 U15323 ( .IN1(n7842), .IN2(n14764), .QN(n14763) );
  INVX0 U15324 ( .INP(n14765), .ZN(n14762) );
  NOR2X0 U15325 ( .IN1(n14764), .IN2(n7842), .QN(n14765) );
  NOR2X0 U15326 ( .IN1(n14766), .IN2(n14767), .QN(n14764) );
  NOR2X0 U15327 ( .IN1(WX2142), .IN2(n7843), .QN(n14767) );
  INVX0 U15328 ( .INP(n14768), .ZN(n14766) );
  NAND2X0 U15329 ( .IN1(n7843), .IN2(WX2142), .QN(n14768) );
  NAND2X0 U15330 ( .IN1(n9104), .IN2(n8663), .QN(n14760) );
  NAND2X0 U15331 ( .IN1(n255), .IN2(n9287), .QN(n14739) );
  NOR2X0 U15332 ( .IN1(n9226), .IN2(n9027), .QN(n255) );
  NAND2X0 U15333 ( .IN1(test_so21), .IN2(n9315), .QN(n14738) );
  NAND4X0 U15334 ( .IN1(n14769), .IN2(n14770), .IN3(n14771), .IN4(n14772), 
        .QN(WX1947) );
  NAND2X0 U15335 ( .IN1(n14773), .IN2(n11869), .QN(n14772) );
  NAND2X0 U15336 ( .IN1(n14774), .IN2(n11873), .QN(n11869) );
  NAND2X0 U15337 ( .IN1(n14775), .IN2(n14776), .QN(n14774) );
  NAND2X0 U15338 ( .IN1(n16312), .IN2(n9122), .QN(n14776) );
  NAND2X0 U15339 ( .IN1(TM1), .IN2(n8664), .QN(n14775) );
  NAND2X0 U15340 ( .IN1(n14777), .IN2(n14778), .QN(n14773) );
  NAND2X0 U15341 ( .IN1(n9104), .IN2(n11873), .QN(n14778) );
  NAND2X0 U15342 ( .IN1(n14779), .IN2(n14780), .QN(n11873) );
  NAND2X0 U15343 ( .IN1(n7844), .IN2(n14781), .QN(n14780) );
  INVX0 U15344 ( .INP(n14782), .ZN(n14779) );
  NOR2X0 U15345 ( .IN1(n14781), .IN2(n7844), .QN(n14782) );
  NOR2X0 U15346 ( .IN1(n14783), .IN2(n14784), .QN(n14781) );
  NOR2X0 U15347 ( .IN1(WX2140), .IN2(n7845), .QN(n14784) );
  INVX0 U15348 ( .INP(n14785), .ZN(n14783) );
  NAND2X0 U15349 ( .IN1(n7845), .IN2(WX2140), .QN(n14785) );
  NAND2X0 U15350 ( .IN1(n9103), .IN2(n8664), .QN(n14777) );
  NAND2X0 U15351 ( .IN1(n13872), .IN2(n9336), .QN(n14771) );
  NOR2X0 U15352 ( .IN1(n14786), .IN2(n14787), .QN(n13872) );
  INVX0 U15353 ( .INP(n14788), .ZN(n14787) );
  NAND2X0 U15354 ( .IN1(n14789), .IN2(n14790), .QN(n14788) );
  NOR2X0 U15355 ( .IN1(n14790), .IN2(n14789), .QN(n14786) );
  NAND2X0 U15356 ( .IN1(n14791), .IN2(n14792), .QN(n14789) );
  NAND2X0 U15357 ( .IN1(n8476), .IN2(n14793), .QN(n14792) );
  INVX0 U15358 ( .INP(n14794), .ZN(n14793) );
  NAND2X0 U15359 ( .IN1(n14794), .IN2(WX3433), .QN(n14791) );
  NAND2X0 U15360 ( .IN1(n14795), .IN2(n14796), .QN(n14794) );
  INVX0 U15361 ( .INP(n14797), .ZN(n14796) );
  NOR2X0 U15362 ( .IN1(n8816), .IN2(n16327), .QN(n14797) );
  NAND2X0 U15363 ( .IN1(n16327), .IN2(n8816), .QN(n14795) );
  NOR2X0 U15364 ( .IN1(n14798), .IN2(n14799), .QN(n14790) );
  INVX0 U15365 ( .INP(n14800), .ZN(n14799) );
  NAND2X0 U15366 ( .IN1(n7817), .IN2(n9122), .QN(n14800) );
  NOR2X0 U15367 ( .IN1(n9118), .IN2(n7817), .QN(n14798) );
  NAND2X0 U15368 ( .IN1(n254), .IN2(n9287), .QN(n14770) );
  NOR2X0 U15369 ( .IN1(n9074), .IN2(n9162), .QN(n254) );
  NAND2X0 U15370 ( .IN1(n9300), .IN2(CRC_OUT_8_26), .QN(n14769) );
  NAND4X0 U15371 ( .IN1(n14801), .IN2(n14802), .IN3(n14803), .IN4(n14804), 
        .QN(WX1945) );
  NAND2X0 U15372 ( .IN1(n14805), .IN2(n13892), .QN(n14804) );
  NAND2X0 U15373 ( .IN1(n14806), .IN2(n13895), .QN(n13892) );
  NAND2X0 U15374 ( .IN1(n14807), .IN2(n14808), .QN(n14806) );
  NAND2X0 U15375 ( .IN1(n16326), .IN2(n9122), .QN(n14808) );
  NAND2X0 U15376 ( .IN1(TM1), .IN2(n8607), .QN(n14807) );
  NAND3X0 U15377 ( .IN1(n14809), .IN2(n14810), .IN3(n14811), .QN(n14805) );
  NAND2X0 U15378 ( .IN1(n9328), .IN2(n13895), .QN(n14811) );
  NAND2X0 U15379 ( .IN1(n14812), .IN2(n14813), .QN(n13895) );
  NAND2X0 U15380 ( .IN1(n7818), .IN2(n14814), .QN(n14813) );
  INVX0 U15381 ( .INP(n14815), .ZN(n14812) );
  NOR2X0 U15382 ( .IN1(n14814), .IN2(n7818), .QN(n14815) );
  NOR2X0 U15383 ( .IN1(n14816), .IN2(n14817), .QN(n14814) );
  NOR2X0 U15384 ( .IN1(WX3431), .IN2(n7819), .QN(n14817) );
  INVX0 U15385 ( .INP(n14818), .ZN(n14816) );
  NAND2X0 U15386 ( .IN1(n7819), .IN2(WX3431), .QN(n14818) );
  NAND2X0 U15387 ( .IN1(n9082), .IN2(n8607), .QN(n14810) );
  NAND2X0 U15388 ( .IN1(n16326), .IN2(n9078), .QN(n14809) );
  NAND2X0 U15389 ( .IN1(n14819), .IN2(n11880), .QN(n14803) );
  NAND2X0 U15390 ( .IN1(n14820), .IN2(n11884), .QN(n11880) );
  NAND2X0 U15391 ( .IN1(n14821), .IN2(n14822), .QN(n14820) );
  NAND2X0 U15392 ( .IN1(n16311), .IN2(n9122), .QN(n14822) );
  NAND2X0 U15393 ( .IN1(TM1), .IN2(n8665), .QN(n14821) );
  NAND2X0 U15394 ( .IN1(n14823), .IN2(n14824), .QN(n14819) );
  NAND2X0 U15395 ( .IN1(n9103), .IN2(n11884), .QN(n14824) );
  NAND2X0 U15396 ( .IN1(n14825), .IN2(n14826), .QN(n11884) );
  NAND2X0 U15397 ( .IN1(n7846), .IN2(n14827), .QN(n14826) );
  INVX0 U15398 ( .INP(n14828), .ZN(n14825) );
  NOR2X0 U15399 ( .IN1(n14827), .IN2(n7846), .QN(n14828) );
  NOR2X0 U15400 ( .IN1(n14829), .IN2(n14830), .QN(n14827) );
  NOR2X0 U15401 ( .IN1(WX2138), .IN2(n7847), .QN(n14830) );
  INVX0 U15402 ( .INP(n14831), .ZN(n14829) );
  NAND2X0 U15403 ( .IN1(n7847), .IN2(WX2138), .QN(n14831) );
  NAND2X0 U15404 ( .IN1(n9103), .IN2(n8665), .QN(n14823) );
  NAND2X0 U15405 ( .IN1(n253), .IN2(n9287), .QN(n14802) );
  NOR2X0 U15406 ( .IN1(n9226), .IN2(n9028), .QN(n253) );
  NAND2X0 U15407 ( .IN1(n9300), .IN2(CRC_OUT_8_27), .QN(n14801) );
  NAND4X0 U15408 ( .IN1(n14832), .IN2(n14833), .IN3(n14834), .IN4(n14835), 
        .QN(WX1943) );
  NAND2X0 U15409 ( .IN1(n14836), .IN2(n13901), .QN(n14835) );
  NAND2X0 U15410 ( .IN1(n14837), .IN2(n13904), .QN(n13901) );
  NAND2X0 U15411 ( .IN1(n14838), .IN2(n14839), .QN(n14837) );
  NAND2X0 U15412 ( .IN1(n16325), .IN2(n9122), .QN(n14839) );
  NAND2X0 U15413 ( .IN1(TM1), .IN2(n8608), .QN(n14838) );
  NAND3X0 U15414 ( .IN1(n14840), .IN2(n14841), .IN3(n14842), .QN(n14836) );
  NAND2X0 U15415 ( .IN1(n9328), .IN2(n13904), .QN(n14842) );
  NAND2X0 U15416 ( .IN1(n14843), .IN2(n14844), .QN(n13904) );
  NAND2X0 U15417 ( .IN1(n7820), .IN2(n14845), .QN(n14844) );
  INVX0 U15418 ( .INP(n14846), .ZN(n14843) );
  NOR2X0 U15419 ( .IN1(n14845), .IN2(n7820), .QN(n14846) );
  NOR2X0 U15420 ( .IN1(n14847), .IN2(n14848), .QN(n14845) );
  NOR2X0 U15421 ( .IN1(WX3429), .IN2(n7821), .QN(n14848) );
  INVX0 U15422 ( .INP(n14849), .ZN(n14847) );
  NAND2X0 U15423 ( .IN1(n7821), .IN2(WX3429), .QN(n14849) );
  NAND2X0 U15424 ( .IN1(n10068), .IN2(n8608), .QN(n14841) );
  NAND2X0 U15425 ( .IN1(n16325), .IN2(n10069), .QN(n14840) );
  NAND2X0 U15426 ( .IN1(n11890), .IN2(n9111), .QN(n14834) );
  NOR2X0 U15427 ( .IN1(n14850), .IN2(n14851), .QN(n11890) );
  INVX0 U15428 ( .INP(n14852), .ZN(n14851) );
  NAND2X0 U15429 ( .IN1(n14853), .IN2(n14854), .QN(n14852) );
  NOR2X0 U15430 ( .IN1(n14854), .IN2(n14853), .QN(n14850) );
  NAND2X0 U15431 ( .IN1(n14855), .IN2(n14856), .QN(n14853) );
  NAND2X0 U15432 ( .IN1(n14857), .IN2(WX2072), .QN(n14856) );
  NAND2X0 U15433 ( .IN1(n14858), .IN2(n14859), .QN(n14857) );
  NAND3X0 U15434 ( .IN1(n14858), .IN2(n14859), .IN3(n7849), .QN(n14855) );
  NAND2X0 U15435 ( .IN1(test_so18), .IN2(WX2008), .QN(n14859) );
  NAND2X0 U15436 ( .IN1(n7848), .IN2(n8803), .QN(n14858) );
  NOR2X0 U15437 ( .IN1(n14860), .IN2(n14861), .QN(n14854) );
  INVX0 U15438 ( .INP(n14862), .ZN(n14861) );
  NAND2X0 U15439 ( .IN1(n16310), .IN2(n9123), .QN(n14862) );
  NOR2X0 U15440 ( .IN1(n9118), .IN2(n16310), .QN(n14860) );
  NAND2X0 U15441 ( .IN1(n252), .IN2(n9287), .QN(n14833) );
  NOR2X0 U15442 ( .IN1(n9226), .IN2(n9029), .QN(n252) );
  NAND2X0 U15443 ( .IN1(n9300), .IN2(CRC_OUT_8_28), .QN(n14832) );
  NAND4X0 U15444 ( .IN1(n14863), .IN2(n14864), .IN3(n14865), .IN4(n14866), 
        .QN(WX1941) );
  NAND2X0 U15445 ( .IN1(n14867), .IN2(n13937), .QN(n14866) );
  NAND2X0 U15446 ( .IN1(n14868), .IN2(n13940), .QN(n13937) );
  NAND2X0 U15447 ( .IN1(n14869), .IN2(n14870), .QN(n14868) );
  NAND2X0 U15448 ( .IN1(n16324), .IN2(n9123), .QN(n14870) );
  NAND2X0 U15449 ( .IN1(TM1), .IN2(n8609), .QN(n14869) );
  NAND3X0 U15450 ( .IN1(n14871), .IN2(n14872), .IN3(n14873), .QN(n14867) );
  NAND2X0 U15451 ( .IN1(n9328), .IN2(n13940), .QN(n14873) );
  NAND2X0 U15452 ( .IN1(n14874), .IN2(n14875), .QN(n13940) );
  NAND2X0 U15453 ( .IN1(n7822), .IN2(n14876), .QN(n14875) );
  INVX0 U15454 ( .INP(n14877), .ZN(n14874) );
  NOR2X0 U15455 ( .IN1(n14876), .IN2(n7822), .QN(n14877) );
  NOR2X0 U15456 ( .IN1(n14878), .IN2(n14879), .QN(n14876) );
  NOR2X0 U15457 ( .IN1(WX3427), .IN2(n7823), .QN(n14879) );
  INVX0 U15458 ( .INP(n14880), .ZN(n14878) );
  NAND2X0 U15459 ( .IN1(n7823), .IN2(WX3427), .QN(n14880) );
  NAND2X0 U15460 ( .IN1(n9084), .IN2(n8609), .QN(n14872) );
  NAND2X0 U15461 ( .IN1(n16324), .IN2(n9080), .QN(n14871) );
  NAND2X0 U15462 ( .IN1(n14881), .IN2(n11919), .QN(n14865) );
  NAND2X0 U15463 ( .IN1(n14882), .IN2(n11923), .QN(n11919) );
  NAND2X0 U15464 ( .IN1(n14883), .IN2(n14884), .QN(n14882) );
  NAND2X0 U15465 ( .IN1(n16309), .IN2(n9123), .QN(n14884) );
  NAND2X0 U15466 ( .IN1(TM1), .IN2(n8667), .QN(n14883) );
  NAND2X0 U15467 ( .IN1(n14885), .IN2(n14886), .QN(n14881) );
  NAND2X0 U15468 ( .IN1(n9103), .IN2(n11923), .QN(n14886) );
  NAND2X0 U15469 ( .IN1(n14887), .IN2(n14888), .QN(n11923) );
  NAND2X0 U15470 ( .IN1(n7850), .IN2(n14889), .QN(n14888) );
  INVX0 U15471 ( .INP(n14890), .ZN(n14887) );
  NOR2X0 U15472 ( .IN1(n14889), .IN2(n7850), .QN(n14890) );
  NOR2X0 U15473 ( .IN1(n14891), .IN2(n14892), .QN(n14889) );
  NOR2X0 U15474 ( .IN1(WX2134), .IN2(n7851), .QN(n14892) );
  INVX0 U15475 ( .INP(n14893), .ZN(n14891) );
  NAND2X0 U15476 ( .IN1(n7851), .IN2(WX2134), .QN(n14893) );
  NAND2X0 U15477 ( .IN1(n9103), .IN2(n8667), .QN(n14885) );
  NAND2X0 U15478 ( .IN1(n251), .IN2(n9287), .QN(n14864) );
  NOR2X0 U15479 ( .IN1(n9226), .IN2(n9030), .QN(n251) );
  NAND2X0 U15480 ( .IN1(n9300), .IN2(CRC_OUT_8_29), .QN(n14863) );
  NAND4X0 U15481 ( .IN1(n14894), .IN2(n14895), .IN3(n14896), .IN4(n14897), 
        .QN(WX1939) );
  NAND2X0 U15482 ( .IN1(n14898), .IN2(n11955), .QN(n14897) );
  NAND2X0 U15483 ( .IN1(n14899), .IN2(n11959), .QN(n11955) );
  NAND2X0 U15484 ( .IN1(n14900), .IN2(n14901), .QN(n14899) );
  NAND2X0 U15485 ( .IN1(n16308), .IN2(n9123), .QN(n14901) );
  NAND2X0 U15486 ( .IN1(TM1), .IN2(n8668), .QN(n14900) );
  NAND2X0 U15487 ( .IN1(n14902), .IN2(n14903), .QN(n14898) );
  NAND2X0 U15488 ( .IN1(n9103), .IN2(n11959), .QN(n14903) );
  NAND2X0 U15489 ( .IN1(n14904), .IN2(n14905), .QN(n11959) );
  NAND2X0 U15490 ( .IN1(n7852), .IN2(n14906), .QN(n14905) );
  INVX0 U15491 ( .INP(n14907), .ZN(n14904) );
  NOR2X0 U15492 ( .IN1(n14906), .IN2(n7852), .QN(n14907) );
  NOR2X0 U15493 ( .IN1(n14908), .IN2(n14909), .QN(n14906) );
  NOR2X0 U15494 ( .IN1(WX2132), .IN2(n7853), .QN(n14909) );
  INVX0 U15495 ( .INP(n14910), .ZN(n14908) );
  NAND2X0 U15496 ( .IN1(n7853), .IN2(WX2132), .QN(n14910) );
  NAND2X0 U15497 ( .IN1(n9103), .IN2(n8668), .QN(n14902) );
  NAND2X0 U15498 ( .IN1(n13960), .IN2(n9336), .QN(n14896) );
  NOR2X0 U15499 ( .IN1(n14911), .IN2(n14912), .QN(n13960) );
  INVX0 U15500 ( .INP(n14913), .ZN(n14912) );
  NAND2X0 U15501 ( .IN1(n14914), .IN2(n14915), .QN(n14913) );
  NOR2X0 U15502 ( .IN1(n14915), .IN2(n14914), .QN(n14911) );
  NAND2X0 U15503 ( .IN1(n14916), .IN2(n14917), .QN(n14914) );
  NAND2X0 U15504 ( .IN1(n8472), .IN2(n14918), .QN(n14917) );
  INVX0 U15505 ( .INP(n14919), .ZN(n14918) );
  NAND2X0 U15506 ( .IN1(n14919), .IN2(WX3425), .QN(n14916) );
  NAND2X0 U15507 ( .IN1(n14920), .IN2(n14921), .QN(n14919) );
  INVX0 U15508 ( .INP(n14922), .ZN(n14921) );
  NOR2X0 U15509 ( .IN1(n8817), .IN2(n16323), .QN(n14922) );
  NAND2X0 U15510 ( .IN1(n16323), .IN2(n8817), .QN(n14920) );
  NOR2X0 U15511 ( .IN1(n14923), .IN2(n14924), .QN(n14915) );
  INVX0 U15512 ( .INP(n14925), .ZN(n14924) );
  NAND2X0 U15513 ( .IN1(n7824), .IN2(n9123), .QN(n14925) );
  NOR2X0 U15514 ( .IN1(n9117), .IN2(n7824), .QN(n14923) );
  NAND2X0 U15515 ( .IN1(n250), .IN2(n9287), .QN(n14895) );
  NOR2X0 U15516 ( .IN1(n9226), .IN2(n9031), .QN(n250) );
  NAND2X0 U15517 ( .IN1(n9300), .IN2(CRC_OUT_8_30), .QN(n14894) );
  NAND4X0 U15518 ( .IN1(n14926), .IN2(n14927), .IN3(n14928), .IN4(n14929), 
        .QN(WX1937) );
  NAND2X0 U15519 ( .IN1(n14930), .IN2(n11996), .QN(n14929) );
  NAND2X0 U15520 ( .IN1(n14931), .IN2(n12000), .QN(n11996) );
  NAND2X0 U15521 ( .IN1(n14932), .IN2(n14933), .QN(n14931) );
  NAND2X0 U15522 ( .IN1(n16307), .IN2(n9123), .QN(n14933) );
  NAND2X0 U15523 ( .IN1(TM1), .IN2(n8669), .QN(n14932) );
  NAND2X0 U15524 ( .IN1(n14934), .IN2(n14935), .QN(n14930) );
  NAND2X0 U15525 ( .IN1(n9103), .IN2(n12000), .QN(n14935) );
  NAND2X0 U15526 ( .IN1(n14936), .IN2(n14937), .QN(n12000) );
  NAND2X0 U15527 ( .IN1(n7626), .IN2(n14938), .QN(n14937) );
  INVX0 U15528 ( .INP(n14939), .ZN(n14936) );
  NOR2X0 U15529 ( .IN1(n14938), .IN2(n7626), .QN(n14939) );
  NOR2X0 U15530 ( .IN1(n14940), .IN2(n14941), .QN(n14938) );
  NOR2X0 U15531 ( .IN1(WX2130), .IN2(n7627), .QN(n14941) );
  INVX0 U15532 ( .INP(n14942), .ZN(n14940) );
  NAND2X0 U15533 ( .IN1(n7627), .IN2(WX2130), .QN(n14942) );
  NAND2X0 U15534 ( .IN1(n9103), .IN2(n8669), .QN(n14934) );
  NAND2X0 U15535 ( .IN1(n14943), .IN2(n13980), .QN(n14928) );
  NAND2X0 U15536 ( .IN1(n14944), .IN2(n13983), .QN(n13980) );
  NAND2X0 U15537 ( .IN1(n14945), .IN2(n14946), .QN(n14944) );
  NAND2X0 U15538 ( .IN1(n16322), .IN2(n9123), .QN(n14946) );
  NAND2X0 U15539 ( .IN1(TM1), .IN2(n8611), .QN(n14945) );
  NAND3X0 U15540 ( .IN1(n14947), .IN2(n14948), .IN3(n14949), .QN(n14943) );
  NAND2X0 U15541 ( .IN1(n9328), .IN2(n13983), .QN(n14949) );
  NAND2X0 U15542 ( .IN1(n14950), .IN2(n14951), .QN(n13983) );
  NAND2X0 U15543 ( .IN1(n7624), .IN2(n14952), .QN(n14951) );
  INVX0 U15544 ( .INP(n14953), .ZN(n14950) );
  NOR2X0 U15545 ( .IN1(n14952), .IN2(n7624), .QN(n14953) );
  NOR2X0 U15546 ( .IN1(n14954), .IN2(n14955), .QN(n14952) );
  NOR2X0 U15547 ( .IN1(WX3423), .IN2(n7625), .QN(n14955) );
  INVX0 U15548 ( .INP(n14956), .ZN(n14954) );
  NAND2X0 U15549 ( .IN1(n7625), .IN2(WX3423), .QN(n14956) );
  NAND2X0 U15550 ( .IN1(n9083), .IN2(n8611), .QN(n14948) );
  NOR2X0 U15551 ( .IN1(n9337), .IN2(n9116), .QN(n10068) );
  NAND2X0 U15552 ( .IN1(n16322), .IN2(n9079), .QN(n14947) );
  NOR2X0 U15553 ( .IN1(n9337), .IN2(TM1), .QN(n10069) );
  NAND2X0 U15554 ( .IN1(n9301), .IN2(CRC_OUT_8_31), .QN(n14927) );
  NAND2X0 U15555 ( .IN1(n2245), .IN2(WX1778), .QN(n14926) );
  NOR2X0 U15556 ( .IN1(n9226), .IN2(WX1778), .QN(WX1839) );
  NOR3X0 U15557 ( .IN1(n9151), .IN2(n14957), .IN3(n14958), .QN(WX1326) );
  NOR2X0 U15558 ( .IN1(n8775), .IN2(CRC_OUT_9_30), .QN(n14958) );
  NOR2X0 U15559 ( .IN1(DFF_190_n1), .IN2(WX837), .QN(n14957) );
  NOR3X0 U15560 ( .IN1(n9151), .IN2(n14959), .IN3(n14960), .QN(WX1324) );
  NOR2X0 U15561 ( .IN1(n8697), .IN2(CRC_OUT_9_29), .QN(n14960) );
  NOR2X0 U15562 ( .IN1(DFF_189_n1), .IN2(WX839), .QN(n14959) );
  NOR3X0 U15563 ( .IN1(n9151), .IN2(n14961), .IN3(n14962), .QN(WX1322) );
  NOR2X0 U15564 ( .IN1(n8709), .IN2(CRC_OUT_9_28), .QN(n14962) );
  NOR2X0 U15565 ( .IN1(DFF_188_n1), .IN2(WX841), .QN(n14961) );
  NOR3X0 U15566 ( .IN1(n9151), .IN2(n14963), .IN3(n14964), .QN(WX1320) );
  NOR2X0 U15567 ( .IN1(n8718), .IN2(CRC_OUT_9_27), .QN(n14964) );
  NOR2X0 U15568 ( .IN1(DFF_187_n1), .IN2(WX843), .QN(n14963) );
  NOR3X0 U15569 ( .IN1(n9151), .IN2(n14965), .IN3(n14966), .QN(WX1318) );
  NOR2X0 U15570 ( .IN1(n8724), .IN2(CRC_OUT_9_26), .QN(n14966) );
  NOR2X0 U15571 ( .IN1(DFF_186_n1), .IN2(WX845), .QN(n14965) );
  NOR3X0 U15572 ( .IN1(n9151), .IN2(n14967), .IN3(n14968), .QN(WX1316) );
  NOR2X0 U15573 ( .IN1(n8727), .IN2(CRC_OUT_9_25), .QN(n14968) );
  NOR2X0 U15574 ( .IN1(DFF_185_n1), .IN2(WX847), .QN(n14967) );
  NOR3X0 U15575 ( .IN1(n9151), .IN2(n14969), .IN3(n14970), .QN(WX1314) );
  NOR2X0 U15576 ( .IN1(n8736), .IN2(CRC_OUT_9_24), .QN(n14970) );
  NOR2X0 U15577 ( .IN1(DFF_184_n1), .IN2(WX849), .QN(n14969) );
  NOR3X0 U15578 ( .IN1(n9151), .IN2(n14971), .IN3(n14972), .QN(WX1312) );
  NOR2X0 U15579 ( .IN1(n8745), .IN2(CRC_OUT_9_23), .QN(n14972) );
  NOR2X0 U15580 ( .IN1(DFF_183_n1), .IN2(WX851), .QN(n14971) );
  NOR3X0 U15581 ( .IN1(n9151), .IN2(n14973), .IN3(n14974), .QN(WX1310) );
  NOR2X0 U15582 ( .IN1(n8747), .IN2(CRC_OUT_9_22), .QN(n14974) );
  NOR2X0 U15583 ( .IN1(DFF_182_n1), .IN2(WX853), .QN(n14973) );
  NOR3X0 U15584 ( .IN1(n9151), .IN2(n14975), .IN3(n14976), .QN(WX1308) );
  NOR2X0 U15585 ( .IN1(n8762), .IN2(CRC_OUT_9_21), .QN(n14976) );
  NOR2X0 U15586 ( .IN1(DFF_181_n1), .IN2(WX855), .QN(n14975) );
  NOR3X0 U15587 ( .IN1(n9151), .IN2(n14977), .IN3(n14978), .QN(WX1306) );
  NOR2X0 U15588 ( .IN1(n8768), .IN2(CRC_OUT_9_20), .QN(n14978) );
  NOR2X0 U15589 ( .IN1(DFF_180_n1), .IN2(WX857), .QN(n14977) );
  NOR2X0 U15590 ( .IN1(n9226), .IN2(n14979), .QN(WX1304) );
  NOR2X0 U15591 ( .IN1(n14980), .IN2(n14981), .QN(n14979) );
  NOR2X0 U15592 ( .IN1(test_so10), .IN2(WX859), .QN(n14981) );
  INVX0 U15593 ( .INP(n14982), .ZN(n14980) );
  NAND2X0 U15594 ( .IN1(WX859), .IN2(test_so10), .QN(n14982) );
  NOR3X0 U15595 ( .IN1(n9151), .IN2(n14983), .IN3(n14984), .QN(WX1302) );
  NOR2X0 U15596 ( .IN1(n8706), .IN2(CRC_OUT_9_18), .QN(n14984) );
  NOR2X0 U15597 ( .IN1(DFF_178_n1), .IN2(WX861), .QN(n14983) );
  NOR3X0 U15598 ( .IN1(n9150), .IN2(n14985), .IN3(n14986), .QN(WX1300) );
  NOR2X0 U15599 ( .IN1(n8721), .IN2(CRC_OUT_9_17), .QN(n14986) );
  NOR2X0 U15600 ( .IN1(DFF_177_n1), .IN2(WX863), .QN(n14985) );
  NOR3X0 U15601 ( .IN1(n9150), .IN2(n14987), .IN3(n14988), .QN(WX1298) );
  NOR2X0 U15602 ( .IN1(n8733), .IN2(CRC_OUT_9_16), .QN(n14988) );
  NOR2X0 U15603 ( .IN1(DFF_176_n1), .IN2(WX865), .QN(n14987) );
  NOR3X0 U15604 ( .IN1(n9150), .IN2(n14989), .IN3(n14990), .QN(WX1296) );
  INVX0 U15605 ( .INP(n14991), .ZN(n14990) );
  NAND2X0 U15606 ( .IN1(CRC_OUT_9_15), .IN2(n14992), .QN(n14991) );
  NOR2X0 U15607 ( .IN1(n14992), .IN2(CRC_OUT_9_15), .QN(n14989) );
  NAND2X0 U15608 ( .IN1(n14993), .IN2(n14994), .QN(n14992) );
  NAND2X0 U15609 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .QN(n14994) );
  NAND2X0 U15610 ( .IN1(DFF_191_n1), .IN2(n8798), .QN(n14993) );
  NOR3X0 U15611 ( .IN1(n9150), .IN2(n14995), .IN3(n14996), .QN(WX1294) );
  NOR2X0 U15612 ( .IN1(n8765), .IN2(CRC_OUT_9_14), .QN(n14996) );
  NOR2X0 U15613 ( .IN1(DFF_174_n1), .IN2(WX869), .QN(n14995) );
  NOR3X0 U15614 ( .IN1(n9150), .IN2(n14997), .IN3(n14998), .QN(WX1292) );
  NOR2X0 U15615 ( .IN1(n8777), .IN2(CRC_OUT_9_13), .QN(n14998) );
  NOR2X0 U15616 ( .IN1(DFF_173_n1), .IN2(WX871), .QN(n14997) );
  NOR3X0 U15617 ( .IN1(n9150), .IN2(n14999), .IN3(n15000), .QN(WX1290) );
  NOR2X0 U15618 ( .IN1(n8712), .IN2(CRC_OUT_9_12), .QN(n15000) );
  NOR2X0 U15619 ( .IN1(DFF_172_n1), .IN2(WX873), .QN(n14999) );
  NOR3X0 U15620 ( .IN1(n9150), .IN2(n15001), .IN3(n15002), .QN(WX1288) );
  NOR2X0 U15621 ( .IN1(n8739), .IN2(CRC_OUT_9_11), .QN(n15002) );
  NOR2X0 U15622 ( .IN1(DFF_171_n1), .IN2(WX875), .QN(n15001) );
  NOR2X0 U15623 ( .IN1(n9225), .IN2(n15003), .QN(WX1286) );
  NOR2X0 U15624 ( .IN1(n15004), .IN2(n15005), .QN(n15003) );
  INVX0 U15625 ( .INP(n15006), .ZN(n15005) );
  NAND2X0 U15626 ( .IN1(CRC_OUT_9_10), .IN2(n15007), .QN(n15006) );
  NOR2X0 U15627 ( .IN1(n15007), .IN2(CRC_OUT_9_10), .QN(n15004) );
  NAND2X0 U15628 ( .IN1(n15008), .IN2(n15009), .QN(n15007) );
  NAND2X0 U15629 ( .IN1(n8785), .IN2(CRC_OUT_9_31), .QN(n15009) );
  NAND2X0 U15630 ( .IN1(DFF_191_n1), .IN2(WX877), .QN(n15008) );
  NOR3X0 U15631 ( .IN1(n9150), .IN2(n15010), .IN3(n15011), .QN(WX1284) );
  NOR2X0 U15632 ( .IN1(n8730), .IN2(CRC_OUT_9_9), .QN(n15011) );
  NOR2X0 U15633 ( .IN1(DFF_169_n1), .IN2(WX879), .QN(n15010) );
  NOR3X0 U15634 ( .IN1(n9150), .IN2(n15012), .IN3(n15013), .QN(WX1282) );
  NOR2X0 U15635 ( .IN1(n8743), .IN2(CRC_OUT_9_8), .QN(n15013) );
  NOR2X0 U15636 ( .IN1(DFF_168_n1), .IN2(WX881), .QN(n15012) );
  NOR3X0 U15637 ( .IN1(n9150), .IN2(n15014), .IN3(n15015), .QN(WX1280) );
  NOR2X0 U15638 ( .IN1(n8752), .IN2(CRC_OUT_9_7), .QN(n15015) );
  NOR2X0 U15639 ( .IN1(DFF_167_n1), .IN2(WX883), .QN(n15014) );
  NOR3X0 U15640 ( .IN1(n9150), .IN2(n15016), .IN3(n15017), .QN(WX1278) );
  NOR2X0 U15641 ( .IN1(n8783), .IN2(CRC_OUT_9_6), .QN(n15017) );
  NOR2X0 U15642 ( .IN1(DFF_166_n1), .IN2(WX885), .QN(n15016) );
  NOR3X0 U15643 ( .IN1(n9150), .IN2(n15018), .IN3(n15019), .QN(WX1276) );
  NOR2X0 U15644 ( .IN1(n8770), .IN2(CRC_OUT_9_5), .QN(n15019) );
  NOR2X0 U15645 ( .IN1(DFF_165_n1), .IN2(WX887), .QN(n15018) );
  NOR3X0 U15646 ( .IN1(n9149), .IN2(n15020), .IN3(n15021), .QN(WX1274) );
  NOR2X0 U15647 ( .IN1(n8755), .IN2(CRC_OUT_9_4), .QN(n15021) );
  NOR2X0 U15648 ( .IN1(DFF_164_n1), .IN2(WX889), .QN(n15020) );
  NOR2X0 U15649 ( .IN1(n9225), .IN2(n15022), .QN(WX1272) );
  NOR2X0 U15650 ( .IN1(n15023), .IN2(n15024), .QN(n15022) );
  INVX0 U15651 ( .INP(n15025), .ZN(n15024) );
  NAND2X0 U15652 ( .IN1(CRC_OUT_9_3), .IN2(n15026), .QN(n15025) );
  NOR2X0 U15653 ( .IN1(n15026), .IN2(CRC_OUT_9_3), .QN(n15023) );
  NAND2X0 U15654 ( .IN1(n15027), .IN2(n15028), .QN(n15026) );
  NAND2X0 U15655 ( .IN1(n8758), .IN2(CRC_OUT_9_31), .QN(n15028) );
  NAND2X0 U15656 ( .IN1(DFF_191_n1), .IN2(WX891), .QN(n15027) );
  NOR3X0 U15657 ( .IN1(n9149), .IN2(n15029), .IN3(n15030), .QN(WX1270) );
  NOR2X0 U15658 ( .IN1(n8703), .IN2(CRC_OUT_9_2), .QN(n15030) );
  NOR2X0 U15659 ( .IN1(DFF_162_n1), .IN2(WX893), .QN(n15029) );
  NOR2X0 U15660 ( .IN1(n9225), .IN2(n15031), .QN(WX1268) );
  NOR2X0 U15661 ( .IN1(n15032), .IN2(n15033), .QN(n15031) );
  NOR2X0 U15662 ( .IN1(test_so9), .IN2(WX895), .QN(n15033) );
  INVX0 U15663 ( .INP(n15034), .ZN(n15032) );
  NAND2X0 U15664 ( .IN1(WX895), .IN2(test_so9), .QN(n15034) );
  NOR3X0 U15665 ( .IN1(n9149), .IN2(n15035), .IN3(n15036), .QN(WX1266) );
  NOR2X0 U15666 ( .IN1(n8714), .IN2(CRC_OUT_9_0), .QN(n15036) );
  NOR2X0 U15667 ( .IN1(DFF_160_n1), .IN2(WX897), .QN(n15035) );
  NOR3X0 U15668 ( .IN1(n9149), .IN2(n15037), .IN3(n15038), .QN(WX1264) );
  NOR2X0 U15669 ( .IN1(n8789), .IN2(CRC_OUT_9_31), .QN(n15038) );
  NOR2X0 U15670 ( .IN1(DFF_191_n1), .IN2(WX899), .QN(n15037) );
  NOR3X0 U15671 ( .IN1(n9147), .IN2(n15039), .IN3(n15040), .QN(WX11670) );
  NOR2X0 U15672 ( .IN1(n8134), .IN2(CRC_OUT_1_30), .QN(n15040) );
  NOR2X0 U15673 ( .IN1(DFF_1726_n1), .IN2(WX11181), .QN(n15039) );
  NOR3X0 U15674 ( .IN1(n9149), .IN2(n15041), .IN3(n15042), .QN(WX11668) );
  NOR2X0 U15675 ( .IN1(n8135), .IN2(CRC_OUT_1_29), .QN(n15042) );
  NOR2X0 U15676 ( .IN1(DFF_1725_n1), .IN2(WX11183), .QN(n15041) );
  NOR3X0 U15677 ( .IN1(n9149), .IN2(n15043), .IN3(n15044), .QN(WX11666) );
  NOR2X0 U15678 ( .IN1(n8136), .IN2(CRC_OUT_1_28), .QN(n15044) );
  NOR2X0 U15679 ( .IN1(DFF_1724_n1), .IN2(WX11185), .QN(n15043) );
  NOR3X0 U15680 ( .IN1(n9149), .IN2(n15045), .IN3(n15046), .QN(WX11664) );
  NOR2X0 U15681 ( .IN1(n8137), .IN2(CRC_OUT_1_27), .QN(n15046) );
  NOR2X0 U15682 ( .IN1(DFF_1723_n1), .IN2(WX11187), .QN(n15045) );
  NOR3X0 U15683 ( .IN1(n9149), .IN2(n15047), .IN3(n15048), .QN(WX11662) );
  NOR2X0 U15684 ( .IN1(n8138), .IN2(CRC_OUT_1_26), .QN(n15048) );
  NOR2X0 U15685 ( .IN1(DFF_1722_n1), .IN2(WX11189), .QN(n15047) );
  NOR3X0 U15686 ( .IN1(n9149), .IN2(n15049), .IN3(n15050), .QN(WX11660) );
  NOR2X0 U15687 ( .IN1(n8139), .IN2(CRC_OUT_1_25), .QN(n15050) );
  NOR2X0 U15688 ( .IN1(DFF_1721_n1), .IN2(WX11191), .QN(n15049) );
  NOR3X0 U15689 ( .IN1(n9149), .IN2(n15051), .IN3(n15052), .QN(WX11658) );
  NOR2X0 U15690 ( .IN1(n8140), .IN2(CRC_OUT_1_24), .QN(n15052) );
  NOR2X0 U15691 ( .IN1(DFF_1720_n1), .IN2(WX11193), .QN(n15051) );
  NOR3X0 U15692 ( .IN1(n9149), .IN2(n15053), .IN3(n15054), .QN(WX11656) );
  NOR2X0 U15693 ( .IN1(n8141), .IN2(CRC_OUT_1_23), .QN(n15054) );
  NOR2X0 U15694 ( .IN1(DFF_1719_n1), .IN2(WX11195), .QN(n15053) );
  NOR3X0 U15695 ( .IN1(n9149), .IN2(n15055), .IN3(n15056), .QN(WX11654) );
  NOR2X0 U15696 ( .IN1(n8142), .IN2(CRC_OUT_1_22), .QN(n15056) );
  NOR2X0 U15697 ( .IN1(DFF_1718_n1), .IN2(WX11197), .QN(n15055) );
  NOR3X0 U15698 ( .IN1(n9148), .IN2(n15057), .IN3(n15058), .QN(WX11652) );
  NOR2X0 U15699 ( .IN1(n8143), .IN2(CRC_OUT_1_21), .QN(n15058) );
  NOR2X0 U15700 ( .IN1(DFF_1717_n1), .IN2(WX11199), .QN(n15057) );
  NOR3X0 U15701 ( .IN1(n9148), .IN2(n15059), .IN3(n15060), .QN(WX11650) );
  NOR2X0 U15702 ( .IN1(n8144), .IN2(CRC_OUT_1_20), .QN(n15060) );
  NOR2X0 U15703 ( .IN1(DFF_1716_n1), .IN2(WX11201), .QN(n15059) );
  NOR3X0 U15704 ( .IN1(n9148), .IN2(n15061), .IN3(n15062), .QN(WX11648) );
  NOR2X0 U15705 ( .IN1(n8145), .IN2(CRC_OUT_1_19), .QN(n15062) );
  NOR2X0 U15706 ( .IN1(DFF_1715_n1), .IN2(WX11203), .QN(n15061) );
  NOR2X0 U15707 ( .IN1(n9224), .IN2(n15063), .QN(WX11646) );
  NOR2X0 U15708 ( .IN1(n15064), .IN2(n15065), .QN(n15063) );
  NOR2X0 U15709 ( .IN1(test_so97), .IN2(CRC_OUT_1_18), .QN(n15065) );
  NOR2X0 U15710 ( .IN1(DFF_1714_n1), .IN2(n8804), .QN(n15064) );
  NOR3X0 U15711 ( .IN1(n9148), .IN2(n15066), .IN3(n15067), .QN(WX11644) );
  NOR2X0 U15712 ( .IN1(n8146), .IN2(CRC_OUT_1_17), .QN(n15067) );
  NOR2X0 U15713 ( .IN1(DFF_1713_n1), .IN2(WX11207), .QN(n15066) );
  NOR3X0 U15714 ( .IN1(n9148), .IN2(n15068), .IN3(n15069), .QN(WX11642) );
  NOR2X0 U15715 ( .IN1(n8147), .IN2(CRC_OUT_1_16), .QN(n15069) );
  NOR2X0 U15716 ( .IN1(DFF_1712_n1), .IN2(WX11209), .QN(n15068) );
  NOR3X0 U15717 ( .IN1(n9148), .IN2(n15070), .IN3(n15071), .QN(WX11640) );
  INVX0 U15718 ( .INP(n15072), .ZN(n15071) );
  NAND2X0 U15719 ( .IN1(CRC_OUT_1_15), .IN2(n15073), .QN(n15072) );
  NOR2X0 U15720 ( .IN1(n15073), .IN2(CRC_OUT_1_15), .QN(n15070) );
  NAND2X0 U15721 ( .IN1(n15074), .IN2(n15075), .QN(n15073) );
  NAND2X0 U15722 ( .IN1(test_so100), .IN2(WX11211), .QN(n15075) );
  NAND2X0 U15723 ( .IN1(n8105), .IN2(n8790), .QN(n15074) );
  NOR2X0 U15724 ( .IN1(n9227), .IN2(n15076), .QN(WX11638) );
  NOR2X0 U15725 ( .IN1(n15077), .IN2(n15078), .QN(n15076) );
  NOR2X0 U15726 ( .IN1(test_so99), .IN2(WX11213), .QN(n15078) );
  INVX0 U15727 ( .INP(n15079), .ZN(n15077) );
  NAND2X0 U15728 ( .IN1(WX11213), .IN2(test_so99), .QN(n15079) );
  NOR3X0 U15729 ( .IN1(n9148), .IN2(n15080), .IN3(n15081), .QN(WX11636) );
  NOR2X0 U15730 ( .IN1(n8149), .IN2(CRC_OUT_1_13), .QN(n15081) );
  NOR2X0 U15731 ( .IN1(DFF_1709_n1), .IN2(WX11215), .QN(n15080) );
  NOR3X0 U15732 ( .IN1(n9148), .IN2(n15082), .IN3(n15083), .QN(WX11634) );
  NOR2X0 U15733 ( .IN1(n8150), .IN2(CRC_OUT_1_12), .QN(n15083) );
  NOR2X0 U15734 ( .IN1(DFF_1708_n1), .IN2(WX11217), .QN(n15082) );
  NOR3X0 U15735 ( .IN1(n9148), .IN2(n15084), .IN3(n15085), .QN(WX11632) );
  NOR2X0 U15736 ( .IN1(n8151), .IN2(CRC_OUT_1_11), .QN(n15085) );
  NOR2X0 U15737 ( .IN1(DFF_1707_n1), .IN2(WX11219), .QN(n15084) );
  NOR3X0 U15738 ( .IN1(n9148), .IN2(n15086), .IN3(n15087), .QN(WX11630) );
  INVX0 U15739 ( .INP(n15088), .ZN(n15087) );
  NAND2X0 U15740 ( .IN1(CRC_OUT_1_10), .IN2(n15089), .QN(n15088) );
  NOR2X0 U15741 ( .IN1(n15089), .IN2(CRC_OUT_1_10), .QN(n15086) );
  NAND2X0 U15742 ( .IN1(n15090), .IN2(n15091), .QN(n15089) );
  NAND2X0 U15743 ( .IN1(test_so100), .IN2(WX11221), .QN(n15091) );
  NAND2X0 U15744 ( .IN1(n8106), .IN2(n8790), .QN(n15090) );
  NOR3X0 U15745 ( .IN1(n9147), .IN2(n15092), .IN3(n15093), .QN(WX11628) );
  NOR2X0 U15746 ( .IN1(n8152), .IN2(CRC_OUT_1_9), .QN(n15093) );
  NOR2X0 U15747 ( .IN1(DFF_1705_n1), .IN2(WX11223), .QN(n15092) );
  NOR3X0 U15748 ( .IN1(n9152), .IN2(n15094), .IN3(n15095), .QN(WX11626) );
  NOR2X0 U15749 ( .IN1(n8153), .IN2(CRC_OUT_1_8), .QN(n15095) );
  NOR2X0 U15750 ( .IN1(DFF_1704_n1), .IN2(WX11225), .QN(n15094) );
  NOR3X0 U15751 ( .IN1(n9147), .IN2(n15096), .IN3(n15097), .QN(WX11624) );
  NOR2X0 U15752 ( .IN1(n8154), .IN2(CRC_OUT_1_7), .QN(n15097) );
  NOR2X0 U15753 ( .IN1(DFF_1703_n1), .IN2(WX11227), .QN(n15096) );
  NOR3X0 U15754 ( .IN1(n9147), .IN2(n15098), .IN3(n15099), .QN(WX11622) );
  NOR2X0 U15755 ( .IN1(n8155), .IN2(CRC_OUT_1_6), .QN(n15099) );
  NOR2X0 U15756 ( .IN1(DFF_1702_n1), .IN2(WX11229), .QN(n15098) );
  NOR3X0 U15757 ( .IN1(n9147), .IN2(n15100), .IN3(n15101), .QN(WX11620) );
  NOR2X0 U15758 ( .IN1(n8156), .IN2(CRC_OUT_1_5), .QN(n15101) );
  NOR2X0 U15759 ( .IN1(DFF_1701_n1), .IN2(WX11231), .QN(n15100) );
  NOR3X0 U15760 ( .IN1(n9147), .IN2(n15102), .IN3(n15103), .QN(WX11618) );
  NOR2X0 U15761 ( .IN1(n8157), .IN2(CRC_OUT_1_4), .QN(n15103) );
  NOR2X0 U15762 ( .IN1(DFF_1700_n1), .IN2(WX11233), .QN(n15102) );
  NOR3X0 U15763 ( .IN1(n9147), .IN2(n15104), .IN3(n15105), .QN(WX11616) );
  INVX0 U15764 ( .INP(n15106), .ZN(n15105) );
  NAND2X0 U15765 ( .IN1(CRC_OUT_1_3), .IN2(n15107), .QN(n15106) );
  NOR2X0 U15766 ( .IN1(n15107), .IN2(CRC_OUT_1_3), .QN(n15104) );
  NAND2X0 U15767 ( .IN1(n15108), .IN2(n15109), .QN(n15107) );
  NAND2X0 U15768 ( .IN1(test_so100), .IN2(WX11235), .QN(n15109) );
  NAND2X0 U15769 ( .IN1(n8107), .IN2(n8790), .QN(n15108) );
  NOR3X0 U15770 ( .IN1(n9148), .IN2(n15110), .IN3(n15111), .QN(WX11614) );
  NOR2X0 U15771 ( .IN1(n8158), .IN2(CRC_OUT_1_2), .QN(n15111) );
  NOR2X0 U15772 ( .IN1(DFF_1698_n1), .IN2(WX11237), .QN(n15110) );
  NOR2X0 U15773 ( .IN1(n9227), .IN2(n15112), .QN(WX11612) );
  NOR2X0 U15774 ( .IN1(n15113), .IN2(n15114), .QN(n15112) );
  NOR2X0 U15775 ( .IN1(test_so98), .IN2(CRC_OUT_1_1), .QN(n15114) );
  NOR2X0 U15776 ( .IN1(DFF_1697_n1), .IN2(n8794), .QN(n15113) );
  NOR3X0 U15777 ( .IN1(n9148), .IN2(n15115), .IN3(n15116), .QN(WX11610) );
  NOR2X0 U15778 ( .IN1(n8159), .IN2(CRC_OUT_1_0), .QN(n15116) );
  NOR2X0 U15779 ( .IN1(DFF_1696_n1), .IN2(WX11241), .QN(n15115) );
  NOR2X0 U15780 ( .IN1(n9227), .IN2(n15117), .QN(WX11608) );
  NOR2X0 U15781 ( .IN1(n15118), .IN2(n15119), .QN(n15117) );
  NOR2X0 U15782 ( .IN1(test_so100), .IN2(WX11243), .QN(n15119) );
  NOR2X0 U15783 ( .IN1(n8126), .IN2(n8790), .QN(n15118) );
  NOR2X0 U15784 ( .IN1(n16427), .IN2(n9159), .QN(WX11082) );
  NOR2X0 U15785 ( .IN1(n16426), .IN2(n9158), .QN(WX11080) );
  NOR2X0 U15786 ( .IN1(n16425), .IN2(n9158), .QN(WX11078) );
  NOR2X0 U15787 ( .IN1(n16424), .IN2(n9158), .QN(WX11076) );
  NOR2X0 U15788 ( .IN1(n16423), .IN2(n9158), .QN(WX11074) );
  NOR2X0 U15789 ( .IN1(n16422), .IN2(n9158), .QN(WX11072) );
  NOR2X0 U15790 ( .IN1(n16421), .IN2(n9158), .QN(WX11070) );
  NOR2X0 U15791 ( .IN1(n16420), .IN2(n9158), .QN(WX11068) );
  NOR2X0 U15792 ( .IN1(n16419), .IN2(n9158), .QN(WX11066) );
  NOR2X0 U15793 ( .IN1(n9228), .IN2(n8826), .QN(WX11064) );
  NOR2X0 U15794 ( .IN1(n16418), .IN2(n9158), .QN(WX11062) );
  NOR2X0 U15795 ( .IN1(n16417), .IN2(n9157), .QN(WX11060) );
  NOR2X0 U15796 ( .IN1(n16416), .IN2(n9156), .QN(WX11058) );
  NOR2X0 U15797 ( .IN1(n16415), .IN2(n9156), .QN(WX11056) );
  NOR2X0 U15798 ( .IN1(n16414), .IN2(n9157), .QN(WX11054) );
  NOR2X0 U15799 ( .IN1(n16413), .IN2(n9156), .QN(WX11052) );
  NAND4X0 U15800 ( .IN1(n15120), .IN2(n15121), .IN3(n15122), .IN4(n15123), 
        .QN(WX11050) );
  NAND2X0 U15801 ( .IN1(n9103), .IN2(n9960), .QN(n15123) );
  NAND2X0 U15802 ( .IN1(n15124), .IN2(n15125), .QN(n9960) );
  INVX0 U15803 ( .INP(n15126), .ZN(n15125) );
  NOR2X0 U15804 ( .IN1(n15127), .IN2(n15128), .QN(n15126) );
  NAND2X0 U15805 ( .IN1(n15128), .IN2(n15127), .QN(n15124) );
  NOR2X0 U15806 ( .IN1(n15129), .IN2(n15130), .QN(n15127) );
  NOR2X0 U15807 ( .IN1(WX11243), .IN2(n7855), .QN(n15130) );
  INVX0 U15808 ( .INP(n15131), .ZN(n15129) );
  NAND2X0 U15809 ( .IN1(n7855), .IN2(WX11243), .QN(n15131) );
  NAND2X0 U15810 ( .IN1(n15132), .IN2(n15133), .QN(n15128) );
  NAND2X0 U15811 ( .IN1(n7854), .IN2(WX11115), .QN(n15133) );
  INVX0 U15812 ( .INP(n15134), .ZN(n15132) );
  NOR2X0 U15813 ( .IN1(WX11115), .IN2(n7854), .QN(n15134) );
  NAND2X0 U15814 ( .IN1(n1969), .IN2(n9287), .QN(n15122) );
  NOR2X0 U15815 ( .IN1(n9228), .IN2(n9032), .QN(n1969) );
  NAND2X0 U15816 ( .IN1(DATA_0_0), .IN2(n9336), .QN(n15121) );
  NAND2X0 U15817 ( .IN1(n9301), .IN2(CRC_OUT_1_0), .QN(n15120) );
  NAND4X0 U15818 ( .IN1(n15135), .IN2(n15136), .IN3(n15137), .IN4(n15138), 
        .QN(WX11048) );
  NAND2X0 U15819 ( .IN1(n9103), .IN2(n9967), .QN(n15138) );
  NAND2X0 U15820 ( .IN1(n15139), .IN2(n15140), .QN(n9967) );
  INVX0 U15821 ( .INP(n15141), .ZN(n15140) );
  NOR2X0 U15822 ( .IN1(n15142), .IN2(n15143), .QN(n15141) );
  NAND2X0 U15823 ( .IN1(n15143), .IN2(n15142), .QN(n15139) );
  NOR2X0 U15824 ( .IN1(n15144), .IN2(n15145), .QN(n15142) );
  NOR2X0 U15825 ( .IN1(WX11241), .IN2(n7857), .QN(n15145) );
  INVX0 U15826 ( .INP(n15146), .ZN(n15144) );
  NAND2X0 U15827 ( .IN1(n7857), .IN2(WX11241), .QN(n15146) );
  NAND2X0 U15828 ( .IN1(n15147), .IN2(n15148), .QN(n15143) );
  NAND2X0 U15829 ( .IN1(n7856), .IN2(WX11113), .QN(n15148) );
  INVX0 U15830 ( .INP(n15149), .ZN(n15147) );
  NOR2X0 U15831 ( .IN1(WX11113), .IN2(n7856), .QN(n15149) );
  NAND2X0 U15832 ( .IN1(n1968), .IN2(n9287), .QN(n15137) );
  NOR2X0 U15833 ( .IN1(n9228), .IN2(n9033), .QN(n1968) );
  NAND2X0 U15834 ( .IN1(DATA_0_1), .IN2(n9336), .QN(n15136) );
  NAND2X0 U15835 ( .IN1(n9301), .IN2(CRC_OUT_1_1), .QN(n15135) );
  NAND4X0 U15836 ( .IN1(n15150), .IN2(n15151), .IN3(n15152), .IN4(n15153), 
        .QN(WX11046) );
  NAND3X0 U15837 ( .IN1(n9972), .IN2(n9973), .IN3(n9092), .QN(n15153) );
  NAND3X0 U15838 ( .IN1(n15154), .IN2(n15155), .IN3(n15156), .QN(n9973) );
  INVX0 U15839 ( .INP(n15157), .ZN(n15156) );
  NAND2X0 U15840 ( .IN1(n15157), .IN2(n15158), .QN(n9972) );
  NAND2X0 U15841 ( .IN1(n15154), .IN2(n15155), .QN(n15158) );
  NAND2X0 U15842 ( .IN1(n7859), .IN2(WX11111), .QN(n15155) );
  NAND2X0 U15843 ( .IN1(n3535), .IN2(WX11175), .QN(n15154) );
  NOR2X0 U15844 ( .IN1(n15159), .IN2(n15160), .QN(n15157) );
  NOR2X0 U15845 ( .IN1(n8794), .IN2(n7858), .QN(n15160) );
  INVX0 U15846 ( .INP(n15161), .ZN(n15159) );
  NAND2X0 U15847 ( .IN1(n7858), .IN2(n8794), .QN(n15161) );
  NAND2X0 U15848 ( .IN1(n1967), .IN2(n9287), .QN(n15152) );
  NOR2X0 U15849 ( .IN1(n9228), .IN2(n9034), .QN(n1967) );
  NAND2X0 U15850 ( .IN1(DATA_0_2), .IN2(n9336), .QN(n15151) );
  NAND2X0 U15851 ( .IN1(n9301), .IN2(CRC_OUT_1_2), .QN(n15150) );
  NAND4X0 U15852 ( .IN1(n15162), .IN2(n15163), .IN3(n15164), .IN4(n15165), 
        .QN(WX11044) );
  NAND2X0 U15853 ( .IN1(n9103), .IN2(n9981), .QN(n15165) );
  NAND2X0 U15854 ( .IN1(n15166), .IN2(n15167), .QN(n9981) );
  INVX0 U15855 ( .INP(n15168), .ZN(n15167) );
  NOR2X0 U15856 ( .IN1(n15169), .IN2(n15170), .QN(n15168) );
  NAND2X0 U15857 ( .IN1(n15170), .IN2(n15169), .QN(n15166) );
  NOR2X0 U15858 ( .IN1(n15171), .IN2(n15172), .QN(n15169) );
  NOR2X0 U15859 ( .IN1(WX11237), .IN2(n7861), .QN(n15172) );
  INVX0 U15860 ( .INP(n15173), .ZN(n15171) );
  NAND2X0 U15861 ( .IN1(n7861), .IN2(WX11237), .QN(n15173) );
  NAND2X0 U15862 ( .IN1(n15174), .IN2(n15175), .QN(n15170) );
  NAND2X0 U15863 ( .IN1(n7860), .IN2(WX11109), .QN(n15175) );
  INVX0 U15864 ( .INP(n15176), .ZN(n15174) );
  NOR2X0 U15865 ( .IN1(WX11109), .IN2(n7860), .QN(n15176) );
  NAND2X0 U15866 ( .IN1(n1966), .IN2(n9287), .QN(n15164) );
  NOR2X0 U15867 ( .IN1(n9228), .IN2(n9035), .QN(n1966) );
  NAND2X0 U15868 ( .IN1(DATA_0_3), .IN2(n9336), .QN(n15163) );
  NAND2X0 U15869 ( .IN1(n9301), .IN2(CRC_OUT_1_3), .QN(n15162) );
  NAND4X0 U15870 ( .IN1(n15177), .IN2(n15178), .IN3(n15179), .IN4(n15180), 
        .QN(WX11042) );
  NAND3X0 U15871 ( .IN1(n9986), .IN2(n9987), .IN3(n9092), .QN(n15180) );
  NAND3X0 U15872 ( .IN1(n15181), .IN2(n15182), .IN3(n15183), .QN(n9987) );
  INVX0 U15873 ( .INP(n15184), .ZN(n15183) );
  NAND2X0 U15874 ( .IN1(n15184), .IN2(n15185), .QN(n9986) );
  NAND2X0 U15875 ( .IN1(n15181), .IN2(n15182), .QN(n15185) );
  NAND2X0 U15876 ( .IN1(n8107), .IN2(WX11107), .QN(n15182) );
  NAND2X0 U15877 ( .IN1(n3539), .IN2(WX11235), .QN(n15181) );
  NOR2X0 U15878 ( .IN1(n15186), .IN2(n15187), .QN(n15184) );
  INVX0 U15879 ( .INP(n15188), .ZN(n15187) );
  NAND2X0 U15880 ( .IN1(test_so96), .IN2(WX11043), .QN(n15188) );
  NOR2X0 U15881 ( .IN1(WX11043), .IN2(test_so96), .QN(n15186) );
  NAND2X0 U15882 ( .IN1(n1965), .IN2(n9287), .QN(n15179) );
  NOR2X0 U15883 ( .IN1(n9228), .IN2(n9036), .QN(n1965) );
  NAND2X0 U15884 ( .IN1(DATA_0_4), .IN2(n9336), .QN(n15178) );
  NAND2X0 U15885 ( .IN1(n9301), .IN2(CRC_OUT_1_4), .QN(n15177) );
  NAND4X0 U15886 ( .IN1(n15189), .IN2(n15190), .IN3(n15191), .IN4(n15192), 
        .QN(WX11040) );
  NAND2X0 U15887 ( .IN1(n9103), .IN2(n9994), .QN(n15192) );
  NAND2X0 U15888 ( .IN1(n15193), .IN2(n15194), .QN(n9994) );
  INVX0 U15889 ( .INP(n15195), .ZN(n15194) );
  NOR2X0 U15890 ( .IN1(n15196), .IN2(n15197), .QN(n15195) );
  NAND2X0 U15891 ( .IN1(n15197), .IN2(n15196), .QN(n15193) );
  NOR2X0 U15892 ( .IN1(n15198), .IN2(n15199), .QN(n15196) );
  NOR2X0 U15893 ( .IN1(WX11233), .IN2(n7864), .QN(n15199) );
  INVX0 U15894 ( .INP(n15200), .ZN(n15198) );
  NAND2X0 U15895 ( .IN1(n7864), .IN2(WX11233), .QN(n15200) );
  NAND2X0 U15896 ( .IN1(n15201), .IN2(n15202), .QN(n15197) );
  NAND2X0 U15897 ( .IN1(n7863), .IN2(WX11105), .QN(n15202) );
  INVX0 U15898 ( .INP(n15203), .ZN(n15201) );
  NOR2X0 U15899 ( .IN1(WX11105), .IN2(n7863), .QN(n15203) );
  NAND2X0 U15900 ( .IN1(n1964), .IN2(n9287), .QN(n15191) );
  NOR2X0 U15901 ( .IN1(n9228), .IN2(n9037), .QN(n1964) );
  NAND2X0 U15902 ( .IN1(DATA_0_5), .IN2(n9336), .QN(n15190) );
  NAND2X0 U15903 ( .IN1(n9301), .IN2(CRC_OUT_1_5), .QN(n15189) );
  NAND4X0 U15904 ( .IN1(n15204), .IN2(n15205), .IN3(n15206), .IN4(n15207), 
        .QN(WX11038) );
  NAND3X0 U15905 ( .IN1(n9999), .IN2(n10000), .IN3(n9091), .QN(n15207) );
  NAND3X0 U15906 ( .IN1(n15208), .IN2(n15209), .IN3(n15210), .QN(n10000) );
  INVX0 U15907 ( .INP(n15211), .ZN(n15210) );
  NAND2X0 U15908 ( .IN1(n15211), .IN2(n15212), .QN(n9999) );
  NAND2X0 U15909 ( .IN1(n15208), .IN2(n15209), .QN(n15212) );
  NAND2X0 U15910 ( .IN1(n8156), .IN2(WX11167), .QN(n15209) );
  NAND2X0 U15911 ( .IN1(n7866), .IN2(WX11231), .QN(n15208) );
  NOR2X0 U15912 ( .IN1(n15213), .IN2(n15214), .QN(n15211) );
  INVX0 U15913 ( .INP(n15215), .ZN(n15214) );
  NAND2X0 U15914 ( .IN1(test_so94), .IN2(WX11039), .QN(n15215) );
  NOR2X0 U15915 ( .IN1(WX11039), .IN2(test_so94), .QN(n15213) );
  NAND2X0 U15916 ( .IN1(n1963), .IN2(n9288), .QN(n15206) );
  NOR2X0 U15917 ( .IN1(n9228), .IN2(n9038), .QN(n1963) );
  NAND2X0 U15918 ( .IN1(DATA_0_6), .IN2(n9335), .QN(n15205) );
  NAND2X0 U15919 ( .IN1(n9301), .IN2(CRC_OUT_1_6), .QN(n15204) );
  NAND4X0 U15920 ( .IN1(n15216), .IN2(n15217), .IN3(n15218), .IN4(n15219), 
        .QN(WX11036) );
  NAND2X0 U15921 ( .IN1(n9103), .IN2(n10007), .QN(n15219) );
  NAND2X0 U15922 ( .IN1(n15220), .IN2(n15221), .QN(n10007) );
  INVX0 U15923 ( .INP(n15222), .ZN(n15221) );
  NOR2X0 U15924 ( .IN1(n15223), .IN2(n15224), .QN(n15222) );
  NAND2X0 U15925 ( .IN1(n15224), .IN2(n15223), .QN(n15220) );
  NOR2X0 U15926 ( .IN1(n15225), .IN2(n15226), .QN(n15223) );
  NOR2X0 U15927 ( .IN1(WX11229), .IN2(n7868), .QN(n15226) );
  INVX0 U15928 ( .INP(n15227), .ZN(n15225) );
  NAND2X0 U15929 ( .IN1(n7868), .IN2(WX11229), .QN(n15227) );
  NAND2X0 U15930 ( .IN1(n15228), .IN2(n15229), .QN(n15224) );
  NAND2X0 U15931 ( .IN1(n7867), .IN2(WX11101), .QN(n15229) );
  INVX0 U15932 ( .INP(n15230), .ZN(n15228) );
  NOR2X0 U15933 ( .IN1(WX11101), .IN2(n7867), .QN(n15230) );
  NAND2X0 U15934 ( .IN1(n1962), .IN2(n9288), .QN(n15218) );
  NOR2X0 U15935 ( .IN1(n9228), .IN2(n9039), .QN(n1962) );
  NAND2X0 U15936 ( .IN1(DATA_0_7), .IN2(n9336), .QN(n15217) );
  NAND2X0 U15937 ( .IN1(n9301), .IN2(CRC_OUT_1_7), .QN(n15216) );
  NAND4X0 U15938 ( .IN1(n15231), .IN2(n15232), .IN3(n15233), .IN4(n15234), 
        .QN(WX11034) );
  NAND3X0 U15939 ( .IN1(n10012), .IN2(n10013), .IN3(n9091), .QN(n15234) );
  NAND3X0 U15940 ( .IN1(n15235), .IN2(n15236), .IN3(n15237), .QN(n10013) );
  INVX0 U15941 ( .INP(n15238), .ZN(n15237) );
  NAND2X0 U15942 ( .IN1(n15238), .IN2(n15239), .QN(n10012) );
  NAND2X0 U15943 ( .IN1(n15235), .IN2(n15236), .QN(n15239) );
  NAND2X0 U15944 ( .IN1(n8154), .IN2(WX11099), .QN(n15236) );
  NAND2X0 U15945 ( .IN1(n3547), .IN2(WX11227), .QN(n15235) );
  NOR2X0 U15946 ( .IN1(n15240), .IN2(n15241), .QN(n15238) );
  INVX0 U15947 ( .INP(n15242), .ZN(n15241) );
  NAND2X0 U15948 ( .IN1(test_so92), .IN2(WX11163), .QN(n15242) );
  NOR2X0 U15949 ( .IN1(WX11163), .IN2(test_so92), .QN(n15240) );
  NAND2X0 U15950 ( .IN1(n1961), .IN2(n9288), .QN(n15233) );
  NOR2X0 U15951 ( .IN1(n9228), .IN2(n9040), .QN(n1961) );
  NAND2X0 U15952 ( .IN1(DATA_0_8), .IN2(n9335), .QN(n15232) );
  NAND2X0 U15953 ( .IN1(n9301), .IN2(CRC_OUT_1_8), .QN(n15231) );
  NAND4X0 U15954 ( .IN1(n15243), .IN2(n15244), .IN3(n15245), .IN4(n15246), 
        .QN(WX11032) );
  NAND2X0 U15955 ( .IN1(n9103), .IN2(n10020), .QN(n15246) );
  NAND2X0 U15956 ( .IN1(n15247), .IN2(n15248), .QN(n10020) );
  INVX0 U15957 ( .INP(n15249), .ZN(n15248) );
  NOR2X0 U15958 ( .IN1(n15250), .IN2(n15251), .QN(n15249) );
  NAND2X0 U15959 ( .IN1(n15251), .IN2(n15250), .QN(n15247) );
  NOR2X0 U15960 ( .IN1(n15252), .IN2(n15253), .QN(n15250) );
  NOR2X0 U15961 ( .IN1(WX11225), .IN2(n7871), .QN(n15253) );
  INVX0 U15962 ( .INP(n15254), .ZN(n15252) );
  NAND2X0 U15963 ( .IN1(n7871), .IN2(WX11225), .QN(n15254) );
  NAND2X0 U15964 ( .IN1(n15255), .IN2(n15256), .QN(n15251) );
  NAND2X0 U15965 ( .IN1(n7870), .IN2(WX11097), .QN(n15256) );
  INVX0 U15966 ( .INP(n15257), .ZN(n15255) );
  NOR2X0 U15967 ( .IN1(WX11097), .IN2(n7870), .QN(n15257) );
  NAND2X0 U15968 ( .IN1(n1960), .IN2(n9288), .QN(n15245) );
  NOR2X0 U15969 ( .IN1(n9229), .IN2(n9041), .QN(n1960) );
  NAND2X0 U15970 ( .IN1(DATA_0_9), .IN2(n9335), .QN(n15244) );
  NAND2X0 U15971 ( .IN1(n9301), .IN2(CRC_OUT_1_9), .QN(n15243) );
  NAND4X0 U15972 ( .IN1(n15258), .IN2(n15259), .IN3(n15260), .IN4(n15261), 
        .QN(WX11030) );
  NAND2X0 U15973 ( .IN1(n9103), .IN2(n10026), .QN(n15261) );
  NAND2X0 U15974 ( .IN1(n15262), .IN2(n15263), .QN(n10026) );
  INVX0 U15975 ( .INP(n15264), .ZN(n15263) );
  NOR2X0 U15976 ( .IN1(n15265), .IN2(n15266), .QN(n15264) );
  NAND2X0 U15977 ( .IN1(n15266), .IN2(n15265), .QN(n15262) );
  NOR2X0 U15978 ( .IN1(n15267), .IN2(n15268), .QN(n15265) );
  NOR2X0 U15979 ( .IN1(WX11223), .IN2(n7873), .QN(n15268) );
  INVX0 U15980 ( .INP(n15269), .ZN(n15267) );
  NAND2X0 U15981 ( .IN1(n7873), .IN2(WX11223), .QN(n15269) );
  NAND2X0 U15982 ( .IN1(n15270), .IN2(n15271), .QN(n15266) );
  NAND2X0 U15983 ( .IN1(n7872), .IN2(WX11095), .QN(n15271) );
  INVX0 U15984 ( .INP(n15272), .ZN(n15270) );
  NOR2X0 U15985 ( .IN1(WX11095), .IN2(n7872), .QN(n15272) );
  NAND2X0 U15986 ( .IN1(n1959), .IN2(n9288), .QN(n15260) );
  NOR2X0 U15987 ( .IN1(n9075), .IN2(n9156), .QN(n1959) );
  NAND2X0 U15988 ( .IN1(DATA_0_10), .IN2(n9335), .QN(n15259) );
  NAND2X0 U15989 ( .IN1(n9301), .IN2(CRC_OUT_1_10), .QN(n15258) );
  NAND4X0 U15990 ( .IN1(n15273), .IN2(n15274), .IN3(n15275), .IN4(n15276), 
        .QN(WX11028) );
  NAND2X0 U15991 ( .IN1(n9103), .IN2(n10032), .QN(n15276) );
  NAND2X0 U15992 ( .IN1(n15277), .IN2(n15278), .QN(n10032) );
  INVX0 U15993 ( .INP(n15279), .ZN(n15278) );
  NOR2X0 U15994 ( .IN1(n15280), .IN2(n15281), .QN(n15279) );
  NAND2X0 U15995 ( .IN1(n15281), .IN2(n15280), .QN(n15277) );
  NOR2X0 U15996 ( .IN1(n15282), .IN2(n15283), .QN(n15280) );
  NOR2X0 U15997 ( .IN1(WX11221), .IN2(n7875), .QN(n15283) );
  INVX0 U15998 ( .INP(n15284), .ZN(n15282) );
  NAND2X0 U15999 ( .IN1(n7875), .IN2(WX11221), .QN(n15284) );
  NAND2X0 U16000 ( .IN1(n15285), .IN2(n15286), .QN(n15281) );
  NAND2X0 U16001 ( .IN1(n7874), .IN2(WX11093), .QN(n15286) );
  INVX0 U16002 ( .INP(n15287), .ZN(n15285) );
  NOR2X0 U16003 ( .IN1(WX11093), .IN2(n7874), .QN(n15287) );
  NAND2X0 U16004 ( .IN1(n1958), .IN2(n9288), .QN(n15275) );
  NOR2X0 U16005 ( .IN1(n9229), .IN2(n9042), .QN(n1958) );
  NAND2X0 U16006 ( .IN1(DATA_0_11), .IN2(n9335), .QN(n15274) );
  NAND2X0 U16007 ( .IN1(n9302), .IN2(CRC_OUT_1_11), .QN(n15273) );
  NAND4X0 U16008 ( .IN1(n15288), .IN2(n15289), .IN3(n15290), .IN4(n15291), 
        .QN(WX11026) );
  NAND2X0 U16009 ( .IN1(n9103), .IN2(n10038), .QN(n15291) );
  NAND2X0 U16010 ( .IN1(n15292), .IN2(n15293), .QN(n10038) );
  INVX0 U16011 ( .INP(n15294), .ZN(n15293) );
  NOR2X0 U16012 ( .IN1(n15295), .IN2(n15296), .QN(n15294) );
  NAND2X0 U16013 ( .IN1(n15296), .IN2(n15295), .QN(n15292) );
  NOR2X0 U16014 ( .IN1(n15297), .IN2(n15298), .QN(n15295) );
  NOR2X0 U16015 ( .IN1(WX11219), .IN2(n7877), .QN(n15298) );
  INVX0 U16016 ( .INP(n15299), .ZN(n15297) );
  NAND2X0 U16017 ( .IN1(n7877), .IN2(WX11219), .QN(n15299) );
  NAND2X0 U16018 ( .IN1(n15300), .IN2(n15301), .QN(n15296) );
  NAND2X0 U16019 ( .IN1(n7876), .IN2(WX11091), .QN(n15301) );
  INVX0 U16020 ( .INP(n15302), .ZN(n15300) );
  NOR2X0 U16021 ( .IN1(WX11091), .IN2(n7876), .QN(n15302) );
  NAND2X0 U16022 ( .IN1(n1957), .IN2(n9288), .QN(n15290) );
  NOR2X0 U16023 ( .IN1(n9229), .IN2(n9043), .QN(n1957) );
  NAND2X0 U16024 ( .IN1(DATA_0_12), .IN2(n9335), .QN(n15289) );
  NAND2X0 U16025 ( .IN1(n9302), .IN2(CRC_OUT_1_12), .QN(n15288) );
  NAND4X0 U16026 ( .IN1(n15303), .IN2(n15304), .IN3(n15305), .IN4(n15306), 
        .QN(WX11024) );
  NAND2X0 U16027 ( .IN1(n9102), .IN2(n10044), .QN(n15306) );
  NAND2X0 U16028 ( .IN1(n15307), .IN2(n15308), .QN(n10044) );
  INVX0 U16029 ( .INP(n15309), .ZN(n15308) );
  NOR2X0 U16030 ( .IN1(n15310), .IN2(n15311), .QN(n15309) );
  NAND2X0 U16031 ( .IN1(n15311), .IN2(n15310), .QN(n15307) );
  NOR2X0 U16032 ( .IN1(n15312), .IN2(n15313), .QN(n15310) );
  NOR2X0 U16033 ( .IN1(WX11217), .IN2(n7879), .QN(n15313) );
  INVX0 U16034 ( .INP(n15314), .ZN(n15312) );
  NAND2X0 U16035 ( .IN1(n7879), .IN2(WX11217), .QN(n15314) );
  NAND2X0 U16036 ( .IN1(n15315), .IN2(n15316), .QN(n15311) );
  NAND2X0 U16037 ( .IN1(n7878), .IN2(WX11089), .QN(n15316) );
  INVX0 U16038 ( .INP(n15317), .ZN(n15315) );
  NOR2X0 U16039 ( .IN1(WX11089), .IN2(n7878), .QN(n15317) );
  NAND2X0 U16040 ( .IN1(n1956), .IN2(n9288), .QN(n15305) );
  NOR2X0 U16041 ( .IN1(n9229), .IN2(n9044), .QN(n1956) );
  NAND2X0 U16042 ( .IN1(DATA_0_13), .IN2(n9335), .QN(n15304) );
  NAND2X0 U16043 ( .IN1(n9302), .IN2(CRC_OUT_1_13), .QN(n15303) );
  NAND4X0 U16044 ( .IN1(n15318), .IN2(n15319), .IN3(n15320), .IN4(n15321), 
        .QN(WX11022) );
  NAND2X0 U16045 ( .IN1(n9102), .IN2(n10051), .QN(n15321) );
  NAND2X0 U16046 ( .IN1(n15322), .IN2(n15323), .QN(n10051) );
  INVX0 U16047 ( .INP(n15324), .ZN(n15323) );
  NOR2X0 U16048 ( .IN1(n15325), .IN2(n15326), .QN(n15324) );
  NAND2X0 U16049 ( .IN1(n15326), .IN2(n15325), .QN(n15322) );
  NOR2X0 U16050 ( .IN1(n15327), .IN2(n15328), .QN(n15325) );
  NOR2X0 U16051 ( .IN1(WX11215), .IN2(n7881), .QN(n15328) );
  INVX0 U16052 ( .INP(n15329), .ZN(n15327) );
  NAND2X0 U16053 ( .IN1(n7881), .IN2(WX11215), .QN(n15329) );
  NAND2X0 U16054 ( .IN1(n15330), .IN2(n15331), .QN(n15326) );
  NAND2X0 U16055 ( .IN1(n7880), .IN2(WX11087), .QN(n15331) );
  INVX0 U16056 ( .INP(n15332), .ZN(n15330) );
  NOR2X0 U16057 ( .IN1(WX11087), .IN2(n7880), .QN(n15332) );
  NAND2X0 U16058 ( .IN1(n1955), .IN2(n9288), .QN(n15320) );
  NOR2X0 U16059 ( .IN1(n9229), .IN2(n9045), .QN(n1955) );
  NAND2X0 U16060 ( .IN1(DATA_0_14), .IN2(n9335), .QN(n15319) );
  NAND2X0 U16061 ( .IN1(test_so99), .IN2(n9314), .QN(n15318) );
  NAND4X0 U16062 ( .IN1(n15333), .IN2(n15334), .IN3(n15335), .IN4(n15336), 
        .QN(WX11020) );
  NAND2X0 U16063 ( .IN1(n9102), .IN2(n10057), .QN(n15336) );
  NAND2X0 U16064 ( .IN1(n15337), .IN2(n15338), .QN(n10057) );
  INVX0 U16065 ( .INP(n15339), .ZN(n15338) );
  NOR2X0 U16066 ( .IN1(n15340), .IN2(n15341), .QN(n15339) );
  NAND2X0 U16067 ( .IN1(n15341), .IN2(n15340), .QN(n15337) );
  NOR2X0 U16068 ( .IN1(n15342), .IN2(n15343), .QN(n15340) );
  NOR2X0 U16069 ( .IN1(WX11213), .IN2(n7883), .QN(n15343) );
  INVX0 U16070 ( .INP(n15344), .ZN(n15342) );
  NAND2X0 U16071 ( .IN1(n7883), .IN2(WX11213), .QN(n15344) );
  NAND2X0 U16072 ( .IN1(n15345), .IN2(n15346), .QN(n15341) );
  NAND2X0 U16073 ( .IN1(n7882), .IN2(WX11085), .QN(n15346) );
  INVX0 U16074 ( .INP(n15347), .ZN(n15345) );
  NOR2X0 U16075 ( .IN1(WX11085), .IN2(n7882), .QN(n15347) );
  NAND2X0 U16076 ( .IN1(n1954), .IN2(n9288), .QN(n15335) );
  NOR2X0 U16077 ( .IN1(n9229), .IN2(n9046), .QN(n1954) );
  NAND2X0 U16078 ( .IN1(DATA_0_15), .IN2(n9335), .QN(n15334) );
  NAND2X0 U16079 ( .IN1(n9302), .IN2(CRC_OUT_1_15), .QN(n15333) );
  NAND4X0 U16080 ( .IN1(n15348), .IN2(n15349), .IN3(n15350), .IN4(n15351), 
        .QN(WX11018) );
  NAND2X0 U16081 ( .IN1(n15352), .IN2(n10063), .QN(n15351) );
  NAND2X0 U16082 ( .IN1(n15353), .IN2(n10067), .QN(n10063) );
  NAND2X0 U16083 ( .IN1(n15354), .IN2(n15355), .QN(n15353) );
  NAND2X0 U16084 ( .IN1(n16427), .IN2(n9123), .QN(n15355) );
  NAND2X0 U16085 ( .IN1(TM1), .IN2(n8246), .QN(n15354) );
  NAND2X0 U16086 ( .IN1(n15356), .IN2(n15357), .QN(n15352) );
  NAND2X0 U16087 ( .IN1(n9102), .IN2(n10067), .QN(n15357) );
  NAND2X0 U16088 ( .IN1(n15358), .IN2(n15359), .QN(n10067) );
  NAND2X0 U16089 ( .IN1(n7628), .IN2(n15360), .QN(n15359) );
  INVX0 U16090 ( .INP(n15361), .ZN(n15358) );
  NOR2X0 U16091 ( .IN1(n15360), .IN2(n7628), .QN(n15361) );
  NOR2X0 U16092 ( .IN1(n15362), .IN2(n15363), .QN(n15360) );
  NOR2X0 U16093 ( .IN1(WX11211), .IN2(n7629), .QN(n15363) );
  INVX0 U16094 ( .INP(n15364), .ZN(n15362) );
  NAND2X0 U16095 ( .IN1(n7629), .IN2(WX11211), .QN(n15364) );
  NAND2X0 U16096 ( .IN1(n9102), .IN2(n8246), .QN(n15356) );
  NAND2X0 U16097 ( .IN1(n1953), .IN2(n9288), .QN(n15350) );
  NOR2X0 U16098 ( .IN1(n9229), .IN2(n9047), .QN(n1953) );
  NAND2X0 U16099 ( .IN1(DATA_0_16), .IN2(n9335), .QN(n15349) );
  NAND2X0 U16100 ( .IN1(n9302), .IN2(CRC_OUT_1_16), .QN(n15348) );
  NAND4X0 U16101 ( .IN1(n15365), .IN2(n15366), .IN3(n15367), .IN4(n15368), 
        .QN(WX11016) );
  NAND2X0 U16102 ( .IN1(n15369), .IN2(n10081), .QN(n15368) );
  NAND2X0 U16103 ( .IN1(n15370), .IN2(n10085), .QN(n10081) );
  NAND2X0 U16104 ( .IN1(n15371), .IN2(n15372), .QN(n15370) );
  NAND2X0 U16105 ( .IN1(n16426), .IN2(n9123), .QN(n15372) );
  NAND2X0 U16106 ( .IN1(TM1), .IN2(n8247), .QN(n15371) );
  NAND2X0 U16107 ( .IN1(n15373), .IN2(n15374), .QN(n15369) );
  NAND2X0 U16108 ( .IN1(n9102), .IN2(n10085), .QN(n15374) );
  NAND2X0 U16109 ( .IN1(n15375), .IN2(n15376), .QN(n10085) );
  NAND2X0 U16110 ( .IN1(n7630), .IN2(n15377), .QN(n15376) );
  INVX0 U16111 ( .INP(n15378), .ZN(n15375) );
  NOR2X0 U16112 ( .IN1(n15377), .IN2(n7630), .QN(n15378) );
  NOR2X0 U16113 ( .IN1(n15379), .IN2(n15380), .QN(n15377) );
  NOR2X0 U16114 ( .IN1(WX11209), .IN2(n7631), .QN(n15380) );
  INVX0 U16115 ( .INP(n15381), .ZN(n15379) );
  NAND2X0 U16116 ( .IN1(n7631), .IN2(WX11209), .QN(n15381) );
  NAND2X0 U16117 ( .IN1(n9102), .IN2(n8247), .QN(n15373) );
  NAND2X0 U16118 ( .IN1(n1952), .IN2(n9288), .QN(n15367) );
  NOR2X0 U16119 ( .IN1(n9229), .IN2(n9048), .QN(n1952) );
  NAND2X0 U16120 ( .IN1(DATA_0_17), .IN2(n9335), .QN(n15366) );
  NAND2X0 U16121 ( .IN1(n9302), .IN2(CRC_OUT_1_17), .QN(n15365) );
  NAND4X0 U16122 ( .IN1(n15382), .IN2(n15383), .IN3(n15384), .IN4(n15385), 
        .QN(WX11014) );
  NAND2X0 U16123 ( .IN1(n15386), .IN2(n10091), .QN(n15385) );
  NAND2X0 U16124 ( .IN1(n15387), .IN2(n10095), .QN(n10091) );
  NAND2X0 U16125 ( .IN1(n15388), .IN2(n15389), .QN(n15387) );
  NAND2X0 U16126 ( .IN1(n16425), .IN2(n9123), .QN(n15389) );
  NAND2X0 U16127 ( .IN1(TM1), .IN2(n8248), .QN(n15388) );
  NAND2X0 U16128 ( .IN1(n15390), .IN2(n15391), .QN(n15386) );
  NAND2X0 U16129 ( .IN1(n9102), .IN2(n10095), .QN(n15391) );
  NAND2X0 U16130 ( .IN1(n15392), .IN2(n15393), .QN(n10095) );
  NAND2X0 U16131 ( .IN1(n7632), .IN2(n15394), .QN(n15393) );
  INVX0 U16132 ( .INP(n15395), .ZN(n15392) );
  NOR2X0 U16133 ( .IN1(n15394), .IN2(n7632), .QN(n15395) );
  NOR2X0 U16134 ( .IN1(n15396), .IN2(n15397), .QN(n15394) );
  NOR2X0 U16135 ( .IN1(WX11207), .IN2(n7633), .QN(n15397) );
  INVX0 U16136 ( .INP(n15398), .ZN(n15396) );
  NAND2X0 U16137 ( .IN1(n7633), .IN2(WX11207), .QN(n15398) );
  NAND2X0 U16138 ( .IN1(n9106), .IN2(n8248), .QN(n15390) );
  NAND2X0 U16139 ( .IN1(n1951), .IN2(n9288), .QN(n15384) );
  NOR2X0 U16140 ( .IN1(n9229), .IN2(n9049), .QN(n1951) );
  NAND2X0 U16141 ( .IN1(DATA_0_18), .IN2(n9335), .QN(n15383) );
  NAND2X0 U16142 ( .IN1(n9302), .IN2(CRC_OUT_1_18), .QN(n15382) );
  NAND4X0 U16143 ( .IN1(n15399), .IN2(n15400), .IN3(n15401), .IN4(n15402), 
        .QN(WX11012) );
  NAND2X0 U16144 ( .IN1(n10106), .IN2(n9111), .QN(n15402) );
  NOR2X0 U16145 ( .IN1(n15403), .IN2(n15404), .QN(n10106) );
  INVX0 U16146 ( .INP(n15405), .ZN(n15404) );
  NAND2X0 U16147 ( .IN1(n15406), .IN2(n15407), .QN(n15405) );
  NOR2X0 U16148 ( .IN1(n15407), .IN2(n15406), .QN(n15403) );
  NAND2X0 U16149 ( .IN1(n15408), .IN2(n15409), .QN(n15406) );
  NAND2X0 U16150 ( .IN1(n15410), .IN2(WX11141), .QN(n15409) );
  NAND2X0 U16151 ( .IN1(n15411), .IN2(n15412), .QN(n15410) );
  NAND3X0 U16152 ( .IN1(n15411), .IN2(n15412), .IN3(n7635), .QN(n15408) );
  NAND2X0 U16153 ( .IN1(test_so97), .IN2(WX11077), .QN(n15412) );
  NAND2X0 U16154 ( .IN1(n7634), .IN2(n8804), .QN(n15411) );
  NOR2X0 U16155 ( .IN1(n15413), .IN2(n15414), .QN(n15407) );
  INVX0 U16156 ( .INP(n15415), .ZN(n15414) );
  NAND2X0 U16157 ( .IN1(n16424), .IN2(n9123), .QN(n15415) );
  NOR2X0 U16158 ( .IN1(n9117), .IN2(n16424), .QN(n15413) );
  NAND2X0 U16159 ( .IN1(n1950), .IN2(n9288), .QN(n15401) );
  NOR2X0 U16160 ( .IN1(n9229), .IN2(n9050), .QN(n1950) );
  NAND2X0 U16161 ( .IN1(DATA_0_19), .IN2(n9335), .QN(n15400) );
  NAND2X0 U16162 ( .IN1(n9302), .IN2(CRC_OUT_1_19), .QN(n15399) );
  NAND4X0 U16163 ( .IN1(n15416), .IN2(n15417), .IN3(n15418), .IN4(n15419), 
        .QN(WX11010) );
  NAND2X0 U16164 ( .IN1(n15420), .IN2(n10117), .QN(n15419) );
  NAND2X0 U16165 ( .IN1(n15421), .IN2(n10121), .QN(n10117) );
  NAND2X0 U16166 ( .IN1(n15422), .IN2(n15423), .QN(n15421) );
  NAND2X0 U16167 ( .IN1(n16423), .IN2(n9123), .QN(n15423) );
  NAND2X0 U16168 ( .IN1(TM1), .IN2(n8250), .QN(n15422) );
  NAND2X0 U16169 ( .IN1(n15424), .IN2(n15425), .QN(n15420) );
  NAND2X0 U16170 ( .IN1(n9102), .IN2(n10121), .QN(n15425) );
  NAND2X0 U16171 ( .IN1(n15426), .IN2(n15427), .QN(n10121) );
  NAND2X0 U16172 ( .IN1(n7636), .IN2(n15428), .QN(n15427) );
  INVX0 U16173 ( .INP(n15429), .ZN(n15426) );
  NOR2X0 U16174 ( .IN1(n15428), .IN2(n7636), .QN(n15429) );
  NOR2X0 U16175 ( .IN1(n15430), .IN2(n15431), .QN(n15428) );
  NOR2X0 U16176 ( .IN1(WX11203), .IN2(n7637), .QN(n15431) );
  INVX0 U16177 ( .INP(n15432), .ZN(n15430) );
  NAND2X0 U16178 ( .IN1(n7637), .IN2(WX11203), .QN(n15432) );
  NAND2X0 U16179 ( .IN1(n9102), .IN2(n8250), .QN(n15424) );
  NAND2X0 U16180 ( .IN1(n1949), .IN2(n9288), .QN(n15418) );
  NOR2X0 U16181 ( .IN1(n9229), .IN2(n9051), .QN(n1949) );
  NAND2X0 U16182 ( .IN1(DATA_0_20), .IN2(n9335), .QN(n15417) );
  NAND2X0 U16183 ( .IN1(n9302), .IN2(CRC_OUT_1_20), .QN(n15416) );
  NAND4X0 U16184 ( .IN1(n15433), .IN2(n15434), .IN3(n15435), .IN4(n15436), 
        .QN(WX11008) );
  NAND2X0 U16185 ( .IN1(n10131), .IN2(n9111), .QN(n15436) );
  NOR2X0 U16186 ( .IN1(n15437), .IN2(n15438), .QN(n10131) );
  INVX0 U16187 ( .INP(n15439), .ZN(n15438) );
  NAND2X0 U16188 ( .IN1(n15440), .IN2(n15441), .QN(n15439) );
  NOR2X0 U16189 ( .IN1(n15441), .IN2(n15440), .QN(n15437) );
  NAND2X0 U16190 ( .IN1(n15442), .IN2(n15443), .QN(n15440) );
  NAND2X0 U16191 ( .IN1(n8144), .IN2(n15444), .QN(n15443) );
  INVX0 U16192 ( .INP(n15445), .ZN(n15444) );
  NAND2X0 U16193 ( .IN1(n15445), .IN2(WX11201), .QN(n15442) );
  NAND2X0 U16194 ( .IN1(n15446), .IN2(n15447), .QN(n15445) );
  INVX0 U16195 ( .INP(n15448), .ZN(n15447) );
  NOR2X0 U16196 ( .IN1(n8818), .IN2(n16422), .QN(n15448) );
  NAND2X0 U16197 ( .IN1(n16422), .IN2(n8818), .QN(n15446) );
  NOR2X0 U16198 ( .IN1(n15449), .IN2(n15450), .QN(n15441) );
  INVX0 U16199 ( .INP(n15451), .ZN(n15450) );
  NAND2X0 U16200 ( .IN1(n7638), .IN2(n9123), .QN(n15451) );
  NOR2X0 U16201 ( .IN1(n9118), .IN2(n7638), .QN(n15449) );
  NAND2X0 U16202 ( .IN1(n1948), .IN2(n9288), .QN(n15435) );
  NOR2X0 U16203 ( .IN1(n9229), .IN2(n9052), .QN(n1948) );
  NAND2X0 U16204 ( .IN1(DATA_0_21), .IN2(n9335), .QN(n15434) );
  NAND2X0 U16205 ( .IN1(n9302), .IN2(CRC_OUT_1_21), .QN(n15433) );
  NAND4X0 U16206 ( .IN1(n15452), .IN2(n15453), .IN3(n15454), .IN4(n15455), 
        .QN(WX11006) );
  NAND2X0 U16207 ( .IN1(n15456), .IN2(n10142), .QN(n15455) );
  NAND2X0 U16208 ( .IN1(n15457), .IN2(n10146), .QN(n10142) );
  NAND2X0 U16209 ( .IN1(n15458), .IN2(n15459), .QN(n15457) );
  NAND2X0 U16210 ( .IN1(n16421), .IN2(n9123), .QN(n15459) );
  NAND2X0 U16211 ( .IN1(TM1), .IN2(n8252), .QN(n15458) );
  NAND2X0 U16212 ( .IN1(n15460), .IN2(n15461), .QN(n15456) );
  NAND2X0 U16213 ( .IN1(n9102), .IN2(n10146), .QN(n15461) );
  NAND2X0 U16214 ( .IN1(n15462), .IN2(n15463), .QN(n10146) );
  NAND2X0 U16215 ( .IN1(n7639), .IN2(n15464), .QN(n15463) );
  INVX0 U16216 ( .INP(n15465), .ZN(n15462) );
  NOR2X0 U16217 ( .IN1(n15464), .IN2(n7639), .QN(n15465) );
  NOR2X0 U16218 ( .IN1(n15466), .IN2(n15467), .QN(n15464) );
  NOR2X0 U16219 ( .IN1(WX11199), .IN2(n7640), .QN(n15467) );
  INVX0 U16220 ( .INP(n15468), .ZN(n15466) );
  NAND2X0 U16221 ( .IN1(n7640), .IN2(WX11199), .QN(n15468) );
  NAND2X0 U16222 ( .IN1(n9102), .IN2(n8252), .QN(n15460) );
  NAND2X0 U16223 ( .IN1(n1947), .IN2(n9288), .QN(n15454) );
  NOR2X0 U16224 ( .IN1(n9229), .IN2(n9053), .QN(n1947) );
  NAND2X0 U16225 ( .IN1(DATA_0_22), .IN2(n9335), .QN(n15453) );
  NAND2X0 U16226 ( .IN1(n9302), .IN2(CRC_OUT_1_22), .QN(n15452) );
  NAND4X0 U16227 ( .IN1(n15469), .IN2(n15470), .IN3(n15471), .IN4(n15472), 
        .QN(WX11004) );
  NAND2X0 U16228 ( .IN1(n10156), .IN2(n9112), .QN(n15472) );
  NOR2X0 U16229 ( .IN1(n15473), .IN2(n15474), .QN(n10156) );
  INVX0 U16230 ( .INP(n15475), .ZN(n15474) );
  NAND2X0 U16231 ( .IN1(n15476), .IN2(n15477), .QN(n15475) );
  NOR2X0 U16232 ( .IN1(n15477), .IN2(n15476), .QN(n15473) );
  NAND2X0 U16233 ( .IN1(n15478), .IN2(n15479), .QN(n15476) );
  NAND2X0 U16234 ( .IN1(n8142), .IN2(n15480), .QN(n15479) );
  INVX0 U16235 ( .INP(n15481), .ZN(n15480) );
  NAND2X0 U16236 ( .IN1(n15481), .IN2(WX11197), .QN(n15478) );
  NAND2X0 U16237 ( .IN1(n15482), .IN2(n15483), .QN(n15481) );
  INVX0 U16238 ( .INP(n15484), .ZN(n15483) );
  NOR2X0 U16239 ( .IN1(n8819), .IN2(n16420), .QN(n15484) );
  NAND2X0 U16240 ( .IN1(n16420), .IN2(n8819), .QN(n15482) );
  NOR2X0 U16241 ( .IN1(n15485), .IN2(n15486), .QN(n15477) );
  INVX0 U16242 ( .INP(n15487), .ZN(n15486) );
  NAND2X0 U16243 ( .IN1(n7641), .IN2(n9123), .QN(n15487) );
  NOR2X0 U16244 ( .IN1(n9117), .IN2(n7641), .QN(n15485) );
  NAND2X0 U16245 ( .IN1(n1946), .IN2(n9289), .QN(n15471) );
  NOR2X0 U16246 ( .IN1(n9229), .IN2(n9054), .QN(n1946) );
  NAND2X0 U16247 ( .IN1(DATA_0_23), .IN2(n9335), .QN(n15470) );
  NAND2X0 U16248 ( .IN1(n9302), .IN2(CRC_OUT_1_23), .QN(n15469) );
  NAND4X0 U16249 ( .IN1(n15488), .IN2(n15489), .IN3(n15490), .IN4(n15491), 
        .QN(WX11002) );
  NAND2X0 U16250 ( .IN1(n15492), .IN2(n10167), .QN(n15491) );
  NAND2X0 U16251 ( .IN1(n15493), .IN2(n10171), .QN(n10167) );
  NAND2X0 U16252 ( .IN1(n15494), .IN2(n15495), .QN(n15493) );
  NAND2X0 U16253 ( .IN1(n16419), .IN2(n9123), .QN(n15495) );
  NAND2X0 U16254 ( .IN1(TM1), .IN2(n8254), .QN(n15494) );
  NAND2X0 U16255 ( .IN1(n15496), .IN2(n15497), .QN(n15492) );
  NAND2X0 U16256 ( .IN1(n9102), .IN2(n10171), .QN(n15497) );
  NAND2X0 U16257 ( .IN1(n15498), .IN2(n15499), .QN(n10171) );
  NAND2X0 U16258 ( .IN1(n7642), .IN2(n15500), .QN(n15499) );
  INVX0 U16259 ( .INP(n15501), .ZN(n15498) );
  NOR2X0 U16260 ( .IN1(n15500), .IN2(n7642), .QN(n15501) );
  NOR2X0 U16261 ( .IN1(n15502), .IN2(n15503), .QN(n15500) );
  NOR2X0 U16262 ( .IN1(WX11195), .IN2(n7643), .QN(n15503) );
  INVX0 U16263 ( .INP(n15504), .ZN(n15502) );
  NAND2X0 U16264 ( .IN1(n7643), .IN2(WX11195), .QN(n15504) );
  NAND2X0 U16265 ( .IN1(n9102), .IN2(n8254), .QN(n15496) );
  NAND2X0 U16266 ( .IN1(n1945), .IN2(n9289), .QN(n15490) );
  NOR2X0 U16267 ( .IN1(n9229), .IN2(n9055), .QN(n1945) );
  NAND2X0 U16268 ( .IN1(DATA_0_24), .IN2(n9335), .QN(n15489) );
  NAND2X0 U16269 ( .IN1(n9303), .IN2(CRC_OUT_1_24), .QN(n15488) );
  NAND4X0 U16270 ( .IN1(n15505), .IN2(n15506), .IN3(n15507), .IN4(n15508), 
        .QN(WX11000) );
  NAND2X0 U16271 ( .IN1(n15509), .IN2(n10182), .QN(n15508) );
  NAND3X0 U16272 ( .IN1(n15510), .IN2(n15511), .IN3(n10186), .QN(n10182) );
  NAND2X0 U16273 ( .IN1(n8140), .IN2(n9123), .QN(n15511) );
  NAND2X0 U16274 ( .IN1(TM1), .IN2(WX11193), .QN(n15510) );
  NAND2X0 U16275 ( .IN1(n15512), .IN2(n15513), .QN(n15509) );
  NAND2X0 U16276 ( .IN1(n9102), .IN2(n10186), .QN(n15513) );
  NAND2X0 U16277 ( .IN1(n15514), .IN2(n15515), .QN(n10186) );
  NAND2X0 U16278 ( .IN1(n15516), .IN2(WX11129), .QN(n15515) );
  NAND2X0 U16279 ( .IN1(n15517), .IN2(n15518), .QN(n15516) );
  NAND3X0 U16280 ( .IN1(n15517), .IN2(n15518), .IN3(n7645), .QN(n15514) );
  NAND2X0 U16281 ( .IN1(test_so91), .IN2(WX11065), .QN(n15518) );
  NAND2X0 U16282 ( .IN1(n7644), .IN2(n8826), .QN(n15517) );
  NAND2X0 U16283 ( .IN1(n8140), .IN2(n9112), .QN(n15512) );
  NAND2X0 U16284 ( .IN1(n1944), .IN2(n9289), .QN(n15507) );
  NOR2X0 U16285 ( .IN1(n9230), .IN2(n9056), .QN(n1944) );
  NAND2X0 U16286 ( .IN1(DATA_0_25), .IN2(n9334), .QN(n15506) );
  NAND2X0 U16287 ( .IN1(n9303), .IN2(CRC_OUT_1_25), .QN(n15505) );
  NAND4X0 U16288 ( .IN1(n15519), .IN2(n15520), .IN3(n15521), .IN4(n15522), 
        .QN(WX10998) );
  NAND2X0 U16289 ( .IN1(n15523), .IN2(n10197), .QN(n15522) );
  NAND2X0 U16290 ( .IN1(n15524), .IN2(n10201), .QN(n10197) );
  NAND2X0 U16291 ( .IN1(n15525), .IN2(n15526), .QN(n15524) );
  NAND2X0 U16292 ( .IN1(n16418), .IN2(n9123), .QN(n15526) );
  NAND2X0 U16293 ( .IN1(TM1), .IN2(n8257), .QN(n15525) );
  NAND2X0 U16294 ( .IN1(n15527), .IN2(n15528), .QN(n15523) );
  NAND2X0 U16295 ( .IN1(n9102), .IN2(n10201), .QN(n15528) );
  NAND2X0 U16296 ( .IN1(n15529), .IN2(n15530), .QN(n10201) );
  NAND2X0 U16297 ( .IN1(n7646), .IN2(n15531), .QN(n15530) );
  INVX0 U16298 ( .INP(n15532), .ZN(n15529) );
  NOR2X0 U16299 ( .IN1(n15531), .IN2(n7646), .QN(n15532) );
  NOR2X0 U16300 ( .IN1(n15533), .IN2(n15534), .QN(n15531) );
  NOR2X0 U16301 ( .IN1(WX11191), .IN2(n7647), .QN(n15534) );
  INVX0 U16302 ( .INP(n15535), .ZN(n15533) );
  NAND2X0 U16303 ( .IN1(n7647), .IN2(WX11191), .QN(n15535) );
  NAND2X0 U16304 ( .IN1(n9102), .IN2(n8257), .QN(n15527) );
  NAND2X0 U16305 ( .IN1(n1943), .IN2(n9289), .QN(n15521) );
  NOR2X0 U16306 ( .IN1(n9230), .IN2(n9057), .QN(n1943) );
  NAND2X0 U16307 ( .IN1(DATA_0_26), .IN2(n9334), .QN(n15520) );
  NAND2X0 U16308 ( .IN1(n9303), .IN2(CRC_OUT_1_26), .QN(n15519) );
  NAND4X0 U16309 ( .IN1(n15536), .IN2(n15537), .IN3(n15538), .IN4(n15539), 
        .QN(WX10996) );
  NAND2X0 U16310 ( .IN1(n15540), .IN2(n10212), .QN(n15539) );
  NAND2X0 U16311 ( .IN1(n15541), .IN2(n10216), .QN(n10212) );
  NAND2X0 U16312 ( .IN1(n15542), .IN2(n15543), .QN(n15541) );
  NAND2X0 U16313 ( .IN1(n16417), .IN2(n9123), .QN(n15543) );
  NAND2X0 U16314 ( .IN1(TM1), .IN2(n8258), .QN(n15542) );
  NAND2X0 U16315 ( .IN1(n15544), .IN2(n15545), .QN(n15540) );
  NAND2X0 U16316 ( .IN1(n9101), .IN2(n10216), .QN(n15545) );
  NAND2X0 U16317 ( .IN1(n15546), .IN2(n15547), .QN(n10216) );
  NAND2X0 U16318 ( .IN1(n7648), .IN2(n15548), .QN(n15547) );
  INVX0 U16319 ( .INP(n15549), .ZN(n15546) );
  NOR2X0 U16320 ( .IN1(n15548), .IN2(n7648), .QN(n15549) );
  NOR2X0 U16321 ( .IN1(n15550), .IN2(n15551), .QN(n15548) );
  NOR2X0 U16322 ( .IN1(WX11189), .IN2(n7649), .QN(n15551) );
  INVX0 U16323 ( .INP(n15552), .ZN(n15550) );
  NAND2X0 U16324 ( .IN1(n7649), .IN2(WX11189), .QN(n15552) );
  NAND2X0 U16325 ( .IN1(n9101), .IN2(n8258), .QN(n15544) );
  NAND2X0 U16326 ( .IN1(n1942), .IN2(n9289), .QN(n15538) );
  NOR2X0 U16327 ( .IN1(n9076), .IN2(n9157), .QN(n1942) );
  NAND2X0 U16328 ( .IN1(DATA_0_27), .IN2(n9335), .QN(n15537) );
  NAND2X0 U16329 ( .IN1(n9303), .IN2(CRC_OUT_1_27), .QN(n15536) );
  NAND4X0 U16330 ( .IN1(n15553), .IN2(n15554), .IN3(n15555), .IN4(n15556), 
        .QN(WX10994) );
  NAND2X0 U16331 ( .IN1(n15557), .IN2(n10227), .QN(n15556) );
  NAND2X0 U16332 ( .IN1(n15558), .IN2(n10231), .QN(n10227) );
  NAND2X0 U16333 ( .IN1(n15559), .IN2(n15560), .QN(n15558) );
  NAND2X0 U16334 ( .IN1(n16416), .IN2(n9123), .QN(n15560) );
  NAND2X0 U16335 ( .IN1(TM1), .IN2(n8259), .QN(n15559) );
  NAND2X0 U16336 ( .IN1(n15561), .IN2(n15562), .QN(n15557) );
  NAND2X0 U16337 ( .IN1(n9101), .IN2(n10231), .QN(n15562) );
  NAND2X0 U16338 ( .IN1(n15563), .IN2(n15564), .QN(n10231) );
  NAND2X0 U16339 ( .IN1(n7650), .IN2(n15565), .QN(n15564) );
  INVX0 U16340 ( .INP(n15566), .ZN(n15563) );
  NOR2X0 U16341 ( .IN1(n15565), .IN2(n7650), .QN(n15566) );
  NOR2X0 U16342 ( .IN1(n15567), .IN2(n15568), .QN(n15565) );
  NOR2X0 U16343 ( .IN1(WX11187), .IN2(n7651), .QN(n15568) );
  INVX0 U16344 ( .INP(n15569), .ZN(n15567) );
  NAND2X0 U16345 ( .IN1(n7651), .IN2(WX11187), .QN(n15569) );
  NAND2X0 U16346 ( .IN1(n9101), .IN2(n8259), .QN(n15561) );
  NAND2X0 U16347 ( .IN1(n1941), .IN2(n9289), .QN(n15555) );
  NOR2X0 U16348 ( .IN1(n9230), .IN2(n9058), .QN(n1941) );
  NAND2X0 U16349 ( .IN1(DATA_0_28), .IN2(n9334), .QN(n15554) );
  NAND2X0 U16350 ( .IN1(n9303), .IN2(CRC_OUT_1_28), .QN(n15553) );
  NAND4X0 U16351 ( .IN1(n15570), .IN2(n15571), .IN3(n15572), .IN4(n15573), 
        .QN(WX10992) );
  NAND2X0 U16352 ( .IN1(n15574), .IN2(n10242), .QN(n15573) );
  NAND2X0 U16353 ( .IN1(n15575), .IN2(n10246), .QN(n10242) );
  NAND2X0 U16354 ( .IN1(n15576), .IN2(n15577), .QN(n15575) );
  NAND2X0 U16355 ( .IN1(n16415), .IN2(n9123), .QN(n15577) );
  NAND2X0 U16356 ( .IN1(TM1), .IN2(n8260), .QN(n15576) );
  NAND2X0 U16357 ( .IN1(n15578), .IN2(n15579), .QN(n15574) );
  NAND2X0 U16358 ( .IN1(n9101), .IN2(n10246), .QN(n15579) );
  NAND2X0 U16359 ( .IN1(n15580), .IN2(n15581), .QN(n10246) );
  NAND2X0 U16360 ( .IN1(n7652), .IN2(n15582), .QN(n15581) );
  INVX0 U16361 ( .INP(n15583), .ZN(n15580) );
  NOR2X0 U16362 ( .IN1(n15582), .IN2(n7652), .QN(n15583) );
  NOR2X0 U16363 ( .IN1(n15584), .IN2(n15585), .QN(n15582) );
  NOR2X0 U16364 ( .IN1(WX11185), .IN2(n7653), .QN(n15585) );
  INVX0 U16365 ( .INP(n15586), .ZN(n15584) );
  NAND2X0 U16366 ( .IN1(n7653), .IN2(WX11185), .QN(n15586) );
  NAND2X0 U16367 ( .IN1(n9101), .IN2(n8260), .QN(n15578) );
  NAND2X0 U16368 ( .IN1(n1940), .IN2(n9289), .QN(n15572) );
  NOR2X0 U16369 ( .IN1(n9230), .IN2(n9059), .QN(n1940) );
  NAND2X0 U16370 ( .IN1(DATA_0_29), .IN2(n9334), .QN(n15571) );
  NAND2X0 U16371 ( .IN1(n9303), .IN2(CRC_OUT_1_29), .QN(n15570) );
  NAND4X0 U16372 ( .IN1(n15587), .IN2(n15588), .IN3(n15589), .IN4(n15590), 
        .QN(WX10990) );
  NAND2X0 U16373 ( .IN1(n15591), .IN2(n10257), .QN(n15590) );
  NAND2X0 U16374 ( .IN1(n15592), .IN2(n10261), .QN(n10257) );
  NAND2X0 U16375 ( .IN1(n15593), .IN2(n15594), .QN(n15592) );
  NAND2X0 U16376 ( .IN1(n16414), .IN2(n9123), .QN(n15594) );
  NAND2X0 U16377 ( .IN1(TM1), .IN2(n8261), .QN(n15593) );
  NAND2X0 U16378 ( .IN1(n15595), .IN2(n15596), .QN(n15591) );
  NAND2X0 U16379 ( .IN1(n9101), .IN2(n10261), .QN(n15596) );
  NAND2X0 U16380 ( .IN1(n15597), .IN2(n15598), .QN(n10261) );
  NAND2X0 U16381 ( .IN1(n7654), .IN2(n15599), .QN(n15598) );
  INVX0 U16382 ( .INP(n15600), .ZN(n15597) );
  NOR2X0 U16383 ( .IN1(n15599), .IN2(n7654), .QN(n15600) );
  NOR2X0 U16384 ( .IN1(n15601), .IN2(n15602), .QN(n15599) );
  NOR2X0 U16385 ( .IN1(WX11183), .IN2(n7655), .QN(n15602) );
  INVX0 U16386 ( .INP(n15603), .ZN(n15601) );
  NAND2X0 U16387 ( .IN1(n7655), .IN2(WX11183), .QN(n15603) );
  NAND2X0 U16388 ( .IN1(n9101), .IN2(n8261), .QN(n15595) );
  NAND2X0 U16389 ( .IN1(n1939), .IN2(n9289), .QN(n15589) );
  NOR2X0 U16390 ( .IN1(n9117), .IN2(n2183), .QN(n2148) );
  NOR2X0 U16391 ( .IN1(n9230), .IN2(n9060), .QN(n1939) );
  NAND2X0 U16392 ( .IN1(DATA_0_30), .IN2(n9334), .QN(n15588) );
  NAND2X0 U16393 ( .IN1(n9303), .IN2(CRC_OUT_1_30), .QN(n15587) );
  NAND4X0 U16394 ( .IN1(n15604), .IN2(n15605), .IN3(n15606), .IN4(n15607), 
        .QN(WX10988) );
  NAND2X0 U16395 ( .IN1(n15608), .IN2(n10267), .QN(n15607) );
  NAND2X0 U16396 ( .IN1(n15609), .IN2(n10271), .QN(n10267) );
  NAND2X0 U16397 ( .IN1(n15610), .IN2(n15611), .QN(n15609) );
  NAND2X0 U16398 ( .IN1(n16413), .IN2(n9123), .QN(n15611) );
  NAND2X0 U16399 ( .IN1(TM1), .IN2(n8262), .QN(n15610) );
  NAND2X0 U16400 ( .IN1(n15612), .IN2(n15613), .QN(n15608) );
  NAND2X0 U16401 ( .IN1(n9102), .IN2(n10271), .QN(n15613) );
  NAND2X0 U16402 ( .IN1(n15614), .IN2(n15615), .QN(n10271) );
  NAND2X0 U16403 ( .IN1(n7612), .IN2(n15616), .QN(n15615) );
  INVX0 U16404 ( .INP(n15617), .ZN(n15614) );
  NOR2X0 U16405 ( .IN1(n15616), .IN2(n7612), .QN(n15617) );
  NOR2X0 U16406 ( .IN1(n15618), .IN2(n15619), .QN(n15616) );
  NOR2X0 U16407 ( .IN1(WX11181), .IN2(n7613), .QN(n15619) );
  INVX0 U16408 ( .INP(n15620), .ZN(n15618) );
  NAND2X0 U16409 ( .IN1(n7613), .IN2(WX11181), .QN(n15620) );
  NAND2X0 U16410 ( .IN1(n9092), .IN2(n8262), .QN(n15612) );
  NOR3X0 U16411 ( .IN1(n9152), .IN2(TM0), .IN3(n9116), .QN(n9958) );
  NAND2X0 U16412 ( .IN1(DATA_0_31), .IN2(n2153), .QN(n15606) );
  NAND2X0 U16413 ( .IN1(test_so100), .IN2(n9315), .QN(n15605) );
  NAND2X0 U16414 ( .IN1(n2245), .IN2(WX10829), .QN(n15604) );
  NOR2X0 U16415 ( .IN1(n9230), .IN2(WX10829), .QN(WX10890) );
  NOR2X0 U16416 ( .IN1(n9230), .IN2(n15621), .QN(WX10377) );
  NOR2X0 U16417 ( .IN1(n15622), .IN2(n15623), .QN(n15621) );
  NOR2X0 U16418 ( .IN1(test_so85), .IN2(CRC_OUT_2_30), .QN(n15623) );
  NOR2X0 U16419 ( .IN1(DFF_1534_n1), .IN2(n8805), .QN(n15622) );
  NOR3X0 U16420 ( .IN1(n9152), .IN2(n15624), .IN3(n15625), .QN(WX10375) );
  NOR2X0 U16421 ( .IN1(n8160), .IN2(CRC_OUT_2_29), .QN(n15625) );
  NOR2X0 U16422 ( .IN1(DFF_1533_n1), .IN2(WX9890), .QN(n15624) );
  NOR3X0 U16423 ( .IN1(n9152), .IN2(n15626), .IN3(n15627), .QN(WX10373) );
  NOR2X0 U16424 ( .IN1(n8161), .IN2(CRC_OUT_2_28), .QN(n15627) );
  NOR2X0 U16425 ( .IN1(DFF_1532_n1), .IN2(WX9892), .QN(n15626) );
  NOR3X0 U16426 ( .IN1(n9152), .IN2(n15628), .IN3(n15629), .QN(WX10371) );
  NOR2X0 U16427 ( .IN1(n8162), .IN2(CRC_OUT_2_27), .QN(n15629) );
  NOR2X0 U16428 ( .IN1(DFF_1531_n1), .IN2(WX9894), .QN(n15628) );
  NOR3X0 U16429 ( .IN1(n9152), .IN2(n15630), .IN3(n15631), .QN(WX10369) );
  NOR2X0 U16430 ( .IN1(n8163), .IN2(CRC_OUT_2_26), .QN(n15631) );
  NOR2X0 U16431 ( .IN1(DFF_1530_n1), .IN2(WX9896), .QN(n15630) );
  NOR3X0 U16432 ( .IN1(n9152), .IN2(n15632), .IN3(n15633), .QN(WX10367) );
  NOR2X0 U16433 ( .IN1(n8164), .IN2(CRC_OUT_2_25), .QN(n15633) );
  NOR2X0 U16434 ( .IN1(DFF_1529_n1), .IN2(WX9898), .QN(n15632) );
  NOR3X0 U16435 ( .IN1(n9152), .IN2(n15634), .IN3(n15635), .QN(WX10365) );
  NOR2X0 U16436 ( .IN1(n8165), .IN2(CRC_OUT_2_24), .QN(n15635) );
  NOR2X0 U16437 ( .IN1(DFF_1528_n1), .IN2(WX9900), .QN(n15634) );
  NOR3X0 U16438 ( .IN1(n9152), .IN2(n15636), .IN3(n15637), .QN(WX10363) );
  NOR2X0 U16439 ( .IN1(n8166), .IN2(CRC_OUT_2_23), .QN(n15637) );
  NOR2X0 U16440 ( .IN1(DFF_1527_n1), .IN2(WX9902), .QN(n15636) );
  NOR3X0 U16441 ( .IN1(n9152), .IN2(n15638), .IN3(n15639), .QN(WX10361) );
  NOR2X0 U16442 ( .IN1(n8167), .IN2(CRC_OUT_2_22), .QN(n15639) );
  NOR2X0 U16443 ( .IN1(DFF_1526_n1), .IN2(WX9904), .QN(n15638) );
  NOR3X0 U16444 ( .IN1(n9152), .IN2(n15640), .IN3(n15641), .QN(WX10359) );
  NOR2X0 U16445 ( .IN1(n8168), .IN2(CRC_OUT_2_21), .QN(n15641) );
  NOR2X0 U16446 ( .IN1(DFF_1525_n1), .IN2(WX9906), .QN(n15640) );
  NOR3X0 U16447 ( .IN1(n9153), .IN2(n15642), .IN3(n15643), .QN(WX10357) );
  NOR2X0 U16448 ( .IN1(n8169), .IN2(CRC_OUT_2_20), .QN(n15643) );
  NOR2X0 U16449 ( .IN1(DFF_1524_n1), .IN2(WX9908), .QN(n15642) );
  NOR2X0 U16450 ( .IN1(n9231), .IN2(n15644), .QN(WX10355) );
  NOR2X0 U16451 ( .IN1(n15645), .IN2(n15646), .QN(n15644) );
  NOR2X0 U16452 ( .IN1(test_so88), .IN2(WX9910), .QN(n15646) );
  INVX0 U16453 ( .INP(n15647), .ZN(n15645) );
  NAND2X0 U16454 ( .IN1(WX9910), .IN2(test_so88), .QN(n15647) );
  NOR3X0 U16455 ( .IN1(n9153), .IN2(n15648), .IN3(n15649), .QN(WX10353) );
  NOR2X0 U16456 ( .IN1(n8171), .IN2(CRC_OUT_2_18), .QN(n15649) );
  NOR2X0 U16457 ( .IN1(DFF_1522_n1), .IN2(WX9912), .QN(n15648) );
  NOR3X0 U16458 ( .IN1(n9152), .IN2(n15650), .IN3(n15651), .QN(WX10351) );
  NOR2X0 U16459 ( .IN1(n8172), .IN2(CRC_OUT_2_17), .QN(n15651) );
  NOR2X0 U16460 ( .IN1(DFF_1521_n1), .IN2(WX9914), .QN(n15650) );
  NOR3X0 U16461 ( .IN1(n9153), .IN2(n15652), .IN3(n15653), .QN(WX10349) );
  NOR2X0 U16462 ( .IN1(n8173), .IN2(CRC_OUT_2_16), .QN(n15653) );
  NOR2X0 U16463 ( .IN1(DFF_1520_n1), .IN2(WX9916), .QN(n15652) );
  NOR2X0 U16464 ( .IN1(n9231), .IN2(n15654), .QN(WX10347) );
  NOR2X0 U16465 ( .IN1(n15655), .IN2(n15656), .QN(n15654) );
  NOR2X0 U16466 ( .IN1(DFF_1519_n1), .IN2(n15657), .QN(n15656) );
  INVX0 U16467 ( .INP(n15658), .ZN(n15655) );
  NAND2X0 U16468 ( .IN1(n15657), .IN2(DFF_1519_n1), .QN(n15658) );
  NOR2X0 U16469 ( .IN1(n15659), .IN2(n15660), .QN(n15657) );
  NOR2X0 U16470 ( .IN1(WX9918), .IN2(DFF_1535_n1), .QN(n15660) );
  NOR2X0 U16471 ( .IN1(CRC_OUT_2_31), .IN2(n8108), .QN(n15659) );
  NOR3X0 U16472 ( .IN1(n9153), .IN2(n15661), .IN3(n15662), .QN(WX10345) );
  NOR2X0 U16473 ( .IN1(n8174), .IN2(CRC_OUT_2_14), .QN(n15662) );
  NOR2X0 U16474 ( .IN1(DFF_1518_n1), .IN2(WX9920), .QN(n15661) );
  NOR2X0 U16475 ( .IN1(n9231), .IN2(n15663), .QN(WX10343) );
  NOR2X0 U16476 ( .IN1(n15664), .IN2(n15665), .QN(n15663) );
  NOR2X0 U16477 ( .IN1(test_so86), .IN2(CRC_OUT_2_13), .QN(n15665) );
  NOR2X0 U16478 ( .IN1(DFF_1517_n1), .IN2(n8795), .QN(n15664) );
  NOR3X0 U16479 ( .IN1(n9153), .IN2(n15666), .IN3(n15667), .QN(WX10341) );
  NOR2X0 U16480 ( .IN1(n8175), .IN2(CRC_OUT_2_12), .QN(n15667) );
  NOR2X0 U16481 ( .IN1(DFF_1516_n1), .IN2(WX9924), .QN(n15666) );
  NOR3X0 U16482 ( .IN1(n9153), .IN2(n15668), .IN3(n15669), .QN(WX10339) );
  NOR2X0 U16483 ( .IN1(n8176), .IN2(CRC_OUT_2_11), .QN(n15669) );
  NOR2X0 U16484 ( .IN1(DFF_1515_n1), .IN2(WX9926), .QN(n15668) );
  NOR2X0 U16485 ( .IN1(n9231), .IN2(n15670), .QN(WX10337) );
  NOR2X0 U16486 ( .IN1(n15671), .IN2(n15672), .QN(n15670) );
  INVX0 U16487 ( .INP(n15673), .ZN(n15672) );
  NAND2X0 U16488 ( .IN1(CRC_OUT_2_10), .IN2(n15674), .QN(n15673) );
  NOR2X0 U16489 ( .IN1(n15674), .IN2(CRC_OUT_2_10), .QN(n15671) );
  NAND2X0 U16490 ( .IN1(n15675), .IN2(n15676), .QN(n15674) );
  NAND2X0 U16491 ( .IN1(n8109), .IN2(CRC_OUT_2_31), .QN(n15676) );
  NAND2X0 U16492 ( .IN1(DFF_1535_n1), .IN2(WX9928), .QN(n15675) );
  NOR3X0 U16493 ( .IN1(n9153), .IN2(n15677), .IN3(n15678), .QN(WX10335) );
  NOR2X0 U16494 ( .IN1(n8177), .IN2(CRC_OUT_2_9), .QN(n15678) );
  NOR2X0 U16495 ( .IN1(DFF_1513_n1), .IN2(WX9930), .QN(n15677) );
  NOR3X0 U16496 ( .IN1(n9153), .IN2(n15679), .IN3(n15680), .QN(WX10333) );
  NOR2X0 U16497 ( .IN1(n8178), .IN2(CRC_OUT_2_8), .QN(n15680) );
  NOR2X0 U16498 ( .IN1(DFF_1512_n1), .IN2(WX9932), .QN(n15679) );
  NOR3X0 U16499 ( .IN1(n9154), .IN2(n15681), .IN3(n15682), .QN(WX10331) );
  NOR2X0 U16500 ( .IN1(n8179), .IN2(CRC_OUT_2_7), .QN(n15682) );
  NOR2X0 U16501 ( .IN1(DFF_1511_n1), .IN2(WX9934), .QN(n15681) );
  NOR3X0 U16502 ( .IN1(n9153), .IN2(n15683), .IN3(n15684), .QN(WX10329) );
  NOR2X0 U16503 ( .IN1(n8180), .IN2(CRC_OUT_2_6), .QN(n15684) );
  NOR2X0 U16504 ( .IN1(DFF_1510_n1), .IN2(WX9936), .QN(n15683) );
  NOR3X0 U16505 ( .IN1(n9154), .IN2(n15685), .IN3(n15686), .QN(WX10327) );
  NOR2X0 U16506 ( .IN1(n8181), .IN2(CRC_OUT_2_5), .QN(n15686) );
  NOR2X0 U16507 ( .IN1(DFF_1509_n1), .IN2(WX9938), .QN(n15685) );
  NOR3X0 U16508 ( .IN1(n9154), .IN2(n15687), .IN3(n15688), .QN(WX10325) );
  NOR2X0 U16509 ( .IN1(n8182), .IN2(CRC_OUT_2_4), .QN(n15688) );
  NOR2X0 U16510 ( .IN1(DFF_1508_n1), .IN2(WX9940), .QN(n15687) );
  NOR2X0 U16511 ( .IN1(n9232), .IN2(n15689), .QN(WX10323) );
  NOR2X0 U16512 ( .IN1(n15690), .IN2(n15691), .QN(n15689) );
  INVX0 U16513 ( .INP(n15692), .ZN(n15691) );
  NAND2X0 U16514 ( .IN1(CRC_OUT_2_3), .IN2(n15693), .QN(n15692) );
  NOR2X0 U16515 ( .IN1(n15693), .IN2(CRC_OUT_2_3), .QN(n15690) );
  NAND2X0 U16516 ( .IN1(n15694), .IN2(n15695), .QN(n15693) );
  NAND2X0 U16517 ( .IN1(n8110), .IN2(CRC_OUT_2_31), .QN(n15695) );
  NAND2X0 U16518 ( .IN1(DFF_1535_n1), .IN2(WX9942), .QN(n15694) );
  NOR2X0 U16519 ( .IN1(n9232), .IN2(n15696), .QN(WX10321) );
  NOR2X0 U16520 ( .IN1(n15697), .IN2(n15698), .QN(n15696) );
  NOR2X0 U16521 ( .IN1(test_so87), .IN2(WX9944), .QN(n15698) );
  INVX0 U16522 ( .INP(n15699), .ZN(n15697) );
  NAND2X0 U16523 ( .IN1(WX9944), .IN2(test_so87), .QN(n15699) );
  NOR3X0 U16524 ( .IN1(n9153), .IN2(n15700), .IN3(n15701), .QN(WX10319) );
  NOR2X0 U16525 ( .IN1(n8184), .IN2(CRC_OUT_2_1), .QN(n15701) );
  NOR2X0 U16526 ( .IN1(DFF_1505_n1), .IN2(WX9946), .QN(n15700) );
  NOR3X0 U16527 ( .IN1(n9154), .IN2(n15702), .IN3(n15703), .QN(WX10317) );
  NOR2X0 U16528 ( .IN1(n8185), .IN2(CRC_OUT_2_0), .QN(n15703) );
  NOR2X0 U16529 ( .IN1(DFF_1504_n1), .IN2(WX9948), .QN(n15702) );
  NOR3X0 U16530 ( .IN1(n9136), .IN2(n15704), .IN3(n15705), .QN(WX10315) );
  NOR2X0 U16531 ( .IN1(n8127), .IN2(CRC_OUT_2_31), .QN(n15705) );
  NOR2X0 U16532 ( .IN1(DFF_1535_n1), .IN2(WX9950), .QN(n15704) );
  INVX0 U16533 ( .INP(RESET), .ZN(n2182) );
  NAND2X0 U16534 ( .IN1(n15706), .IN2(n15707), .QN(DATA_9_9) );
  INVX0 U16535 ( .INP(n15708), .ZN(n15707) );
  NOR2X0 U16536 ( .IN1(n15709), .IN2(n11716), .QN(n15708) );
  NAND2X0 U16537 ( .IN1(n11716), .IN2(n15709), .QN(n15706) );
  NAND2X0 U16538 ( .IN1(TM0), .IN2(WX529), .QN(n15709) );
  NAND2X0 U16539 ( .IN1(n15710), .IN2(n15711), .QN(n11716) );
  NAND2X0 U16540 ( .IN1(n15712), .IN2(n15713), .QN(n15711) );
  INVX0 U16541 ( .INP(n15714), .ZN(n15710) );
  NOR2X0 U16542 ( .IN1(n15713), .IN2(n15712), .QN(n15714) );
  NAND2X0 U16543 ( .IN1(n15715), .IN2(n15716), .QN(n15712) );
  NAND2X0 U16544 ( .IN1(n8741), .IN2(n15717), .QN(n15716) );
  INVX0 U16545 ( .INP(n15718), .ZN(n15715) );
  NOR2X0 U16546 ( .IN1(n15717), .IN2(n8741), .QN(n15718) );
  NOR2X0 U16547 ( .IN1(n15719), .IN2(n15720), .QN(n15717) );
  NOR2X0 U16548 ( .IN1(WX881), .IN2(n8742), .QN(n15720) );
  INVX0 U16549 ( .INP(n15721), .ZN(n15719) );
  NAND2X0 U16550 ( .IN1(n8742), .IN2(WX881), .QN(n15721) );
  NOR2X0 U16551 ( .IN1(n15722), .IN2(n15723), .QN(n15713) );
  INVX0 U16552 ( .INP(n15724), .ZN(n15723) );
  NAND2X0 U16553 ( .IN1(n3485), .IN2(n2183), .QN(n15724) );
  NOR2X0 U16554 ( .IN1(n2183), .IN2(n3485), .QN(n15722) );
  NAND2X0 U16555 ( .IN1(n15725), .IN2(n15726), .QN(DATA_9_8) );
  INVX0 U16556 ( .INP(n15727), .ZN(n15726) );
  NOR2X0 U16557 ( .IN1(n15728), .IN2(n11710), .QN(n15727) );
  NAND2X0 U16558 ( .IN1(n11710), .IN2(n15728), .QN(n15725) );
  NAND2X0 U16559 ( .IN1(TM0), .IN2(WX531), .QN(n15728) );
  NAND2X0 U16560 ( .IN1(n15729), .IN2(n15730), .QN(n11710) );
  NAND2X0 U16561 ( .IN1(n15731), .IN2(n15732), .QN(n15730) );
  INVX0 U16562 ( .INP(n15733), .ZN(n15729) );
  NOR2X0 U16563 ( .IN1(n15732), .IN2(n15731), .QN(n15733) );
  NAND2X0 U16564 ( .IN1(n15734), .IN2(n15735), .QN(n15731) );
  NAND2X0 U16565 ( .IN1(n8751), .IN2(n15736), .QN(n15735) );
  INVX0 U16566 ( .INP(n15737), .ZN(n15734) );
  NOR2X0 U16567 ( .IN1(n15736), .IN2(n8751), .QN(n15737) );
  NOR2X0 U16568 ( .IN1(n15738), .IN2(n15739), .QN(n15736) );
  INVX0 U16569 ( .INP(n15740), .ZN(n15739) );
  NAND2X0 U16570 ( .IN1(n8753), .IN2(WX883), .QN(n15740) );
  NOR2X0 U16571 ( .IN1(WX883), .IN2(n8753), .QN(n15738) );
  NOR2X0 U16572 ( .IN1(n15741), .IN2(n15742), .QN(n15732) );
  INVX0 U16573 ( .INP(n15743), .ZN(n15742) );
  NAND2X0 U16574 ( .IN1(n3483), .IN2(n2183), .QN(n15743) );
  NOR2X0 U16575 ( .IN1(n2183), .IN2(n3483), .QN(n15741) );
  NAND2X0 U16576 ( .IN1(n15744), .IN2(n15745), .QN(DATA_9_7) );
  INVX0 U16577 ( .INP(n15746), .ZN(n15745) );
  NOR2X0 U16578 ( .IN1(n15747), .IN2(n11704), .QN(n15746) );
  NAND2X0 U16579 ( .IN1(n11704), .IN2(n15747), .QN(n15744) );
  NAND2X0 U16580 ( .IN1(TM0), .IN2(WX533), .QN(n15747) );
  NAND2X0 U16581 ( .IN1(n15748), .IN2(n15749), .QN(n11704) );
  NAND2X0 U16582 ( .IN1(n15750), .IN2(n15751), .QN(n15749) );
  INVX0 U16583 ( .INP(n15752), .ZN(n15748) );
  NOR2X0 U16584 ( .IN1(n15751), .IN2(n15750), .QN(n15752) );
  NAND2X0 U16585 ( .IN1(n15753), .IN2(n15754), .QN(n15750) );
  NAND2X0 U16586 ( .IN1(n8781), .IN2(n15755), .QN(n15754) );
  INVX0 U16587 ( .INP(n15756), .ZN(n15753) );
  NOR2X0 U16588 ( .IN1(n15755), .IN2(n8781), .QN(n15756) );
  NOR2X0 U16589 ( .IN1(n15757), .IN2(n15758), .QN(n15755) );
  NOR2X0 U16590 ( .IN1(WX885), .IN2(n8782), .QN(n15758) );
  INVX0 U16591 ( .INP(n15759), .ZN(n15757) );
  NAND2X0 U16592 ( .IN1(n8782), .IN2(WX885), .QN(n15759) );
  NOR2X0 U16593 ( .IN1(n15760), .IN2(n15761), .QN(n15751) );
  INVX0 U16594 ( .INP(n15762), .ZN(n15761) );
  NAND2X0 U16595 ( .IN1(n3481), .IN2(n2183), .QN(n15762) );
  NOR2X0 U16596 ( .IN1(n2183), .IN2(n3481), .QN(n15760) );
  NOR2X0 U16597 ( .IN1(n15763), .IN2(n15764), .QN(DATA_9_6) );
  INVX0 U16598 ( .INP(n15765), .ZN(n15764) );
  NAND2X0 U16599 ( .IN1(n15766), .IN2(n11698), .QN(n15765) );
  NOR2X0 U16600 ( .IN1(n11698), .IN2(n15766), .QN(n15763) );
  NAND2X0 U16601 ( .IN1(TM0), .IN2(WX535), .QN(n15766) );
  NAND2X0 U16602 ( .IN1(n15767), .IN2(n15768), .QN(n11698) );
  NAND2X0 U16603 ( .IN1(n15769), .IN2(n15770), .QN(n15768) );
  NAND2X0 U16604 ( .IN1(n15771), .IN2(n15772), .QN(n15769) );
  NAND3X0 U16605 ( .IN1(n15771), .IN2(n15772), .IN3(n15773), .QN(n15767) );
  INVX0 U16606 ( .INP(n15770), .ZN(n15773) );
  NOR2X0 U16607 ( .IN1(n15774), .IN2(n15775), .QN(n15770) );
  INVX0 U16608 ( .INP(n15776), .ZN(n15775) );
  NAND2X0 U16609 ( .IN1(n8769), .IN2(n15777), .QN(n15776) );
  NOR2X0 U16610 ( .IN1(n15777), .IN2(n8769), .QN(n15774) );
  NOR2X0 U16611 ( .IN1(n15778), .IN2(n15779), .QN(n15777) );
  INVX0 U16612 ( .INP(n15780), .ZN(n15779) );
  NAND2X0 U16613 ( .IN1(test_so5), .IN2(WX887), .QN(n15780) );
  NOR2X0 U16614 ( .IN1(WX887), .IN2(test_so5), .QN(n15778) );
  NAND2X0 U16615 ( .IN1(n3479), .IN2(n2183), .QN(n15772) );
  NAND2X0 U16616 ( .IN1(TM0), .IN2(WX695), .QN(n15771) );
  NAND2X0 U16617 ( .IN1(n15781), .IN2(n15782), .QN(DATA_9_5) );
  INVX0 U16618 ( .INP(n15783), .ZN(n15782) );
  NOR2X0 U16619 ( .IN1(n15784), .IN2(n11691), .QN(n15783) );
  NAND2X0 U16620 ( .IN1(n11691), .IN2(n15784), .QN(n15781) );
  NAND2X0 U16621 ( .IN1(TM0), .IN2(WX537), .QN(n15784) );
  NAND2X0 U16622 ( .IN1(n15785), .IN2(n15786), .QN(n11691) );
  NAND2X0 U16623 ( .IN1(n15787), .IN2(n15788), .QN(n15786) );
  INVX0 U16624 ( .INP(n15789), .ZN(n15785) );
  NOR2X0 U16625 ( .IN1(n15788), .IN2(n15787), .QN(n15789) );
  NAND2X0 U16626 ( .IN1(n15790), .IN2(n15791), .QN(n15787) );
  NAND2X0 U16627 ( .IN1(n8754), .IN2(n15792), .QN(n15791) );
  INVX0 U16628 ( .INP(n15793), .ZN(n15790) );
  NOR2X0 U16629 ( .IN1(n15792), .IN2(n8754), .QN(n15793) );
  NOR2X0 U16630 ( .IN1(n15794), .IN2(n15795), .QN(n15792) );
  INVX0 U16631 ( .INP(n15796), .ZN(n15795) );
  NAND2X0 U16632 ( .IN1(n8756), .IN2(WX889), .QN(n15796) );
  NOR2X0 U16633 ( .IN1(WX889), .IN2(n8756), .QN(n15794) );
  NOR2X0 U16634 ( .IN1(n15797), .IN2(n15798), .QN(n15788) );
  INVX0 U16635 ( .INP(n15799), .ZN(n15798) );
  NAND2X0 U16636 ( .IN1(n3477), .IN2(n2183), .QN(n15799) );
  NOR2X0 U16637 ( .IN1(n2183), .IN2(n3477), .QN(n15797) );
  NAND2X0 U16638 ( .IN1(n15800), .IN2(n15801), .QN(DATA_9_4) );
  INVX0 U16639 ( .INP(n15802), .ZN(n15801) );
  NOR2X0 U16640 ( .IN1(n15803), .IN2(n11685), .QN(n15802) );
  NAND2X0 U16641 ( .IN1(n11685), .IN2(n15803), .QN(n15800) );
  NAND2X0 U16642 ( .IN1(TM0), .IN2(WX539), .QN(n15803) );
  NAND2X0 U16643 ( .IN1(n15804), .IN2(n15805), .QN(n11685) );
  NAND2X0 U16644 ( .IN1(n15806), .IN2(n15807), .QN(n15805) );
  INVX0 U16645 ( .INP(n15808), .ZN(n15804) );
  NOR2X0 U16646 ( .IN1(n15807), .IN2(n15806), .QN(n15808) );
  NAND2X0 U16647 ( .IN1(n15809), .IN2(n15810), .QN(n15806) );
  NAND2X0 U16648 ( .IN1(n8757), .IN2(n15811), .QN(n15810) );
  INVX0 U16649 ( .INP(n15812), .ZN(n15809) );
  NOR2X0 U16650 ( .IN1(n15811), .IN2(n8757), .QN(n15812) );
  NOR2X0 U16651 ( .IN1(n15813), .IN2(n15814), .QN(n15811) );
  INVX0 U16652 ( .INP(n15815), .ZN(n15814) );
  NAND2X0 U16653 ( .IN1(n8759), .IN2(WX891), .QN(n15815) );
  NOR2X0 U16654 ( .IN1(WX891), .IN2(n8759), .QN(n15813) );
  NOR2X0 U16655 ( .IN1(n15816), .IN2(n15817), .QN(n15807) );
  INVX0 U16656 ( .INP(n15818), .ZN(n15817) );
  NAND2X0 U16657 ( .IN1(n3475), .IN2(n2183), .QN(n15818) );
  NOR2X0 U16658 ( .IN1(n2183), .IN2(n3475), .QN(n15816) );
  NAND2X0 U16659 ( .IN1(n15819), .IN2(n15820), .QN(DATA_9_31) );
  INVX0 U16660 ( .INP(n15821), .ZN(n15820) );
  NOR2X0 U16661 ( .IN1(n15822), .IN2(n12001), .QN(n15821) );
  NAND2X0 U16662 ( .IN1(n12001), .IN2(n15822), .QN(n15819) );
  NAND2X0 U16663 ( .IN1(TM0), .IN2(WX485), .QN(n15822) );
  NAND2X0 U16664 ( .IN1(n15823), .IN2(n15824), .QN(n12001) );
  NAND2X0 U16665 ( .IN1(n15825), .IN2(n15826), .QN(n15824) );
  INVX0 U16666 ( .INP(n15827), .ZN(n15823) );
  NOR2X0 U16667 ( .IN1(n15826), .IN2(n15825), .QN(n15827) );
  NAND2X0 U16668 ( .IN1(n15828), .IN2(n15829), .QN(n15825) );
  NAND2X0 U16669 ( .IN1(n8773), .IN2(n15830), .QN(n15829) );
  INVX0 U16670 ( .INP(n15831), .ZN(n15828) );
  NOR2X0 U16671 ( .IN1(n15830), .IN2(n8773), .QN(n15831) );
  NOR2X0 U16672 ( .IN1(n15832), .IN2(n15833), .QN(n15830) );
  NOR2X0 U16673 ( .IN1(WX837), .IN2(n8774), .QN(n15833) );
  INVX0 U16674 ( .INP(n15834), .ZN(n15832) );
  NAND2X0 U16675 ( .IN1(n8774), .IN2(WX837), .QN(n15834) );
  NOR2X0 U16676 ( .IN1(n15835), .IN2(n15836), .QN(n15826) );
  INVX0 U16677 ( .INP(n15837), .ZN(n15836) );
  NAND2X0 U16678 ( .IN1(n3529), .IN2(n9124), .QN(n15837) );
  NOR2X0 U16679 ( .IN1(n9117), .IN2(n3529), .QN(n15835) );
  NAND2X0 U16680 ( .IN1(n15838), .IN2(n15839), .QN(DATA_9_30) );
  INVX0 U16681 ( .INP(n15840), .ZN(n15839) );
  NOR2X0 U16682 ( .IN1(n15841), .IN2(n11960), .QN(n15840) );
  NAND2X0 U16683 ( .IN1(n11960), .IN2(n15841), .QN(n15838) );
  NAND2X0 U16684 ( .IN1(TM0), .IN2(WX487), .QN(n15841) );
  NAND2X0 U16685 ( .IN1(n15842), .IN2(n15843), .QN(n11960) );
  NAND2X0 U16686 ( .IN1(n15844), .IN2(n15845), .QN(n15843) );
  INVX0 U16687 ( .INP(n15846), .ZN(n15842) );
  NOR2X0 U16688 ( .IN1(n15845), .IN2(n15844), .QN(n15846) );
  NAND2X0 U16689 ( .IN1(n15847), .IN2(n15848), .QN(n15844) );
  NAND2X0 U16690 ( .IN1(n8678), .IN2(n15849), .QN(n15848) );
  INVX0 U16691 ( .INP(n15850), .ZN(n15847) );
  NOR2X0 U16692 ( .IN1(n15849), .IN2(n8678), .QN(n15850) );
  NOR2X0 U16693 ( .IN1(n15851), .IN2(n15852), .QN(n15849) );
  NOR2X0 U16694 ( .IN1(WX839), .IN2(n8679), .QN(n15852) );
  INVX0 U16695 ( .INP(n15853), .ZN(n15851) );
  NAND2X0 U16696 ( .IN1(n8679), .IN2(WX839), .QN(n15853) );
  NOR2X0 U16697 ( .IN1(n15854), .IN2(n15855), .QN(n15845) );
  INVX0 U16698 ( .INP(n15856), .ZN(n15855) );
  NAND2X0 U16699 ( .IN1(n3527), .IN2(n9124), .QN(n15856) );
  NOR2X0 U16700 ( .IN1(n9116), .IN2(n3527), .QN(n15854) );
  NAND2X0 U16701 ( .IN1(n15857), .IN2(n15858), .QN(DATA_9_3) );
  INVX0 U16702 ( .INP(n15859), .ZN(n15858) );
  NOR2X0 U16703 ( .IN1(n15860), .IN2(n11678), .QN(n15859) );
  NAND2X0 U16704 ( .IN1(n11678), .IN2(n15860), .QN(n15857) );
  NAND2X0 U16705 ( .IN1(TM0), .IN2(WX541), .QN(n15860) );
  NAND2X0 U16706 ( .IN1(n15861), .IN2(n15862), .QN(n11678) );
  NAND2X0 U16707 ( .IN1(n15863), .IN2(n15864), .QN(n15862) );
  INVX0 U16708 ( .INP(n15865), .ZN(n15861) );
  NOR2X0 U16709 ( .IN1(n15864), .IN2(n15863), .QN(n15865) );
  NAND2X0 U16710 ( .IN1(n15866), .IN2(n15867), .QN(n15863) );
  NAND2X0 U16711 ( .IN1(n8698), .IN2(n15868), .QN(n15867) );
  INVX0 U16712 ( .INP(n15869), .ZN(n15866) );
  NOR2X0 U16713 ( .IN1(n15868), .IN2(n8698), .QN(n15869) );
  NOR2X0 U16714 ( .IN1(n15870), .IN2(n15871), .QN(n15868) );
  INVX0 U16715 ( .INP(n15872), .ZN(n15871) );
  NAND2X0 U16716 ( .IN1(n8704), .IN2(WX893), .QN(n15872) );
  NOR2X0 U16717 ( .IN1(WX893), .IN2(n8704), .QN(n15870) );
  NOR2X0 U16718 ( .IN1(n15873), .IN2(n15874), .QN(n15864) );
  INVX0 U16719 ( .INP(n15875), .ZN(n15874) );
  NAND2X0 U16720 ( .IN1(n3473), .IN2(n2183), .QN(n15875) );
  NOR2X0 U16721 ( .IN1(n2183), .IN2(n3473), .QN(n15873) );
  NAND2X0 U16722 ( .IN1(n15876), .IN2(n15877), .QN(DATA_9_29) );
  INVX0 U16723 ( .INP(n15878), .ZN(n15877) );
  NOR2X0 U16724 ( .IN1(n15879), .IN2(n11924), .QN(n15878) );
  NAND2X0 U16725 ( .IN1(n11924), .IN2(n15879), .QN(n15876) );
  NAND2X0 U16726 ( .IN1(TM0), .IN2(WX489), .QN(n15879) );
  NAND2X0 U16727 ( .IN1(n15880), .IN2(n15881), .QN(n11924) );
  NAND2X0 U16728 ( .IN1(n15882), .IN2(n15883), .QN(n15881) );
  INVX0 U16729 ( .INP(n15884), .ZN(n15880) );
  NOR2X0 U16730 ( .IN1(n15883), .IN2(n15882), .QN(n15884) );
  NAND2X0 U16731 ( .IN1(n15885), .IN2(n15886), .QN(n15882) );
  NAND2X0 U16732 ( .IN1(n8708), .IN2(n15887), .QN(n15886) );
  INVX0 U16733 ( .INP(n15888), .ZN(n15885) );
  NOR2X0 U16734 ( .IN1(n15887), .IN2(n8708), .QN(n15888) );
  NOR2X0 U16735 ( .IN1(n15889), .IN2(n15890), .QN(n15887) );
  INVX0 U16736 ( .INP(n15891), .ZN(n15890) );
  NAND2X0 U16737 ( .IN1(n8710), .IN2(WX841), .QN(n15891) );
  NOR2X0 U16738 ( .IN1(WX841), .IN2(n8710), .QN(n15889) );
  NOR2X0 U16739 ( .IN1(n15892), .IN2(n15893), .QN(n15883) );
  INVX0 U16740 ( .INP(n15894), .ZN(n15893) );
  NAND2X0 U16741 ( .IN1(n3525), .IN2(n9124), .QN(n15894) );
  NOR2X0 U16742 ( .IN1(n9116), .IN2(n3525), .QN(n15892) );
  NOR2X0 U16743 ( .IN1(n15895), .IN2(n15896), .QN(DATA_9_28) );
  INVX0 U16744 ( .INP(n15897), .ZN(n15896) );
  NAND2X0 U16745 ( .IN1(n15898), .IN2(n11892), .QN(n15897) );
  NOR2X0 U16746 ( .IN1(n11892), .IN2(n15898), .QN(n15895) );
  NAND2X0 U16747 ( .IN1(TM0), .IN2(WX491), .QN(n15898) );
  NAND2X0 U16748 ( .IN1(n15899), .IN2(n15900), .QN(n11892) );
  NAND2X0 U16749 ( .IN1(n15901), .IN2(n15902), .QN(n15900) );
  NAND2X0 U16750 ( .IN1(n15903), .IN2(n15904), .QN(n15901) );
  NAND3X0 U16751 ( .IN1(n15903), .IN2(n15904), .IN3(n15905), .QN(n15899) );
  INVX0 U16752 ( .INP(n15902), .ZN(n15905) );
  NOR2X0 U16753 ( .IN1(n15906), .IN2(n15907), .QN(n15902) );
  INVX0 U16754 ( .INP(n15908), .ZN(n15907) );
  NAND2X0 U16755 ( .IN1(n8717), .IN2(n15909), .QN(n15908) );
  NOR2X0 U16756 ( .IN1(n15909), .IN2(n8717), .QN(n15906) );
  NOR2X0 U16757 ( .IN1(n15910), .IN2(n15911), .QN(n15909) );
  INVX0 U16758 ( .INP(n15912), .ZN(n15911) );
  NAND2X0 U16759 ( .IN1(test_so2), .IN2(WX843), .QN(n15912) );
  NOR2X0 U16760 ( .IN1(WX843), .IN2(test_so2), .QN(n15910) );
  NAND2X0 U16761 ( .IN1(n8719), .IN2(n9124), .QN(n15904) );
  NAND2X0 U16762 ( .IN1(TM1), .IN2(WX715), .QN(n15903) );
  NAND2X0 U16763 ( .IN1(n15913), .IN2(n15914), .QN(DATA_9_27) );
  INVX0 U16764 ( .INP(n15915), .ZN(n15914) );
  NOR2X0 U16765 ( .IN1(n15916), .IN2(n11885), .QN(n15915) );
  NAND2X0 U16766 ( .IN1(n11885), .IN2(n15916), .QN(n15913) );
  NAND2X0 U16767 ( .IN1(TM0), .IN2(WX493), .QN(n15916) );
  NAND2X0 U16768 ( .IN1(n15917), .IN2(n15918), .QN(n11885) );
  NAND2X0 U16769 ( .IN1(n15919), .IN2(n15920), .QN(n15918) );
  INVX0 U16770 ( .INP(n15921), .ZN(n15917) );
  NOR2X0 U16771 ( .IN1(n15920), .IN2(n15919), .QN(n15921) );
  NAND2X0 U16772 ( .IN1(n15922), .IN2(n15923), .QN(n15919) );
  NAND2X0 U16773 ( .IN1(n8723), .IN2(n15924), .QN(n15923) );
  INVX0 U16774 ( .INP(n15925), .ZN(n15922) );
  NOR2X0 U16775 ( .IN1(n15924), .IN2(n8723), .QN(n15925) );
  NOR2X0 U16776 ( .IN1(n15926), .IN2(n15927), .QN(n15924) );
  INVX0 U16777 ( .INP(n15928), .ZN(n15927) );
  NAND2X0 U16778 ( .IN1(n8725), .IN2(WX845), .QN(n15928) );
  NOR2X0 U16779 ( .IN1(WX845), .IN2(n8725), .QN(n15926) );
  NOR2X0 U16780 ( .IN1(n15929), .IN2(n15930), .QN(n15920) );
  INVX0 U16781 ( .INP(n15931), .ZN(n15930) );
  NAND2X0 U16782 ( .IN1(n3521), .IN2(n9124), .QN(n15931) );
  NOR2X0 U16783 ( .IN1(n9116), .IN2(n3521), .QN(n15929) );
  NAND2X0 U16784 ( .IN1(n15932), .IN2(n15933), .QN(DATA_9_26) );
  INVX0 U16785 ( .INP(n15934), .ZN(n15933) );
  NOR2X0 U16786 ( .IN1(n15935), .IN2(n11874), .QN(n15934) );
  NAND2X0 U16787 ( .IN1(n11874), .IN2(n15935), .QN(n15932) );
  NAND2X0 U16788 ( .IN1(TM0), .IN2(WX495), .QN(n15935) );
  NAND2X0 U16789 ( .IN1(n15936), .IN2(n15937), .QN(n11874) );
  NAND2X0 U16790 ( .IN1(n15938), .IN2(n15939), .QN(n15937) );
  INVX0 U16791 ( .INP(n15940), .ZN(n15936) );
  NOR2X0 U16792 ( .IN1(n15939), .IN2(n15938), .QN(n15940) );
  NAND2X0 U16793 ( .IN1(n15941), .IN2(n15942), .QN(n15938) );
  NAND2X0 U16794 ( .IN1(n8726), .IN2(n15943), .QN(n15942) );
  INVX0 U16795 ( .INP(n15944), .ZN(n15941) );
  NOR2X0 U16796 ( .IN1(n15943), .IN2(n8726), .QN(n15944) );
  NOR2X0 U16797 ( .IN1(n15945), .IN2(n15946), .QN(n15943) );
  INVX0 U16798 ( .INP(n15947), .ZN(n15946) );
  NAND2X0 U16799 ( .IN1(n8728), .IN2(WX847), .QN(n15947) );
  NOR2X0 U16800 ( .IN1(WX847), .IN2(n8728), .QN(n15945) );
  NOR2X0 U16801 ( .IN1(n15948), .IN2(n15949), .QN(n15939) );
  INVX0 U16802 ( .INP(n15950), .ZN(n15949) );
  NAND2X0 U16803 ( .IN1(n3519), .IN2(n9124), .QN(n15950) );
  NOR2X0 U16804 ( .IN1(n9117), .IN2(n3519), .QN(n15948) );
  NAND2X0 U16805 ( .IN1(n15951), .IN2(n15952), .QN(DATA_9_25) );
  INVX0 U16806 ( .INP(n15953), .ZN(n15952) );
  NOR2X0 U16807 ( .IN1(n15954), .IN2(n11863), .QN(n15953) );
  NAND2X0 U16808 ( .IN1(n11863), .IN2(n15954), .QN(n15951) );
  NAND2X0 U16809 ( .IN1(TM0), .IN2(WX497), .QN(n15954) );
  NAND2X0 U16810 ( .IN1(n15955), .IN2(n15956), .QN(n11863) );
  NAND2X0 U16811 ( .IN1(n15957), .IN2(n15958), .QN(n15956) );
  INVX0 U16812 ( .INP(n15959), .ZN(n15955) );
  NOR2X0 U16813 ( .IN1(n15958), .IN2(n15957), .QN(n15959) );
  NAND2X0 U16814 ( .IN1(n15960), .IN2(n15961), .QN(n15957) );
  NAND2X0 U16815 ( .IN1(n8735), .IN2(n15962), .QN(n15961) );
  INVX0 U16816 ( .INP(n15963), .ZN(n15960) );
  NOR2X0 U16817 ( .IN1(n15962), .IN2(n8735), .QN(n15963) );
  NOR2X0 U16818 ( .IN1(n15964), .IN2(n15965), .QN(n15962) );
  INVX0 U16819 ( .INP(n15966), .ZN(n15965) );
  NAND2X0 U16820 ( .IN1(n8737), .IN2(WX849), .QN(n15966) );
  NOR2X0 U16821 ( .IN1(WX849), .IN2(n8737), .QN(n15964) );
  NOR2X0 U16822 ( .IN1(n15967), .IN2(n15968), .QN(n15958) );
  INVX0 U16823 ( .INP(n15969), .ZN(n15968) );
  NAND2X0 U16824 ( .IN1(n3517), .IN2(n9124), .QN(n15969) );
  NOR2X0 U16825 ( .IN1(n9116), .IN2(n3517), .QN(n15967) );
  NOR2X0 U16826 ( .IN1(n15970), .IN2(n15971), .QN(DATA_9_24) );
  INVX0 U16827 ( .INP(n15972), .ZN(n15971) );
  NAND2X0 U16828 ( .IN1(n15973), .IN2(n11852), .QN(n15972) );
  NOR2X0 U16829 ( .IN1(n11852), .IN2(n15973), .QN(n15970) );
  NAND2X0 U16830 ( .IN1(TM0), .IN2(WX499), .QN(n15973) );
  NAND2X0 U16831 ( .IN1(n15974), .IN2(n15975), .QN(n11852) );
  NAND2X0 U16832 ( .IN1(n15976), .IN2(n15977), .QN(n15975) );
  NAND2X0 U16833 ( .IN1(n15978), .IN2(n15979), .QN(n15976) );
  NAND3X0 U16834 ( .IN1(n15978), .IN2(n15979), .IN3(n15980), .QN(n15974) );
  INVX0 U16835 ( .INP(n15977), .ZN(n15980) );
  NOR2X0 U16836 ( .IN1(n15981), .IN2(n15982), .QN(n15977) );
  INVX0 U16837 ( .INP(n15983), .ZN(n15982) );
  NAND2X0 U16838 ( .IN1(n8744), .IN2(n15984), .QN(n15983) );
  NOR2X0 U16839 ( .IN1(n15984), .IN2(n8744), .QN(n15981) );
  NOR2X0 U16840 ( .IN1(n15985), .IN2(n15986), .QN(n15984) );
  INVX0 U16841 ( .INP(n15987), .ZN(n15986) );
  NAND2X0 U16842 ( .IN1(test_so4), .IN2(WX851), .QN(n15987) );
  NOR2X0 U16843 ( .IN1(WX851), .IN2(test_so4), .QN(n15985) );
  NAND2X0 U16844 ( .IN1(n3515), .IN2(n9124), .QN(n15979) );
  NAND2X0 U16845 ( .IN1(TM1), .IN2(WX659), .QN(n15978) );
  NAND2X0 U16846 ( .IN1(n15988), .IN2(n15989), .QN(DATA_9_23) );
  INVX0 U16847 ( .INP(n15990), .ZN(n15989) );
  NOR2X0 U16848 ( .IN1(n15991), .IN2(n11840), .QN(n15990) );
  NAND2X0 U16849 ( .IN1(n11840), .IN2(n15991), .QN(n15988) );
  NAND2X0 U16850 ( .IN1(TM0), .IN2(WX501), .QN(n15991) );
  NAND2X0 U16851 ( .IN1(n15992), .IN2(n15993), .QN(n11840) );
  NAND2X0 U16852 ( .IN1(n15994), .IN2(n15995), .QN(n15993) );
  INVX0 U16853 ( .INP(n15996), .ZN(n15992) );
  NOR2X0 U16854 ( .IN1(n15995), .IN2(n15994), .QN(n15996) );
  NAND2X0 U16855 ( .IN1(n15997), .IN2(n15998), .QN(n15994) );
  NAND2X0 U16856 ( .IN1(n8746), .IN2(n15999), .QN(n15998) );
  INVX0 U16857 ( .INP(n16000), .ZN(n15997) );
  NOR2X0 U16858 ( .IN1(n15999), .IN2(n8746), .QN(n16000) );
  NOR2X0 U16859 ( .IN1(n16001), .IN2(n16002), .QN(n15999) );
  INVX0 U16860 ( .INP(n16003), .ZN(n16002) );
  NAND2X0 U16861 ( .IN1(n8748), .IN2(WX853), .QN(n16003) );
  NOR2X0 U16862 ( .IN1(WX853), .IN2(n8748), .QN(n16001) );
  NOR2X0 U16863 ( .IN1(n16004), .IN2(n16005), .QN(n15995) );
  INVX0 U16864 ( .INP(n16006), .ZN(n16005) );
  NAND2X0 U16865 ( .IN1(n3513), .IN2(n9124), .QN(n16006) );
  NOR2X0 U16866 ( .IN1(n9116), .IN2(n3513), .QN(n16004) );
  NAND2X0 U16867 ( .IN1(n16007), .IN2(n16008), .QN(DATA_9_22) );
  INVX0 U16868 ( .INP(n16009), .ZN(n16008) );
  NOR2X0 U16869 ( .IN1(n16010), .IN2(n11829), .QN(n16009) );
  NAND2X0 U16870 ( .IN1(n11829), .IN2(n16010), .QN(n16007) );
  NAND2X0 U16871 ( .IN1(TM0), .IN2(WX503), .QN(n16010) );
  NAND2X0 U16872 ( .IN1(n16011), .IN2(n16012), .QN(n11829) );
  NAND2X0 U16873 ( .IN1(n16013), .IN2(n16014), .QN(n16012) );
  INVX0 U16874 ( .INP(n16015), .ZN(n16011) );
  NOR2X0 U16875 ( .IN1(n16014), .IN2(n16013), .QN(n16015) );
  NAND2X0 U16876 ( .IN1(n16016), .IN2(n16017), .QN(n16013) );
  NAND2X0 U16877 ( .IN1(n8760), .IN2(n16018), .QN(n16017) );
  INVX0 U16878 ( .INP(n16019), .ZN(n16016) );
  NOR2X0 U16879 ( .IN1(n16018), .IN2(n8760), .QN(n16019) );
  NOR2X0 U16880 ( .IN1(n16020), .IN2(n16021), .QN(n16018) );
  NOR2X0 U16881 ( .IN1(WX855), .IN2(n8761), .QN(n16021) );
  INVX0 U16882 ( .INP(n16022), .ZN(n16020) );
  NAND2X0 U16883 ( .IN1(n8761), .IN2(WX855), .QN(n16022) );
  NOR2X0 U16884 ( .IN1(n16023), .IN2(n16024), .QN(n16014) );
  INVX0 U16885 ( .INP(n16025), .ZN(n16024) );
  NAND2X0 U16886 ( .IN1(n3511), .IN2(n9124), .QN(n16025) );
  NOR2X0 U16887 ( .IN1(n9116), .IN2(n3511), .QN(n16023) );
  NAND2X0 U16888 ( .IN1(n16026), .IN2(n16027), .QN(DATA_9_21) );
  INVX0 U16889 ( .INP(n16028), .ZN(n16027) );
  NOR2X0 U16890 ( .IN1(n16029), .IN2(n11818), .QN(n16028) );
  NAND2X0 U16891 ( .IN1(n11818), .IN2(n16029), .QN(n16026) );
  NAND2X0 U16892 ( .IN1(TM0), .IN2(WX505), .QN(n16029) );
  NAND2X0 U16893 ( .IN1(n16030), .IN2(n16031), .QN(n11818) );
  NAND2X0 U16894 ( .IN1(n16032), .IN2(n16033), .QN(n16031) );
  INVX0 U16895 ( .INP(n16034), .ZN(n16030) );
  NOR2X0 U16896 ( .IN1(n16033), .IN2(n16032), .QN(n16034) );
  NAND2X0 U16897 ( .IN1(n16035), .IN2(n16036), .QN(n16032) );
  NAND2X0 U16898 ( .IN1(n8766), .IN2(n16037), .QN(n16036) );
  INVX0 U16899 ( .INP(n16038), .ZN(n16035) );
  NOR2X0 U16900 ( .IN1(n16037), .IN2(n8766), .QN(n16038) );
  NOR2X0 U16901 ( .IN1(n16039), .IN2(n16040), .QN(n16037) );
  NOR2X0 U16902 ( .IN1(WX857), .IN2(n8767), .QN(n16040) );
  INVX0 U16903 ( .INP(n16041), .ZN(n16039) );
  NAND2X0 U16904 ( .IN1(n8767), .IN2(WX857), .QN(n16041) );
  NOR2X0 U16905 ( .IN1(n16042), .IN2(n16043), .QN(n16033) );
  INVX0 U16906 ( .INP(n16044), .ZN(n16043) );
  NAND2X0 U16907 ( .IN1(n3509), .IN2(n9124), .QN(n16044) );
  NOR2X0 U16908 ( .IN1(n9116), .IN2(n3509), .QN(n16042) );
  NOR2X0 U16909 ( .IN1(n16045), .IN2(n16046), .QN(DATA_9_20) );
  INVX0 U16910 ( .INP(n16047), .ZN(n16046) );
  NAND2X0 U16911 ( .IN1(n16048), .IN2(n11807), .QN(n16047) );
  NOR2X0 U16912 ( .IN1(n11807), .IN2(n16048), .QN(n16045) );
  NAND2X0 U16913 ( .IN1(TM0), .IN2(WX507), .QN(n16048) );
  NAND2X0 U16914 ( .IN1(n16049), .IN2(n16050), .QN(n11807) );
  NAND2X0 U16915 ( .IN1(n16051), .IN2(n16052), .QN(n16050) );
  NAND2X0 U16916 ( .IN1(n16053), .IN2(n16054), .QN(n16051) );
  NAND3X0 U16917 ( .IN1(n16053), .IN2(n16054), .IN3(n16055), .QN(n16049) );
  INVX0 U16918 ( .INP(n16052), .ZN(n16055) );
  NOR2X0 U16919 ( .IN1(n16056), .IN2(n16057), .QN(n16052) );
  INVX0 U16920 ( .INP(n16058), .ZN(n16057) );
  NAND2X0 U16921 ( .IN1(n8771), .IN2(n16059), .QN(n16058) );
  NOR2X0 U16922 ( .IN1(n16059), .IN2(n8771), .QN(n16056) );
  NOR2X0 U16923 ( .IN1(n16060), .IN2(n16061), .QN(n16059) );
  INVX0 U16924 ( .INP(n16062), .ZN(n16061) );
  NAND2X0 U16925 ( .IN1(test_so6), .IN2(WX731), .QN(n16062) );
  NOR2X0 U16926 ( .IN1(WX731), .IN2(test_so6), .QN(n16060) );
  NAND2X0 U16927 ( .IN1(n3507), .IN2(n9124), .QN(n16054) );
  NAND2X0 U16928 ( .IN1(TM1), .IN2(WX667), .QN(n16053) );
  NOR2X0 U16929 ( .IN1(n16063), .IN2(n16064), .QN(DATA_9_2) );
  INVX0 U16930 ( .INP(n16065), .ZN(n16064) );
  NAND2X0 U16931 ( .IN1(n16066), .IN2(n11672), .QN(n16065) );
  NOR2X0 U16932 ( .IN1(n11672), .IN2(n16066), .QN(n16063) );
  NAND2X0 U16933 ( .IN1(TM0), .IN2(WX543), .QN(n16066) );
  NAND2X0 U16934 ( .IN1(n16067), .IN2(n16068), .QN(n11672) );
  NAND2X0 U16935 ( .IN1(n16069), .IN2(n16070), .QN(n16068) );
  NAND2X0 U16936 ( .IN1(n16071), .IN2(n16072), .QN(n16069) );
  NAND3X0 U16937 ( .IN1(n16071), .IN2(n16072), .IN3(n16073), .QN(n16067) );
  INVX0 U16938 ( .INP(n16070), .ZN(n16073) );
  NOR2X0 U16939 ( .IN1(n16074), .IN2(n16075), .QN(n16070) );
  INVX0 U16940 ( .INP(n16076), .ZN(n16075) );
  NAND2X0 U16941 ( .IN1(n8779), .IN2(n16077), .QN(n16076) );
  NOR2X0 U16942 ( .IN1(n16077), .IN2(n8779), .QN(n16074) );
  NOR2X0 U16943 ( .IN1(n16078), .IN2(n16079), .QN(n16077) );
  INVX0 U16944 ( .INP(n16080), .ZN(n16079) );
  NAND2X0 U16945 ( .IN1(test_so7), .IN2(WX895), .QN(n16080) );
  NOR2X0 U16946 ( .IN1(WX895), .IN2(test_so7), .QN(n16078) );
  NAND2X0 U16947 ( .IN1(n3471), .IN2(n2183), .QN(n16072) );
  NAND2X0 U16948 ( .IN1(TM0), .IN2(WX703), .QN(n16071) );
  NAND2X0 U16949 ( .IN1(n16081), .IN2(n16082), .QN(DATA_9_19) );
  INVX0 U16950 ( .INP(n16083), .ZN(n16082) );
  NOR2X0 U16951 ( .IN1(n16084), .IN2(n11795), .QN(n16083) );
  NAND2X0 U16952 ( .IN1(n11795), .IN2(n16084), .QN(n16081) );
  NAND2X0 U16953 ( .IN1(TM0), .IN2(WX509), .QN(n16084) );
  NAND2X0 U16954 ( .IN1(n16085), .IN2(n16086), .QN(n11795) );
  NAND2X0 U16955 ( .IN1(n16087), .IN2(n16088), .QN(n16086) );
  INVX0 U16956 ( .INP(n16089), .ZN(n16085) );
  NOR2X0 U16957 ( .IN1(n16088), .IN2(n16087), .QN(n16089) );
  NAND2X0 U16958 ( .IN1(n16090), .IN2(n16091), .QN(n16087) );
  NAND2X0 U16959 ( .IN1(n8705), .IN2(n16092), .QN(n16091) );
  INVX0 U16960 ( .INP(n16093), .ZN(n16090) );
  NOR2X0 U16961 ( .IN1(n16092), .IN2(n8705), .QN(n16093) );
  NOR2X0 U16962 ( .IN1(n16094), .IN2(n16095), .QN(n16092) );
  INVX0 U16963 ( .INP(n16096), .ZN(n16095) );
  NAND2X0 U16964 ( .IN1(n8707), .IN2(WX861), .QN(n16096) );
  NOR2X0 U16965 ( .IN1(WX861), .IN2(n8707), .QN(n16094) );
  NOR2X0 U16966 ( .IN1(n16097), .IN2(n16098), .QN(n16088) );
  INVX0 U16967 ( .INP(n16099), .ZN(n16098) );
  NAND2X0 U16968 ( .IN1(n3505), .IN2(n9124), .QN(n16099) );
  NOR2X0 U16969 ( .IN1(n9116), .IN2(n3505), .QN(n16097) );
  NAND2X0 U16970 ( .IN1(n16100), .IN2(n16101), .QN(DATA_9_18) );
  INVX0 U16971 ( .INP(n16102), .ZN(n16101) );
  NOR2X0 U16972 ( .IN1(n16103), .IN2(n11784), .QN(n16102) );
  NAND2X0 U16973 ( .IN1(n11784), .IN2(n16103), .QN(n16100) );
  NAND2X0 U16974 ( .IN1(TM0), .IN2(WX511), .QN(n16103) );
  NAND2X0 U16975 ( .IN1(n16104), .IN2(n16105), .QN(n11784) );
  NAND2X0 U16976 ( .IN1(n16106), .IN2(n16107), .QN(n16105) );
  INVX0 U16977 ( .INP(n16108), .ZN(n16104) );
  NOR2X0 U16978 ( .IN1(n16107), .IN2(n16106), .QN(n16108) );
  NAND2X0 U16979 ( .IN1(n16109), .IN2(n16110), .QN(n16106) );
  NAND2X0 U16980 ( .IN1(n8720), .IN2(n16111), .QN(n16110) );
  INVX0 U16981 ( .INP(n16112), .ZN(n16109) );
  NOR2X0 U16982 ( .IN1(n16111), .IN2(n8720), .QN(n16112) );
  NOR2X0 U16983 ( .IN1(n16113), .IN2(n16114), .QN(n16111) );
  INVX0 U16984 ( .INP(n16115), .ZN(n16114) );
  NAND2X0 U16985 ( .IN1(n8722), .IN2(WX863), .QN(n16115) );
  NOR2X0 U16986 ( .IN1(WX863), .IN2(n8722), .QN(n16113) );
  NOR2X0 U16987 ( .IN1(n16116), .IN2(n16117), .QN(n16107) );
  INVX0 U16988 ( .INP(n16118), .ZN(n16117) );
  NAND2X0 U16989 ( .IN1(n3503), .IN2(n9124), .QN(n16118) );
  NOR2X0 U16990 ( .IN1(n9116), .IN2(n3503), .QN(n16116) );
  NAND2X0 U16991 ( .IN1(n16119), .IN2(n16120), .QN(DATA_9_17) );
  INVX0 U16992 ( .INP(n16121), .ZN(n16120) );
  NOR2X0 U16993 ( .IN1(n16122), .IN2(n11778), .QN(n16121) );
  NAND2X0 U16994 ( .IN1(n11778), .IN2(n16122), .QN(n16119) );
  NAND2X0 U16995 ( .IN1(TM0), .IN2(WX513), .QN(n16122) );
  NAND2X0 U16996 ( .IN1(n16123), .IN2(n16124), .QN(n11778) );
  NAND2X0 U16997 ( .IN1(n16125), .IN2(n16126), .QN(n16124) );
  INVX0 U16998 ( .INP(n16127), .ZN(n16123) );
  NOR2X0 U16999 ( .IN1(n16126), .IN2(n16125), .QN(n16127) );
  NAND2X0 U17000 ( .IN1(n16128), .IN2(n16129), .QN(n16125) );
  NAND2X0 U17001 ( .IN1(n8732), .IN2(n16130), .QN(n16129) );
  INVX0 U17002 ( .INP(n16131), .ZN(n16128) );
  NOR2X0 U17003 ( .IN1(n16130), .IN2(n8732), .QN(n16131) );
  NOR2X0 U17004 ( .IN1(n16132), .IN2(n16133), .QN(n16130) );
  INVX0 U17005 ( .INP(n16134), .ZN(n16133) );
  NAND2X0 U17006 ( .IN1(n8734), .IN2(WX865), .QN(n16134) );
  NOR2X0 U17007 ( .IN1(WX865), .IN2(n8734), .QN(n16132) );
  NOR2X0 U17008 ( .IN1(n16135), .IN2(n16136), .QN(n16126) );
  INVX0 U17009 ( .INP(n16137), .ZN(n16136) );
  NAND2X0 U17010 ( .IN1(n3501), .IN2(n9124), .QN(n16137) );
  NOR2X0 U17011 ( .IN1(n9116), .IN2(n3501), .QN(n16135) );
  NOR2X0 U17012 ( .IN1(n16138), .IN2(n16139), .QN(DATA_9_16) );
  INVX0 U17013 ( .INP(n16140), .ZN(n16139) );
  NAND2X0 U17014 ( .IN1(n16141), .IN2(n11767), .QN(n16140) );
  NOR2X0 U17015 ( .IN1(n11767), .IN2(n16141), .QN(n16138) );
  NAND2X0 U17016 ( .IN1(TM0), .IN2(WX515), .QN(n16141) );
  NAND2X0 U17017 ( .IN1(n16142), .IN2(n16143), .QN(n11767) );
  NAND2X0 U17018 ( .IN1(n16144), .IN2(n16145), .QN(n16143) );
  NAND2X0 U17019 ( .IN1(n16146), .IN2(n16147), .QN(n16144) );
  NAND3X0 U17020 ( .IN1(n16146), .IN2(n16147), .IN3(n16148), .QN(n16142) );
  INVX0 U17021 ( .INP(n16145), .ZN(n16148) );
  NOR2X0 U17022 ( .IN1(n16149), .IN2(n16150), .QN(n16145) );
  INVX0 U17023 ( .INP(n16151), .ZN(n16150) );
  NAND2X0 U17024 ( .IN1(n8749), .IN2(n16152), .QN(n16151) );
  NOR2X0 U17025 ( .IN1(n16152), .IN2(n8749), .QN(n16149) );
  NOR2X0 U17026 ( .IN1(n16153), .IN2(n16154), .QN(n16152) );
  NOR2X0 U17027 ( .IN1(n8798), .IN2(n8750), .QN(n16154) );
  INVX0 U17028 ( .INP(n16155), .ZN(n16153) );
  NAND2X0 U17029 ( .IN1(n8750), .IN2(n8798), .QN(n16155) );
  NAND2X0 U17030 ( .IN1(n3499), .IN2(n9118), .QN(n16147) );
  INVX0 U17031 ( .INP(TM1), .ZN(n10633) );
  NAND2X0 U17032 ( .IN1(TM1), .IN2(WX675), .QN(n16146) );
  NAND2X0 U17033 ( .IN1(n16156), .IN2(n16157), .QN(DATA_9_15) );
  INVX0 U17034 ( .INP(n16158), .ZN(n16157) );
  NOR2X0 U17035 ( .IN1(n16159), .IN2(n11755), .QN(n16158) );
  NAND2X0 U17036 ( .IN1(n11755), .IN2(n16159), .QN(n16156) );
  NAND2X0 U17037 ( .IN1(TM0), .IN2(WX517), .QN(n16159) );
  NAND2X0 U17038 ( .IN1(n16160), .IN2(n16161), .QN(n11755) );
  NAND2X0 U17039 ( .IN1(n16162), .IN2(n16163), .QN(n16161) );
  INVX0 U17040 ( .INP(n16164), .ZN(n16160) );
  NOR2X0 U17041 ( .IN1(n16163), .IN2(n16162), .QN(n16164) );
  NAND2X0 U17042 ( .IN1(n16165), .IN2(n16166), .QN(n16162) );
  NAND2X0 U17043 ( .IN1(n8763), .IN2(n16167), .QN(n16166) );
  INVX0 U17044 ( .INP(n16168), .ZN(n16165) );
  NOR2X0 U17045 ( .IN1(n16167), .IN2(n8763), .QN(n16168) );
  NOR2X0 U17046 ( .IN1(n16169), .IN2(n16170), .QN(n16167) );
  NOR2X0 U17047 ( .IN1(WX869), .IN2(n8764), .QN(n16170) );
  INVX0 U17048 ( .INP(n16171), .ZN(n16169) );
  NAND2X0 U17049 ( .IN1(n8764), .IN2(WX869), .QN(n16171) );
  NOR2X0 U17050 ( .IN1(n16172), .IN2(n16173), .QN(n16163) );
  INVX0 U17051 ( .INP(n16174), .ZN(n16173) );
  NAND2X0 U17052 ( .IN1(n3497), .IN2(n2183), .QN(n16174) );
  NOR2X0 U17053 ( .IN1(n2183), .IN2(n3497), .QN(n16172) );
  NAND2X0 U17054 ( .IN1(n16175), .IN2(n16176), .QN(DATA_9_14) );
  INVX0 U17055 ( .INP(n16177), .ZN(n16176) );
  NOR2X0 U17056 ( .IN1(n16178), .IN2(n11749), .QN(n16177) );
  NAND2X0 U17057 ( .IN1(n11749), .IN2(n16178), .QN(n16175) );
  NAND2X0 U17058 ( .IN1(test_so1), .IN2(TM0), .QN(n16178) );
  NAND2X0 U17059 ( .IN1(n16179), .IN2(n16180), .QN(n11749) );
  NAND2X0 U17060 ( .IN1(n16181), .IN2(n16182), .QN(n16180) );
  INVX0 U17061 ( .INP(n16183), .ZN(n16179) );
  NOR2X0 U17062 ( .IN1(n16182), .IN2(n16181), .QN(n16183) );
  NAND2X0 U17063 ( .IN1(n16184), .IN2(n16185), .QN(n16181) );
  NAND2X0 U17064 ( .IN1(n8776), .IN2(n16186), .QN(n16185) );
  INVX0 U17065 ( .INP(n16187), .ZN(n16184) );
  NOR2X0 U17066 ( .IN1(n16186), .IN2(n8776), .QN(n16187) );
  NOR2X0 U17067 ( .IN1(n16188), .IN2(n16189), .QN(n16186) );
  INVX0 U17068 ( .INP(n16190), .ZN(n16189) );
  NAND2X0 U17069 ( .IN1(n8778), .IN2(WX871), .QN(n16190) );
  NOR2X0 U17070 ( .IN1(WX871), .IN2(n8778), .QN(n16188) );
  NOR2X0 U17071 ( .IN1(n16191), .IN2(n16192), .QN(n16182) );
  INVX0 U17072 ( .INP(n16193), .ZN(n16192) );
  NAND2X0 U17073 ( .IN1(n3495), .IN2(n2183), .QN(n16193) );
  NOR2X0 U17074 ( .IN1(n2183), .IN2(n3495), .QN(n16191) );
  NAND2X0 U17075 ( .IN1(n16194), .IN2(n16195), .QN(DATA_9_13) );
  INVX0 U17076 ( .INP(n16196), .ZN(n16195) );
  NOR2X0 U17077 ( .IN1(n16197), .IN2(n11742), .QN(n16196) );
  NAND2X0 U17078 ( .IN1(n11742), .IN2(n16197), .QN(n16194) );
  NAND2X0 U17079 ( .IN1(TM0), .IN2(WX521), .QN(n16197) );
  NAND2X0 U17080 ( .IN1(n16198), .IN2(n16199), .QN(n11742) );
  NAND2X0 U17081 ( .IN1(n16200), .IN2(n16201), .QN(n16199) );
  INVX0 U17082 ( .INP(n16202), .ZN(n16198) );
  NOR2X0 U17083 ( .IN1(n16201), .IN2(n16200), .QN(n16202) );
  NAND2X0 U17084 ( .IN1(n16203), .IN2(n16204), .QN(n16200) );
  NAND2X0 U17085 ( .IN1(n8711), .IN2(n16205), .QN(n16204) );
  INVX0 U17086 ( .INP(n16206), .ZN(n16203) );
  NOR2X0 U17087 ( .IN1(n16205), .IN2(n8711), .QN(n16206) );
  NOR2X0 U17088 ( .IN1(n16207), .IN2(n16208), .QN(n16205) );
  INVX0 U17089 ( .INP(n16209), .ZN(n16208) );
  NAND2X0 U17090 ( .IN1(n8713), .IN2(WX873), .QN(n16209) );
  NOR2X0 U17091 ( .IN1(WX873), .IN2(n8713), .QN(n16207) );
  NOR2X0 U17092 ( .IN1(n16210), .IN2(n16211), .QN(n16201) );
  INVX0 U17093 ( .INP(n16212), .ZN(n16211) );
  NAND2X0 U17094 ( .IN1(n3493), .IN2(n2183), .QN(n16212) );
  NOR2X0 U17095 ( .IN1(n2183), .IN2(n3493), .QN(n16210) );
  NAND2X0 U17096 ( .IN1(n16213), .IN2(n16214), .QN(DATA_9_12) );
  INVX0 U17097 ( .INP(n16215), .ZN(n16214) );
  NOR2X0 U17098 ( .IN1(n16216), .IN2(n11736), .QN(n16215) );
  NAND2X0 U17099 ( .IN1(n11736), .IN2(n16216), .QN(n16213) );
  NAND2X0 U17100 ( .IN1(TM0), .IN2(WX523), .QN(n16216) );
  NAND2X0 U17101 ( .IN1(n16217), .IN2(n16218), .QN(n11736) );
  NAND2X0 U17102 ( .IN1(n16219), .IN2(n16220), .QN(n16218) );
  INVX0 U17103 ( .INP(n16221), .ZN(n16217) );
  NOR2X0 U17104 ( .IN1(n16220), .IN2(n16219), .QN(n16221) );
  NAND2X0 U17105 ( .IN1(n16222), .IN2(n16223), .QN(n16219) );
  NAND2X0 U17106 ( .IN1(n8738), .IN2(n16224), .QN(n16223) );
  INVX0 U17107 ( .INP(n16225), .ZN(n16222) );
  NOR2X0 U17108 ( .IN1(n16224), .IN2(n8738), .QN(n16225) );
  NOR2X0 U17109 ( .IN1(n16226), .IN2(n16227), .QN(n16224) );
  INVX0 U17110 ( .INP(n16228), .ZN(n16227) );
  NAND2X0 U17111 ( .IN1(n8740), .IN2(WX875), .QN(n16228) );
  NOR2X0 U17112 ( .IN1(WX875), .IN2(n8740), .QN(n16226) );
  NOR2X0 U17113 ( .IN1(n16229), .IN2(n16230), .QN(n16220) );
  INVX0 U17114 ( .INP(n16231), .ZN(n16230) );
  NAND2X0 U17115 ( .IN1(n3491), .IN2(n2183), .QN(n16231) );
  NOR2X0 U17116 ( .IN1(n2183), .IN2(n3491), .QN(n16229) );
  NAND2X0 U17117 ( .IN1(n16232), .IN2(n16233), .QN(DATA_9_11) );
  INVX0 U17118 ( .INP(n16234), .ZN(n16233) );
  NOR2X0 U17119 ( .IN1(n16235), .IN2(n11730), .QN(n16234) );
  NAND2X0 U17120 ( .IN1(n11730), .IN2(n16235), .QN(n16232) );
  NAND2X0 U17121 ( .IN1(TM0), .IN2(WX525), .QN(n16235) );
  NAND2X0 U17122 ( .IN1(n16236), .IN2(n16237), .QN(n11730) );
  NAND2X0 U17123 ( .IN1(n16238), .IN2(n16239), .QN(n16237) );
  INVX0 U17124 ( .INP(n16240), .ZN(n16236) );
  NOR2X0 U17125 ( .IN1(n16239), .IN2(n16238), .QN(n16240) );
  NAND2X0 U17126 ( .IN1(n16241), .IN2(n16242), .QN(n16238) );
  NAND2X0 U17127 ( .IN1(n8784), .IN2(n16243), .QN(n16242) );
  INVX0 U17128 ( .INP(n16244), .ZN(n16241) );
  NOR2X0 U17129 ( .IN1(n16243), .IN2(n8784), .QN(n16244) );
  NOR2X0 U17130 ( .IN1(n16245), .IN2(n16246), .QN(n16243) );
  INVX0 U17131 ( .INP(n16247), .ZN(n16246) );
  NAND2X0 U17132 ( .IN1(n8786), .IN2(WX877), .QN(n16247) );
  NOR2X0 U17133 ( .IN1(WX877), .IN2(n8786), .QN(n16245) );
  NOR2X0 U17134 ( .IN1(n16248), .IN2(n16249), .QN(n16239) );
  INVX0 U17135 ( .INP(n16250), .ZN(n16249) );
  NAND2X0 U17136 ( .IN1(n3489), .IN2(n2183), .QN(n16250) );
  NOR2X0 U17137 ( .IN1(n2183), .IN2(n3489), .QN(n16248) );
  NOR2X0 U17138 ( .IN1(n16251), .IN2(n16252), .QN(DATA_9_10) );
  INVX0 U17139 ( .INP(n16253), .ZN(n16252) );
  NAND2X0 U17140 ( .IN1(n16254), .IN2(n11724), .QN(n16253) );
  NOR2X0 U17141 ( .IN1(n11724), .IN2(n16254), .QN(n16251) );
  NAND2X0 U17142 ( .IN1(TM0), .IN2(WX527), .QN(n16254) );
  NAND2X0 U17143 ( .IN1(n16255), .IN2(n16256), .QN(n11724) );
  NAND2X0 U17144 ( .IN1(n16257), .IN2(n16258), .QN(n16256) );
  NAND2X0 U17145 ( .IN1(n16259), .IN2(n16260), .QN(n16257) );
  NAND3X0 U17146 ( .IN1(n16259), .IN2(n16260), .IN3(n16261), .QN(n16255) );
  INVX0 U17147 ( .INP(n16258), .ZN(n16261) );
  NOR2X0 U17148 ( .IN1(n16262), .IN2(n16263), .QN(n16258) );
  INVX0 U17149 ( .INP(n16264), .ZN(n16263) );
  NAND2X0 U17150 ( .IN1(n8729), .IN2(n16265), .QN(n16264) );
  NOR2X0 U17151 ( .IN1(n16265), .IN2(n8729), .QN(n16262) );
  NOR2X0 U17152 ( .IN1(n16266), .IN2(n16267), .QN(n16265) );
  INVX0 U17153 ( .INP(n16268), .ZN(n16267) );
  NAND2X0 U17154 ( .IN1(test_so3), .IN2(WX879), .QN(n16268) );
  NOR2X0 U17155 ( .IN1(WX879), .IN2(test_so3), .QN(n16266) );
  NAND2X0 U17156 ( .IN1(n8731), .IN2(n2183), .QN(n16260) );
  NAND2X0 U17157 ( .IN1(TM0), .IN2(WX751), .QN(n16259) );
  NAND2X0 U17158 ( .IN1(n16269), .IN2(n16270), .QN(DATA_9_1) );
  INVX0 U17159 ( .INP(n16271), .ZN(n16270) );
  NOR2X0 U17160 ( .IN1(n16272), .IN2(n11665), .QN(n16271) );
  NAND2X0 U17161 ( .IN1(n11665), .IN2(n16272), .QN(n16269) );
  NAND2X0 U17162 ( .IN1(TM0), .IN2(WX545), .QN(n16272) );
  NAND2X0 U17163 ( .IN1(n16273), .IN2(n16274), .QN(n11665) );
  NAND2X0 U17164 ( .IN1(n16275), .IN2(n16276), .QN(n16274) );
  INVX0 U17165 ( .INP(n16277), .ZN(n16273) );
  NOR2X0 U17166 ( .IN1(n16276), .IN2(n16275), .QN(n16277) );
  NAND2X0 U17167 ( .IN1(n16278), .IN2(n16279), .QN(n16275) );
  NAND2X0 U17168 ( .IN1(n8714), .IN2(n16280), .QN(n16279) );
  INVX0 U17169 ( .INP(n16281), .ZN(n16280) );
  NAND2X0 U17170 ( .IN1(n16281), .IN2(WX897), .QN(n16278) );
  NAND2X0 U17171 ( .IN1(n16282), .IN2(n16283), .QN(n16281) );
  INVX0 U17172 ( .INP(n16284), .ZN(n16283) );
  NOR2X0 U17173 ( .IN1(WX833), .IN2(n8715), .QN(n16284) );
  NAND2X0 U17174 ( .IN1(n8715), .IN2(WX833), .QN(n16282) );
  NOR2X0 U17175 ( .IN1(n16285), .IN2(n16286), .QN(n16276) );
  INVX0 U17176 ( .INP(n16287), .ZN(n16286) );
  NAND2X0 U17177 ( .IN1(n3469), .IN2(n2183), .QN(n16287) );
  NOR2X0 U17178 ( .IN1(n2183), .IN2(n3469), .QN(n16285) );
  NAND2X0 U17179 ( .IN1(n16288), .IN2(n16289), .QN(DATA_9_0) );
  INVX0 U17180 ( .INP(n16290), .ZN(n16289) );
  NOR2X0 U17181 ( .IN1(n16291), .IN2(n11659), .QN(n16290) );
  NAND2X0 U17182 ( .IN1(n11659), .IN2(n16291), .QN(n16288) );
  NAND2X0 U17183 ( .IN1(TM0), .IN2(WX547), .QN(n16291) );
  NAND2X0 U17184 ( .IN1(n16292), .IN2(n16293), .QN(n11659) );
  NAND2X0 U17185 ( .IN1(n16294), .IN2(n16295), .QN(n16293) );
  INVX0 U17186 ( .INP(n16296), .ZN(n16292) );
  NOR2X0 U17187 ( .IN1(n16295), .IN2(n16294), .QN(n16296) );
  NAND2X0 U17188 ( .IN1(n16297), .IN2(n16298), .QN(n16294) );
  NAND2X0 U17189 ( .IN1(n8787), .IN2(n16299), .QN(n16298) );
  INVX0 U17190 ( .INP(n16300), .ZN(n16297) );
  NOR2X0 U17191 ( .IN1(n16299), .IN2(n8787), .QN(n16300) );
  NOR2X0 U17192 ( .IN1(n16301), .IN2(n16302), .QN(n16299) );
  NOR2X0 U17193 ( .IN1(WX899), .IN2(n8788), .QN(n16302) );
  INVX0 U17194 ( .INP(n16303), .ZN(n16301) );
  NAND2X0 U17195 ( .IN1(n8788), .IN2(WX899), .QN(n16303) );
  NOR2X0 U17196 ( .IN1(n16304), .IN2(n16305), .QN(n16295) );
  INVX0 U17197 ( .INP(n16306), .ZN(n16305) );
  NAND2X0 U17198 ( .IN1(n3467), .IN2(n2183), .QN(n16306) );
  NOR2X0 U17199 ( .IN1(n2183), .IN2(n3467), .QN(n16304) );
  INVX0 U17200 ( .INP(TM0), .ZN(n2183) );
  NOR2X0 U3558_U2 ( .IN1(n9180), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n9273), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n2183), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n9180), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n9180), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n9204), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n9198), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n9192), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n9192), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n9192), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n9192), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n9192), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n9192), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n9192), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n9192), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n9193), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n9193), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n9193), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n9193), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n9193), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n9193), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n9193), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n9193), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n9193), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n9193), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n9193), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n9193), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n9193), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n9194), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n9194), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n9194), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n9194), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n9194), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n9194), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n9194), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n9194), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n9194), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n9194), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n9194), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n9194), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n9194), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n9195), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n9195), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n9195), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n9195), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n9195), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n9195), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n9195), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n9195), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n9195), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n9195), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n9195), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n9195), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n9195), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n9196), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n9196), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n9196), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n9196), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n9196), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n9196), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n9196), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n9196), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n9196), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n9196), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n9196), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n9196), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n9196), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n9197), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n9197), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n9197), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n9197), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n9197), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n9197), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n9197), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n9197), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n9197), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n9197), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n9197), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n9197), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n9197), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n9198), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n9198), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n9198), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n9198), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n9198), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n9198), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n9198), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n9198), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n9198), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n9198), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n9198), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n9198), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n9199), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n9199), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n9199), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n9199), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n9199), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n9199), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n9199), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n9199), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n9199), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n9199), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n9199), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n9199), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n9199), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n9200), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n9200), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n9200), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n9200), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n9200), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n9200), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n9200), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n9200), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n9200), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n9200), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n9200), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n9200), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n9200), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n9201), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n9201), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n9201), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n9201), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n9201), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n9201), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n9201), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n9201), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n9201), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n9201), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n9201), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n9201), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n9201), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n9202), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n9202), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n9202), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n9202), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n9202), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n9202), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n9202), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n9202), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n9202), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n9202), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n9202), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n9202), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n9202), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n9203), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n9203), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n9203), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n9203), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n9203), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n9203), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n9203), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n9203), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n9203), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n9203), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n9203), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n9203), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n9203), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n9204), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n9204), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n9204), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n9204), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n9204), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n9204), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n9186), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n9180), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n9180), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n9180), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n9180), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n9180), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n9180), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n9180), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n9180), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n9180), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n9180), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n9181), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n9181), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n9181), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n9181), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n9181), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n9181), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n9181), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n9181), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n9181), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n9181), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n9181), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n9181), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n9181), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n9182), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n9182), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n9182), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n9182), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n9182), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n9182), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n9182), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n9182), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n9182), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n9182), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n9182), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n9182), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n9182), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n9183), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n9183), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n9183), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n9183), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n9183), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n9183), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n9183), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n9183), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n9183), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n9183), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n9183), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n9183), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n9183), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n9184), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n9184), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n9184), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n9184), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n9184), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n9184), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n9184), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n9184), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n9184), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n9184), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n9184), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n9184), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n9184), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n9185), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n9185), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n9185), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n9185), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n9185), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n9185), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n9185), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n9185), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n9185), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n9185), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n9185), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n9185), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n9185), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n9186), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n9186), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n9186), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n9186), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n9186), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n9186), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n9186), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n9186), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n9186), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n9186), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n9186), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n9186), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n9187), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n9187), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n9187), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n9187), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n9187), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n9187), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n9187), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n9187), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n9187), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n9187), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n9187), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n9187), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n9187), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n9188), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n9188), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n9188), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n9188), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n9188), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n9188), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n9188), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n9188), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n9188), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n9188), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n9188), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n9188), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n9188), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n9189), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n9189), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n9189), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n9189), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n9189), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n9189), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n9189), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n9189), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n9189), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n9189), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n9189), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n9189), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n9189), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n9190), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n9190), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n9190), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n9190), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n9190), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n9190), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n9190), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n9190), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n9190), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n9190), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n9190), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n9190), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n9190), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n9191), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n9191), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n9191), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n9191), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n9191), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n9191), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n9191), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n9191), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n9191), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n9191), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n9191), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n9191), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n9191), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n9192), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n9192), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n9192), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n9192), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n9192), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n9222), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n9224), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n9223), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n9222), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n9222), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n9223), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n9223), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n9222), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n9221), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n9221), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n9221), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n9221), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n9221), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n9220), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n9220), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n9221), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n9220), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n9220), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n9223), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n9223), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n9223), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n9223), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n9223), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n9223), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n9223), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n9222), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n9222), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n9223), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n9222), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n9222), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n9220), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n9221), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n9221), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n9221), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n9220), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n9222), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n9222), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n9221), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n9222), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n9222), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n9221), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n9223), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n9222), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n9224), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n9223), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n9221), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n9221), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n9220), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n9220), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n9220), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n9220), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n9219), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n9220), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n9220), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n9220), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n9219), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n9212), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n9204), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n9204), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n9204), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n9204), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n9204), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n9204), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n9205), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n9205), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n9205), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n9205), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n9205), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n9205), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n9205), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n9205), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n9205), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n9205), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n9205), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n9205), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n9205), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n9206), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n9206), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n9206), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n9206), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n9206), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n9206), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n9206), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n9206), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n9206), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n9206), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n9206), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n9206), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n9206), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n9207), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n9207), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n9207), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n9207), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n9207), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n9219), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n9207), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n9207), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n9207), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n9207), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n9207), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n9207), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n9207), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n9208), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n9208), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n9208), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n9208), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n9208), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n9208), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n9208), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n9208), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n9208), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n9208), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n9208), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n9208), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n9208), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n9209), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n9209), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n9209), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n9209), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n9209), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n9209), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n9209), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n9209), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n9209), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n9209), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n9209), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n9209), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n9209), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n9210), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n9210), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n9210), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n9210), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n9210), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n9210), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n9210), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n9210), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n9210), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n9210), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n9210), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n9210), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n9210), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n9211), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n9211), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n9211), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n9211), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n9211), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n9211), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n9211), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n9211), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n9211), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n9211), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n9211), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n9211), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n9211), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n9212), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n9219), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n9219), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n9219), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n9219), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n9219), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n9219), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n9219), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n9219), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n9219), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n9219), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n9218), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n9218), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n9218), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n9218), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n9218), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n9218), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n9218), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n9218), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n9218), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n9218), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n9218), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n9218), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n9218), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n9217), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n9217), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n9217), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n9217), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n9217), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n9217), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n9217), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n9217), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n9217), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n9217), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n9217), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n9217), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n9217), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n9216), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n9216), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n9216), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n9216), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n9216), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n9216), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n9216), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n9216), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n9216), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n9216), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n9216), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n9216), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n9216), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n9215), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n9215), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n9215), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n9215), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n9215), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n9215), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n9215), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n9215), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n9215), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n9215), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n9215), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n9215), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n9214), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n9214), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n9214), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n9214), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n9214), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n9214), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n9214), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n9214), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n9214), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n9214), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n9214), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n9214), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n9214), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n9213), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n9213), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n9213), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n9213), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n9213), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n9213), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n9213), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n9213), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n9213), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n9213), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n9213), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n9213), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n9213), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n9212), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n9212), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n9212), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n9212), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n9212), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n9212), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n9212), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n9212), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n9212), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n9212), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n9212), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n9215), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n9207), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n9165), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n9172), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n9172), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n9172), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n9172), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n9172), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n9172), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n9172), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n9171), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n9171), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n9171), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n9171), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n9171), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n9171), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n9171), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n9171), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n9171), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n9171), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n9171), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n9171), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n9171), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n9170), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n9170), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n9170), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n9170), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n9170), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n9170), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n9170), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n9170), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n9170), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n9170), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n9170), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n9170), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n9170), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n9169), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n9169), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n9169), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n9169), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n9169), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n9169), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n9169), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n9169), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n9169), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n9169), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n9169), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n9169), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n9169), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n9168), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n9168), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n9168), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n9168), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n9168), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n9168), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n9168), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n9168), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n9168), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n9168), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n9168), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n9168), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n9167), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n9167), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n9167), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n9167), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n9167), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n9167), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n9167), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n9167), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n9167), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n9167), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n9167), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n9172), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n9167), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n9166), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n9167), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n9166), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n9166), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n9166), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n9166), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n9166), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n9166), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n9166), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n9166), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n9166), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n9166), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n9166), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n9166), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n9165), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n9165), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n9165), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n9165), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n9165), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n9165), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n9165), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n9165), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n9165), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n9165), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n9165), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n9168), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n9172), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n9172), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n9172), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n9172), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n9172), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n9173), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n9173), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n9173), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n9173), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n9173), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n9173), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n9173), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n9173), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n9173), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n9173), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n9173), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n9173), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n9173), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n9174), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n9174), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n9174), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n9174), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n9174), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n9174), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n9174), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n9174), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n9174), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n9174), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n9174), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n9174), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n9174), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n9175), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n9175), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n9175), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n9175), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n9175), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n9175), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n9175), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n9175), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n9175), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n9175), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n9175), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n9175), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n9175), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n9176), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n9176), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n9176), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n9176), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n9176), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n9176), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n9176), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n9176), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n9176), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n9176), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n9176), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n9176), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n9176), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n9177), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n9177), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n9177), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n9177), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n9177), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n9177), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n9177), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n9177), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n9177), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n9177), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n9177), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n9177), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n9177), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n9178), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n9178), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n9178), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n9178), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n9178), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n9178), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n9178), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n9178), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n9178), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n9178), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n9178), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n9178), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n9178), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n9179), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n9179), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n9179), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n9179), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n9179), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n9179), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n9179), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n9179), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n9179), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n9179), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n9179), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n9179), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n9179), .IN2(U6482_n1), .QN(WX708) );
endmodule

