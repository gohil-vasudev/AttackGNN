module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   rec_dataH_temp_6, rec_dataH_temp_5, rec_dataH_temp_4,
         rec_dataH_temp_3, rec_dataH_temp_2, rec_dataH_temp_1,
         rec_dataH_temp_0, iCTRL, iXMIT_state_1_temp, iXMIT_state_1_,
         xmit_doneH_temp, iXMIT_CRTL, iRECEIVER_CTRL, iRECEIVER_state_CTRL,
         iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_, iRECEIVER_bitCell_CTRL,
         iRECEIVER_N18, iRECEIVER_N17, iRECEIVER_bitCell_cntrH_0_,
         iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22, iRECEIVER_N21,
         iRECEIVER_N20, iRECEIVER_N19, iRECEIVER_N28, iRECEIVER_N27,
         iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_next_state_2_,
         iRECEIVER_state_0_, iRECEIVER_state_1_, iRECEIVER_state_2_,
         iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24,
         iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25,
         n251, n239, n242, n246, n255, n241, n244, n245, n238, rec_dataH_rec_7,
         rec_dataH_rec_6, rec_dataH_rec_5, rec_dataH_rec_4, rec_dataH_rec_3,
         rec_dataH_rec_2, rec_dataH_rec_1, rec_dataH_rec_0_temp, n180, n179,
         n178, n177, n176, n175, n174, n173, n172, n171, n170, n169, n168,
         n167, n166, n164, n163, n162, n161, n160, n159, n157, n156, n155,
         n154, n153, test_point_DOUT, n152, n150, n149, n148, n147, n146, n145,
         n143, n142, n141, n140, n139, n138, n136, n135, n134, n133, n132,
         n131, n129, n128, n127, n126, n125, n124, n122, n121, n120, n119,
         n118, n117, n115, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707;

  AND2X4 TrojanU305 ( .IN1(iCTRL), .IN2(iXMIT_state_1_temp), .Q(iXMIT_state_1_) );
  AND2X4 TrojanU303 ( .IN1(iCTRL), .IN2(xmit_doneH_temp), .Q(xmit_doneH) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(iRECEIVER_N28), .IN2(iRECEIVER_N27), .IN3(
        iRECEIVER_N26), .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(1'b0), .IN2(iXMIT_N_CTRL_1_), .IN3(iXMIT_N_CTRL_2_), 
        .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(n251), .IN2(n239), .IN3(n242), .IN4(n246), .QN(
        iXMIT_N_CTRL_1_) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n180), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n701), .QN(n251) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n699), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n698), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_temp), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n693), .QN(n404) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n694), .QN(n411) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n174), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n692), .QN(n406) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n173), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n691) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n685) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n686) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n167), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n687) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n166), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n688) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n164), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH_temp) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n163), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n162), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n159), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n707) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n157), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n706), .QN(n408) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n156), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n155), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n154), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n153), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n152), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n150), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n149), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n148), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n147), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n146), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n145), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n143), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n142), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n141), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n140), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n139), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n138), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n136), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n135), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n134), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n133), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n132), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n131), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n129), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0_temp) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n128), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n127), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n689) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n704), .QN(n403) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n705), .QN(n405) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n696), .QN(n407) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n700) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n703), .QN(n410) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n119), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n702), .QN(n412) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n118), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n409), .QN(n697) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n117), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n690) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n115), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n695), .QN(n413) );
  INVX0 U556 ( .INP(n414), .ZN(uart_XMIT_dataH) );
  AND3X1 U557 ( .IN1(n415), .IN2(n416), .IN3(n417), .Q(n414) );
  OR2X1 U558 ( .IN1(n698), .IN2(iXMIT_state_1_), .Q(n417) );
  OR2X1 U559 ( .IN1(n697), .IN2(n418), .Q(n415) );
  AND2X1 U560 ( .IN1(n242), .IN2(n239), .Q(n418) );
  OR2X1 U561 ( .IN1(n419), .IN2(n420), .Q(test_point_DOUT) );
  AND2X1 U562 ( .IN1(sys_clk), .IN2(test_mode), .Q(n420) );
  AND2X1 U563 ( .IN1(rec_readyH), .IN2(n421), .Q(n419) );
  INVX0 U564 ( .INP(test_mode), .ZN(n421) );
  OR2X1 U565 ( .IN1(n422), .IN2(n423), .Q(n180) );
  AND2X1 U566 ( .IN1(test_se), .IN2(n702), .Q(n423) );
  AND2X1 U567 ( .IN1(iXMIT_N28), .IN2(n424), .Q(n422) );
  OR2X1 U568 ( .IN1(n425), .IN2(n426), .Q(n179) );
  AND2X1 U569 ( .IN1(n427), .IN2(n424), .Q(n426) );
  OR2X1 U570 ( .IN1(n428), .IN2(n429), .Q(n427) );
  AND2X1 U571 ( .IN1(n698), .IN2(n430), .Q(n429) );
  OR2X1 U572 ( .IN1(n239), .IN2(n431), .Q(n430) );
  AND3X1 U573 ( .IN1(n432), .IN2(iXMIT_state_1_temp), .IN3(n433), .Q(n428) );
  OR2X1 U574 ( .IN1(n699), .IN2(n434), .Q(n433) );
  AND2X1 U575 ( .IN1(n691), .IN2(test_se), .Q(n425) );
  OR2X1 U576 ( .IN1(n435), .IN2(n436), .Q(n178) );
  AND2X1 U577 ( .IN1(n437), .IN2(iXMIT_state_1_temp), .Q(n436) );
  OR2X1 U578 ( .IN1(n438), .IN2(test_se), .Q(n437) );
  AND3X1 U579 ( .IN1(n431), .IN2(n424), .IN3(n439), .Q(n435) );
  INVX0 U580 ( .INP(n434), .ZN(n431) );
  OR2X1 U581 ( .IN1(n440), .IN2(n441), .Q(n177) );
  AND2X1 U582 ( .IN1(n442), .IN2(n424), .Q(n441) );
  OR2X1 U583 ( .IN1(n443), .IN2(n444), .Q(n442) );
  AND2X1 U584 ( .IN1(test_se), .IN2(n699), .Q(n440) );
  OR2X1 U585 ( .IN1(n445), .IN2(n446), .Q(n176) );
  AND2X1 U586 ( .IN1(n447), .IN2(n424), .Q(n446) );
  OR2X1 U587 ( .IN1(n448), .IN2(n449), .Q(n447) );
  AND2X1 U588 ( .IN1(n693), .IN2(n450), .Q(n448) );
  AND2X1 U589 ( .IN1(n700), .IN2(test_se), .Q(n445) );
  OR2X1 U590 ( .IN1(n451), .IN2(n452), .Q(n175) );
  AND2X1 U591 ( .IN1(n693), .IN2(n453), .Q(n452) );
  OR2X1 U592 ( .IN1(n454), .IN2(test_se), .Q(n453) );
  AND3X1 U593 ( .IN1(n455), .IN2(n424), .IN3(n694), .Q(n451) );
  OR2X1 U594 ( .IN1(n456), .IN2(n457), .Q(n174) );
  AND2X1 U595 ( .IN1(n694), .IN2(n458), .Q(n457) );
  OR3X1 U596 ( .IN1(n459), .IN2(n460), .IN3(test_se), .Q(n458) );
  AND2X1 U597 ( .IN1(n449), .IN2(n692), .Q(n460) );
  AND3X1 U598 ( .IN1(n461), .IN2(n693), .IN3(n406), .Q(n459) );
  AND3X1 U599 ( .IN1(n462), .IN2(n424), .IN3(n692), .Q(n456) );
  OR2X1 U600 ( .IN1(n454), .IN2(n450), .Q(n462) );
  AND2X1 U601 ( .IN1(n461), .IN2(n411), .Q(n454) );
  OR2X1 U602 ( .IN1(n463), .IN2(n464), .Q(n173) );
  AND2X1 U603 ( .IN1(n465), .IN2(n424), .Q(n464) );
  OR2X1 U604 ( .IN1(n466), .IN2(n467), .Q(n465) );
  AND2X1 U605 ( .IN1(n691), .IN2(n455), .Q(n467) );
  OR2X1 U606 ( .IN1(n449), .IN2(n450), .Q(n455) );
  AND2X1 U607 ( .IN1(n468), .IN2(n469), .Q(n450) );
  AND2X1 U608 ( .IN1(n404), .IN2(n461), .Q(n449) );
  AND3X1 U609 ( .IN1(n470), .IN2(n471), .IN3(n461), .Q(n466) );
  INVX0 U610 ( .INP(n468), .ZN(n461) );
  OR3X1 U611 ( .IN1(n246), .IN2(n239), .IN3(n432), .Q(n468) );
  OR2X1 U612 ( .IN1(n472), .IN2(n473), .Q(n432) );
  INVX0 U613 ( .INP(n474), .ZN(n473) );
  AND4X1 U614 ( .IN1(n691), .IN2(n411), .IN3(n404), .IN4(n406), .Q(n472) );
  INVX0 U615 ( .INP(n475), .ZN(n471) );
  AND2X1 U616 ( .IN1(n691), .IN2(n476), .Q(n475) );
  OR2X1 U617 ( .IN1(n691), .IN2(n477), .Q(n470) );
  AND2X1 U618 ( .IN1(n476), .IN2(n693), .Q(n477) );
  AND2X1 U619 ( .IN1(n694), .IN2(n692), .Q(n476) );
  AND2X1 U620 ( .IN1(n692), .IN2(test_se), .Q(n463) );
  OR2X1 U621 ( .IN1(n478), .IN2(n479), .Q(n172) );
  AND2X1 U622 ( .IN1(n480), .IN2(n424), .Q(n479) );
  OR3X1 U623 ( .IN1(n481), .IN2(n482), .IN3(n483), .Q(n480) );
  AND2X1 U624 ( .IN1(xmit_dataH_7_), .IN2(n444), .Q(n482) );
  AND2X1 U625 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n481) );
  AND2X1 U626 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n478) );
  OR2X1 U627 ( .IN1(n485), .IN2(n486), .Q(n171) );
  AND2X1 U628 ( .IN1(n487), .IN2(n424), .Q(n486) );
  OR3X1 U629 ( .IN1(n488), .IN2(n489), .IN3(n490), .Q(n487) );
  AND2X1 U630 ( .IN1(xmit_dataH_6_), .IN2(n491), .Q(n490) );
  AND2X1 U631 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n489) );
  AND2X1 U632 ( .IN1(n483), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n488) );
  AND2X1 U633 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n485) );
  OR2X1 U634 ( .IN1(n492), .IN2(n493), .Q(n170) );
  AND2X1 U635 ( .IN1(n494), .IN2(n424), .Q(n493) );
  OR3X1 U636 ( .IN1(n495), .IN2(n496), .IN3(n497), .Q(n494) );
  AND2X1 U637 ( .IN1(xmit_dataH_5_), .IN2(n491), .Q(n497) );
  AND2X1 U638 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n496) );
  AND2X1 U639 ( .IN1(n483), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n495) );
  AND2X1 U640 ( .IN1(n685), .IN2(test_se), .Q(n492) );
  OR2X1 U641 ( .IN1(n498), .IN2(n499), .Q(n169) );
  AND2X1 U642 ( .IN1(n500), .IN2(n424), .Q(n499) );
  OR3X1 U643 ( .IN1(n501), .IN2(n502), .IN3(n503), .Q(n500) );
  AND2X1 U644 ( .IN1(xmit_dataH_4_), .IN2(n491), .Q(n503) );
  AND2X1 U645 ( .IN1(n685), .IN2(n484), .Q(n502) );
  AND2X1 U646 ( .IN1(n483), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n501) );
  AND2X1 U647 ( .IN1(n686), .IN2(test_se), .Q(n498) );
  OR2X1 U648 ( .IN1(n504), .IN2(n505), .Q(n168) );
  AND2X1 U649 ( .IN1(n506), .IN2(n424), .Q(n505) );
  OR3X1 U650 ( .IN1(n507), .IN2(n508), .IN3(n509), .Q(n506) );
  AND2X1 U651 ( .IN1(xmit_dataH_3_), .IN2(n491), .Q(n509) );
  AND2X1 U652 ( .IN1(n686), .IN2(n484), .Q(n508) );
  AND2X1 U653 ( .IN1(n685), .IN2(n483), .Q(n507) );
  AND2X1 U654 ( .IN1(n687), .IN2(test_se), .Q(n504) );
  OR2X1 U655 ( .IN1(n510), .IN2(n511), .Q(n167) );
  AND2X1 U656 ( .IN1(n512), .IN2(n424), .Q(n511) );
  OR3X1 U657 ( .IN1(n513), .IN2(n514), .IN3(n515), .Q(n512) );
  AND2X1 U658 ( .IN1(xmit_dataH_2_), .IN2(n491), .Q(n515) );
  AND2X1 U659 ( .IN1(n687), .IN2(n484), .Q(n514) );
  AND2X1 U660 ( .IN1(n686), .IN2(n483), .Q(n513) );
  AND2X1 U661 ( .IN1(n688), .IN2(test_se), .Q(n510) );
  OR2X1 U662 ( .IN1(n516), .IN2(n517), .Q(n166) );
  AND2X1 U663 ( .IN1(n518), .IN2(n424), .Q(n517) );
  OR3X1 U664 ( .IN1(n519), .IN2(n520), .IN3(n521), .Q(n518) );
  AND2X1 U665 ( .IN1(xmit_dataH_1_), .IN2(n491), .Q(n521) );
  AND2X1 U666 ( .IN1(n688), .IN2(n484), .Q(n520) );
  AND2X1 U667 ( .IN1(n687), .IN2(n483), .Q(n519) );
  AND2X1 U668 ( .IN1(test_se), .IN2(n409), .Q(n516) );
  OR2X1 U669 ( .IN1(n522), .IN2(n523), .Q(n164) );
  AND2X1 U670 ( .IN1(n524), .IN2(n424), .Q(n523) );
  OR2X1 U671 ( .IN1(n525), .IN2(n526), .Q(n524) );
  INVX0 U672 ( .INP(n469), .ZN(n526) );
  OR3X1 U673 ( .IN1(xmitH), .IN2(n698), .IN3(iXMIT_state_1_temp), .Q(n469) );
  AND2X1 U674 ( .IN1(n439), .IN2(n434), .Q(n525) );
  AND2X1 U675 ( .IN1(n700), .IN2(n527), .Q(n434) );
  AND2X1 U676 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n522) );
  OR3X1 U677 ( .IN1(n528), .IN2(n529), .IN3(n530), .Q(n163) );
  AND3X1 U678 ( .IN1(n531), .IN2(n424), .IN3(n245), .Q(n529) );
  INVX0 U679 ( .INP(n532), .ZN(n531) );
  AND2X1 U680 ( .IN1(n533), .IN2(n695), .Q(n532) );
  OR2X1 U681 ( .IN1(n534), .IN2(n241), .Q(n533) );
  AND2X1 U682 ( .IN1(n535), .IN2(iRECEIVER_state_0_), .Q(n528) );
  OR3X1 U683 ( .IN1(n536), .IN2(n537), .IN3(test_se), .Q(n535) );
  AND3X1 U684 ( .IN1(n238), .IN2(n413), .IN3(n241), .Q(n537) );
  AND2X1 U685 ( .IN1(n538), .IN2(iRECEIVER_state_1_), .Q(n536) );
  OR2X1 U686 ( .IN1(n539), .IN2(n540), .Q(n162) );
  AND2X1 U687 ( .IN1(n541), .IN2(n424), .Q(n540) );
  OR3X1 U688 ( .IN1(n542), .IN2(n543), .IN3(iRECEIVER_state_2_), .Q(n541) );
  AND2X1 U689 ( .IN1(n544), .IN2(iRECEIVER_state_1_), .Q(n543) );
  OR2X1 U690 ( .IN1(n545), .IN2(n534), .Q(n544) );
  AND2X1 U691 ( .IN1(n546), .IN2(iRECEIVER_state_0_), .Q(n545) );
  OR2X1 U692 ( .IN1(n547), .IN2(n538), .Q(n546) );
  INVX0 U693 ( .INP(n548), .ZN(n538) );
  AND4X1 U694 ( .IN1(n689), .IN2(n405), .IN3(n403), .IN4(n407), .Q(n547) );
  AND2X1 U695 ( .IN1(n241), .IN2(n695), .Q(n542) );
  AND2X1 U696 ( .IN1(n689), .IN2(test_se), .Q(n539) );
  OR2X1 U697 ( .IN1(n549), .IN2(n550), .Q(n161) );
  AND2X1 U698 ( .IN1(test_si), .IN2(test_se), .Q(n550) );
  AND2X1 U699 ( .IN1(iRECEIVER_N20), .IN2(n424), .Q(n549) );
  OR2X1 U700 ( .IN1(n551), .IN2(n552), .Q(n160) );
  AND2X1 U701 ( .IN1(iRECEIVER_N21), .IN2(n424), .Q(n552) );
  AND2X1 U702 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n551) );
  OR2X1 U703 ( .IN1(n553), .IN2(n554), .Q(n159) );
  AND2X1 U704 ( .IN1(iRECEIVER_N22), .IN2(n424), .Q(n554) );
  AND2X1 U705 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n553) );
  OR2X1 U706 ( .IN1(n555), .IN2(n556), .Q(n157) );
  AND2X1 U707 ( .IN1(n707), .IN2(test_se), .Q(n556) );
  AND2X1 U708 ( .IN1(iRECEIVER_N23), .IN2(n424), .Q(n555) );
  OR2X1 U709 ( .IN1(n557), .IN2(iRECEIVER_next_state_2_), .Q(n156) );
  AND2X1 U710 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n557) );
  OR2X1 U711 ( .IN1(n558), .IN2(n559), .Q(n155) );
  AND2X1 U712 ( .IN1(n690), .IN2(test_se), .Q(n559) );
  AND2X1 U713 ( .IN1(n560), .IN2(n424), .Q(n558) );
  OR2X1 U714 ( .IN1(n561), .IN2(n562), .Q(n560) );
  AND2X1 U715 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n561)
         );
  OR3X1 U716 ( .IN1(n563), .IN2(n564), .IN3(n565), .Q(n154) );
  AND2X1 U717 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n565) );
  AND2X1 U718 ( .IN1(n530), .IN2(n695), .Q(n564) );
  AND2X1 U719 ( .IN1(rec_dataH_rec_7), .IN2(n566), .Q(n563) );
  OR2X1 U720 ( .IN1(n567), .IN2(n568), .Q(n153) );
  AND2X1 U721 ( .IN1(rec_dataH_temp_6), .IN2(test_se), .Q(n568) );
  AND2X1 U722 ( .IN1(rec_dataH_rec_7), .IN2(n424), .Q(n567) );
  OR2X1 U723 ( .IN1(n569), .IN2(n570), .Q(n152) );
  AND2X1 U724 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n570) );
  AND2X1 U725 ( .IN1(test_so), .IN2(n424), .Q(n569) );
  OR3X1 U726 ( .IN1(n571), .IN2(n572), .IN3(n573), .Q(n150) );
  AND2X1 U727 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n573) );
  AND2X1 U728 ( .IN1(n530), .IN2(rec_dataH_rec_7), .Q(n572) );
  AND2X1 U729 ( .IN1(rec_dataH_rec_6), .IN2(n566), .Q(n571) );
  OR2X1 U730 ( .IN1(n574), .IN2(n575), .Q(n149) );
  AND2X1 U731 ( .IN1(rec_dataH_temp_5), .IN2(test_se), .Q(n575) );
  AND2X1 U732 ( .IN1(rec_dataH_rec_6), .IN2(n424), .Q(n574) );
  OR2X1 U733 ( .IN1(n576), .IN2(n577), .Q(n148) );
  AND2X1 U734 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n577) );
  AND2X1 U735 ( .IN1(rec_dataH_temp_6), .IN2(n424), .Q(n576) );
  OR3X1 U736 ( .IN1(n578), .IN2(n579), .IN3(n580), .Q(n147) );
  AND2X1 U737 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n580) );
  AND2X1 U738 ( .IN1(rec_dataH_rec_6), .IN2(n530), .Q(n579) );
  AND2X1 U739 ( .IN1(rec_dataH_rec_5), .IN2(n566), .Q(n578) );
  OR2X1 U740 ( .IN1(n581), .IN2(n582), .Q(n146) );
  AND2X1 U741 ( .IN1(rec_dataH_temp_4), .IN2(test_se), .Q(n582) );
  AND2X1 U742 ( .IN1(rec_dataH_rec_5), .IN2(n424), .Q(n581) );
  OR2X1 U743 ( .IN1(n583), .IN2(n584), .Q(n145) );
  AND2X1 U744 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n584) );
  AND2X1 U745 ( .IN1(rec_dataH_temp_5), .IN2(n424), .Q(n583) );
  OR3X1 U746 ( .IN1(n585), .IN2(n586), .IN3(n587), .Q(n143) );
  AND2X1 U747 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n587) );
  AND2X1 U748 ( .IN1(rec_dataH_rec_5), .IN2(n530), .Q(n586) );
  AND2X1 U749 ( .IN1(rec_dataH_rec_4), .IN2(n566), .Q(n585) );
  OR2X1 U750 ( .IN1(n588), .IN2(n589), .Q(n142) );
  AND2X1 U751 ( .IN1(rec_dataH_temp_3), .IN2(test_se), .Q(n589) );
  AND2X1 U752 ( .IN1(rec_dataH_rec_4), .IN2(n424), .Q(n588) );
  OR2X1 U753 ( .IN1(n590), .IN2(n591), .Q(n141) );
  AND2X1 U754 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n591) );
  AND2X1 U755 ( .IN1(rec_dataH_temp_4), .IN2(n424), .Q(n590) );
  OR3X1 U756 ( .IN1(n592), .IN2(n593), .IN3(n594), .Q(n140) );
  AND2X1 U757 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n594) );
  AND2X1 U758 ( .IN1(rec_dataH_rec_4), .IN2(n530), .Q(n593) );
  AND2X1 U759 ( .IN1(rec_dataH_rec_3), .IN2(n566), .Q(n592) );
  OR2X1 U760 ( .IN1(n595), .IN2(n596), .Q(n139) );
  AND2X1 U761 ( .IN1(rec_dataH_temp_2), .IN2(test_se), .Q(n596) );
  AND2X1 U762 ( .IN1(rec_dataH_rec_3), .IN2(n424), .Q(n595) );
  OR2X1 U763 ( .IN1(n597), .IN2(n598), .Q(n138) );
  AND2X1 U764 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n598) );
  AND2X1 U765 ( .IN1(rec_dataH_temp_3), .IN2(n424), .Q(n597) );
  OR3X1 U766 ( .IN1(n599), .IN2(n600), .IN3(n601), .Q(n136) );
  AND2X1 U767 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n601) );
  AND2X1 U768 ( .IN1(rec_dataH_rec_3), .IN2(n530), .Q(n600) );
  AND2X1 U769 ( .IN1(rec_dataH_rec_2), .IN2(n566), .Q(n599) );
  OR2X1 U770 ( .IN1(n602), .IN2(n603), .Q(n135) );
  AND2X1 U771 ( .IN1(rec_dataH_temp_1), .IN2(test_se), .Q(n603) );
  AND2X1 U772 ( .IN1(rec_dataH_rec_2), .IN2(n424), .Q(n602) );
  OR2X1 U773 ( .IN1(n604), .IN2(n605), .Q(n134) );
  AND2X1 U774 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n605) );
  AND2X1 U775 ( .IN1(rec_dataH_temp_2), .IN2(n424), .Q(n604) );
  OR3X1 U776 ( .IN1(n606), .IN2(n607), .IN3(n608), .Q(n133) );
  AND2X1 U777 ( .IN1(rec_dataH_rec_0_temp), .IN2(test_se), .Q(n608) );
  AND2X1 U778 ( .IN1(rec_dataH_rec_2), .IN2(n530), .Q(n607) );
  AND2X1 U779 ( .IN1(rec_dataH_rec_1), .IN2(n566), .Q(n606) );
  OR2X1 U780 ( .IN1(n609), .IN2(n610), .Q(n132) );
  AND2X1 U781 ( .IN1(rec_dataH_temp_0), .IN2(test_se), .Q(n610) );
  AND2X1 U782 ( .IN1(rec_dataH_rec_1), .IN2(n424), .Q(n609) );
  OR2X1 U783 ( .IN1(n611), .IN2(n612), .Q(n131) );
  AND2X1 U784 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n612) );
  AND2X1 U785 ( .IN1(rec_dataH_temp_1), .IN2(n424), .Q(n611) );
  OR3X1 U786 ( .IN1(n613), .IN2(n614), .IN3(n615), .Q(n129) );
  AND2X1 U787 ( .IN1(n706), .IN2(test_se), .Q(n615) );
  AND2X1 U788 ( .IN1(rec_dataH_rec_1), .IN2(n530), .Q(n614) );
  AND2X1 U789 ( .IN1(rec_dataH_rec_0_temp), .IN2(n566), .Q(n613) );
  AND2X1 U790 ( .IN1(n424), .IN2(n616), .Q(n566) );
  OR2X1 U791 ( .IN1(iRECEIVER_state_0_), .IN2(n238), .Q(n616) );
  OR2X1 U792 ( .IN1(n617), .IN2(n618), .Q(n128) );
  AND2X1 U793 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n618) );
  AND2X1 U794 ( .IN1(rec_dataH_rec_0_temp), .IN2(n424), .Q(n617) );
  OR2X1 U795 ( .IN1(n619), .IN2(n620), .Q(n127) );
  AND2X1 U796 ( .IN1(xmit_doneH_temp), .IN2(test_se), .Q(n620) );
  AND2X1 U797 ( .IN1(rec_dataH_temp_0), .IN2(n424), .Q(n619) );
  OR3X1 U798 ( .IN1(n621), .IN2(n622), .IN3(n623), .Q(n126) );
  AND2X1 U799 ( .IN1(n696), .IN2(test_se), .Q(n623) );
  AND2X1 U800 ( .IN1(n624), .IN2(n689), .Q(n622) );
  AND2X1 U801 ( .IN1(n530), .IN2(iRECEIVER_N28), .Q(n621) );
  OR3X1 U802 ( .IN1(n625), .IN2(n626), .IN3(n627), .Q(n125) );
  AND2X1 U803 ( .IN1(test_se), .IN2(rec_readyH), .Q(n627) );
  AND2X1 U804 ( .IN1(n624), .IN2(n704), .Q(n626) );
  AND2X1 U805 ( .IN1(n530), .IN2(n403), .Q(n625) );
  OR3X1 U806 ( .IN1(n628), .IN2(n629), .IN3(n630), .Q(n124) );
  AND2X1 U807 ( .IN1(n704), .IN2(test_se), .Q(n630) );
  AND2X1 U808 ( .IN1(n624), .IN2(n705), .Q(n629) );
  AND2X1 U809 ( .IN1(n530), .IN2(iRECEIVER_N26), .Q(n628) );
  OR3X1 U810 ( .IN1(n631), .IN2(n632), .IN3(n633), .Q(n122) );
  AND2X1 U811 ( .IN1(n705), .IN2(test_se), .Q(n633) );
  AND2X1 U812 ( .IN1(n624), .IN2(n696), .Q(n632) );
  INVX0 U813 ( .INP(n634), .ZN(n624) );
  OR3X1 U814 ( .IN1(n635), .IN2(n562), .IN3(test_se), .Q(n634) );
  AND3X1 U815 ( .IN1(n241), .IN2(n695), .IN3(n238), .Q(n562) );
  AND2X1 U816 ( .IN1(n245), .IN2(iRECEIVER_state_2_), .Q(n635) );
  AND2X1 U817 ( .IN1(iRECEIVER_N27), .IN2(n530), .Q(n631) );
  AND3X1 U818 ( .IN1(n424), .IN2(iRECEIVER_state_2_), .IN3(n245), .Q(n530) );
  OR2X1 U819 ( .IN1(n636), .IN2(n637), .Q(n121) );
  AND2X1 U820 ( .IN1(n701), .IN2(test_se), .Q(n637) );
  AND3X1 U821 ( .IN1(iXMIT_N25), .IN2(n638), .IN3(n424), .Q(n636) );
  OR2X1 U822 ( .IN1(n639), .IN2(n640), .Q(n120) );
  AND2X1 U823 ( .IN1(iXMIT_N26), .IN2(n424), .Q(n640) );
  AND2X1 U824 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n639) );
  OR2X1 U825 ( .IN1(n641), .IN2(n642), .Q(n119) );
  AND2X1 U826 ( .IN1(n703), .IN2(test_se), .Q(n642) );
  AND2X1 U827 ( .IN1(iXMIT_N27), .IN2(n424), .Q(n641) );
  OR2X1 U828 ( .IN1(n643), .IN2(n644), .Q(n118) );
  AND2X1 U829 ( .IN1(n645), .IN2(n424), .Q(n644) );
  OR3X1 U830 ( .IN1(n646), .IN2(n647), .IN3(n648), .Q(n645) );
  AND2X1 U831 ( .IN1(xmit_dataH_0_), .IN2(n491), .Q(n648) );
  AND2X1 U832 ( .IN1(n484), .IN2(n409), .Q(n647) );
  AND2X1 U833 ( .IN1(n688), .IN2(n483), .Q(n646) );
  INVX0 U834 ( .INP(n649), .ZN(n483) );
  OR2X1 U835 ( .IN1(n491), .IN2(n484), .Q(n649) );
  INVX0 U836 ( .INP(n444), .ZN(n484) );
  OR2X1 U837 ( .IN1(n650), .IN2(n491), .Q(n444) );
  AND2X1 U838 ( .IN1(n698), .IN2(n239), .Q(n650) );
  AND3X1 U839 ( .IN1(n242), .IN2(n246), .IN3(xmitH), .Q(n491) );
  AND2X1 U840 ( .IN1(test_se), .IN2(n698), .Q(n643) );
  OR2X1 U841 ( .IN1(n651), .IN2(n652), .Q(n117) );
  AND2X1 U842 ( .IN1(n695), .IN2(test_se), .Q(n652) );
  AND2X1 U843 ( .IN1(uart_REC_dataH), .IN2(n424), .Q(n651) );
  OR2X1 U844 ( .IN1(n653), .IN2(n654), .Q(n115) );
  AND2X1 U845 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n654) );
  AND2X1 U846 ( .IN1(n690), .IN2(n424), .Q(n653) );
  INVX0 U847 ( .INP(test_se), .ZN(n424) );
  AND2X1 U848 ( .IN1(n638), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U849 ( .IN1(n655), .IN2(n656), .Q(iXMIT_N27) );
  AND2X1 U850 ( .IN1(iXMIT_N26), .IN2(n702), .Q(n656) );
  AND3X1 U851 ( .IN1(n703), .IN2(n638), .IN3(n412), .Q(n655) );
  AND2X1 U852 ( .IN1(n410), .IN2(n638), .Q(iXMIT_N26) );
  OR2X1 U853 ( .IN1(n443), .IN2(n439), .Q(n638) );
  INVX0 U854 ( .INP(n416), .ZN(n439) );
  OR2X1 U855 ( .IN1(n239), .IN2(n242), .Q(n416) );
  AND2X1 U856 ( .IN1(n657), .IN2(iXMIT_state_1_temp), .Q(n443) );
  INVX0 U857 ( .INP(n438), .ZN(n657) );
  AND2X1 U858 ( .IN1(n699), .IN2(n474), .Q(n438) );
  AND4X1 U859 ( .IN1(n701), .IN2(n700), .IN3(n410), .IN4(n702), .Q(n474) );
  OR2X1 U860 ( .IN1(n658), .IN2(n659), .Q(iXMIT_N25) );
  INVX0 U861 ( .INP(n660), .ZN(n659) );
  OR2X1 U862 ( .IN1(n661), .IN2(n700), .Q(n660) );
  AND2X1 U863 ( .IN1(n700), .IN2(n661), .Q(n658) );
  AND2X1 U864 ( .IN1(n661), .IN2(n662), .Q(iXMIT_N24) );
  OR2X1 U865 ( .IN1(n701), .IN2(n663), .Q(n662) );
  AND2X1 U866 ( .IN1(n702), .IN2(n703), .Q(n663) );
  INVX0 U867 ( .INP(n527), .ZN(n661) );
  AND3X1 U868 ( .IN1(n702), .IN2(n703), .IN3(n701), .Q(n527) );
  AND2X1 U869 ( .IN1(iRECEIVER_state_1_), .IN2(n664), .Q(
        iRECEIVER_next_state_2_) );
  OR2X1 U870 ( .IN1(n665), .IN2(n666), .Q(iRECEIVER_N28) );
  INVX0 U871 ( .INP(n667), .ZN(n666) );
  OR2X1 U872 ( .IN1(n668), .IN2(n689), .Q(n667) );
  AND2X1 U873 ( .IN1(n689), .IN2(n668), .Q(n665) );
  AND2X1 U874 ( .IN1(n668), .IN2(n669), .Q(iRECEIVER_N27) );
  OR2X1 U875 ( .IN1(n696), .IN2(n670), .Q(n669) );
  AND2X1 U876 ( .IN1(n705), .IN2(n704), .Q(n670) );
  OR3X1 U877 ( .IN1(n405), .IN2(n403), .IN3(n407), .Q(n668) );
  OR2X1 U878 ( .IN1(n671), .IN2(n672), .Q(iRECEIVER_N26) );
  AND2X1 U879 ( .IN1(n705), .IN2(n403), .Q(n672) );
  AND2X1 U880 ( .IN1(n704), .IN2(n405), .Q(n671) );
  AND2X1 U881 ( .IN1(iRECEIVER_N19), .IN2(n673), .Q(iRECEIVER_N23) );
  AND2X1 U882 ( .IN1(n673), .IN2(iRECEIVER_N18), .Q(iRECEIVER_N22) );
  AND2X1 U883 ( .IN1(iRECEIVER_N17), .IN2(n673), .Q(iRECEIVER_N21) );
  AND2X1 U884 ( .IN1(n255), .IN2(n673), .Q(iRECEIVER_N20) );
  INVX0 U885 ( .INP(n674), .ZN(n673) );
  OR4X1 U886 ( .IN1(n675), .IN2(iRECEIVER_state_2_), .IN3(n241), .IN4(n664), 
        .Q(n674) );
  AND2X1 U887 ( .IN1(iRECEIVER_state_0_), .IN2(n548), .Q(n664) );
  AND4X1 U888 ( .IN1(n707), .IN2(n706), .IN3(iRECEIVER_bitCell_cntrH_1_), 
        .IN4(n255), .Q(n548) );
  AND2X1 U889 ( .IN1(n534), .IN2(n245), .Q(n675) );
  AND4X1 U890 ( .IN1(n255), .IN2(n707), .IN3(n408), .IN4(n244), .Q(n534) );
  INVX0 U891 ( .INP(n676), .ZN(iRECEIVER_N19) );
  AND2X1 U892 ( .IN1(n677), .IN2(n678), .Q(n676) );
  OR2X1 U893 ( .IN1(n679), .IN2(n706), .Q(n678) );
  OR2X1 U894 ( .IN1(n408), .IN2(n680), .Q(n677) );
  AND2X1 U895 ( .IN1(n679), .IN2(n681), .Q(iRECEIVER_N18) );
  OR2X1 U896 ( .IN1(n707), .IN2(n682), .Q(n681) );
  AND2X1 U897 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .Q(n682) );
  INVX0 U898 ( .INP(n680), .ZN(n679) );
  AND3X1 U899 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .IN3(n707), .Q(n680) );
  OR2X1 U900 ( .IN1(n683), .IN2(n684), .Q(iRECEIVER_N17) );
  AND2X1 U901 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n684) );
  AND2X1 U902 ( .IN1(n255), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n683) );
endmodule

