module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n716_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n705_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n269_, new_n512_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n151_, keyIn_0_3 );
nand g001 ( new_n152_, N29, N42, N75 );
nand g002 ( new_n153_, new_n152_, new_n151_ );
nand g003 ( new_n154_, keyIn_0_3, N29, N42, N75 );
nand g004 ( N388, new_n153_, new_n154_ );
nand g005 ( new_n156_, N29, N36, N80 );
not g006 ( N389, new_n156_ );
not g007 ( new_n158_, keyIn_0_4 );
nand g008 ( new_n159_, N29, N36, N42 );
not g009 ( new_n160_, new_n159_ );
nand g010 ( new_n161_, new_n160_, new_n158_ );
nand g011 ( new_n162_, new_n159_, keyIn_0_4 );
nand g012 ( N390, new_n161_, new_n162_ );
nand g013 ( new_n164_, N85, N86 );
not g014 ( N391, new_n164_ );
not g015 ( new_n166_, keyIn_0_0 );
nand g016 ( new_n167_, N1, N8 );
not g017 ( new_n168_, new_n167_ );
nand g018 ( new_n169_, new_n168_, N13, N17 );
nand g019 ( new_n170_, new_n169_, new_n166_ );
not g020 ( new_n171_, new_n170_ );
nor g021 ( new_n172_, new_n169_, new_n166_ );
nor g022 ( N418, new_n171_, new_n172_ );
not g023 ( new_n174_, keyIn_0_1 );
nand g024 ( new_n175_, new_n160_, new_n174_ );
nand g025 ( new_n176_, new_n159_, keyIn_0_1 );
nand g026 ( new_n177_, new_n175_, new_n176_ );
nand g027 ( new_n178_, N1, N26 );
nand g028 ( new_n179_, N13, N17 );
nor g029 ( new_n180_, new_n178_, new_n179_ );
nand g030 ( N419, new_n177_, new_n180_ );
nand g031 ( N420, N59, N75, N80 );
nand g032 ( N421, N36, N59, N80 );
nand g033 ( new_n184_, N36, N42, N59 );
nand g034 ( new_n185_, new_n184_, keyIn_0_5 );
not g035 ( new_n186_, keyIn_0_5 );
nand g036 ( new_n187_, new_n186_, N36, N42, N59 );
nand g037 ( new_n188_, new_n185_, new_n187_ );
not g038 ( N422, new_n188_ );
not g039 ( new_n190_, N90 );
nor g040 ( new_n191_, N87, N88 );
nor g041 ( N423, new_n191_, new_n190_ );
nand g042 ( N446, new_n175_, new_n176_, new_n180_ );
not g043 ( new_n194_, keyIn_0_2 );
nand g044 ( new_n195_, N1, N26, N51 );
nand g045 ( new_n196_, new_n195_, new_n194_ );
nand g046 ( new_n197_, keyIn_0_2, N1, N26, N51 );
nand g047 ( new_n198_, new_n196_, new_n197_ );
not g048 ( N447, new_n198_ );
nand g049 ( new_n200_, new_n168_, N13, N55 );
nand g050 ( new_n201_, N29, N68 );
nor g051 ( N448, new_n200_, new_n201_ );
not g052 ( new_n203_, keyIn_0_12 );
not g053 ( new_n204_, new_n200_ );
nand g054 ( new_n205_, N59, N68 );
not g055 ( new_n206_, new_n205_ );
nand g056 ( new_n207_, new_n204_, N74, new_n206_ );
not g057 ( new_n208_, new_n207_ );
nor g058 ( new_n209_, new_n208_, new_n203_ );
nor g059 ( new_n210_, new_n207_, keyIn_0_12 );
nor g060 ( N449, new_n209_, new_n210_ );
not g061 ( new_n212_, keyIn_0_9 );
not g062 ( new_n213_, new_n191_ );
nand g063 ( new_n214_, new_n213_, N89 );
nand g064 ( new_n215_, new_n214_, new_n212_ );
nand g065 ( new_n216_, new_n213_, keyIn_0_9, N89 );
nand g066 ( N450, new_n215_, new_n216_ );
not g067 ( new_n218_, keyIn_0_19 );
not g068 ( new_n219_, N135 );
nor g069 ( new_n220_, N111, N116 );
nor g070 ( new_n221_, new_n220_, keyIn_0_6 );
not g071 ( new_n222_, keyIn_0_6 );
nor g072 ( new_n223_, new_n222_, N111, N116 );
nor g073 ( new_n224_, new_n221_, new_n223_ );
nand g074 ( new_n225_, N111, N116 );
not g075 ( new_n226_, new_n225_ );
nor g076 ( new_n227_, new_n224_, new_n226_ );
nand g077 ( new_n228_, N121, N126 );
not g078 ( new_n229_, new_n228_ );
nor g079 ( new_n230_, N121, N126 );
nor g080 ( new_n231_, new_n229_, new_n230_ );
nor g081 ( new_n232_, new_n227_, new_n231_ );
nand g082 ( new_n233_, new_n227_, new_n231_ );
not g083 ( new_n234_, new_n233_ );
nor g084 ( new_n235_, new_n234_, new_n232_ );
not g085 ( new_n236_, new_n235_ );
nand g086 ( new_n237_, new_n236_, new_n218_, new_n219_ );
nand g087 ( new_n238_, new_n235_, N135 );
nand g088 ( new_n239_, new_n236_, new_n219_ );
nand g089 ( new_n240_, new_n239_, keyIn_0_19 );
nand g090 ( new_n241_, new_n240_, new_n237_, new_n238_ );
not g091 ( new_n242_, new_n241_ );
not g092 ( new_n243_, N130 );
not g093 ( new_n244_, N91 );
not g094 ( new_n245_, N96 );
nand g095 ( new_n246_, new_n244_, new_n245_ );
nand g096 ( new_n247_, N91, N96 );
nand g097 ( new_n248_, new_n246_, new_n247_ );
not g098 ( new_n249_, N101 );
not g099 ( new_n250_, N106 );
nand g100 ( new_n251_, new_n249_, new_n250_ );
nand g101 ( new_n252_, N101, N106 );
nand g102 ( new_n253_, new_n251_, new_n252_ );
nand g103 ( new_n254_, new_n248_, new_n253_ );
nand g104 ( new_n255_, new_n246_, new_n251_, new_n247_, new_n252_ );
nand g105 ( new_n256_, new_n254_, new_n255_ );
nand g106 ( new_n257_, new_n256_, new_n243_ );
nand g107 ( new_n258_, new_n254_, N130, new_n255_ );
nand g108 ( new_n259_, new_n242_, new_n257_, new_n258_ );
nor g109 ( new_n260_, new_n259_, keyIn_0_32 );
nand g110 ( new_n261_, new_n259_, keyIn_0_32 );
nand g111 ( new_n262_, new_n257_, new_n258_ );
nand g112 ( new_n263_, new_n241_, new_n262_ );
nand g113 ( new_n264_, new_n261_, new_n263_ );
nor g114 ( N767, new_n264_, new_n260_ );
not g115 ( new_n266_, keyIn_0_25 );
nand g116 ( new_n267_, N171, N177 );
not g117 ( new_n268_, new_n267_ );
nor g118 ( new_n269_, N171, N177 );
nor g119 ( new_n270_, new_n268_, new_n269_ );
not g120 ( new_n271_, keyIn_0_13 );
not g121 ( new_n272_, N159 );
not g122 ( new_n273_, N165 );
nand g123 ( new_n274_, new_n272_, new_n273_ );
nand g124 ( new_n275_, N159, N165 );
nand g125 ( new_n276_, new_n274_, new_n271_, new_n275_ );
nand g126 ( new_n277_, new_n276_, new_n270_ );
not g127 ( new_n278_, new_n270_ );
nand g128 ( new_n279_, new_n278_, new_n271_, new_n274_, new_n275_ );
nand g129 ( new_n280_, new_n279_, new_n266_, new_n243_, new_n277_ );
nand g130 ( new_n281_, new_n279_, new_n277_, new_n243_ );
nand g131 ( new_n282_, new_n281_, keyIn_0_25 );
nand g132 ( new_n283_, new_n279_, new_n277_ );
nand g133 ( new_n284_, new_n283_, N130 );
nand g134 ( new_n285_, new_n282_, new_n284_, keyIn_0_31, new_n280_ );
not g135 ( new_n286_, new_n285_ );
not g136 ( new_n287_, keyIn_0_26 );
not g137 ( new_n288_, N207 );
not g138 ( new_n289_, N183 );
not g139 ( new_n290_, N189 );
nand g140 ( new_n291_, new_n289_, new_n290_ );
nand g141 ( new_n292_, N183, N189 );
nand g142 ( new_n293_, new_n291_, new_n292_ );
not g143 ( new_n294_, N195 );
not g144 ( new_n295_, N201 );
nand g145 ( new_n296_, new_n294_, new_n295_ );
nand g146 ( new_n297_, N195, N201 );
nand g147 ( new_n298_, new_n296_, new_n297_ );
nand g148 ( new_n299_, new_n293_, new_n298_ );
nand g149 ( new_n300_, new_n291_, new_n296_, new_n292_, new_n297_ );
nand g150 ( new_n301_, new_n299_, new_n300_ );
nand g151 ( new_n302_, new_n301_, new_n288_ );
nand g152 ( new_n303_, new_n302_, new_n287_ );
nand g153 ( new_n304_, new_n301_, keyIn_0_26, new_n288_ );
nand g154 ( new_n305_, new_n303_, new_n304_ );
nand g155 ( new_n306_, new_n299_, N207, new_n300_ );
nand g156 ( new_n307_, new_n305_, new_n306_ );
nand g157 ( new_n308_, new_n286_, new_n307_ );
nand g158 ( new_n309_, new_n285_, new_n305_, new_n306_ );
nand g159 ( N768, new_n308_, new_n309_ );
not g160 ( new_n311_, keyIn_0_52 );
not g161 ( new_n312_, keyIn_0_37 );
nand g162 ( new_n313_, N59, N156 );
not g163 ( new_n314_, new_n313_ );
nand g164 ( new_n315_, N17, N42 );
not g165 ( new_n316_, new_n315_ );
nor g166 ( new_n317_, N17, N42 );
nor g167 ( new_n318_, new_n316_, new_n317_ );
nand g168 ( new_n319_, new_n318_, new_n196_, new_n197_, new_n314_ );
nand g169 ( new_n320_, N42, N59, N75 );
nand g170 ( new_n321_, new_n168_, N17, N51, new_n320_ );
nand g171 ( new_n322_, new_n319_, new_n321_ );
nand g172 ( new_n323_, new_n322_, N126 );
nand g173 ( new_n324_, new_n323_, keyIn_0_24 );
not g174 ( new_n325_, keyIn_0_24 );
nand g175 ( new_n326_, new_n322_, new_n325_, N126 );
nand g176 ( new_n327_, new_n324_, new_n326_ );
not g177 ( new_n328_, keyIn_0_15 );
nand g178 ( new_n329_, N29, N55, N75, N80 );
not g179 ( new_n330_, new_n329_ );
nand g180 ( new_n331_, new_n330_, new_n196_, new_n197_ );
nand g181 ( new_n332_, new_n331_, new_n328_ );
nand g182 ( new_n333_, new_n330_, new_n196_, keyIn_0_15, new_n197_ );
nand g183 ( new_n334_, new_n332_, new_n333_ );
nand g184 ( new_n335_, keyIn_0_10, N268 );
not g185 ( new_n336_, new_n335_ );
nor g186 ( new_n337_, keyIn_0_10, N268 );
nor g187 ( new_n338_, new_n336_, new_n337_ );
nand g188 ( new_n339_, new_n334_, new_n338_ );
nand g189 ( new_n340_, new_n196_, N17, new_n197_, new_n313_ );
nand g190 ( new_n341_, new_n340_, N1 );
nand g191 ( new_n342_, new_n341_, N153 );
nand g192 ( new_n343_, new_n339_, new_n342_ );
not g193 ( new_n344_, new_n343_ );
nand g194 ( new_n345_, new_n344_, new_n327_ );
nand g195 ( new_n346_, new_n345_, N201 );
nand g196 ( new_n347_, new_n346_, new_n312_ );
nand g197 ( new_n348_, new_n345_, keyIn_0_37, N201 );
nand g198 ( new_n349_, new_n347_, new_n348_ );
not g199 ( new_n350_, new_n349_ );
not g200 ( new_n351_, keyIn_0_38 );
nand g201 ( new_n352_, new_n344_, new_n327_, new_n295_ );
nand g202 ( new_n353_, new_n352_, new_n351_ );
nand g203 ( new_n354_, new_n344_, new_n327_, keyIn_0_38, new_n295_ );
nand g204 ( new_n355_, new_n353_, new_n354_ );
nand g205 ( new_n356_, new_n350_, new_n355_ );
not g206 ( new_n357_, new_n356_ );
nand g207 ( new_n358_, new_n357_, N261 );
not g208 ( new_n359_, N261 );
nand g209 ( new_n360_, new_n356_, new_n359_ );
nand g210 ( new_n361_, new_n358_, new_n311_, new_n360_ );
nand g211 ( new_n362_, new_n358_, new_n360_ );
nand g212 ( new_n363_, new_n362_, keyIn_0_52 );
nand g213 ( new_n364_, new_n363_, N219, new_n361_ );
nand g214 ( new_n365_, N121, N210 );
nand g215 ( new_n366_, new_n364_, new_n365_ );
nand g216 ( new_n367_, new_n366_, keyIn_0_56 );
not g217 ( new_n368_, keyIn_0_56 );
nand g218 ( new_n369_, new_n364_, new_n368_, new_n365_ );
nand g219 ( new_n370_, new_n367_, new_n369_ );
not g220 ( new_n371_, keyIn_0_16 );
not g221 ( new_n372_, keyIn_0_14 );
nand g222 ( new_n373_, new_n204_, N42, N72, new_n206_ );
not g223 ( new_n374_, new_n373_ );
nand g224 ( new_n375_, new_n374_, keyIn_0_8 );
not g225 ( new_n376_, keyIn_0_8 );
nand g226 ( new_n377_, new_n373_, new_n376_ );
nand g227 ( new_n378_, new_n375_, N73, new_n377_ );
nand g228 ( new_n379_, new_n378_, keyIn_0_11 );
not g229 ( new_n380_, keyIn_0_11 );
nand g230 ( new_n381_, new_n375_, new_n380_, N73, new_n377_ );
nand g231 ( new_n382_, new_n379_, new_n381_ );
nand g232 ( new_n383_, new_n382_, new_n372_ );
nand g233 ( new_n384_, new_n379_, keyIn_0_14, new_n381_ );
nand g234 ( new_n385_, new_n383_, new_n384_ );
nand g235 ( new_n386_, new_n385_, new_n371_ );
nand g236 ( new_n387_, new_n383_, keyIn_0_16, new_n384_ );
nand g237 ( new_n388_, new_n386_, new_n387_ );
nand g238 ( new_n389_, new_n388_, N201 );
nand g239 ( new_n390_, new_n389_, keyIn_0_28 );
not g240 ( new_n391_, keyIn_0_28 );
nand g241 ( new_n392_, new_n388_, new_n391_, N201 );
nand g242 ( new_n393_, new_n390_, new_n392_ );
nand g243 ( new_n394_, new_n357_, N228 );
nand g244 ( new_n395_, N255, N267 );
nand g245 ( new_n396_, new_n345_, N246 );
nand g246 ( new_n397_, new_n394_, new_n395_, new_n396_ );
nand g247 ( new_n398_, new_n349_, N237 );
nand g248 ( new_n399_, new_n398_, keyIn_0_50 );
not g249 ( new_n400_, keyIn_0_50 );
nand g250 ( new_n401_, new_n349_, new_n400_, N237 );
nand g251 ( new_n402_, new_n399_, new_n401_ );
nor g252 ( new_n403_, new_n397_, new_n402_ );
nand g253 ( N850, new_n370_, new_n393_, new_n403_ );
not g254 ( new_n405_, keyIn_0_51 );
nand g255 ( new_n406_, new_n341_, N146 );
nand g256 ( new_n407_, new_n322_, keyIn_0_23, N116 );
not g257 ( new_n408_, keyIn_0_23 );
nand g258 ( new_n409_, new_n322_, N116 );
nand g259 ( new_n410_, new_n409_, new_n408_ );
nand g260 ( new_n411_, new_n410_, new_n339_, new_n406_, new_n407_ );
nand g261 ( new_n412_, new_n411_, keyIn_0_30 );
not g262 ( new_n413_, keyIn_0_30 );
nand g263 ( new_n414_, new_n407_, new_n406_ );
not g264 ( new_n415_, new_n414_ );
nand g265 ( new_n416_, new_n415_, new_n413_, new_n339_, new_n410_ );
nand g266 ( new_n417_, new_n416_, new_n412_ );
nand g267 ( new_n418_, new_n417_, new_n290_ );
nand g268 ( new_n419_, new_n341_, N149 );
nand g269 ( new_n420_, new_n322_, N121 );
nand g270 ( new_n421_, new_n339_, new_n420_, new_n294_, new_n419_ );
nand g271 ( new_n422_, new_n349_, new_n418_, new_n421_ );
nand g272 ( new_n423_, new_n422_, new_n405_ );
nand g273 ( new_n424_, new_n349_, keyIn_0_51, new_n418_, new_n421_ );
nand g274 ( new_n425_, new_n423_, new_n424_ );
not g275 ( new_n426_, keyIn_0_42 );
nand g276 ( new_n427_, new_n355_, N261 );
not g277 ( new_n428_, new_n427_ );
nand g278 ( new_n429_, new_n428_, new_n426_, new_n418_, new_n421_ );
nand g279 ( new_n430_, new_n418_, new_n355_, N261, new_n421_ );
nand g280 ( new_n431_, new_n430_, keyIn_0_42 );
nand g281 ( new_n432_, new_n339_, new_n419_, new_n420_ );
nand g282 ( new_n433_, new_n432_, N195 );
not g283 ( new_n434_, new_n433_ );
nand g284 ( new_n435_, new_n418_, new_n434_ );
not g285 ( new_n436_, new_n417_ );
nand g286 ( new_n437_, new_n436_, N189 );
nand g287 ( new_n438_, new_n435_, new_n437_ );
not g288 ( new_n439_, new_n438_ );
nand g289 ( new_n440_, new_n425_, new_n429_, new_n431_, new_n439_ );
not g290 ( new_n441_, new_n440_ );
not g291 ( new_n442_, keyIn_0_36 );
not g292 ( new_n443_, keyIn_0_29 );
not g293 ( new_n444_, keyIn_0_22 );
nand g294 ( new_n445_, new_n322_, N111 );
nand g295 ( new_n446_, new_n445_, new_n444_ );
nand g296 ( new_n447_, new_n322_, keyIn_0_22, N111 );
nand g297 ( new_n448_, new_n446_, new_n447_ );
nand g298 ( new_n449_, new_n341_, N143 );
nand g299 ( new_n450_, new_n339_, new_n449_ );
not g300 ( new_n451_, new_n450_ );
nand g301 ( new_n452_, new_n451_, new_n448_ );
nand g302 ( new_n453_, new_n452_, new_n443_ );
nand g303 ( new_n454_, new_n451_, new_n448_, keyIn_0_29 );
nand g304 ( new_n455_, new_n453_, new_n454_ );
nand g305 ( new_n456_, new_n455_, N183 );
nand g306 ( new_n457_, new_n456_, new_n442_ );
nand g307 ( new_n458_, new_n455_, keyIn_0_36, N183 );
nand g308 ( new_n459_, new_n457_, new_n458_ );
nand g309 ( new_n460_, new_n453_, new_n289_, new_n454_ );
nand g310 ( new_n461_, new_n459_, new_n460_ );
nor g311 ( new_n462_, new_n441_, new_n461_ );
nand g312 ( new_n463_, new_n462_, keyIn_0_53 );
nand g313 ( new_n464_, new_n441_, new_n461_ );
not g314 ( new_n465_, keyIn_0_53 );
not g315 ( new_n466_, new_n462_ );
nand g316 ( new_n467_, new_n466_, new_n465_ );
nand g317 ( new_n468_, new_n467_, keyIn_0_55, new_n463_, new_n464_ );
not g318 ( new_n469_, keyIn_0_55 );
nand g319 ( new_n470_, new_n467_, new_n463_, new_n464_ );
nand g320 ( new_n471_, new_n470_, new_n469_ );
nand g321 ( new_n472_, new_n471_, N219, new_n468_ );
not g322 ( new_n473_, keyIn_0_47 );
not g323 ( new_n474_, new_n461_ );
nand g324 ( new_n475_, new_n474_, N228 );
nand g325 ( new_n476_, new_n475_, new_n473_ );
nand g326 ( new_n477_, new_n388_, N183 );
nand g327 ( new_n478_, new_n477_, keyIn_0_27 );
not g328 ( new_n479_, keyIn_0_27 );
nand g329 ( new_n480_, new_n388_, new_n479_, N183 );
nand g330 ( new_n481_, new_n478_, new_n480_ );
nand g331 ( new_n482_, new_n455_, N246 );
nand g332 ( new_n483_, N106, N210 );
nand g333 ( new_n484_, new_n481_, new_n482_, new_n483_ );
not g334 ( new_n485_, new_n484_ );
nand g335 ( new_n486_, new_n474_, keyIn_0_47, N228 );
nand g336 ( new_n487_, new_n459_, keyIn_0_40 );
not g337 ( new_n488_, keyIn_0_40 );
nand g338 ( new_n489_, new_n457_, new_n488_, new_n458_ );
nand g339 ( new_n490_, new_n487_, N237, new_n489_ );
nand g340 ( new_n491_, new_n485_, new_n476_, new_n486_, new_n490_ );
not g341 ( new_n492_, new_n491_ );
nand g342 ( N863, new_n472_, new_n492_ );
nand g343 ( new_n494_, new_n437_, new_n418_ );
nor g344 ( new_n495_, new_n428_, new_n349_ );
not g345 ( new_n496_, new_n495_ );
nand g346 ( new_n497_, new_n496_, new_n421_ );
nand g347 ( new_n498_, new_n434_, keyIn_0_49 );
not g348 ( new_n499_, keyIn_0_49 );
nand g349 ( new_n500_, new_n433_, new_n499_ );
nand g350 ( new_n501_, new_n498_, new_n500_ );
not g351 ( new_n502_, new_n501_ );
nand g352 ( new_n503_, new_n497_, new_n494_, new_n502_ );
not g353 ( new_n504_, new_n494_ );
nand g354 ( new_n505_, new_n497_, new_n502_ );
nand g355 ( new_n506_, new_n505_, new_n504_ );
nand g356 ( new_n507_, new_n506_, N219, new_n503_ );
nand g357 ( new_n508_, new_n436_, N189, N237 );
nand g358 ( new_n509_, N111, N210 );
nand g359 ( new_n510_, new_n388_, N189 );
nand g360 ( new_n511_, new_n510_, new_n508_, new_n509_ );
not g361 ( new_n512_, keyIn_0_41 );
nand g362 ( new_n513_, new_n436_, N246 );
nand g363 ( new_n514_, N255, N259 );
nand g364 ( new_n515_, new_n513_, new_n514_ );
nand g365 ( new_n516_, new_n515_, new_n512_ );
nand g366 ( new_n517_, new_n513_, keyIn_0_41, new_n514_ );
nand g367 ( new_n518_, new_n516_, new_n517_ );
nor g368 ( new_n519_, new_n511_, new_n518_ );
not g369 ( new_n520_, keyIn_0_48 );
nand g370 ( new_n521_, new_n504_, N228 );
nand g371 ( new_n522_, new_n521_, new_n520_ );
nand g372 ( new_n523_, new_n504_, keyIn_0_48, N228 );
nand g373 ( N864, new_n507_, new_n519_, new_n522_, new_n523_ );
nand g374 ( new_n525_, new_n433_, new_n421_ );
not g375 ( new_n526_, new_n525_ );
nand g376 ( new_n527_, new_n496_, new_n526_ );
nand g377 ( new_n528_, new_n495_, new_n525_ );
nand g378 ( new_n529_, new_n527_, N219, new_n528_ );
nand g379 ( new_n530_, new_n388_, N195 );
nand g380 ( new_n531_, new_n526_, N228 );
nand g381 ( new_n532_, new_n434_, N237 );
nand g382 ( new_n533_, new_n432_, N246 );
nand g383 ( new_n534_, N255, N260 );
nand g384 ( new_n535_, N116, N210 );
nand g385 ( new_n536_, new_n532_, new_n533_, new_n534_, new_n535_ );
not g386 ( new_n537_, new_n536_ );
nand g387 ( N865, new_n529_, new_n530_, new_n531_, new_n537_ );
nand g388 ( new_n539_, new_n440_, new_n460_ );
not g389 ( new_n540_, keyIn_0_46 );
nand g390 ( new_n541_, new_n487_, new_n489_ );
nand g391 ( new_n542_, new_n541_, new_n540_ );
nand g392 ( new_n543_, new_n487_, keyIn_0_46, new_n489_ );
nand g393 ( new_n544_, new_n539_, new_n542_, new_n543_ );
nand g394 ( new_n545_, new_n544_, keyIn_0_54 );
not g395 ( new_n546_, keyIn_0_54 );
nand g396 ( new_n547_, new_n539_, new_n546_, new_n542_, new_n543_ );
nand g397 ( new_n548_, new_n545_, new_n547_ );
not g398 ( new_n549_, N177 );
not g399 ( new_n550_, keyIn_0_18 );
not g400 ( new_n551_, N268 );
nand g401 ( new_n552_, N29, N75, N80 );
not g402 ( new_n553_, new_n552_ );
nand g403 ( new_n554_, N447, N17, new_n551_, new_n553_ );
nand g404 ( new_n555_, new_n554_, new_n550_ );
not g405 ( new_n556_, new_n554_ );
nand g406 ( new_n557_, new_n556_, keyIn_0_18 );
nand g407 ( new_n558_, new_n557_, new_n555_ );
nand g408 ( new_n559_, new_n322_, N106 );
nand g409 ( new_n560_, N138, N152 );
not g410 ( new_n561_, N55 );
nor g411 ( new_n562_, new_n198_, new_n561_, new_n314_ );
nand g412 ( new_n563_, new_n562_, N153 );
nand g413 ( new_n564_, new_n563_, new_n560_ );
not g414 ( new_n565_, new_n564_ );
nand g415 ( new_n566_, new_n558_, new_n549_, new_n559_, new_n565_ );
nand g416 ( new_n567_, new_n548_, new_n566_ );
nand g417 ( new_n568_, new_n558_, new_n559_, new_n565_ );
nand g418 ( new_n569_, new_n568_, N177 );
nand g419 ( new_n570_, new_n567_, new_n569_ );
not g420 ( new_n571_, N171 );
not g421 ( new_n572_, keyIn_0_17 );
nand g422 ( new_n573_, new_n562_, N149 );
nand g423 ( new_n574_, new_n573_, new_n572_ );
nand g424 ( new_n575_, new_n562_, keyIn_0_17, N149 );
nand g425 ( new_n576_, new_n574_, new_n575_ );
nand g426 ( new_n577_, new_n322_, N101 );
nand g427 ( new_n578_, N17, N138 );
nand g428 ( new_n579_, new_n576_, new_n554_, new_n577_, new_n578_ );
not g429 ( new_n580_, new_n579_ );
nand g430 ( new_n581_, new_n580_, new_n571_ );
nand g431 ( new_n582_, new_n570_, new_n581_ );
not g432 ( new_n583_, keyIn_0_35 );
nand g433 ( new_n584_, new_n579_, N171 );
nand g434 ( new_n585_, new_n584_, new_n583_ );
nand g435 ( new_n586_, new_n579_, keyIn_0_35, N171 );
nand g436 ( new_n587_, new_n585_, new_n586_ );
not g437 ( new_n588_, new_n587_ );
nand g438 ( new_n589_, new_n582_, new_n588_ );
nand g439 ( new_n590_, new_n562_, N146 );
nand g440 ( new_n591_, new_n590_, keyIn_0_21, new_n554_ );
not g441 ( new_n592_, keyIn_0_21 );
nand g442 ( new_n593_, new_n590_, new_n554_ );
nand g443 ( new_n594_, new_n593_, new_n592_ );
nand g444 ( new_n595_, N51, N138 );
nand g445 ( new_n596_, new_n322_, N96 );
nand g446 ( new_n597_, new_n594_, new_n591_, new_n595_, new_n596_ );
nor g447 ( new_n598_, new_n597_, N165 );
not g448 ( new_n599_, new_n598_ );
nand g449 ( new_n600_, new_n589_, new_n599_ );
nand g450 ( new_n601_, new_n597_, N165 );
nand g451 ( new_n602_, new_n600_, new_n601_ );
not g452 ( new_n603_, keyIn_0_20 );
nand g453 ( new_n604_, new_n562_, N143 );
nand g454 ( new_n605_, new_n604_, new_n603_, new_n554_ );
nand g455 ( new_n606_, new_n604_, new_n554_ );
nand g456 ( new_n607_, new_n606_, keyIn_0_20 );
nand g457 ( new_n608_, N8, N138 );
nand g458 ( new_n609_, new_n322_, N91 );
nand g459 ( new_n610_, new_n607_, new_n605_, new_n608_, new_n609_ );
nor g460 ( new_n611_, new_n610_, N159 );
not g461 ( new_n612_, new_n611_ );
nor g462 ( new_n613_, new_n612_, keyIn_0_33 );
nand g463 ( new_n614_, new_n612_, keyIn_0_33 );
not g464 ( new_n615_, new_n614_ );
nor g465 ( new_n616_, new_n615_, new_n613_ );
not g466 ( new_n617_, new_n616_ );
nand g467 ( new_n618_, new_n602_, new_n617_ );
nand g468 ( new_n619_, new_n610_, N159 );
not g469 ( new_n620_, new_n619_ );
nand g470 ( new_n621_, new_n620_, keyIn_0_43 );
not g471 ( new_n622_, keyIn_0_43 );
nand g472 ( new_n623_, new_n619_, new_n622_ );
nand g473 ( new_n624_, new_n621_, new_n623_ );
not g474 ( new_n625_, new_n624_ );
nand g475 ( new_n626_, new_n618_, new_n625_ );
nand g476 ( new_n627_, new_n626_, keyIn_0_59 );
not g477 ( new_n628_, keyIn_0_59 );
nand g478 ( new_n629_, new_n618_, new_n628_, new_n625_ );
nand g479 ( N866, new_n627_, new_n629_ );
not g480 ( new_n631_, keyIn_0_62 );
not g481 ( new_n632_, new_n548_ );
nand g482 ( new_n633_, new_n569_, new_n566_ );
nand g483 ( new_n634_, new_n632_, keyIn_0_57, new_n633_ );
not g484 ( new_n635_, keyIn_0_57 );
nand g485 ( new_n636_, new_n632_, new_n633_ );
nand g486 ( new_n637_, new_n636_, new_n635_ );
not g487 ( new_n638_, new_n633_ );
nand g488 ( new_n639_, new_n548_, new_n638_ );
nand g489 ( new_n640_, new_n637_, N219, new_n634_, new_n639_ );
nand g490 ( new_n641_, new_n388_, N177 );
nand g491 ( new_n642_, new_n638_, N228 );
nand g492 ( new_n643_, new_n568_, N177, N237 );
nand g493 ( new_n644_, new_n568_, N246 );
nand g494 ( new_n645_, N101, N210 );
nand g495 ( new_n646_, new_n643_, new_n644_, new_n645_ );
not g496 ( new_n647_, new_n646_ );
nand g497 ( new_n648_, new_n641_, new_n642_, new_n647_ );
not g498 ( new_n649_, new_n648_ );
nand g499 ( new_n650_, new_n640_, new_n649_ );
nand g500 ( new_n651_, new_n650_, new_n631_ );
nand g501 ( new_n652_, new_n640_, keyIn_0_62, new_n649_ );
nand g502 ( N874, new_n651_, new_n652_ );
nor g503 ( new_n654_, new_n616_, new_n620_ );
nand g504 ( new_n655_, new_n602_, new_n654_ );
not g505 ( new_n656_, new_n654_ );
nand g506 ( new_n657_, new_n600_, new_n601_, new_n656_ );
nand g507 ( new_n658_, new_n655_, N219, new_n657_ );
not g508 ( new_n659_, keyIn_0_39 );
nand g509 ( new_n660_, new_n388_, N159 );
not g510 ( new_n661_, keyIn_0_34 );
nand g511 ( new_n662_, new_n610_, N246 );
nand g512 ( new_n663_, new_n662_, new_n661_ );
nand g513 ( new_n664_, new_n610_, keyIn_0_34, N246 );
nand g514 ( new_n665_, new_n663_, new_n664_ );
nand g515 ( new_n666_, new_n660_, new_n665_ );
nand g516 ( new_n667_, new_n666_, new_n659_ );
nand g517 ( new_n668_, new_n660_, keyIn_0_39, new_n665_ );
nand g518 ( new_n669_, new_n667_, new_n668_ );
nand g519 ( new_n670_, new_n654_, N228 );
not g520 ( new_n671_, new_n338_ );
nand g521 ( new_n672_, new_n671_, N210 );
nand g522 ( new_n673_, new_n620_, N237 );
nand g523 ( new_n674_, new_n673_, new_n672_ );
not g524 ( new_n675_, new_n674_ );
nand g525 ( N878, new_n658_, new_n669_, new_n670_, new_n675_ );
not g526 ( new_n677_, keyIn_0_60 );
not g527 ( new_n678_, new_n601_ );
nor g528 ( new_n679_, new_n678_, new_n598_ );
not g529 ( new_n680_, new_n679_ );
not g530 ( new_n681_, keyIn_0_44 );
nand g531 ( new_n682_, new_n588_, new_n681_ );
nand g532 ( new_n683_, new_n587_, keyIn_0_44 );
nand g533 ( new_n684_, new_n682_, new_n683_ );
not g534 ( new_n685_, new_n684_ );
nand g535 ( new_n686_, new_n582_, new_n680_, new_n685_ );
nand g536 ( new_n687_, new_n686_, keyIn_0_58 );
not g537 ( new_n688_, keyIn_0_58 );
nand g538 ( new_n689_, new_n582_, new_n688_, new_n680_, new_n685_ );
nand g539 ( new_n690_, new_n687_, new_n689_ );
nand g540 ( new_n691_, new_n582_, new_n685_ );
nand g541 ( new_n692_, new_n691_, new_n679_ );
nand g542 ( new_n693_, new_n690_, N219, new_n692_ );
not g543 ( new_n694_, keyIn_0_7 );
nand g544 ( new_n695_, N91, N210 );
nand g545 ( new_n696_, new_n695_, new_n694_ );
nand g546 ( new_n697_, keyIn_0_7, N91, N210 );
nand g547 ( new_n698_, new_n696_, new_n697_ );
nand g548 ( new_n699_, new_n693_, new_n698_ );
nand g549 ( new_n700_, new_n699_, new_n677_ );
nand g550 ( new_n701_, new_n693_, keyIn_0_60, new_n698_ );
nand g551 ( new_n702_, new_n700_, new_n701_ );
nand g552 ( new_n703_, new_n388_, N165 );
nand g553 ( new_n704_, new_n679_, N228 );
nand g554 ( new_n705_, new_n678_, N237 );
nand g555 ( new_n706_, new_n597_, N246 );
nand g556 ( new_n707_, new_n703_, new_n704_, new_n705_, new_n706_ );
not g557 ( new_n708_, new_n707_ );
nand g558 ( N879, new_n702_, new_n708_ );
not g559 ( new_n710_, keyIn_0_61 );
nand g560 ( new_n711_, new_n588_, new_n581_ );
not g561 ( new_n712_, new_n711_ );
nand g562 ( new_n713_, new_n570_, new_n712_ );
nand g563 ( new_n714_, new_n567_, new_n569_, new_n711_ );
nand g564 ( new_n715_, new_n713_, N219, new_n714_ );
nand g565 ( new_n716_, N96, N210 );
nand g566 ( new_n717_, new_n715_, new_n716_ );
nand g567 ( new_n718_, new_n717_, new_n710_ );
nand g568 ( new_n719_, new_n715_, keyIn_0_61, new_n716_ );
nand g569 ( new_n720_, new_n718_, new_n719_ );
nand g570 ( new_n721_, new_n587_, N237 );
nand g571 ( new_n722_, new_n721_, keyIn_0_45 );
not g572 ( new_n723_, keyIn_0_45 );
nand g573 ( new_n724_, new_n587_, new_n723_, N237 );
nand g574 ( new_n725_, new_n722_, new_n724_ );
not g575 ( new_n726_, new_n725_ );
nand g576 ( new_n727_, new_n388_, N171 );
nand g577 ( new_n728_, new_n579_, N246 );
nand g578 ( new_n729_, new_n712_, N228 );
nand g579 ( new_n730_, new_n729_, new_n727_, new_n728_ );
nor g580 ( new_n731_, new_n730_, new_n726_ );
nand g581 ( new_n732_, new_n720_, new_n731_ );
nand g582 ( new_n733_, new_n732_, keyIn_0_63 );
not g583 ( new_n734_, keyIn_0_63 );
nand g584 ( new_n735_, new_n720_, new_n734_, new_n731_ );
nand g585 ( N880, new_n733_, new_n735_ );
endmodule