module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n767_, new_n401_, new_n514_, new_n601_, new_n842_, new_n556_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n481_, new_n1073_, new_n902_, new_n449_, new_n580_, new_n639_, new_n484_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n350_, new_n655_, new_n1054_, new_n1083_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n764_, new_n906_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n429_, new_n355_, new_n926_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n398_, new_n646_, new_n395_, new_n538_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n473_, new_n790_, new_n1081_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n347_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n1002_, new_n834_, new_n369_, new_n448_, new_n867_, new_n1032_, new_n901_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1065_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n499_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n377_, new_n539_, new_n905_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n780_, new_n984_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_;

nand g000 ( new_n343_, N29, N42, N75 );
xnor g001 ( N388, new_n343_, keyIn_0_5 );
nand g002 ( new_n345_, N29, N36, N80 );
xnor g003 ( N389, new_n345_, keyIn_0_6 );
nand g004 ( new_n347_, N29, N36, N42 );
not g005 ( N390, new_n347_ );
nand g006 ( new_n349_, N85, N86 );
nand g007 ( new_n350_, new_n349_, keyIn_0_11 );
not g008 ( new_n351_, keyIn_0_11 );
nand g009 ( new_n352_, new_n351_, N85, N86 );
nand g010 ( N391, new_n350_, new_n352_ );
nand g011 ( new_n354_, N1, N8, N13, N17 );
xnor g012 ( new_n355_, new_n354_, keyIn_0_0 );
xor g013 ( N418, new_n355_, keyIn_0_40 );
nand g014 ( new_n357_, N1, N13, N17, N26 );
xor g015 ( new_n358_, new_n357_, keyIn_0_1 );
xnor g016 ( new_n359_, new_n347_, keyIn_0_2 );
not g017 ( new_n360_, new_n359_ );
nand g018 ( N419, new_n358_, new_n360_ );
nand g019 ( new_n362_, N59, N75, N80 );
xnor g020 ( new_n363_, new_n362_, keyIn_0_7 );
xnor g021 ( N420, new_n363_, keyIn_0_46 );
nand g022 ( new_n365_, N36, N59, N80 );
xor g023 ( new_n366_, new_n365_, keyIn_0_9 );
xnor g024 ( N421, new_n366_, keyIn_0_47 );
nand g025 ( new_n368_, N36, N42, N59 );
xor g026 ( new_n369_, new_n368_, keyIn_0_10 );
xnor g027 ( N422, new_n369_, keyIn_0_48 );
or g028 ( new_n371_, N87, N88 );
nand g029 ( new_n372_, new_n371_, keyIn_0_12 );
or g030 ( new_n373_, keyIn_0_12, N87, N88 );
nand g031 ( new_n374_, new_n372_, new_n373_ );
nand g032 ( new_n375_, new_n374_, N90 );
xnor g033 ( N423, new_n375_, keyIn_0_50 );
nand g034 ( new_n377_, new_n359_, keyIn_0_41 );
or g035 ( new_n378_, new_n359_, keyIn_0_41 );
nand g036 ( new_n379_, new_n378_, new_n358_, new_n377_ );
xor g037 ( N446, new_n379_, keyIn_0_58 );
nand g038 ( new_n381_, N1, N26, N51 );
xnor g039 ( new_n382_, new_n381_, keyIn_0_43 );
xnor g040 ( N447, new_n382_, keyIn_0_60 );
and g041 ( new_n384_, N1, N8, N13, N55 );
nand g042 ( new_n385_, new_n384_, N29, N68 );
xnor g043 ( N448, new_n385_, keyIn_0_62 );
nand g044 ( new_n387_, new_n384_, N59, N68, N74 );
xnor g045 ( new_n388_, new_n387_, keyIn_0_45 );
xnor g046 ( N449, new_n388_, keyIn_0_63 );
nand g047 ( new_n390_, new_n374_, N89 );
xor g048 ( N450, new_n390_, keyIn_0_49 );
not g049 ( new_n392_, N135 );
or g050 ( new_n393_, N121, N126 );
nand g051 ( new_n394_, new_n393_, keyIn_0_18 );
nand g052 ( new_n395_, N121, N126 );
or g053 ( new_n396_, new_n393_, keyIn_0_18 );
nand g054 ( new_n397_, new_n396_, new_n394_, new_n395_ );
xnor g055 ( new_n398_, new_n397_, keyIn_0_53 );
xor g056 ( new_n399_, new_n398_, keyIn_0_68 );
nor g057 ( new_n400_, N111, N116 );
xor g058 ( new_n401_, new_n400_, keyIn_0_17 );
nand g059 ( new_n402_, N111, N116 );
xor g060 ( new_n403_, new_n402_, keyIn_0_16 );
nand g061 ( new_n404_, new_n401_, new_n403_ );
xnor g062 ( new_n405_, new_n404_, keyIn_0_52 );
xor g063 ( new_n406_, new_n405_, keyIn_0_67 );
nand g064 ( new_n407_, new_n406_, new_n399_ );
nand g065 ( new_n408_, new_n407_, keyIn_0_78 );
or g066 ( new_n409_, new_n407_, keyIn_0_78 );
nand g067 ( new_n410_, new_n405_, new_n398_ );
xnor g068 ( new_n411_, new_n410_, keyIn_0_69 );
nand g069 ( new_n412_, new_n409_, new_n408_, new_n411_ );
xor g070 ( new_n413_, new_n412_, keyIn_0_87 );
nor g071 ( new_n414_, new_n413_, new_n392_ );
xnor g072 ( new_n415_, new_n414_, keyIn_0_104 );
nand g073 ( new_n416_, new_n413_, new_n392_ );
xnor g074 ( new_n417_, new_n416_, keyIn_0_105 );
nand g075 ( new_n418_, new_n415_, new_n417_ );
xnor g076 ( new_n419_, new_n418_, keyIn_0_123 );
xnor g077 ( new_n420_, new_n419_, keyIn_0_129 );
not g078 ( new_n421_, N130 );
nor g079 ( new_n422_, N91, N96 );
xnor g080 ( new_n423_, new_n422_, keyIn_0_14 );
nand g081 ( new_n424_, N91, N96 );
xnor g082 ( new_n425_, new_n424_, keyIn_0_13 );
nand g083 ( new_n426_, new_n423_, new_n425_ );
xor g084 ( new_n427_, new_n426_, keyIn_0_51 );
or g085 ( new_n428_, new_n427_, keyIn_0_64 );
not g086 ( new_n429_, N101 );
not g087 ( new_n430_, N106 );
nand g088 ( new_n431_, new_n429_, new_n430_ );
nand g089 ( new_n432_, new_n431_, keyIn_0_15 );
nand g090 ( new_n433_, N101, N106 );
or g091 ( new_n434_, new_n431_, keyIn_0_15 );
nand g092 ( new_n435_, new_n434_, new_n432_, new_n433_ );
xor g093 ( new_n436_, new_n435_, keyIn_0_65 );
nand g094 ( new_n437_, new_n427_, keyIn_0_64 );
nand g095 ( new_n438_, new_n428_, new_n436_, new_n437_ );
or g096 ( new_n439_, new_n438_, keyIn_0_77 );
nand g097 ( new_n440_, new_n438_, keyIn_0_77 );
nand g098 ( new_n441_, new_n427_, new_n435_ );
xor g099 ( new_n442_, new_n441_, keyIn_0_66 );
nand g100 ( new_n443_, new_n439_, new_n440_, new_n442_ );
xnor g101 ( new_n444_, new_n443_, keyIn_0_86 );
nor g102 ( new_n445_, new_n444_, new_n421_ );
xnor g103 ( new_n446_, new_n445_, keyIn_0_102 );
nand g104 ( new_n447_, new_n444_, new_n421_ );
xnor g105 ( new_n448_, new_n447_, keyIn_0_103 );
nand g106 ( new_n449_, new_n446_, new_n448_ );
xnor g107 ( new_n450_, new_n449_, keyIn_0_122 );
xnor g108 ( new_n451_, new_n450_, keyIn_0_128 );
and g109 ( new_n452_, new_n420_, new_n451_ );
nand g110 ( new_n453_, new_n452_, keyIn_0_138 );
nand g111 ( new_n454_, new_n419_, new_n450_ );
or g112 ( new_n455_, new_n452_, keyIn_0_138 );
nand g113 ( new_n456_, new_n455_, new_n453_, new_n454_ );
xor g114 ( N767, new_n456_, keyIn_0_156 );
nor g115 ( new_n458_, N171, N177 );
xor g116 ( new_n459_, new_n458_, keyIn_0_28 );
nand g117 ( new_n460_, N171, N177 );
xor g118 ( new_n461_, new_n460_, keyIn_0_27 );
nand g119 ( new_n462_, new_n459_, new_n461_ );
xor g120 ( new_n463_, new_n462_, keyIn_0_72 );
nor g121 ( new_n464_, N159, N165 );
xnor g122 ( new_n465_, new_n464_, keyIn_0_26 );
nand g123 ( new_n466_, N159, N165 );
xnor g124 ( new_n467_, new_n466_, keyIn_0_25 );
nand g125 ( new_n468_, new_n465_, new_n467_ );
xor g126 ( new_n469_, new_n468_, keyIn_0_71 );
nand g127 ( new_n470_, new_n463_, new_n469_ );
xor g128 ( new_n471_, new_n470_, keyIn_0_84 );
nand g129 ( new_n472_, new_n462_, new_n468_ );
nand g130 ( new_n473_, new_n471_, new_n472_ );
xor g131 ( new_n474_, new_n473_, keyIn_0_101 );
nor g132 ( new_n475_, new_n474_, new_n421_ );
xor g133 ( new_n476_, new_n475_, keyIn_0_114 );
nand g134 ( new_n477_, new_n474_, new_n421_ );
xor g135 ( new_n478_, new_n477_, keyIn_0_115 );
nand g136 ( new_n479_, new_n476_, new_n478_ );
or g137 ( new_n480_, new_n479_, keyIn_0_136 );
not g138 ( new_n481_, N207 );
nor g139 ( new_n482_, N195, N201 );
xnor g140 ( new_n483_, new_n482_, keyIn_0_31 );
nand g141 ( new_n484_, N195, N201 );
xnor g142 ( new_n485_, new_n484_, keyIn_0_30 );
nand g143 ( new_n486_, new_n483_, new_n485_ );
xnor g144 ( new_n487_, new_n486_, keyIn_0_57 );
xnor g145 ( new_n488_, new_n487_, keyIn_0_73 );
nor g146 ( new_n489_, keyIn_0_29, N189 );
xnor g147 ( new_n490_, new_n489_, keyIn_0_56 );
not g148 ( new_n491_, N183 );
nand g149 ( new_n492_, keyIn_0_29, N189 );
nand g150 ( new_n493_, new_n492_, new_n491_ );
xor g151 ( new_n494_, new_n490_, new_n493_ );
nand g152 ( new_n495_, new_n488_, new_n494_ );
xor g153 ( new_n496_, new_n495_, keyIn_0_85 );
not g154 ( new_n497_, new_n494_ );
nand g155 ( new_n498_, new_n497_, new_n487_ );
xnor g156 ( new_n499_, new_n498_, keyIn_0_74 );
nand g157 ( new_n500_, new_n496_, new_n499_ );
nor g158 ( new_n501_, new_n500_, new_n481_ );
xnor g159 ( new_n502_, new_n501_, keyIn_0_116 );
nand g160 ( new_n503_, new_n500_, new_n481_ );
nand g161 ( new_n504_, new_n479_, keyIn_0_136 );
nand g162 ( new_n505_, new_n480_, new_n502_, new_n503_, new_n504_ );
xor g163 ( new_n506_, new_n505_, keyIn_0_139 );
nand g164 ( new_n507_, new_n502_, new_n503_ );
nand g165 ( new_n508_, new_n479_, new_n507_ );
xnor g166 ( new_n509_, new_n508_, keyIn_0_137 );
nand g167 ( new_n510_, new_n506_, new_n509_ );
xor g168 ( N768, new_n510_, keyIn_0_157 );
not g169 ( new_n512_, keyIn_0_192 );
not g170 ( new_n513_, N261 );
not g171 ( new_n514_, N201 );
not g172 ( new_n515_, keyIn_0_59 );
not g173 ( new_n516_, keyIn_0_42 );
nand g174 ( new_n517_, new_n381_, new_n516_ );
or g175 ( new_n518_, new_n381_, new_n516_ );
nand g176 ( new_n519_, new_n518_, new_n517_ );
nand g177 ( new_n520_, new_n519_, new_n515_ );
nand g178 ( new_n521_, new_n518_, keyIn_0_59, new_n517_ );
nand g179 ( new_n522_, new_n520_, new_n521_ );
not g180 ( new_n523_, keyIn_0_55 );
not g181 ( new_n524_, N17 );
not g182 ( new_n525_, N42 );
nand g183 ( new_n526_, new_n524_, new_n525_ );
nand g184 ( new_n527_, new_n526_, keyIn_0_23 );
or g185 ( new_n528_, keyIn_0_23, N17, N42 );
nand g186 ( new_n529_, new_n527_, new_n528_ );
not g187 ( new_n530_, keyIn_0_24 );
nand g188 ( new_n531_, N17, N42 );
nand g189 ( new_n532_, new_n531_, new_n530_ );
nand g190 ( new_n533_, keyIn_0_24, N17, N42 );
nand g191 ( new_n534_, new_n532_, new_n533_ );
nand g192 ( new_n535_, new_n529_, new_n523_, new_n534_ );
nand g193 ( new_n536_, N59, N156 );
not g194 ( new_n537_, new_n536_ );
nand g195 ( new_n538_, new_n529_, new_n534_ );
nand g196 ( new_n539_, new_n538_, keyIn_0_55 );
and g197 ( new_n540_, new_n539_, new_n537_ );
nand g198 ( new_n541_, new_n540_, keyIn_0_82, new_n522_, new_n535_ );
not g199 ( new_n542_, keyIn_0_82 );
nand g200 ( new_n543_, new_n522_, new_n539_, new_n535_, new_n537_ );
nand g201 ( new_n544_, new_n543_, new_n542_ );
nand g202 ( new_n545_, new_n541_, new_n544_ );
nand g203 ( new_n546_, N1, N8, N17, N51 );
xnor g204 ( new_n547_, new_n546_, keyIn_0_3 );
nand g205 ( new_n548_, N42, N59, N75 );
xnor g206 ( new_n549_, new_n548_, keyIn_0_8 );
nand g207 ( new_n550_, new_n547_, new_n549_ );
xor g208 ( new_n551_, new_n550_, keyIn_0_70 );
nand g209 ( new_n552_, new_n545_, new_n551_ );
nand g210 ( new_n553_, new_n552_, keyIn_0_88 );
not g211 ( new_n554_, keyIn_0_88 );
nand g212 ( new_n555_, new_n545_, new_n554_, new_n551_ );
nand g213 ( new_n556_, new_n553_, new_n555_ );
nand g214 ( new_n557_, new_n556_, N126 );
not g215 ( new_n558_, keyIn_0_97 );
xor g216 ( new_n559_, new_n536_, keyIn_0_22 );
nand g217 ( new_n560_, new_n522_, keyIn_0_83, N17, new_n559_ );
not g218 ( new_n561_, keyIn_0_83 );
nand g219 ( new_n562_, new_n522_, N17, new_n559_ );
nand g220 ( new_n563_, new_n562_, new_n561_ );
nand g221 ( new_n564_, new_n563_, N1, new_n560_ );
xnor g222 ( new_n565_, new_n564_, new_n558_ );
nand g223 ( new_n566_, new_n565_, N153 );
nand g224 ( new_n567_, new_n557_, keyIn_0_127, new_n566_ );
not g225 ( new_n568_, N55 );
nand g226 ( new_n569_, new_n522_, N29, N75, N80 );
nor g227 ( new_n570_, new_n569_, new_n568_ );
or g228 ( new_n571_, new_n570_, keyIn_0_81 );
xnor g229 ( new_n572_, keyIn_0_19, N268 );
xnor g230 ( new_n573_, new_n572_, keyIn_0_54 );
nand g231 ( new_n574_, new_n570_, keyIn_0_81 );
nand g232 ( new_n575_, new_n571_, new_n573_, new_n574_ );
not g233 ( new_n576_, keyIn_0_127 );
nand g234 ( new_n577_, new_n557_, new_n566_ );
nand g235 ( new_n578_, new_n577_, new_n576_ );
nand g236 ( new_n579_, new_n578_, new_n567_, new_n575_ );
nand g237 ( new_n580_, new_n579_, keyIn_0_135 );
not g238 ( new_n581_, keyIn_0_135 );
nand g239 ( new_n582_, new_n578_, new_n581_, new_n567_, new_n575_ );
nand g240 ( new_n583_, new_n580_, new_n582_ );
nand g241 ( new_n584_, new_n583_, new_n514_ );
nand g242 ( new_n585_, new_n584_, keyIn_0_154 );
not g243 ( new_n586_, keyIn_0_154 );
nand g244 ( new_n587_, new_n583_, new_n586_, new_n514_ );
and g245 ( new_n588_, new_n585_, new_n587_ );
and g246 ( new_n589_, new_n580_, new_n582_ );
nand g247 ( new_n590_, new_n589_, N201 );
nand g248 ( new_n591_, new_n588_, new_n590_ );
nor g249 ( new_n592_, new_n591_, new_n513_ );
or g250 ( new_n593_, new_n592_, new_n512_ );
nand g251 ( new_n594_, new_n591_, new_n513_ );
nand g252 ( new_n595_, new_n592_, new_n512_ );
nand g253 ( new_n596_, new_n593_, new_n594_, new_n595_ );
or g254 ( new_n597_, new_n596_, keyIn_0_209 );
nand g255 ( new_n598_, new_n596_, keyIn_0_209 );
nand g256 ( new_n599_, new_n597_, N219, new_n598_ );
or g257 ( new_n600_, new_n599_, keyIn_0_215 );
nand g258 ( new_n601_, new_n599_, keyIn_0_215 );
not g259 ( new_n602_, keyIn_0_193 );
and g260 ( new_n603_, new_n588_, N228, new_n590_ );
or g261 ( new_n604_, new_n603_, new_n602_ );
nand g262 ( new_n605_, new_n603_, new_n602_ );
xnor g263 ( new_n606_, new_n590_, keyIn_0_172 );
nand g264 ( new_n607_, new_n606_, N237 );
xnor g265 ( new_n608_, new_n607_, keyIn_0_194 );
nand g266 ( new_n609_, new_n608_, new_n604_, new_n605_ );
xnor g267 ( new_n610_, new_n609_, keyIn_0_210 );
not g268 ( new_n611_, N246 );
nor g269 ( new_n612_, new_n583_, new_n611_ );
nand g270 ( new_n613_, new_n612_, keyIn_0_155 );
or g271 ( new_n614_, new_n612_, keyIn_0_155 );
nand g272 ( new_n615_, N255, N267 );
xor g273 ( new_n616_, new_n615_, keyIn_0_39 );
nand g274 ( new_n617_, new_n614_, new_n613_, new_n616_ );
and g275 ( new_n618_, new_n617_, keyIn_0_173 );
nor g276 ( new_n619_, new_n617_, keyIn_0_173 );
nand g277 ( new_n620_, N42, N59, N68, N72 );
not g278 ( new_n621_, new_n620_ );
or g279 ( new_n622_, new_n621_, keyIn_0_4 );
nand g280 ( new_n623_, new_n621_, keyIn_0_4 );
nand g281 ( new_n624_, new_n622_, new_n384_, new_n623_ );
xnor g282 ( new_n625_, new_n624_, keyIn_0_44 );
nand g283 ( new_n626_, new_n625_, N73 );
xnor g284 ( new_n627_, new_n626_, keyIn_0_61 );
xor g285 ( new_n628_, new_n627_, keyIn_0_76 );
and g286 ( new_n629_, new_n628_, N201 );
nand g287 ( new_n630_, N121, N210 );
xnor g288 ( new_n631_, new_n630_, keyIn_0_38 );
nor g289 ( new_n632_, new_n618_, new_n619_, new_n629_, new_n631_ );
nand g290 ( new_n633_, new_n600_, new_n601_, new_n610_, new_n632_ );
xnor g291 ( new_n634_, new_n633_, keyIn_0_223 );
xnor g292 ( new_n635_, new_n634_, keyIn_0_229 );
xnor g293 ( N850, new_n635_, keyIn_0_234 );
not g294 ( new_n637_, keyIn_0_245 );
not g295 ( new_n638_, keyIn_0_233 );
not g296 ( new_n639_, keyIn_0_226 );
not g297 ( new_n640_, keyIn_0_220 );
not g298 ( new_n641_, keyIn_0_165 );
and g299 ( new_n642_, new_n556_, N111 );
nand g300 ( new_n643_, new_n642_, keyIn_0_111 );
nand g301 ( new_n644_, new_n565_, N143 );
or g302 ( new_n645_, new_n642_, keyIn_0_111 );
nand g303 ( new_n646_, new_n645_, new_n643_, new_n644_ );
xnor g304 ( new_n647_, new_n646_, keyIn_0_126 );
xor g305 ( new_n648_, new_n575_, keyIn_0_98 );
nand g306 ( new_n649_, new_n647_, new_n648_ );
xnor g307 ( new_n650_, new_n649_, keyIn_0_132 );
or g308 ( new_n651_, new_n650_, new_n491_ );
xor g309 ( new_n652_, new_n651_, keyIn_0_149 );
nand g310 ( new_n653_, new_n650_, new_n491_ );
xnor g311 ( new_n654_, new_n653_, keyIn_0_150 );
nand g312 ( new_n655_, new_n652_, new_n654_ );
xnor g313 ( new_n656_, new_n655_, new_n641_ );
not g314 ( new_n657_, keyIn_0_204 );
nor g315 ( new_n658_, new_n583_, new_n514_ );
or g316 ( new_n659_, new_n658_, keyIn_0_172 );
nand g317 ( new_n660_, new_n658_, keyIn_0_172 );
nand g318 ( new_n661_, new_n556_, N116 );
xor g319 ( new_n662_, new_n575_, keyIn_0_99 );
nand g320 ( new_n663_, new_n565_, N146 );
nand g321 ( new_n664_, new_n662_, new_n661_, new_n663_ );
xor g322 ( new_n665_, new_n664_, keyIn_0_133 );
nor g323 ( new_n666_, new_n665_, N189 );
not g324 ( new_n667_, new_n666_ );
not g325 ( new_n668_, N195 );
not g326 ( new_n669_, keyIn_0_134 );
nand g327 ( new_n670_, new_n565_, N149 );
nand g328 ( new_n671_, new_n670_, keyIn_0_112 );
not g329 ( new_n672_, keyIn_0_112 );
nand g330 ( new_n673_, new_n565_, new_n672_, N149 );
nand g331 ( new_n674_, new_n671_, new_n673_ );
not g332 ( new_n675_, keyIn_0_113 );
nand g333 ( new_n676_, new_n556_, new_n675_, N121 );
xnor g334 ( new_n677_, new_n575_, keyIn_0_100 );
nand g335 ( new_n678_, new_n556_, N121 );
nand g336 ( new_n679_, new_n678_, keyIn_0_113 );
and g337 ( new_n680_, new_n679_, new_n677_ );
nand g338 ( new_n681_, new_n680_, new_n669_, new_n674_, new_n676_ );
nand g339 ( new_n682_, new_n674_, new_n679_, new_n676_, new_n677_ );
nand g340 ( new_n683_, new_n682_, keyIn_0_134 );
nand g341 ( new_n684_, new_n681_, new_n683_, new_n668_ );
nand g342 ( new_n685_, new_n684_, keyIn_0_152 );
not g343 ( new_n686_, keyIn_0_152 );
nand g344 ( new_n687_, new_n681_, new_n683_, new_n686_, new_n668_ );
nand g345 ( new_n688_, new_n685_, new_n687_ );
nand g346 ( new_n689_, new_n659_, new_n667_, new_n660_, new_n688_ );
nand g347 ( new_n690_, new_n689_, keyIn_0_197 );
nand g348 ( new_n691_, new_n665_, N189 );
and g349 ( new_n692_, new_n690_, new_n691_ );
not g350 ( new_n693_, keyIn_0_169 );
nand g351 ( new_n694_, new_n681_, new_n683_ );
nand g352 ( new_n695_, new_n694_, N195 );
nand g353 ( new_n696_, new_n695_, new_n693_ );
nand g354 ( new_n697_, new_n694_, keyIn_0_169, N195 );
nand g355 ( new_n698_, new_n696_, new_n697_ );
nand g356 ( new_n699_, new_n698_, new_n667_ );
nand g357 ( new_n700_, new_n699_, keyIn_0_196 );
not g358 ( new_n701_, keyIn_0_196 );
nand g359 ( new_n702_, new_n698_, new_n701_, new_n667_ );
nand g360 ( new_n703_, new_n700_, new_n702_ );
not g361 ( new_n704_, keyIn_0_197 );
nand g362 ( new_n705_, new_n606_, new_n704_, new_n667_, new_n688_ );
and g363 ( new_n706_, new_n703_, new_n705_ );
nand g364 ( new_n707_, new_n688_, new_n585_, N261, new_n587_ );
nor g365 ( new_n708_, new_n707_, new_n666_ );
xnor g366 ( new_n709_, new_n708_, keyIn_0_176 );
nand g367 ( new_n710_, new_n709_, new_n706_, new_n692_ );
nand g368 ( new_n711_, new_n710_, new_n657_ );
nand g369 ( new_n712_, new_n709_, new_n706_, keyIn_0_204, new_n692_ );
nand g370 ( new_n713_, new_n711_, new_n712_ );
not g371 ( new_n714_, new_n713_ );
nand g372 ( new_n715_, new_n656_, keyIn_0_211, new_n714_ );
not g373 ( new_n716_, keyIn_0_211 );
nand g374 ( new_n717_, new_n656_, new_n714_ );
nand g375 ( new_n718_, new_n717_, new_n716_ );
not g376 ( new_n719_, new_n656_ );
nand g377 ( new_n720_, new_n719_, new_n713_ );
nand g378 ( new_n721_, new_n718_, new_n715_, new_n720_ );
or g379 ( new_n722_, new_n721_, keyIn_0_216 );
nand g380 ( new_n723_, new_n721_, keyIn_0_216 );
nand g381 ( new_n724_, new_n722_, N219, new_n723_ );
nand g382 ( new_n725_, new_n724_, new_n640_ );
nand g383 ( new_n726_, new_n722_, keyIn_0_220, N219, new_n723_ );
nand g384 ( new_n727_, new_n725_, new_n726_ );
not g385 ( new_n728_, N210 );
nor g386 ( new_n729_, new_n430_, new_n728_ );
or g387 ( new_n730_, new_n729_, keyIn_0_34 );
nand g388 ( new_n731_, keyIn_0_34, N106, N210 );
nand g389 ( new_n732_, new_n730_, new_n731_ );
nand g390 ( new_n733_, new_n727_, new_n639_, new_n732_ );
nand g391 ( new_n734_, new_n727_, new_n732_ );
nand g392 ( new_n735_, new_n734_, keyIn_0_226 );
nand g393 ( new_n736_, new_n719_, N228 );
xnor g394 ( new_n737_, new_n651_, keyIn_0_149 );
nand g395 ( new_n738_, new_n737_, N237 );
xnor g396 ( new_n739_, new_n738_, keyIn_0_186 );
nand g397 ( new_n740_, new_n736_, new_n739_ );
nor g398 ( new_n741_, new_n740_, keyIn_0_205 );
or g399 ( new_n742_, new_n650_, new_n611_ );
nand g400 ( new_n743_, new_n628_, N183 );
xnor g401 ( new_n744_, new_n743_, keyIn_0_121 );
nand g402 ( new_n745_, new_n742_, new_n744_ );
xor g403 ( new_n746_, new_n745_, keyIn_0_166 );
and g404 ( new_n747_, new_n740_, keyIn_0_205 );
nor g405 ( new_n748_, new_n747_, new_n741_, new_n746_ );
nand g406 ( new_n749_, new_n735_, new_n733_, new_n748_ );
nand g407 ( new_n750_, new_n749_, new_n638_ );
nand g408 ( new_n751_, new_n735_, keyIn_0_233, new_n733_, new_n748_ );
nand g409 ( new_n752_, new_n750_, new_n751_ );
nand g410 ( new_n753_, new_n752_, keyIn_0_238 );
not g411 ( new_n754_, keyIn_0_238 );
nand g412 ( new_n755_, new_n750_, new_n754_, new_n751_ );
nand g413 ( new_n756_, new_n753_, new_n755_ );
nand g414 ( new_n757_, new_n756_, new_n637_ );
nand g415 ( new_n758_, new_n753_, keyIn_0_245, new_n755_ );
nand g416 ( N863, new_n757_, new_n758_ );
not g417 ( new_n760_, keyIn_0_221 );
xnor g418 ( new_n761_, new_n707_, keyIn_0_175 );
nand g419 ( new_n762_, new_n606_, keyIn_0_195, new_n688_ );
not g420 ( new_n763_, keyIn_0_195 );
nand g421 ( new_n764_, new_n606_, new_n688_ );
nand g422 ( new_n765_, new_n764_, new_n763_ );
xor g423 ( new_n766_, new_n698_, keyIn_0_189 );
nand g424 ( new_n767_, new_n761_, new_n765_, new_n762_, new_n766_ );
xnor g425 ( new_n768_, new_n767_, keyIn_0_206 );
nand g426 ( new_n769_, new_n667_, new_n691_ );
xnor g427 ( new_n770_, new_n769_, keyIn_0_167 );
and g428 ( new_n771_, new_n768_, new_n770_ );
nand g429 ( new_n772_, new_n771_, keyIn_0_212 );
or g430 ( new_n773_, new_n771_, keyIn_0_212 );
or g431 ( new_n774_, new_n768_, new_n770_ );
nand g432 ( new_n775_, new_n773_, N219, new_n772_, new_n774_ );
nand g433 ( new_n776_, new_n775_, new_n760_ );
or g434 ( new_n777_, new_n775_, new_n760_ );
nand g435 ( new_n778_, N111, N210 );
xor g436 ( new_n779_, new_n778_, keyIn_0_35 );
nand g437 ( new_n780_, new_n777_, new_n776_, new_n779_ );
xnor g438 ( new_n781_, new_n780_, keyIn_0_227 );
nand g439 ( new_n782_, new_n770_, N228 );
not g440 ( new_n783_, new_n782_ );
nor g441 ( new_n784_, new_n783_, keyIn_0_187 );
not g442 ( new_n785_, N237 );
nor g443 ( new_n786_, new_n691_, new_n785_ );
nand g444 ( new_n787_, new_n786_, keyIn_0_188 );
nand g445 ( new_n788_, new_n628_, N189 );
or g446 ( new_n789_, new_n786_, keyIn_0_188 );
nand g447 ( new_n790_, new_n789_, new_n787_, new_n788_ );
nor g448 ( new_n791_, new_n784_, new_n790_ );
nand g449 ( new_n792_, new_n665_, N246 );
xnor g450 ( new_n793_, new_n792_, keyIn_0_151 );
nand g451 ( new_n794_, N255, N259 );
nand g452 ( new_n795_, new_n794_, keyIn_0_36 );
not g453 ( new_n796_, keyIn_0_36 );
nand g454 ( new_n797_, new_n796_, N255, N259 );
nand g455 ( new_n798_, new_n795_, new_n797_ );
nand g456 ( new_n799_, new_n793_, new_n798_ );
xnor g457 ( new_n800_, new_n799_, keyIn_0_168 );
nand g458 ( new_n801_, new_n783_, keyIn_0_187 );
nand g459 ( new_n802_, new_n781_, new_n791_, new_n800_, new_n801_ );
xnor g460 ( new_n803_, new_n802_, keyIn_0_239 );
xor g461 ( N864, new_n803_, keyIn_0_246 );
not g462 ( new_n805_, keyIn_0_228 );
not g463 ( new_n806_, keyIn_0_222 );
not g464 ( new_n807_, keyIn_0_217 );
not g465 ( new_n808_, keyIn_0_213 );
nand g466 ( new_n809_, new_n688_, new_n695_ );
xnor g467 ( new_n810_, new_n809_, keyIn_0_170 );
nand g468 ( new_n811_, new_n588_, N261 );
xnor g469 ( new_n812_, new_n811_, keyIn_0_174 );
nor g470 ( new_n813_, new_n812_, new_n606_ );
xnor g471 ( new_n814_, new_n813_, keyIn_0_207 );
nor g472 ( new_n815_, new_n814_, new_n810_ );
or g473 ( new_n816_, new_n815_, new_n808_ );
nand g474 ( new_n817_, new_n814_, new_n810_ );
nand g475 ( new_n818_, new_n817_, keyIn_0_214 );
or g476 ( new_n819_, new_n817_, keyIn_0_214 );
nand g477 ( new_n820_, new_n815_, new_n808_ );
nand g478 ( new_n821_, new_n816_, new_n819_, new_n818_, new_n820_ );
or g479 ( new_n822_, new_n821_, new_n807_ );
nand g480 ( new_n823_, new_n821_, new_n807_ );
nand g481 ( new_n824_, new_n822_, N219, new_n823_ );
or g482 ( new_n825_, new_n824_, new_n806_ );
nand g483 ( new_n826_, N116, N210 );
nand g484 ( new_n827_, new_n824_, new_n806_ );
nand g485 ( new_n828_, new_n825_, new_n826_, new_n827_ );
or g486 ( new_n829_, new_n828_, new_n805_ );
nand g487 ( new_n830_, new_n828_, new_n805_ );
not g488 ( new_n831_, keyIn_0_208 );
nand g489 ( new_n832_, new_n810_, N228 );
or g490 ( new_n833_, new_n832_, keyIn_0_190 );
nand g491 ( new_n834_, new_n698_, N237 );
xnor g492 ( new_n835_, new_n834_, keyIn_0_191 );
nand g493 ( new_n836_, new_n832_, keyIn_0_190 );
nand g494 ( new_n837_, new_n833_, new_n835_, new_n836_ );
nor g495 ( new_n838_, new_n837_, new_n831_ );
and g496 ( new_n839_, new_n837_, new_n831_ );
and g497 ( new_n840_, new_n694_, N246 );
nand g498 ( new_n841_, new_n840_, keyIn_0_153 );
and g499 ( new_n842_, N255, N260 );
or g500 ( new_n843_, new_n842_, keyIn_0_37 );
nand g501 ( new_n844_, keyIn_0_37, N255, N260 );
nand g502 ( new_n845_, new_n843_, new_n844_ );
or g503 ( new_n846_, new_n840_, keyIn_0_153 );
nand g504 ( new_n847_, new_n846_, new_n841_, new_n845_ );
nor g505 ( new_n848_, new_n847_, keyIn_0_171 );
nand g506 ( new_n849_, new_n628_, N195 );
nand g507 ( new_n850_, new_n847_, keyIn_0_171 );
nand g508 ( new_n851_, new_n850_, new_n849_ );
nor g509 ( new_n852_, new_n839_, new_n838_, new_n848_, new_n851_ );
nand g510 ( new_n853_, new_n829_, new_n830_, new_n852_ );
xor g511 ( new_n854_, new_n853_, keyIn_0_240 );
xnor g512 ( N865, new_n854_, keyIn_0_247 );
not g513 ( new_n856_, keyIn_0_225 );
or g514 ( new_n857_, new_n569_, new_n524_ );
or g515 ( new_n858_, new_n857_, keyIn_0_80 );
nand g516 ( new_n859_, new_n857_, keyIn_0_80 );
nand g517 ( new_n860_, new_n858_, new_n572_, new_n859_ );
xor g518 ( new_n861_, new_n860_, keyIn_0_92 );
nand g519 ( new_n862_, new_n522_, N55, new_n559_ );
xor g520 ( new_n863_, new_n862_, keyIn_0_79 );
nand g521 ( new_n864_, new_n863_, N146 );
xnor g522 ( new_n865_, new_n864_, keyIn_0_91 );
nand g523 ( new_n866_, new_n861_, new_n865_ );
xnor g524 ( new_n867_, new_n866_, keyIn_0_107 );
nand g525 ( new_n868_, new_n556_, N96 );
or g526 ( new_n869_, new_n868_, keyIn_0_106 );
nand g527 ( new_n870_, new_n868_, keyIn_0_106 );
nand g528 ( new_n871_, N51, N138 );
xnor g529 ( new_n872_, new_n871_, keyIn_0_20 );
nand g530 ( new_n873_, new_n867_, new_n869_, new_n870_, new_n872_ );
xnor g531 ( new_n874_, new_n873_, keyIn_0_130 );
nor g532 ( new_n875_, new_n874_, N165 );
xnor g533 ( new_n876_, new_n875_, keyIn_0_144 );
not g534 ( new_n877_, keyIn_0_131 );
nand g535 ( new_n878_, new_n556_, N101 );
and g536 ( new_n879_, N17, N138 );
or g537 ( new_n880_, new_n879_, keyIn_0_21 );
nand g538 ( new_n881_, keyIn_0_21, N17, N138 );
nand g539 ( new_n882_, new_n880_, new_n881_ );
nand g540 ( new_n883_, new_n878_, new_n882_ );
xnor g541 ( new_n884_, new_n883_, keyIn_0_124 );
xor g542 ( new_n885_, new_n860_, keyIn_0_94 );
nand g543 ( new_n886_, new_n863_, N149 );
xnor g544 ( new_n887_, new_n886_, keyIn_0_93 );
nand g545 ( new_n888_, new_n885_, new_n887_ );
xor g546 ( new_n889_, new_n888_, keyIn_0_108 );
nand g547 ( new_n890_, new_n889_, new_n884_ );
xnor g548 ( new_n891_, new_n890_, new_n877_ );
nor g549 ( new_n892_, new_n891_, N171 );
xor g550 ( new_n893_, new_n892_, keyIn_0_145 );
and g551 ( new_n894_, new_n893_, new_n876_ );
nand g552 ( new_n895_, new_n713_, new_n654_ );
xnor g553 ( new_n896_, new_n737_, keyIn_0_185 );
nand g554 ( new_n897_, new_n895_, new_n896_ );
not g555 ( new_n898_, keyIn_0_125 );
and g556 ( new_n899_, new_n556_, N106 );
not g557 ( new_n900_, new_n899_ );
or g558 ( new_n901_, new_n900_, keyIn_0_109 );
nand g559 ( new_n902_, N138, N152 );
nand g560 ( new_n903_, new_n900_, keyIn_0_109 );
nand g561 ( new_n904_, new_n901_, new_n902_, new_n903_ );
or g562 ( new_n905_, new_n904_, new_n898_ );
xnor g563 ( new_n906_, new_n860_, keyIn_0_96 );
nand g564 ( new_n907_, new_n863_, N153 );
xnor g565 ( new_n908_, new_n907_, keyIn_0_95 );
nand g566 ( new_n909_, new_n906_, new_n908_ );
xnor g567 ( new_n910_, new_n909_, keyIn_0_110 );
nand g568 ( new_n911_, new_n904_, new_n898_ );
nand g569 ( new_n912_, new_n905_, new_n910_, new_n911_ );
nor g570 ( new_n913_, new_n912_, N177 );
xor g571 ( new_n914_, new_n913_, keyIn_0_147 );
nand g572 ( new_n915_, new_n897_, new_n856_, new_n894_, new_n914_ );
nand g573 ( new_n916_, new_n897_, new_n894_, new_n914_ );
nand g574 ( new_n917_, new_n916_, keyIn_0_225 );
nand g575 ( new_n918_, new_n912_, N177 );
xnor g576 ( new_n919_, new_n918_, keyIn_0_146 );
xnor g577 ( new_n920_, new_n919_, keyIn_0_162 );
nand g578 ( new_n921_, new_n894_, new_n920_ );
or g579 ( new_n922_, new_n921_, keyIn_0_200 );
nand g580 ( new_n923_, new_n921_, keyIn_0_200 );
and g581 ( new_n924_, new_n891_, N171 );
nand g582 ( new_n925_, new_n876_, new_n924_ );
nor g583 ( new_n926_, new_n925_, keyIn_0_199 );
and g584 ( new_n927_, new_n925_, keyIn_0_199 );
nand g585 ( new_n928_, new_n874_, N165 );
xor g586 ( new_n929_, new_n928_, keyIn_0_143 );
xnor g587 ( new_n930_, new_n929_, keyIn_0_179 );
nor g588 ( new_n931_, new_n930_, new_n927_, new_n926_ );
and g589 ( new_n932_, new_n922_, new_n923_, new_n931_ );
nand g590 ( new_n933_, new_n917_, new_n915_, new_n932_ );
nand g591 ( new_n934_, new_n556_, N91 );
not g592 ( new_n935_, new_n860_ );
or g593 ( new_n936_, new_n935_, keyIn_0_90 );
nand g594 ( new_n937_, N8, N138 );
nand g595 ( new_n938_, new_n863_, N143 );
nand g596 ( new_n939_, new_n938_, keyIn_0_89 );
nand g597 ( new_n940_, new_n935_, keyIn_0_90 );
or g598 ( new_n941_, new_n938_, keyIn_0_89 );
and g599 ( new_n942_, new_n940_, new_n939_, new_n941_ );
nand g600 ( new_n943_, new_n942_, new_n934_, new_n936_, new_n937_ );
nor g601 ( new_n944_, new_n943_, N159 );
xnor g602 ( new_n945_, new_n944_, keyIn_0_141 );
and g603 ( new_n946_, new_n933_, new_n945_ );
nand g604 ( new_n947_, new_n946_, keyIn_0_235 );
nand g605 ( new_n948_, new_n943_, N159 );
xnor g606 ( new_n949_, new_n948_, keyIn_0_140 );
xor g607 ( new_n950_, new_n949_, keyIn_0_177 );
or g608 ( new_n951_, new_n946_, keyIn_0_235 );
nand g609 ( new_n952_, new_n951_, new_n947_, new_n950_ );
xor g610 ( new_n953_, new_n952_, keyIn_0_241 );
xnor g611 ( N866, new_n953_, keyIn_0_248 );
nand g612 ( new_n955_, new_n914_, new_n919_ );
xor g613 ( new_n956_, new_n955_, keyIn_0_163 );
nand g614 ( new_n957_, new_n897_, new_n956_ );
xor g615 ( new_n958_, new_n957_, keyIn_0_219 );
not g616 ( new_n959_, keyIn_0_218 );
or g617 ( new_n960_, new_n897_, new_n956_ );
or g618 ( new_n961_, new_n960_, new_n959_ );
nand g619 ( new_n962_, new_n960_, new_n959_ );
nand g620 ( new_n963_, new_n958_, new_n961_, N219, new_n962_ );
and g621 ( new_n964_, new_n956_, N228 );
nand g622 ( new_n965_, new_n964_, keyIn_0_184 );
or g623 ( new_n966_, new_n964_, keyIn_0_184 );
and g624 ( new_n967_, new_n920_, N237 );
not g625 ( new_n968_, keyIn_0_164 );
and g626 ( new_n969_, new_n912_, N246 );
nand g627 ( new_n970_, new_n969_, keyIn_0_148 );
nand g628 ( new_n971_, new_n628_, N177 );
xnor g629 ( new_n972_, new_n971_, keyIn_0_120 );
or g630 ( new_n973_, new_n969_, keyIn_0_148 );
nand g631 ( new_n974_, new_n973_, new_n970_, new_n972_ );
nor g632 ( new_n975_, new_n974_, new_n968_ );
nor g633 ( new_n976_, new_n429_, new_n728_ );
and g634 ( new_n977_, new_n974_, new_n968_ );
nor g635 ( new_n978_, new_n967_, new_n975_, new_n976_, new_n977_ );
nand g636 ( new_n979_, new_n963_, new_n965_, new_n966_, new_n978_ );
xnor g637 ( new_n980_, new_n979_, keyIn_0_244 );
xnor g638 ( N874, new_n980_, keyIn_0_253 );
not g639 ( new_n982_, keyIn_0_251 );
not g640 ( new_n983_, keyIn_0_249 );
not g641 ( new_n984_, keyIn_0_236 );
not g642 ( new_n985_, new_n949_ );
nand g643 ( new_n986_, new_n985_, new_n945_ );
xor g644 ( new_n987_, new_n986_, keyIn_0_158 );
nand g645 ( new_n988_, new_n933_, new_n987_ );
nand g646 ( new_n989_, new_n988_, keyIn_0_230 );
not g647 ( new_n990_, keyIn_0_230 );
nand g648 ( new_n991_, new_n933_, new_n990_, new_n987_ );
nand g649 ( new_n992_, new_n989_, new_n991_ );
or g650 ( new_n993_, new_n933_, new_n987_ );
nand g651 ( new_n994_, new_n992_, new_n984_, new_n993_ );
nand g652 ( new_n995_, new_n992_, new_n993_ );
nand g653 ( new_n996_, new_n995_, keyIn_0_236 );
nand g654 ( new_n997_, new_n996_, N219, new_n994_ );
nor g655 ( new_n998_, new_n573_, new_n728_ );
xor g656 ( new_n999_, new_n998_, keyIn_0_75 );
nand g657 ( new_n1000_, new_n997_, new_n999_ );
nand g658 ( new_n1001_, new_n1000_, new_n983_ );
nand g659 ( new_n1002_, new_n997_, keyIn_0_249, new_n999_ );
nand g660 ( new_n1003_, new_n1001_, new_n1002_ );
not g661 ( new_n1004_, keyIn_0_201 );
nand g662 ( new_n1005_, new_n987_, N228 );
or g663 ( new_n1006_, new_n1005_, keyIn_0_178 );
nand g664 ( new_n1007_, new_n949_, N237 );
nand g665 ( new_n1008_, new_n1005_, keyIn_0_178 );
nand g666 ( new_n1009_, new_n1006_, new_n1007_, new_n1008_ );
nor g667 ( new_n1010_, new_n1009_, new_n1004_ );
and g668 ( new_n1011_, new_n1009_, new_n1004_ );
and g669 ( new_n1012_, new_n943_, N246 );
nand g670 ( new_n1013_, new_n1012_, keyIn_0_142 );
or g671 ( new_n1014_, new_n1012_, keyIn_0_142 );
nand g672 ( new_n1015_, new_n628_, N159 );
xnor g673 ( new_n1016_, new_n1015_, keyIn_0_117 );
nand g674 ( new_n1017_, new_n1014_, new_n1013_, new_n1016_ );
nor g675 ( new_n1018_, new_n1011_, new_n1010_, new_n1017_ );
nand g676 ( new_n1019_, new_n1003_, new_n1018_ );
nand g677 ( new_n1020_, new_n1019_, new_n982_ );
nand g678 ( new_n1021_, new_n1003_, keyIn_0_251, new_n1018_ );
nand g679 ( new_n1022_, new_n1020_, new_n1021_ );
nand g680 ( new_n1023_, new_n1022_, keyIn_0_254 );
not g681 ( new_n1024_, keyIn_0_254 );
nand g682 ( new_n1025_, new_n1020_, new_n1024_, new_n1021_ );
nand g683 ( N878, new_n1023_, new_n1025_ );
not g684 ( new_n1027_, keyIn_0_255 );
not g685 ( new_n1028_, keyIn_0_224 );
nand g686 ( new_n1029_, new_n897_, new_n893_, new_n914_ );
or g687 ( new_n1030_, new_n1029_, new_n1028_ );
nand g688 ( new_n1031_, new_n1029_, new_n1028_ );
nand g689 ( new_n1032_, new_n893_, new_n920_ );
nor g690 ( new_n1033_, new_n1032_, keyIn_0_198 );
xnor g691 ( new_n1034_, new_n924_, keyIn_0_181 );
and g692 ( new_n1035_, new_n1032_, keyIn_0_198 );
nor g693 ( new_n1036_, new_n1035_, new_n1033_, new_n1034_ );
nand g694 ( new_n1037_, new_n1030_, new_n1031_, new_n1036_ );
nand g695 ( new_n1038_, new_n929_, new_n876_ );
xnor g696 ( new_n1039_, new_n1038_, keyIn_0_159 );
nand g697 ( new_n1040_, new_n1037_, new_n1039_ );
or g698 ( new_n1041_, new_n1037_, new_n1039_ );
nand g699 ( new_n1042_, new_n1041_, N219, new_n1040_ );
xnor g700 ( new_n1043_, new_n1042_, keyIn_0_242 );
and g701 ( new_n1044_, N91, N210 );
or g702 ( new_n1045_, new_n1044_, keyIn_0_32 );
nand g703 ( new_n1046_, keyIn_0_32, N91, N210 );
nand g704 ( new_n1047_, new_n1045_, new_n1046_ );
nand g705 ( new_n1048_, new_n1043_, new_n1047_ );
xor g706 ( new_n1049_, new_n1048_, keyIn_0_250 );
not g707 ( new_n1050_, keyIn_0_202 );
nand g708 ( new_n1051_, new_n1039_, keyIn_0_180, N228 );
or g709 ( new_n1052_, new_n929_, new_n785_ );
not g710 ( new_n1053_, keyIn_0_180 );
nand g711 ( new_n1054_, new_n1039_, N228 );
nand g712 ( new_n1055_, new_n1054_, new_n1053_ );
nand g713 ( new_n1056_, new_n1055_, new_n1051_, new_n1052_ );
nor g714 ( new_n1057_, new_n1056_, new_n1050_ );
and g715 ( new_n1058_, new_n1056_, new_n1050_ );
nand g716 ( new_n1059_, new_n628_, N165 );
xor g717 ( new_n1060_, new_n1059_, keyIn_0_118 );
and g718 ( new_n1061_, new_n874_, N246 );
nor g719 ( new_n1062_, new_n1058_, new_n1057_, new_n1060_, new_n1061_ );
nand g720 ( new_n1063_, new_n1049_, new_n1062_ );
xnor g721 ( N879, new_n1063_, new_n1027_ );
not g722 ( new_n1065_, keyIn_0_237 );
not g723 ( new_n1066_, new_n924_ );
nand g724 ( new_n1067_, new_n893_, new_n1066_ );
xor g725 ( new_n1068_, new_n1067_, keyIn_0_160 );
nand g726 ( new_n1069_, new_n897_, new_n914_ );
xnor g727 ( new_n1070_, new_n920_, keyIn_0_183 );
nand g728 ( new_n1071_, new_n1069_, new_n1070_ );
nor g729 ( new_n1072_, new_n1071_, new_n1068_ );
or g730 ( new_n1073_, new_n1072_, keyIn_0_231 );
nand g731 ( new_n1074_, new_n1071_, new_n1068_ );
nand g732 ( new_n1075_, new_n1074_, keyIn_0_232 );
or g733 ( new_n1076_, new_n1074_, keyIn_0_232 );
nand g734 ( new_n1077_, new_n1072_, keyIn_0_231 );
nand g735 ( new_n1078_, new_n1073_, new_n1076_, new_n1075_, new_n1077_ );
or g736 ( new_n1079_, new_n1078_, new_n1065_ );
nand g737 ( new_n1080_, new_n1078_, new_n1065_ );
nand g738 ( new_n1081_, new_n1079_, N219, new_n1080_ );
or g739 ( new_n1082_, new_n1081_, keyIn_0_243 );
nand g740 ( new_n1083_, new_n1081_, keyIn_0_243 );
nand g741 ( new_n1084_, new_n1068_, N228 );
nand g742 ( new_n1085_, new_n924_, N237 );
xnor g743 ( new_n1086_, new_n1085_, keyIn_0_182 );
and g744 ( new_n1087_, new_n1084_, new_n1086_ );
and g745 ( new_n1088_, new_n1087_, keyIn_0_203 );
nor g746 ( new_n1089_, new_n1087_, keyIn_0_203 );
nand g747 ( new_n1090_, new_n891_, N246 );
nand g748 ( new_n1091_, new_n628_, N171 );
xnor g749 ( new_n1092_, new_n1091_, keyIn_0_119 );
and g750 ( new_n1093_, new_n1090_, new_n1092_ );
nand g751 ( new_n1094_, new_n1093_, keyIn_0_161 );
or g752 ( new_n1095_, new_n1093_, keyIn_0_161 );
nand g753 ( new_n1096_, N96, N210 );
xor g754 ( new_n1097_, new_n1096_, keyIn_0_33 );
nand g755 ( new_n1098_, new_n1095_, new_n1094_, new_n1097_ );
nor g756 ( new_n1099_, new_n1088_, new_n1089_, new_n1098_ );
nand g757 ( new_n1100_, new_n1082_, new_n1083_, new_n1099_ );
xnor g758 ( N880, new_n1100_, keyIn_0_252 );
endmodule