module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n390_, new_n743_, new_n366_, new_n566_, new_n641_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n451_, new_n489_, new_n424_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n552_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n626_, new_n716_, new_n701_, new_n257_, new_n481_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n634_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n498_, new_n492_, new_n496_, new_n650_, new_n708_, new_n750_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n447_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n739_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n696_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n762_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n577_, new_n374_, new_n376_, new_n380_, new_n747_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n407_, new_n666_, new_n480_, new_n625_, new_n736_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n755_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n307_, new_n597_, new_n408_, new_n470_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n760_, new_n627_, new_n704_, new_n567_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n709_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n757_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n536_, new_n464_, new_n573_, new_n405_;

and g000 ( N388, N29, N42, N75 );
and g001 ( N389, N29, N36, N80 );
nand g002 ( new_n217_, N29, N36, N42 );
not g003 ( N390, new_n217_ );
and g004 ( N391, N85, N86 );
and g005 ( N418, N1, N8, N13, N17 );
and g006 ( new_n221_, N1, N13, N17, N26 );
nand g007 ( N419, new_n221_, new_n217_ );
nand g008 ( N420, N59, N75, N80 );
nand g009 ( N421, N36, N59, N80 );
nand g010 ( N422, N36, N42, N59 );
not g011 ( new_n226_, N90 );
nor g012 ( new_n227_, N87, N88 );
nor g013 ( N423, new_n227_, new_n226_ );
nand g014 ( N446, new_n221_, N390 );
not g015 ( new_n230_, keyIn_0_0 );
nand g016 ( new_n231_, new_n230_, N1, N26, N51 );
nand g017 ( new_n232_, N1, N26, N51 );
nand g018 ( new_n233_, new_n232_, keyIn_0_0 );
nand g019 ( N447, new_n233_, new_n231_ );
not g020 ( new_n235_, N29 );
not g021 ( new_n236_, N68 );
nand g022 ( new_n237_, N1, N8, N13, N55 );
nor g023 ( N448, new_n237_, new_n235_, new_n236_ );
not g024 ( new_n239_, N59 );
nor g025 ( new_n240_, new_n237_, new_n239_, new_n236_ );
and g026 ( N449, new_n240_, N74 );
not g027 ( new_n242_, N89 );
nor g028 ( N450, new_n227_, new_n242_ );
xnor g029 ( new_n244_, N101, N106 );
xnor g030 ( new_n245_, new_n244_, keyIn_0_13 );
not g031 ( new_n246_, new_n245_ );
xor g032 ( new_n247_, N91, N96 );
xnor g033 ( new_n248_, new_n247_, keyIn_0_12 );
nor g034 ( new_n249_, new_n246_, new_n248_ );
xnor g035 ( new_n250_, new_n249_, keyIn_0_28 );
nand g036 ( new_n251_, new_n246_, new_n248_ );
xor g037 ( new_n252_, new_n251_, keyIn_0_23 );
nand g038 ( new_n253_, new_n252_, new_n250_ );
xnor g039 ( new_n254_, new_n253_, keyIn_0_37 );
xnor g040 ( new_n255_, new_n254_, N130 );
xor g041 ( new_n256_, N121, N126 );
xnor g042 ( new_n257_, new_n256_, keyIn_0_15 );
xnor g043 ( new_n258_, N111, N116 );
xnor g044 ( new_n259_, new_n258_, keyIn_0_14 );
not g045 ( new_n260_, new_n259_ );
nor g046 ( new_n261_, new_n260_, new_n257_ );
xor g047 ( new_n262_, new_n261_, keyIn_0_29 );
nand g048 ( new_n263_, new_n260_, new_n257_ );
xnor g049 ( new_n264_, new_n263_, keyIn_0_24 );
nand g050 ( new_n265_, new_n262_, new_n264_ );
xnor g051 ( new_n266_, new_n265_, keyIn_0_38 );
xnor g052 ( new_n267_, new_n266_, N135 );
xnor g053 ( N767, new_n267_, new_n255_ );
not g054 ( new_n269_, keyIn_0_27 );
xor g055 ( new_n270_, N183, N189 );
xnor g056 ( new_n271_, new_n270_, keyIn_0_20 );
xnor g057 ( new_n272_, N195, N201 );
xnor g058 ( new_n273_, new_n272_, keyIn_0_21 );
or g059 ( new_n274_, new_n271_, new_n273_ );
or g060 ( new_n275_, new_n274_, new_n269_ );
nand g061 ( new_n276_, new_n271_, new_n273_ );
or g062 ( new_n277_, new_n276_, keyIn_0_36 );
nand g063 ( new_n278_, new_n276_, keyIn_0_36 );
nand g064 ( new_n279_, new_n274_, new_n269_ );
nand g065 ( new_n280_, new_n275_, new_n277_, new_n278_, new_n279_ );
xnor g066 ( new_n281_, new_n280_, keyIn_0_50 );
xnor g067 ( new_n282_, new_n281_, N207 );
xor g068 ( new_n283_, N171, N177 );
xnor g069 ( new_n284_, new_n283_, keyIn_0_19 );
xnor g070 ( new_n285_, N159, N165 );
xnor g071 ( new_n286_, new_n285_, keyIn_0_18 );
nor g072 ( new_n287_, new_n284_, new_n286_ );
xnor g073 ( new_n288_, new_n287_, keyIn_0_35 );
nand g074 ( new_n289_, new_n284_, new_n286_ );
xor g075 ( new_n290_, new_n289_, keyIn_0_26 );
nand g076 ( new_n291_, new_n290_, new_n288_ );
xor g077 ( new_n292_, new_n291_, keyIn_0_49 );
xnor g078 ( new_n293_, new_n292_, N130 );
xnor g079 ( N768, new_n293_, new_n282_ );
not g080 ( new_n295_, keyIn_0_70 );
not g081 ( new_n296_, keyIn_0_61 );
not g082 ( new_n297_, keyIn_0_34 );
not g083 ( new_n298_, keyIn_0_22 );
not g084 ( new_n299_, keyIn_0_8 );
nand g085 ( new_n300_, N447, new_n299_ );
nand g086 ( new_n301_, new_n233_, keyIn_0_8, new_n231_ );
nand g087 ( new_n302_, new_n300_, new_n301_ );
nand g088 ( new_n303_, new_n302_, new_n298_ );
nand g089 ( new_n304_, new_n300_, keyIn_0_22, new_n301_ );
nand g090 ( new_n305_, new_n303_, new_n304_ );
nand g091 ( new_n306_, N59, N156 );
xnor g092 ( new_n307_, new_n306_, keyIn_0_5 );
nand g093 ( new_n308_, new_n305_, new_n297_, N17, new_n307_ );
nand g094 ( new_n309_, new_n305_, N17, new_n307_ );
nand g095 ( new_n310_, new_n309_, keyIn_0_34 );
nand g096 ( new_n311_, new_n310_, new_n308_ );
nand g097 ( new_n312_, new_n311_, keyIn_0_44, N1 );
not g098 ( new_n313_, keyIn_0_44 );
nand g099 ( new_n314_, new_n311_, N1 );
nand g100 ( new_n315_, new_n314_, new_n313_ );
nand g101 ( new_n316_, new_n315_, new_n312_ );
nand g102 ( new_n317_, new_n316_, new_n296_, N153 );
nand g103 ( new_n318_, new_n316_, N153 );
nand g104 ( new_n319_, new_n318_, keyIn_0_61 );
not g105 ( new_n320_, keyIn_0_39 );
not g106 ( new_n321_, new_n306_ );
not g107 ( new_n322_, keyIn_0_17 );
not g108 ( new_n323_, keyIn_0_6 );
nor g109 ( new_n324_, N17, N42 );
xnor g110 ( new_n325_, new_n324_, new_n323_ );
not g111 ( new_n326_, keyIn_0_7 );
nand g112 ( new_n327_, N17, N42 );
xnor g113 ( new_n328_, new_n327_, new_n326_ );
nand g114 ( new_n329_, new_n325_, new_n322_, new_n328_ );
nand g115 ( new_n330_, new_n325_, new_n328_ );
nand g116 ( new_n331_, new_n330_, keyIn_0_17 );
nand g117 ( new_n332_, new_n331_, new_n329_ );
nand g118 ( new_n333_, new_n305_, keyIn_0_33, new_n321_, new_n332_ );
not g119 ( new_n334_, keyIn_0_33 );
nand g120 ( new_n335_, new_n305_, new_n321_, new_n332_ );
nand g121 ( new_n336_, new_n335_, new_n334_ );
not g122 ( new_n337_, keyIn_0_9 );
not g123 ( new_n338_, keyIn_0_1 );
nand g124 ( new_n339_, N1, N8, N17, N51 );
xnor g125 ( new_n340_, new_n339_, new_n338_ );
nand g126 ( new_n341_, new_n340_, new_n337_ );
xnor g127 ( new_n342_, new_n339_, keyIn_0_1 );
nand g128 ( new_n343_, new_n342_, keyIn_0_9 );
nand g129 ( new_n344_, new_n341_, new_n343_ );
not g130 ( new_n345_, keyIn_0_11 );
not g131 ( new_n346_, keyIn_0_3 );
nand g132 ( new_n347_, N42, N59, N75 );
xnor g133 ( new_n348_, new_n347_, new_n346_ );
nand g134 ( new_n349_, new_n348_, new_n345_ );
xnor g135 ( new_n350_, new_n347_, keyIn_0_3 );
nand g136 ( new_n351_, new_n350_, keyIn_0_11 );
nand g137 ( new_n352_, new_n349_, new_n351_ );
nand g138 ( new_n353_, new_n344_, keyIn_0_25, new_n352_ );
not g139 ( new_n354_, keyIn_0_25 );
nand g140 ( new_n355_, new_n344_, new_n352_ );
nand g141 ( new_n356_, new_n355_, new_n354_ );
nand g142 ( new_n357_, new_n356_, new_n353_ );
nand g143 ( new_n358_, new_n336_, new_n357_, new_n320_, new_n333_ );
nand g144 ( new_n359_, new_n336_, new_n357_, new_n333_ );
nand g145 ( new_n360_, new_n359_, keyIn_0_39 );
nand g146 ( new_n361_, new_n360_, new_n358_ );
nand g147 ( new_n362_, new_n361_, keyIn_0_62, N126 );
not g148 ( new_n363_, keyIn_0_62 );
nand g149 ( new_n364_, new_n361_, N126 );
nand g150 ( new_n365_, new_n364_, new_n363_ );
nand g151 ( new_n366_, new_n365_, new_n362_ );
nand g152 ( new_n367_, new_n366_, new_n319_, new_n295_, new_n317_ );
nand g153 ( new_n368_, new_n366_, new_n317_, new_n319_ );
nand g154 ( new_n369_, new_n368_, keyIn_0_70 );
nand g155 ( new_n370_, new_n369_, new_n367_ );
nand g156 ( new_n371_, N29, N75, N80 );
xor g157 ( new_n372_, new_n371_, keyIn_0_2 );
and g158 ( new_n373_, new_n305_, new_n372_ );
nand g159 ( new_n374_, new_n373_, N55 );
xnor g160 ( new_n375_, new_n374_, keyIn_0_32 );
xor g161 ( new_n376_, keyIn_0_4, N268 );
xnor g162 ( new_n377_, new_n376_, keyIn_0_16 );
nand g163 ( new_n378_, new_n375_, new_n377_ );
xnor g164 ( new_n379_, new_n378_, keyIn_0_48 );
nand g165 ( new_n380_, new_n370_, keyIn_0_78, new_n379_ );
not g166 ( new_n381_, keyIn_0_78 );
nand g167 ( new_n382_, new_n370_, new_n379_ );
nand g168 ( new_n383_, new_n382_, new_n381_ );
nand g169 ( new_n384_, new_n383_, keyIn_0_83, N201, new_n380_ );
not g170 ( new_n385_, keyIn_0_83 );
nand g171 ( new_n386_, new_n383_, N201, new_n380_ );
nand g172 ( new_n387_, new_n386_, new_n385_ );
not g173 ( new_n388_, N201 );
nand g174 ( new_n389_, new_n383_, new_n380_ );
nand g175 ( new_n390_, new_n389_, new_n388_ );
nand g176 ( new_n391_, new_n390_, keyIn_0_84 );
not g177 ( new_n392_, keyIn_0_84 );
nand g178 ( new_n393_, new_n389_, new_n392_, new_n388_ );
nand g179 ( new_n394_, new_n391_, new_n393_ );
nand g180 ( new_n395_, new_n394_, new_n384_, new_n387_ );
xor g181 ( new_n396_, new_n395_, keyIn_0_94 );
or g182 ( new_n397_, new_n396_, N261 );
nand g183 ( new_n398_, new_n396_, N261 );
nand g184 ( new_n399_, new_n397_, N219, new_n398_ );
nand g185 ( new_n400_, new_n396_, N228 );
nand g186 ( new_n401_, new_n387_, new_n384_ );
xnor g187 ( new_n402_, new_n401_, keyIn_0_93 );
nand g188 ( new_n403_, new_n402_, N237 );
nand g189 ( new_n404_, new_n383_, N246, new_n380_ );
nand g190 ( new_n405_, new_n240_, N42, N72 );
nand g191 ( new_n406_, new_n405_, keyIn_0_10 );
or g192 ( new_n407_, new_n405_, keyIn_0_10 );
and g193 ( new_n408_, new_n407_, N73, new_n406_ );
nand g194 ( new_n409_, new_n408_, N201 );
nand g195 ( new_n410_, N255, N267 );
nand g196 ( new_n411_, N121, N210 );
and g197 ( new_n412_, new_n404_, new_n409_, new_n410_, new_n411_ );
nand g198 ( new_n413_, new_n399_, new_n400_, new_n403_, new_n412_ );
xor g199 ( N850, new_n413_, keyIn_0_112 );
not g200 ( new_n415_, keyIn_0_103 );
not g201 ( new_n416_, keyIn_0_80 );
not g202 ( new_n417_, N189 );
nand g203 ( new_n418_, new_n316_, N146 );
or g204 ( new_n419_, new_n418_, keyIn_0_57 );
nand g205 ( new_n420_, new_n418_, keyIn_0_57 );
nand g206 ( new_n421_, new_n361_, N116 );
xnor g207 ( new_n422_, new_n421_, keyIn_0_58 );
nand g208 ( new_n423_, new_n422_, new_n419_, keyIn_0_68, new_n420_ );
not g209 ( new_n424_, keyIn_0_68 );
nand g210 ( new_n425_, new_n422_, new_n419_, new_n420_ );
nand g211 ( new_n426_, new_n425_, new_n424_ );
xor g212 ( new_n427_, new_n378_, keyIn_0_46 );
nand g213 ( new_n428_, new_n426_, keyIn_0_76, new_n423_, new_n427_ );
not g214 ( new_n429_, keyIn_0_76 );
nand g215 ( new_n430_, new_n426_, new_n423_, new_n427_ );
nand g216 ( new_n431_, new_n430_, new_n429_ );
nand g217 ( new_n432_, new_n431_, new_n428_ );
nand g218 ( new_n433_, new_n432_, new_n416_, new_n417_ );
nand g219 ( new_n434_, new_n432_, new_n417_ );
nand g220 ( new_n435_, new_n434_, keyIn_0_80 );
and g221 ( new_n436_, new_n435_, new_n433_ );
not g222 ( new_n437_, keyIn_0_59 );
nand g223 ( new_n438_, new_n316_, new_n437_, N149 );
nand g224 ( new_n439_, new_n316_, N149 );
nand g225 ( new_n440_, new_n439_, keyIn_0_59 );
nand g226 ( new_n441_, new_n440_, new_n438_ );
nand g227 ( new_n442_, new_n361_, N121 );
xnor g228 ( new_n443_, new_n442_, keyIn_0_60 );
nand g229 ( new_n444_, new_n441_, new_n443_, keyIn_0_69 );
not g230 ( new_n445_, keyIn_0_69 );
nand g231 ( new_n446_, new_n441_, new_n443_ );
nand g232 ( new_n447_, new_n446_, new_n445_ );
nand g233 ( new_n448_, new_n447_, new_n444_ );
xnor g234 ( new_n449_, new_n378_, keyIn_0_47 );
not g235 ( new_n450_, new_n449_ );
nand g236 ( new_n451_, new_n448_, keyIn_0_77, new_n450_ );
not g237 ( new_n452_, keyIn_0_77 );
nand g238 ( new_n453_, new_n448_, new_n450_ );
nand g239 ( new_n454_, new_n453_, new_n452_ );
nand g240 ( new_n455_, new_n454_, N195, new_n451_ );
xnor g241 ( new_n456_, new_n455_, keyIn_0_81 );
nand g242 ( new_n457_, new_n456_, keyIn_0_91 );
not g243 ( new_n458_, keyIn_0_91 );
nand g244 ( new_n459_, new_n455_, keyIn_0_81 );
or g245 ( new_n460_, new_n455_, keyIn_0_81 );
nand g246 ( new_n461_, new_n460_, new_n458_, new_n459_ );
nand g247 ( new_n462_, new_n457_, new_n436_, new_n461_ );
nand g248 ( new_n463_, new_n462_, keyIn_0_98 );
not g249 ( new_n464_, keyIn_0_98 );
nand g250 ( new_n465_, new_n457_, new_n464_, new_n436_, new_n461_ );
nand g251 ( new_n466_, new_n463_, new_n465_ );
not g252 ( new_n467_, N195 );
nand g253 ( new_n468_, new_n454_, new_n451_ );
nand g254 ( new_n469_, new_n468_, keyIn_0_82, new_n467_ );
not g255 ( new_n470_, keyIn_0_82 );
nand g256 ( new_n471_, new_n468_, new_n467_ );
nand g257 ( new_n472_, new_n471_, new_n470_ );
and g258 ( new_n473_, new_n472_, new_n469_ );
nand g259 ( new_n474_, new_n402_, new_n436_, new_n473_ );
nand g260 ( new_n475_, new_n474_, keyIn_0_99 );
nand g261 ( new_n476_, new_n472_, new_n433_, new_n435_, new_n469_ );
nand g262 ( new_n477_, new_n394_, N261 );
nor g263 ( new_n478_, new_n477_, new_n476_, keyIn_0_96 );
not g264 ( new_n479_, keyIn_0_96 );
nor g265 ( new_n480_, new_n477_, new_n476_ );
nor g266 ( new_n481_, new_n480_, new_n479_ );
nor g267 ( new_n482_, new_n481_, new_n478_ );
nor g268 ( new_n483_, new_n432_, new_n417_ );
xnor g269 ( new_n484_, new_n483_, keyIn_0_79 );
nor g270 ( new_n485_, new_n476_, keyIn_0_99 );
nand g271 ( new_n486_, new_n485_, new_n402_ );
nand g272 ( new_n487_, new_n486_, new_n484_ );
nor g273 ( new_n488_, new_n482_, new_n487_ );
nand g274 ( new_n489_, new_n488_, new_n415_, new_n466_, new_n475_ );
not g275 ( new_n490_, new_n478_ );
or g276 ( new_n491_, new_n477_, new_n476_ );
nand g277 ( new_n492_, new_n491_, keyIn_0_96 );
nand g278 ( new_n493_, new_n492_, new_n490_ );
and g279 ( new_n494_, new_n486_, new_n484_ );
nand g280 ( new_n495_, new_n493_, new_n494_, new_n466_, new_n475_ );
nand g281 ( new_n496_, new_n495_, keyIn_0_103 );
nand g282 ( new_n497_, new_n489_, new_n496_ );
not g283 ( new_n498_, keyIn_0_67 );
nand g284 ( new_n499_, new_n316_, N143 );
or g285 ( new_n500_, new_n499_, keyIn_0_55 );
nand g286 ( new_n501_, new_n361_, N111 );
xnor g287 ( new_n502_, new_n501_, keyIn_0_56 );
nand g288 ( new_n503_, new_n499_, keyIn_0_55 );
nand g289 ( new_n504_, new_n502_, new_n500_, new_n503_ );
or g290 ( new_n505_, new_n504_, new_n498_ );
nand g291 ( new_n506_, new_n504_, new_n498_ );
xnor g292 ( new_n507_, new_n378_, keyIn_0_45 );
nand g293 ( new_n508_, new_n505_, new_n506_, new_n507_ );
xor g294 ( new_n509_, new_n508_, keyIn_0_75 );
nand g295 ( new_n510_, new_n509_, N183 );
or g296 ( new_n511_, new_n509_, N183 );
nand g297 ( new_n512_, new_n511_, new_n510_ );
xnor g298 ( new_n513_, new_n512_, keyIn_0_89 );
not g299 ( new_n514_, new_n513_ );
and g300 ( new_n515_, new_n497_, new_n514_ );
or g301 ( new_n516_, new_n515_, keyIn_0_106 );
nand g302 ( new_n517_, new_n515_, keyIn_0_106 );
nand g303 ( new_n518_, new_n489_, new_n496_, new_n513_ );
nand g304 ( new_n519_, new_n516_, N219, new_n517_, new_n518_ );
nand g305 ( new_n520_, new_n514_, N228 );
nand g306 ( new_n521_, new_n509_, N183, N237 );
nand g307 ( new_n522_, new_n509_, N246 );
nand g308 ( new_n523_, new_n408_, N183 );
nand g309 ( new_n524_, N106, N210 );
and g310 ( new_n525_, new_n521_, new_n522_, new_n523_, new_n524_ );
nand g311 ( new_n526_, new_n519_, new_n520_, new_n525_ );
xor g312 ( N863, new_n526_, keyIn_0_121 );
nand g313 ( new_n528_, new_n457_, new_n461_ );
not g314 ( new_n529_, keyIn_0_95 );
not g315 ( new_n530_, new_n473_ );
nor g316 ( new_n531_, new_n530_, new_n477_ );
or g317 ( new_n532_, new_n531_, new_n529_ );
nand g318 ( new_n533_, new_n531_, new_n529_ );
not g319 ( new_n534_, new_n402_ );
nor g320 ( new_n535_, new_n534_, new_n530_ );
xor g321 ( new_n536_, new_n535_, keyIn_0_97 );
nand g322 ( new_n537_, new_n536_, new_n528_, new_n532_, new_n533_ );
xnor g323 ( new_n538_, new_n537_, keyIn_0_104 );
nand g324 ( new_n539_, new_n484_, new_n436_ );
xnor g325 ( new_n540_, new_n539_, keyIn_0_90 );
nand g326 ( new_n541_, new_n538_, new_n540_ );
or g327 ( new_n542_, new_n541_, keyIn_0_107 );
nand g328 ( new_n543_, new_n541_, keyIn_0_107 );
or g329 ( new_n544_, new_n538_, new_n540_ );
nand g330 ( new_n545_, new_n542_, N219, new_n543_, new_n544_ );
nand g331 ( new_n546_, new_n540_, N228 );
not g332 ( new_n547_, N237 );
or g333 ( new_n548_, new_n484_, new_n547_ );
nand g334 ( new_n549_, new_n431_, N246, new_n428_ );
nand g335 ( new_n550_, new_n408_, N189 );
nand g336 ( new_n551_, N255, N259 );
nand g337 ( new_n552_, N111, N210 );
and g338 ( new_n553_, new_n549_, new_n550_, new_n551_, new_n552_ );
nand g339 ( new_n554_, new_n545_, new_n546_, new_n548_, new_n553_ );
xnor g340 ( N864, new_n554_, keyIn_0_122 );
not g341 ( new_n556_, keyIn_0_108 );
nand g342 ( new_n557_, new_n534_, new_n477_ );
xnor g343 ( new_n558_, new_n557_, keyIn_0_105 );
nand g344 ( new_n559_, new_n473_, new_n456_ );
xnor g345 ( new_n560_, new_n559_, keyIn_0_92 );
or g346 ( new_n561_, new_n558_, new_n560_ );
or g347 ( new_n562_, new_n561_, new_n556_ );
nand g348 ( new_n563_, new_n561_, new_n556_ );
nand g349 ( new_n564_, new_n558_, new_n560_ );
nand g350 ( new_n565_, new_n562_, N219, new_n563_, new_n564_ );
not g351 ( new_n566_, N228 );
nor g352 ( new_n567_, new_n560_, new_n566_ );
nor g353 ( new_n568_, new_n528_, new_n547_ );
and g354 ( new_n569_, new_n454_, N246, new_n451_ );
nand g355 ( new_n570_, new_n408_, N195 );
nand g356 ( new_n571_, N116, N210 );
nand g357 ( new_n572_, N255, N260 );
nand g358 ( new_n573_, new_n570_, new_n571_, new_n572_ );
nor g359 ( new_n574_, new_n567_, new_n568_, new_n569_, new_n573_ );
nand g360 ( new_n575_, new_n565_, new_n574_ );
xnor g361 ( N865, new_n575_, keyIn_0_123 );
not g362 ( new_n577_, keyIn_0_115 );
not g363 ( new_n578_, keyIn_0_110 );
nand g364 ( new_n579_, new_n497_, keyIn_0_109, new_n511_ );
not g365 ( new_n580_, keyIn_0_109 );
nand g366 ( new_n581_, new_n497_, new_n511_ );
nand g367 ( new_n582_, new_n581_, new_n580_ );
nand g368 ( new_n583_, new_n582_, new_n579_ );
nand g369 ( new_n584_, new_n583_, new_n578_, new_n510_ );
nand g370 ( new_n585_, new_n583_, new_n510_ );
nand g371 ( new_n586_, new_n585_, keyIn_0_110 );
nand g372 ( new_n587_, new_n586_, new_n584_ );
not g373 ( new_n588_, N177 );
nand g374 ( new_n589_, new_n361_, N106 );
nand g375 ( new_n590_, N138, N152 );
nand g376 ( new_n591_, new_n589_, new_n590_ );
xnor g377 ( new_n592_, new_n591_, keyIn_0_66 );
nand g378 ( new_n593_, new_n373_, N17 );
xor g379 ( new_n594_, new_n593_, keyIn_0_31 );
nand g380 ( new_n595_, new_n594_, new_n376_ );
xnor g381 ( new_n596_, new_n595_, keyIn_0_43 );
nand g382 ( new_n597_, new_n305_, N55, new_n307_ );
xor g383 ( new_n598_, new_n597_, keyIn_0_30 );
nand g384 ( new_n599_, new_n598_, N153 );
nand g385 ( new_n600_, new_n596_, new_n599_ );
xor g386 ( new_n601_, new_n600_, keyIn_0_54 );
nand g387 ( new_n602_, new_n601_, new_n592_ );
xor g388 ( new_n603_, new_n602_, keyIn_0_74 );
not g389 ( new_n604_, new_n603_ );
nand g390 ( new_n605_, new_n604_, new_n588_ );
nand g391 ( new_n606_, new_n361_, N96 );
nand g392 ( new_n607_, N51, N138 );
nand g393 ( new_n608_, new_n606_, new_n607_ );
xor g394 ( new_n609_, new_n608_, keyIn_0_64 );
xor g395 ( new_n610_, new_n595_, keyIn_0_41 );
nand g396 ( new_n611_, new_n598_, N146 );
nand g397 ( new_n612_, new_n610_, new_n611_ );
xnor g398 ( new_n613_, new_n612_, keyIn_0_52 );
nand g399 ( new_n614_, new_n613_, new_n609_ );
xor g400 ( new_n615_, new_n614_, keyIn_0_72 );
or g401 ( new_n616_, new_n615_, N165 );
not g402 ( new_n617_, N171 );
nand g403 ( new_n618_, new_n361_, N101 );
nand g404 ( new_n619_, N17, N138 );
nand g405 ( new_n620_, new_n618_, new_n619_ );
xnor g406 ( new_n621_, new_n620_, keyIn_0_65 );
xnor g407 ( new_n622_, new_n595_, keyIn_0_42 );
nand g408 ( new_n623_, new_n598_, N149 );
nand g409 ( new_n624_, new_n622_, new_n623_ );
xor g410 ( new_n625_, new_n624_, keyIn_0_53 );
nand g411 ( new_n626_, new_n625_, new_n621_ );
or g412 ( new_n627_, new_n626_, keyIn_0_73 );
nand g413 ( new_n628_, new_n626_, keyIn_0_73 );
nand g414 ( new_n629_, new_n627_, new_n628_ );
nand g415 ( new_n630_, new_n629_, new_n617_ );
and g416 ( new_n631_, new_n616_, new_n630_ );
nand g417 ( new_n632_, new_n587_, new_n605_, new_n631_ );
xnor g418 ( new_n633_, new_n632_, new_n577_ );
nor g419 ( new_n634_, new_n604_, new_n588_ );
nand g420 ( new_n635_, new_n631_, new_n634_ );
xnor g421 ( new_n636_, new_n635_, keyIn_0_102 );
nor g422 ( new_n637_, new_n629_, new_n617_ );
nand g423 ( new_n638_, new_n616_, new_n637_ );
or g424 ( new_n639_, new_n638_, keyIn_0_101 );
nand g425 ( new_n640_, new_n638_, keyIn_0_101 );
nand g426 ( new_n641_, new_n615_, N165 );
and g427 ( new_n642_, new_n636_, new_n639_, new_n640_, new_n641_ );
nand g428 ( new_n643_, new_n633_, keyIn_0_116, new_n642_ );
not g429 ( new_n644_, keyIn_0_116 );
nand g430 ( new_n645_, new_n633_, new_n642_ );
nand g431 ( new_n646_, new_n645_, new_n644_ );
nand g432 ( new_n647_, new_n646_, new_n643_ );
nand g433 ( new_n648_, new_n361_, N91 );
nand g434 ( new_n649_, N8, N138 );
nand g435 ( new_n650_, new_n648_, new_n649_ );
xor g436 ( new_n651_, new_n650_, keyIn_0_63 );
xor g437 ( new_n652_, new_n595_, keyIn_0_40 );
nand g438 ( new_n653_, new_n598_, N143 );
nand g439 ( new_n654_, new_n652_, new_n653_ );
xnor g440 ( new_n655_, new_n654_, keyIn_0_51 );
nand g441 ( new_n656_, new_n655_, new_n651_ );
xnor g442 ( new_n657_, new_n656_, keyIn_0_71 );
nor g443 ( new_n658_, new_n657_, N159 );
not g444 ( new_n659_, new_n658_ );
nand g445 ( new_n660_, new_n647_, new_n659_ );
nand g446 ( new_n661_, new_n657_, N159 );
nand g447 ( N866, new_n660_, new_n661_ );
not g448 ( new_n663_, new_n634_ );
nand g449 ( new_n664_, new_n663_, new_n605_ );
xnor g450 ( new_n665_, new_n664_, keyIn_0_88 );
nand g451 ( new_n666_, new_n587_, new_n665_ );
or g452 ( new_n667_, new_n666_, keyIn_0_111 );
nand g453 ( new_n668_, new_n666_, keyIn_0_111 );
or g454 ( new_n669_, new_n587_, new_n665_ );
nand g455 ( new_n670_, new_n667_, N219, new_n668_, new_n669_ );
nand g456 ( new_n671_, new_n665_, N228 );
nand g457 ( new_n672_, new_n634_, N237 );
nand g458 ( new_n673_, new_n603_, N246 );
nand g459 ( new_n674_, new_n408_, N177 );
nand g460 ( new_n675_, N101, N210 );
and g461 ( new_n676_, new_n672_, new_n673_, new_n674_, new_n675_ );
nand g462 ( new_n677_, new_n670_, new_n671_, new_n676_ );
xor g463 ( N874, new_n677_, keyIn_0_124 );
not g464 ( new_n679_, keyIn_0_125 );
nand g465 ( new_n680_, new_n659_, new_n661_ );
xnor g466 ( new_n681_, new_n680_, keyIn_0_85 );
nand g467 ( new_n682_, new_n646_, new_n643_, new_n681_ );
not g468 ( new_n683_, new_n681_ );
nand g469 ( new_n684_, new_n647_, new_n683_ );
nand g470 ( new_n685_, new_n684_, N219, new_n682_ );
nor g471 ( new_n686_, new_n681_, new_n566_ );
nor g472 ( new_n687_, new_n661_, new_n547_ );
nand g473 ( new_n688_, new_n657_, N246 );
nand g474 ( new_n689_, new_n408_, N159 );
not g475 ( new_n690_, N210 );
or g476 ( new_n691_, new_n377_, new_n690_ );
nand g477 ( new_n692_, new_n688_, new_n689_, new_n691_ );
nor g478 ( new_n693_, new_n686_, new_n687_, new_n692_ );
nand g479 ( new_n694_, new_n685_, new_n679_, new_n693_ );
nand g480 ( new_n695_, new_n685_, new_n693_ );
nand g481 ( new_n696_, new_n695_, keyIn_0_125 );
nand g482 ( N878, new_n696_, new_n694_ );
not g483 ( new_n698_, keyIn_0_126 );
not g484 ( new_n699_, keyIn_0_117 );
nand g485 ( new_n700_, new_n587_, keyIn_0_114, new_n605_, new_n630_ );
not g486 ( new_n701_, keyIn_0_114 );
nand g487 ( new_n702_, new_n587_, new_n605_, new_n630_ );
nand g488 ( new_n703_, new_n702_, new_n701_ );
nand g489 ( new_n704_, new_n634_, new_n630_ );
and g490 ( new_n705_, new_n704_, keyIn_0_100 );
nor g491 ( new_n706_, new_n704_, keyIn_0_100 );
nor g492 ( new_n707_, new_n705_, new_n706_, new_n637_ );
nand g493 ( new_n708_, new_n703_, new_n699_, new_n700_, new_n707_ );
nand g494 ( new_n709_, new_n703_, new_n700_, new_n707_ );
nand g495 ( new_n710_, new_n709_, keyIn_0_117 );
nand g496 ( new_n711_, new_n710_, new_n708_ );
nand g497 ( new_n712_, new_n616_, new_n641_ );
xor g498 ( new_n713_, new_n712_, keyIn_0_86 );
nand g499 ( new_n714_, new_n711_, keyIn_0_119, new_n713_ );
not g500 ( new_n715_, keyIn_0_119 );
nand g501 ( new_n716_, new_n711_, new_n713_ );
nand g502 ( new_n717_, new_n716_, new_n715_ );
or g503 ( new_n718_, new_n711_, new_n713_ );
nand g504 ( new_n719_, new_n717_, new_n718_, N219, new_n714_ );
and g505 ( new_n720_, new_n713_, N228 );
nor g506 ( new_n721_, new_n641_, new_n547_ );
nand g507 ( new_n722_, new_n615_, N246 );
nand g508 ( new_n723_, new_n408_, N165 );
nand g509 ( new_n724_, N91, N210 );
nand g510 ( new_n725_, new_n722_, new_n723_, new_n724_ );
nor g511 ( new_n726_, new_n720_, new_n721_, new_n725_ );
nand g512 ( new_n727_, new_n719_, new_n726_ );
nand g513 ( new_n728_, new_n727_, new_n698_ );
nand g514 ( new_n729_, new_n719_, keyIn_0_126, new_n726_ );
nand g515 ( N879, new_n728_, new_n729_ );
not g516 ( new_n731_, keyIn_0_127 );
not g517 ( new_n732_, keyIn_0_120 );
not g518 ( new_n733_, keyIn_0_118 );
not g519 ( new_n734_, keyIn_0_113 );
nand g520 ( new_n735_, new_n587_, new_n734_, new_n605_ );
nand g521 ( new_n736_, new_n587_, new_n605_ );
nand g522 ( new_n737_, new_n736_, keyIn_0_113 );
nand g523 ( new_n738_, new_n737_, new_n735_ );
nand g524 ( new_n739_, new_n738_, new_n733_, new_n663_ );
nand g525 ( new_n740_, new_n738_, new_n663_ );
nand g526 ( new_n741_, new_n740_, keyIn_0_118 );
nand g527 ( new_n742_, new_n741_, new_n739_ );
not g528 ( new_n743_, new_n637_ );
nand g529 ( new_n744_, new_n743_, new_n630_ );
xor g530 ( new_n745_, new_n744_, keyIn_0_87 );
nand g531 ( new_n746_, new_n742_, new_n732_, new_n745_ );
nand g532 ( new_n747_, new_n742_, new_n745_ );
nand g533 ( new_n748_, new_n747_, keyIn_0_120 );
not g534 ( new_n749_, new_n745_ );
nand g535 ( new_n750_, new_n741_, new_n739_, new_n749_ );
and g536 ( new_n751_, new_n750_, N219 );
nand g537 ( new_n752_, new_n748_, new_n751_, new_n746_ );
nor g538 ( new_n753_, new_n749_, new_n566_ );
nor g539 ( new_n754_, new_n743_, new_n547_ );
nand g540 ( new_n755_, new_n627_, N246, new_n628_ );
nand g541 ( new_n756_, new_n408_, N171 );
nand g542 ( new_n757_, N96, N210 );
nand g543 ( new_n758_, new_n755_, new_n756_, new_n757_ );
nor g544 ( new_n759_, new_n753_, new_n754_, new_n758_ );
nand g545 ( new_n760_, new_n752_, new_n759_ );
nand g546 ( new_n761_, new_n760_, new_n731_ );
nand g547 ( new_n762_, new_n752_, keyIn_0_127, new_n759_ );
nand g548 ( N880, new_n761_, new_n762_ );
endmodule