module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g33533, g34435, g34788, g34839, g36, g44, g53,
         g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
         g6751, g6753, g84, g90, g91, g92, g99, test_so10, test_so26,
         test_so35, test_so39, test_so42, test_so44, test_so46, test_so80,
         test_so86, test_so92, test_so100, g34783, n2730, n4896, n4895, n4837,
         n4921, n4920, n5045, g559, n4959, g33046, g5057, n5615, g34441, g2771,
         n5544, g33982, g1882, g34007, g2299, g24276, g4040, n5530, g30381,
         g2547, n5782, g30405, g3243, g25604, g452, g30416, g3542, g30466,
         g5232, g25736, g5813, g34617, g33974, g1744, g30505, g5909, g33554,
         g1802, n5536, g30432, g3554, g33064, g6219, n5385, g34881, g807,
         n5479, g6031, g24216, g847, n5709, g24232, n9367, DFF_24_n1, g34733,
         g4172, n5493, g34882, g4372, g33026, g3512, g31867, n5471, g25668,
         g3490, n5454, g24344, n5432, g4235, g33966, g1600, g33550, g1714,
         n5460, g30393, g3155, n5366, g29248, g2236, g4571, g4555, g24274,
         g3698, g33973, g1736, g30360, g1968, n5664, g34460, g30494, g5607,
         g30384, g2657, n5316, g24340, n5439, g29223, g490, n5708, g26881,
         g311, n5317, g34252, g772, n5334, g30489, g5587, g29301, g6177, n5874,
         g6377, g33022, g3167, n5652, g30496, g5615, g33043, g4567, g29263,
         g30533, g6287, g24256, n5302, g34015, g2563, g34031, g4776, n5707,
         g34452, g4593, n5303, g34646, g6199, n5644, g34001, g2295, g25633,
         g1384, g24259, g1339, g33049, g5180, n5384, g34609, g2844, g31869,
         g1024, g30490, g30427, g3598, g21894, g4264, g33965, g767, n5333,
         g34645, g5853, n5499, g33571, g2089, g34267, g4933, g26971, g4521,
         n5752, g34644, g5507, n5643, g30534, g6291, g33535, g294, n5680,
         g30498, g25728, g25743, g25684, g3813, g25613, g562, g34438, g608,
         n5475, g24244, g1205, n5547, g30439, g3909, g30541, g6259, g30519,
         g5905, g25621, g921, g34807, g2955, g25599, g203, g24235, g34036,
         g4878, n5283, g30476, g5204, g30429, g3606, g32997, g1926, n5510,
         g33063, g6215, n5651, g30424, g3586, g32977, g291, n5679, g34026,
         g4674, n5440, g30420, g3570, g33560, g29226, g676, n5751, g25619,
         g843, g34455, g4332, n5540, g30457, g4153, g33625, g6336, g34790,
         g622, n5672, g30414, g3506, n5576, g26966, g4558, g25656, g3111,
         g30390, g25688, g34727, g939, n5415, g278, n5627, g26963, g4492,
         g34034, g4864, n5318, g33541, g1036, g28093, g24236, g1178, g30404,
         g3239, g28051, g718, g29303, g6195, g26917, g1135, n5328, g33624,
         g6395, n5396, g24337, g34911, g554, g33963, g496, g34627, g3853,
         n5641, g29282, g5134, n5807, g25676, g33013, g2485, n5509, g32981,
         g925, n5725, g34976, n9357, DFF_150_n1, g30483, g5555, g32994, g1798,
         n5833, g28070, g34806, g2941, g30453, g3905, g33539, g763, n5332,
         g30526, g6255, g4375, g34035, g4871, n5443, g34636, g4722, n5345,
         g32978, g590, n5472, g30348, g1632, n5836, g24336, n5438, g3100,
         g24250, g29236, g1437, g29298, g6154, n5747, g1579, g30499, g5567,
         g33976, g1752, g32996, g1917, g30335, g744, n5470, g34637, g4737,
         n5867, g25694, DFF_178_n1, g30528, g6267, g24251, g1442, g30521,
         g26960, g4477, n5849, g24239, g34259, g4643, n5382, g30474, g5264,
         n5703, g33016, g2610, g34643, g5160, n5498, g30510, g5933, g29239,
         g1454, g26897, g753, g34729, g1296, g34625, g3151, n5495, g24353,
         g6727, n5531, g33029, g3530, n5569, g33615, g4104, g24253, g1532,
         g24281, g33997, n9352, g34971, n9351, DFF_206_n1, g34263, g4754,
         n5877, g24237, g1189, n5642, g33584, g2287, n5353, g24280, g4273,
         n5764, g26920, g1389, g33548, g29296, g5835, n5663, g30338, g1171,
         n5363, g21895, g4269, n5763, g33588, g2399, n5762, g34041, g4983,
         n5367, g30495, g5611, g29279, g4572, g25655, g3143, n5882, g34795,
         g2898, g24269, g3343, g30403, g3235, g33042, g30419, g3566, g34023,
         n9348, DFF_228_n1, g28090, g4961, n5770, g34642, g4927, n5879, g30370,
         g2259, n5419, g34448, g2819, n5609, g26946, g5802, g34610, g2852,
         g24209, g417, n5358, g28047, g681, g24206, g437, g26891, g30504,
         g5901, g34798, g2886, g25669, g3494, n5889, g30480, g5511, n5575,
         g33027, g3518, n5645, g33972, g1604, g25697, g5092, g28099, g4831,
         g26947, g4382, n5714, g24350, g6386, g24210, g479, g30455, g3965,
         g28084, g33993, g2008, g736, g30444, g3933, g33537, g222, g25650,
         g3050, n5998, g25625, g1052, g30366, g2122, n5784, g33593, g2465,
         n5523, g30502, g5889, g33036, g4495, g25595, g34462, g33024, g3179,
         n5390, g33552, g1728, n5352, g34014, g2433, g29273, g3835, n5662,
         g25748, g6187, n5453, g34638, g4917, n5408, g30341, g1070, g26899,
         g822, n5422, g30336, g914, n5560, g5339, g26940, g4164, g25622,
         g34447, g2807, n5379, g33613, g4054, n5395, g25749, g6191, n5888,
         g25704, g5077, n5455, g33053, g5523, n5647, g3680, g30555, g6637,
         g25601, g174, n5402, g33971, g1682, g26892, g355, g1087, g26915,
         g1105, n5478, g33008, g30538, g6307, g3802, g25750, g6159, g30369,
         g2255, n5414, g34446, g2815, n5404, g29230, g911, n5559, g43, g33975,
         g1748, g30497, g5551, g30418, g3558, g25721, g5499, n5885, g34622,
         g30438, g3901, g34266, g4888, n5863, g30540, g6251, g32986, g1373,
         g25648, g33960, g157, n5678, g34442, g2783, n5403, g4281, g30421,
         g3574, g33573, g2112, g34730, g1283, n5635, g24205, g10122_Tj, g4297,
         n5698, g32979, g758, n5331, g4639, n5727, g25763, g6537, n5884,
         g30481, g5543, g30517, g5961, g30539, g6243, g34880, n9340, g24242,
         n5654, g30436, g29265, g3476, n5786, g32990, g1664, g24245, g1246,
         n5756, g30553, g6629, g26907, g246, n6008, g24278, g4049, g26955,
         g24282, g2932, g4575, g31894, g4098, n5350, g33037, g4498, g26894,
         g528, n5327, g34977, n5477, g25654, g3139, n5447, g33962, g34451,
         g4584, n5539, g34250, g142, n5724, g29295, g5831, g26905, g239,
         g25629, g1216, n5442, g34792, g2848, g25703, g5022, g32983, g1030,
         g30402, g3231, g25757, g1430, n9336, g33999, g2241, g24262, g1564,
         g25729, g6148, g30558, g6649, g34781, g110, g26901, g225, n5597,
         g26961, g33039, g4504, g33059, g5873, n5388, g31899, g5037, n5611,
         g33007, g2319, n5375, g25720, g5495, n5446, g21891, g30462, g5208,
         g30487, g5579, g33058, g5869, n5649, g24261, g1589, n5755, g25730,
         g5752, n5996, g30531, g6279, g30506, g34804, g2975, n5750, g25747,
         g6167, n5430, n5701, g33601, g2599, n5524, g26922, g1448, n5343,
         g29250, g2370, g30459, g5164, n5570, g1333, n5616, g33534, g153,
         n5677, g30543, g6549, n5571, g29275, g4087, n5480, g34030, g34980,
         g2984, n5842, g30451, g3961, g25627, g962, n5630, g34657, g101,
         g30552, g6625, g34979, n9332, DFF_420_n1, g30337, g1018, g24254,
         g24277, g4045, g29237, g1467, g30378, g2461, n5840, g33019, n5300,
         g33623, g5990, g29235, g1256, n5558, g31902, g5029, n5601, g29306,
         g6519, n5806, g25689, g4169, n5729, g33978, g1816, g26970, g4369,
         g4578, g34253, g4459, n5765, g29272, g3831, n5872, g33595, g2514,
         g33610, g3288, n5400, g33589, g34605, g2145, n5307, g30350, g1700,
         n5417, g25611, g513, n5548, g2841, n5963, g33619, g5297, n5588,
         g34022, g2763, g34033, g4793, n5368, g34726, g952, g31870, g1263,
         n5674, g33985, g1950, g29283, g5138, n5871, g34003, g2307, g25677,
         g34463, g4664, g33006, g2223, g29292, g5808, n5749, g30557, g6645,
         g33989, g2016, g33033, g3873, n5387, n5699, g34005, g2315, g26932,
         g2811, g30516, g5957, g33575, g2047, g33032, g30486, g5575, g34974,
         n9327, DFF_477_n1, g25678, g3752, n5994, g30440, g3917, g1585, n5757,
         g26949, g4388, g30530, g6275, g30542, g6311, g25624, g1041, g30383,
         g33597, g2537, g34598, g26957, g4430, g26967, n9325, g28102, g4826,
         g30524, g6239, g26903, g232, g30475, g5268, g34647, g6545, n5497,
         g30377, n9324, g33553, g1772, n5504, g31903, g5052, n5607, g25715,
         g33984, g1890, g33602, g2629, n5521, g28045, g572, n5337, g34603,
         g2130, n5487, g33035, g4108, n5715, g4308, g24208, g475, g990, n5622,
         g31, n5469, g34970, n9322, DFF_514_n1, g33614, g3990, n5594, g33060,
         g30362, g1992, g33023, g3171, n5603, g26898, g812, n5733, g25618,
         g832, g30518, g5897, g4570, n5702, g26959, g4455, g34801, g2902,
         g26884, g333, g25600, g168, n5606, g26933, g28066, g3684, g33612,
         g3639, n5591, g24268, g3338, n5527, g25716, g5406, n5992, g26906,
         g269, g24203, g401, g24346, g6040, g24207, g441, g25701, n5690,
         g29269, g3808, n5745, g9, n5468, g34255, g30450, g3957, g30456, g4093,
         n5340, g32991, g1760, n5602, g24348, n5437, g34249, g160, n5843,
         g30371, g2279, n5778, g29268, g3498, g29224, g586, n5336, g33017,
         g2619, n5508, g30339, g1183, n5599, g33967, g1608, g33559, g1779,
         g29255, g2652, g30368, g2193, n5839, g30375, g2393, n5421, g28052,
         g661, g28089, g4950, n5772, g33055, g5535, n5566, g30392, g2834,
         g30343, g1361, g30523, g6235, g24233, g1146, n5851, g33018, g32976,
         g150, n5676, g30349, g1696, n5628, g33067, g6555, g26900, g33034,
         g3881, n5564, g30551, g6621, g25667, g3470, n5424, g30452, g3897,
         g34719, g518, g538, g33607, g2606, g26923, g1472, n5290, g24211,
         g33050, g5188, n5567, g24341, g5689, n5529, g24201, g405, g30463,
         g5216, g6494, g34464, g4669, g996, g24335, g4531, g34611, g2860,
         g34262, g4743, g30546, g6593, g25591, g4411, g30347, g1413, g30556,
         g6641, g6, g33562, g1936, n5534, g55, g25610, g504, n5519, g33015,
         g2587, n5372, g31896, g4480, g34004, n9314, g30428, g30485, g5571,
         g30422, g3578, g25714, g29294, g5827, n5809, g30423, g3582, g30529,
         g6271, g34028, g4688, n5656, g33587, g2380, g30460, g5196, g30401,
         g3227, g33990, n9312, g29309, g6541, g30411, g3203, g33546, g1668,
         n5598, g28085, g4760, n5775, g26904, g262, g33556, g1840, n5451,
         g25722, g5467, g25605, g460, g33062, g6209, g26893, n5704, g28050,
         g655, g34626, g33583, g2204, n5620, g30472, g5256, g34454, g4608,
         n5274, g34850, g794, n5291, g4423, g24272, g3689, n5532, g5685,
         g24214, g703, n5821, g26909, g862, n5682, g30406, g3247, g33569,
         g2040, n5505, DFF_672_n1, g34628, g4146, n5981, g34458, g4633, n5844,
         g24240, n5304, g34634, g4732, n5296, g25700, n5689, g29293, g5817,
         g33009, g2351, n5511, g33603, g2648, g24355, g6736, g34268, g4944,
         n5875, g25691, g4072, g26890, g29264, g3466, g28072, g4116, g31900,
         g5041, n5605, g26956, g4434, g29271, g3827, n5808, g29304, g6500,
         n5748, g29261, g3133, n5661, g28063, g3333, g979, n5320, g34027,
         g4681, g33961, g298, n5675, g33604, g32995, g1894, n5374, g34624,
         g2988, g30415, g3538, g33536, g301, g26888, n9306, DFF_709_n1, g28055,
         g827, n5728, g24238, g33600, g2555, n5351, g28105, g5011, g34721,
         g199, g29307, g6523, n5870, g30345, g34453, g4601, n5365, g32980,
         g854, g29238, g1484, n5865, g34639, g4922, n5346, g25695, g5080,
         n5893, g33057, g5863, g26969, g4581, n5670, g29253, g2518, g34021,
         g2567, g26895, g568, n5335, g30413, g3263, g30549, g6613, g24347,
         g25758, g6444, n5990, g34808, g2965, g30501, g5857, n5573, g33969,
         n9303, g34440, g890, n5305, g30433, g3562, g21900, g26921, g1404,
         g29270, g3817, n9302, n6010, g33038, g4501, g31865, g26926, g2724,
         n5301, g28083, g4704, n5771, g34797, g22, g2878, g30478, g5220,
         g34724, g617, n5339, g24212, g26883, g316, g32985, g1277, g25761,
         g6513, n5426, g26886, g336, n5824, g34796, g2882, g32982, g33561,
         g1906, n5503, g26880, g305, n5282, g34975, g8, g26931, g2799, g34641,
         g4912, n5297, g34629, g4157, n5983, g33598, g2541, n5461, g33576,
         g2153, n5356, g34720, g550, g26902, g255, g29244, g30468, g5240,
         g26924, g1478, n5289, g33031, g3863, g29245, g1959, g29266, g3480,
         n5868, g30559, g6653, g34794, g2864, g28087, g4894, n5774, g30435,
         g3857, n5572, g25609, g28057, g1002, g34439, g776, n5330, g28, n5324,
         g1236, g34260, g4646, n5712, g33012, g2476, g32989, g1657, n5525,
         g34006, g2375, g63, g358, g26910, g896, n5431, g28043, g33021, g3161,
         g29251, g2384, n5700, g34456, g4616, n5608, g26968, g4561, g33991,
         g2024, g3451, g26930, g2795, g34599, g613, n5474, g28082, g4527,
         g33557, g1844, g30511, g5937, g33045, g30379, g2523, n5281, g24267,
         n5436, g34020, g2643, g24249, g1489, n5850, g25592, g30382, n9295,
         g29285, g5156, n5526, n9294, DFF_829_n1, g25662, g21896, g33563,
         g1955, g33622, g33582, g2273, n5458, g28086, g4771, n5769, g25744,
         g6098, n5988, g29262, g3147, g24270, g3347, g33581, g2269, g191,
         g24266, g2712, g34849, g626, n5288, g33618, g2729, g5357, n5393,
         g34038, g34032, g4709, n5518, g34803, g2927, g34459, g4340, n5653,
         g30509, g5929, g34640, g4907, n5295, g28069, g4035, g21899, g2946,
         g31868, g918, n5673, g26938, g4082, g25756, g30363, g30334, g577,
         n5294, g33970, g1620, g30391, g2831, g25615, g667, g33540, g930,
         n5731, g30445, g3937, g25617, g817, n5822, g24247, g1249, g24215,
         g837, n5562, g33964, g599, n5550, g25719, g5475, n5425, g29228,
         g30514, g5949, g33627, g6682, n5590, g24231, g904, g34615, g2873,
         n5488, g30356, g1854, n5785, g25696, g5084, n5681, g30493, g5603,
         n5726, g33594, g2495, n5522, g34009, g2437, g30365, g2102, n5666,
         g33004, g2208, g34018, g25685, g4064, n5416, g34040, g4899, n5517,
         g25639, g2719, n5465, g34029, g4785, n5361, g30488, g5583, g34600,
         g781, n5551, g29300, g6173, n5810, g34802, g2917, g25614, g686,
         g28058, g1252, n5554, g29225, g671, g33580, g30532, g6283, g33054,
         g5527, n5389, g26962, g4489, g33564, g1974, n5450, g32984, g1270,
         n5716, g34039, g4966, n5706, g33065, g6227, n5568, g30443, g3929,
         g29291, g5503, g24279, g30508, g5925, g29232, g1124, g34269, g4955,
         n5614, g30464, g5224, g33988, g2012, g30522, g6203, n5574, g25708,
         g5120, g30374, g2389, n5631, g26953, g4438, g34008, g2429, g34444,
         g2787, n5610, g34731, g33606, g2675, n5457, g24334, n5541, g34265,
         g4836, n5713, g30340, g1199, g24257, n5401, g30482, g5547, g34604,
         g2138, n5275, g33591, g2338, g30525, g6247, g26929, g2791, g30448,
         g34602, g1291, n2549, g30513, g5945, g30469, g5244, g33608, g2759,
         g33626, g6741, n5398, g34725, g785, n5293, g30342, g1259, n5553,
         g29267, g3484, n5668, g25593, g209, n5595, g30548, g6609, g33052,
         g5517, g34012, g2449, g34017, n9281, g24263, g2715, n5299, g26912,
         g936, n5557, g30364, g2098, n5280, g34254, g4462, n5671, g34251, g604,
         n5473, g30560, g6589, g33983, n9280, g24204, g429, g33980, g1870,
         g34631, g29243, g1825, g25623, g1008, n5321, g26950, g4392, n5710,
         g30431, g3546, g30467, g5236, g30353, g1768, n5834, g34467, g4854,
         g30442, g3925, g29305, g6509, g25616, g732, n5732, g29252, g2504,
         g4519, g4520, g33003, g2185, n5376, g34613, g37, g4031, g33570, g2070,
         n5535, g34734, g4176, n5494, g24275, n5435, g4405, g872, g29302,
         g6181, n5667, g24349, g34264, g4765, n5613, g30484, g5563, g25634,
         g1395, g33567, g1913, g33585, g2331, n5513, g30527, g6263, g34978,
         n9276, DFF_1012_n1, g30447, g3945, g347, n5860, g34256, g4473, g25630,
         g1266, g29290, g5489, n5660, g29227, g31872, g2748, n5516, g29287,
         g5471, g31897, g4540, g6723, g30562, g6605, g34011, n9274, g33996,
         g2173, g21898, g33014, g2491, g34465, g4849, g33995, g2169, g30372,
         n9273, g30545, g30389, g33590, g2407, n5459, g34616, g2868, g26927,
         g2767, g32992, g1783, n5596, g25631, g1312, n5466, g30477, g5212,
         g34632, g4245, n5640, g28046, g645, g4291, g26896, g25602, g26916,
         g1129, n5329, g33578, g2227, n5538, g33579, g2246, g30354, g1830,
         n5413, g30425, g3590, g24200, g392, g33544, g1592, n5362, g25764,
         g6505, g24246, g1221, g30507, g5921, g26889, g30333, g218, g32998,
         g1932, g32987, g1624, n5370, g25702, g5062, g29286, g5462, n5744,
         g34606, g2689, n5347, g33070, g6573, n5563, g29240, g1677, g32999,
         g2028, n5371, g33605, g2671, g24255, g26945, g33558, g1848, n5464,
         g25699, n5669, g29289, g5485, n5869, g30388, g2741, n5349, g29254,
         g2638, g28074, g4122, g34450, g4322, n5506, g30512, g5941, g33572,
         g2108, n5452, g25, g33551, g33538, g595, n5476, g33005, g2217, n5512,
         g24248, n9267, DFF_1092_n1, g33002, g2066, n5832, g24234, g1152,
         n5618, g30471, g5252, g34000, g2165, g34016, g2571, g33048, g5176,
         n5650, g25628, g26934, g2827, g34468, g4859, g24202, g424, g33542,
         g1274, n5730, n9265, g34445, g2803, n5545, g33555, g1821, g34013,
         g2509, g28091, g5073, g26919, n5556, g30554, g6633, g29281, g5124,
         g30537, g6303, g28092, g5069, g34732, g2994, n5634, g28049, g650,
         g33545, g1636, n5549, g30441, g3921, g29247, g24354, g6732, g25636,
         g1306, n5796, g26914, g1061, g25670, g3462, g33998, g2181, g25626,
         g956, n5341, g33977, g1756, g29297, g5849, g28071, g4112, g30387,
         n9262, g33577, g2197, n5514, g33592, g26913, g1046, g28044, g482,
         n5820, g26948, g4401, g30344, g1514, n5364, g26885, g329, n5766,
         g33069, g6565, n5386, g34621, g2950, g28059, g1345, g25762, g6533,
         n5445, g34633, g4727, n5312, g24352, g26925, g1536, g30446, g3941,
         g25597, g370, g24342, g5694, g30357, g1858, n5892, g26908, g446,
         g30399, g3219, g29242, g1811, g30547, g6601, g34010, g2441, g33986,
         g1874, g34257, g30544, g6581, g30561, g6597, g5008, n5637, g30430,
         g3610, g34799, g2890, g33565, g1978, g33968, g1612, g34843, g112,
         g34793, g2856, g33566, g1982, n5462, g30465, g28073, g4119, g24351,
         g6390, g30346, g1542, g21893, g4258, g4818, n5636, g31904, g5033,
         g34635, g4717, n5344, g25637, g1554, n5768, g29274, g3849, g30396,
         g3199, g25735, g34037, g4975, n5360, g34791, g790, n5292, g30520,
         g5913, g30358, g1902, n5837, g29299, g6163, g25690, g4125, g28096,
         g4821, g28088, g4939, n5776, g24241, n5392, g30397, g3207, g4483,
         g30409, g29284, g5142, n5658, g30470, g5248, g30367, g2126, g24273,
         g3694, g29288, g5481, n5805, g30359, g1964, n5315, g25698, g5097,
         n5753, g30398, g3215, n9255, g26952, g4427, g26928, g2779, n5694,
         g26954, DFF_1225_n1, g30351, g1720, n5780, g31871, g1367, g5112, g19,
         g26939, g4145, g33994, g2161, g25596, g376, n5633, g33586, g2361,
         n5537, g21901, g31866, g582, n5552, g33000, g2051, g26918, g1193,
         g30373, g2327, n5841, g28056, g907, n5555, g34601, g947, n5286,
         g30355, g1834, n5665, g30426, g3594, g34805, g2999, g34002, g2303,
         g28053, g29229, g723, n5826, g33620, g5703, n5397, g34722, g546,
         n5492, g33599, g2472, n5619, g30515, g5953, g25649, g33979, g1740,
         g30417, g3550, g25683, g3845, n5886, g33574, g2116, n5463, g30410,
         g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777, g33596,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g4417,
         g33068, g6561, n5646, g29233, g1141, n5691, g24258, n5655, g30376,
         g33549, g1710, g29308, g6527, n5659, g30408, g3255, g29241, g1691,
         g34620, g2936, g33621, g5644, g25707, g5152, n5883, g24339, g5352,
         g34443, g2775, n5378, g34619, g2922, g29234, g30503, g5893, g30550,
         g6617, g33001, g2060, n5507, g33040, g4512, g30492, g5599, g25664,
         g3401, n5986, g26944, g4366, g34614, n5342, g29260, g3129, n5861,
         g33047, g5170, g24298, g25733, g5821, n5429, g30536, g6299, g29246,
         g2079, g34261, g4698, n5862, g33611, g3703, n5399, g25638, g1559,
         n5441, g34728, n9247, g29222, g411, n5629, g25742, g30449, g3953,
         g34608, g2704, n5377, g24345, g6035, n5528, n9245, g25635, g1300,
         n5483, g25686, g4057, n5711, g30461, g5200, g34466, g4843, g31901,
         g5046, n5578, g29249, g2250, g26882, n5456, g33041, g33011, g2453,
         n5373, g25734, g5841, n5449, n5705, g34618, g2912, g33010, g2357,
         g31864, g164, n5561, g34630, g4253, n5484, g31898, g5016, n5369,
         g25653, g3119, n5423, g25632, g1351, n5322, g32988, g33616, g29280,
         g5115, n5743, g33609, g3352, n5604, g30563, g6657, g33044, g4552,
         g30437, g3893, g30412, g3211, g30491, g5595, g30434, g3614, g34612,
         g29259, g3125, n5781, g25681, g3821, n5428, g25687, g4141, n5612,
         g33617, g30479, g5272, g29256, g2735, n5600, g28054, g728, g30535,
         g6295, g30385, g2661, n5418, g30361, g1988, n5783, g25705, g24260,
         g1548, n5546, g29257, g3106, n5742, g34461, g4659, g34258, g4358,
         n5348, g32993, g1792, n5359, g33992, g2084, g30394, g3187, g34449,
         g4311, n5323, g34019, g2583, g18597, n9240, DFF_1381_n1, g29231,
         g1094, g25682, g21897, g4284, g30395, g3191, g21892, g4239, g4180,
         n5380, g28048, g691, n5520, g34723, g534, n5490, g25598, g385, n5632,
         g33987, g2004, g30380, g2527, n5420, g5456, g26965, n6007, g25706,
         g30458, g4507, n5846, g24338, g5348, g30400, g3223, g34623, g2970,
         g24343, g5698, g30473, g5260, g24252, g1521, g33028, g3522, n5383,
         g29258, g3115, g30407, g3251, g26958, g34457, g33568, g1996, n5355,
         g25663, g26964, g4515, g34735, g4300, n5639, g30352, n9236, g33543,
         g1379, g24271, n5433, g33981, g1878, g30500, g5619, g34649, g71,
         g29277, g25612, n5287, g28060, n2505, n2499, n2461, n2396, n2668,
         n3141, n3122, g72, n5960, n4689, n5961, n4708, n3593, n3589, n3595,
         n3574, n3570, n3576, n3517, n3513, n3519, n3628, n3624, n3630, n3555,
         n3551, n3557, n3646, n3642, n3648, n3536, n3532, n3538, n3611, n3607,
         n3613, n3006, n3765, n3505, n3525, n3635, n4888, n3550, n2595, n2527,
         n3524, n3005, n3623, n3549, n3003, n3007, n3569, n3606, n3588, n3165,
         n3799, n3033, n3622, n3587, n3586, n3605, n3604, n3568, n3567, n3548,
         n3512, n3511, n3531, n3530, n3641, n3640, n3131, n3111, n4537, n4201,
         n3745, n3684, n3274, n2982, n2706, n2649, n2556, n2509, n2487, n2427,
         n2423, n2421, n4172, n4173, n4190, n4191, n4388, n4210, n3951, n3774,
         n3842, n3808, n3908, n3984, n3875, n4015, n3914, n3780, n3957, n3848,
         n3990, n3814, n3881, n4022, n4027, n3785, n3962, n3853, n3886, n3819,
         n3995, n3919, n3682, n3272, n2980, n2704, n2647, n2554, n2507, n2485,
         n2425, n2419, n2405, n2760, n2552, n4946, n4198, n2404, n3653, n4962,
         n4948, n2726, n2727, n3195, n2774, n3116, n4945, n4525, n4518, n3281,
         n3277, n3276, n2989, n2991, n2710, n2707, n3174, n3362, n3676, n2644,
         n3146, n3115, n3833, n3023, n3933, n3729, n2601, n3664, n3662, n3673,
         n3671, n2607, n3506, n2790, n4490, n4178, n4514, n4196, n3736, n3741,
         n2598, n4814, n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145,
         n3164, n2422, n4037, n4034, n4039, n3972, n3969, n3929, n3926, n3863,
         n3860, n4003, n4002, n4032, n4035, n3797, n3792, n3790, n3795, n3891,
         n3893, n3827, n3826, n3896, n4007, n3931, n3793, n3924, n3831, n3829,
         n3927, n3974, n3898, n3970, n4000, n3865, n3861, n3824, n3894, n3967,
         n3858, n4005, n3395, n4956, n5026, n3941, n3733, n4798, n4805, n4175,
         n4193, n3738, n4721, n4523, n4524, n4526, n2573, n2577, n2563, n2567,
         n4938, n4913, n4714, n4516, n4517, n5111, n4819, n3730, n3121, n3180,
         n4305, n4283, n2608, n4447, n4448, n4402, n4403, n4425, n4436, n4437,
         n4391, n4392, n4379, n4380, n4414, n4415, n4458, n4459, n5016, n5014,
         n3064, n3065, n4535, n5112, n3675, counter_31, counter_30, counter_29,
         counter_28, counter_27, counter_26, counter_25, counter_24,
         counter_23, counter_22, counter_21, counter_20, counter_19,
         counter_18, counter_17, counter_16, counter_15, counter_14,
         counter_13, counter_12, counter_11, counter_10, counter_9, counter_8,
         counter_7, counter_6, counter_5, counter_4, counter_3, counter_2,
         counter_1, counter_0, carry_31, carry_30, carry_29, carry_28,
         carry_27, carry_26, carry_25, carry_24, carry_23, carry_22, carry_21,
         carry_20, carry_19, carry_18, carry_17, carry_16, carry_15, carry_14,
         carry_13, carry_12, carry_11, carry_10, carry_9, carry_8, carry_7,
         carry_6, carry_5, carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16,
         N17, N18, N19, N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87,
         n73, n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74,
         n58, n59, n60, n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68,
         n69, n70, n71, n72, n5, n42, n44, n46, n51, n53, n55, n56, n99, n100,
         n101, n112, n113, n114, g33959, n192, n198, n199, n205, n207, n209,
         n214, n279, n335, n411, n422, n424, n429, n431, n433, n438, n468,
         n494, n495, n496, n503, n526, n527, n528, n530, n542, n543, n631,
         n686, n700, n712, n714, n716, n720, n744, n745, n746, n750, n751,
         n752, n807, n811, n826, n828, n830, n835, n853, n935, n936, n937,
         n939, g25259, n1009, n1010, n1011, n1073, n1074, n1075, n1135, n1136,
         n1137, g25167, n1161, n1220, n1242, n1249, n1376, n1401, n1403, n1405,
         n1409, n1411, n1415, n1526, n1680, n1721, n1782, n8045, n8048, n8051,
         n8052, n8054, n8055, n8070, n8071, n8072, n8073, n8074, n8079, n8080,
         n8083, n8084, n8086, n8087, n8088, n8090, n8091, n8095, n8096, n8097,
         n8099, n8100, n8102, n8103, n8104, n8105, n8106, n8111, n8117, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8137, n8138, n8139, n8140,
         n8142, n8144, n8148, n8150, n8151, n8152, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8177, n8179, n8180, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8192, n8193,
         n8194, n8196, n8197, n8198, n8201, n8202, n8204, n8205, n8207, n8208,
         n8209, n8212, n8213, n8215, n8216, n8218, n8220, n8221, n8223, n8225,
         n8227, n8229, n8230, n8231, n8232, n8266, n8268, n8270, n8272, n8274,
         n8276, n8278, n8279, n8281, n8283, n8285, n8287, n8288, n8290, n8292,
         n8294, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8312, n8313, n8318, n8321,
         n8324, n8327, n8330, n8333, n8336, n8339, n8351, n8365, n8366, n8367,
         n8368, n8370, n8371, n8372, n8373, n8375, n8377, n8380, n8382, n8384,
         n8385, n8386, n8387, n8389, n8390, n8391, n8392, n8394, n8395, n8396,
         n8397, n8399, n8401, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8448, n8449, n8450, n8451, n8452, n8455, n8458, n8459,
         n8460, n8461, n8462, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8475, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8498, n8499, n8501, n8502, n8504, n8505, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8532, n8533, n8536, n8537, n8538, n8539, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8554, n8555,
         n8556, n8557, n8560, n8561, n8562, n8566, n8567, n8568, n8569, n8570,
         g32975, n8572, n8573, n8574, n8575, n8576, n8577, g31860, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9241,
         n9242, n9243, n9244, n9246, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9256, n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9266,
         n9268, n9269, n9270, n9271, n9272, n9275, n9277, n9278, n9279, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9296, n9297, n9298, n9299, n9300, n9301, n9304, n9305, n9307,
         n9308, n9309, n9310, n9311, n9313, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9323, n9326, n9328, n9329, n9330, n9331, n9333, n9334,
         n9335, n9337, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9349, n9350, n9353, n9354, n9355, n9356, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, U5116_n1, U5126_n1, U5127_n1, U5128_n1, U5129_n1,
         U5353_n1, U5355_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1,
         U5966_n1, U5967_n1, U5968_n1, U6100_n1, U6211_n1, U6212_n1, U6213_n1,
         U6214_n1, U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6279_n1, U6280_n1,
         U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1,
         U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6338_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6417_n1,
         U6446_n1, U6465_n1, U6497_n1, U6523_n1, U6542_n1, U6552_n1, U6553_n1,
         U6554_n1, U6555_n1, U6556_n1, U6559_n1, U6560_n1, U6561_n1, U6570_n1,
         U6911_n1, U6912_n1, U6917_n1, U6926_n1, U6927_n1, U6929_n1, U6931_n1,
         U6932_n1, U6933_n1, U6934_n1, U6935_n1, U6936_n1, U6937_n1, U6938_n1,
         U6939_n1, U6940_n1, U6941_n1, U6944_n1, U6950_n1, U6954_n1, U6955_n1,
         U6956_n1, U6957_n1, U7174_n1, U7248_n1, U7249_n1, U7402_n1, U7405_n1,
         U7413_n1, U7416_n1, U7427_n1, U7438_n1, U7449_n1, U7455_n1, U7464_n1,
         U7467_n1, U7482_n1, U7492_n1, U7513_n1, U7516_n1, U7549_n1, U7561_n1,
         U7574_n1, U7577_n1, U7585_n1, U7595_n1, U7614_n1, U7621_n1, U7629_n1,
         U7636_n1, U7639_n1, U7649_n1, U7652_n1, U7668_n1, U7673_n1, U7690_n1,
         U7707_n1, U7712_n1, U7792_n1, U7794_n1, U7895_n1, U7897_n1, U7977_n1,
         U8034_n1, U8036_n1, U8050_n1, U8055_n1, U8060_n1, U8070_n1, U8074_n1,
         U8088_n1, U8112_n1, U8113_n1, U8147_n1, U8165_n1, U8185_n1, U8192_n1,
         U8210_n1, U8223_n1, U8224_n1, U8281_n1, U8307_n1, U8974_n1, U8975_n1,
         U9065_n1, U9070_n1, U9075_n1, U9076_n1, U9080_n1, U9084_n1, U9085_n1,
         U9086_n1, U9090_n1, U9098_n1, U9099_n1, U9101_n1, U9107_n1, U9111_n1,
         U9116_n1, U9120_n1, U9124_n1, U9128_n1, U9132_n1, U9136_n1, U9315_n1,
         U9453_n1, U9825_n1, U9886_n1, U9927_n1, U9953_n1, U9957_n1, U9958_n1,
         U9968_n1, U9972_n1, U9992_n1, U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g27831 = g33533;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g31862 = g25259;
  assign g31863 = g25167;
  assign g26801 = g32975;
  assign g25114 = g31860;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n8641), .CLK(n9056), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n8651), .CLK(n9066), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n8696), .CLK(n9111), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n8711), .CLK(n9126), .Q(
        g2299) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n8743), .CLK(n9158), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n8674), .CLK(n9089), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n8730), .CLK(n9145), .Q(g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n8695), .CLK(n9110), .Q(
        g3243) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n8653), .CLK(n9068), .Q(
        g452), .QN(n8313) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n8720), .CLK(n9135), .Q(
        g3542), .QN(n8207) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n8655), .CLK(n9070), .Q(
        g5232) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n8727), .CLK(n9142), .Q(
        g5813), .QN(n8139) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n8681), .CLK(n9096), .Q(
        test_so1), .QN(n8616) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n8650), .CLK(n9065), 
        .Q(g1744) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n8729), .CLK(n9144), .Q(
        g5909), .QN(n8324) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n8666), .CLK(n9081), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n8730), .CLK(n9145), .Q(
        g3554), .QN(n8397) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n8731), .CLK(n9146), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n8676), .CLK(n9091), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n8676), .CLK(n9091), .Q(
        g6031), .QN(n8406) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n8707), .CLK(n9122), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n8695), .CLK(n9110), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n8685), .CLK(n9100), .Q(
        g4172), .QN(n5493) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n8686), .CLK(n9101), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n8686), .CLK(n9101), .Q(
        g3512), .QN(n8490) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n8675), .CLK(n9090), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n8716), .CLK(n9131), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n8688), .CLK(n9103), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n8738), .CLK(n9153), .Q(
        g4235), .QN(n8232) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n8703), .CLK(n9118), .Q(
        g1600) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n8647), .CLK(n9062), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n8728), .CLK(n9143), .Q(
        g14451) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n8728), .CLK(n9143), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n8670), .CLK(n9085), .Q(
        g2236) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n8708), .CLK(n9123), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n8733), .CLK(n9148), .Q(
        g3698), .QN(n8301) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n8650), .CLK(n9065), .Q(
        g1736) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n8694), .CLK(n9109), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n8705), .CLK(n9120), .Q(
        test_so3), .QN(n8605) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n8645), .CLK(n9060), 
        .Q(g5607) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n8646), .CLK(n9061), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n8667), .CLK(n9082), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n8715), .CLK(n9130), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n8715), .CLK(n9130), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n8676), .CLK(n9091), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n8645), .CLK(n9060), .Q(
        g5587) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n8679), .CLK(n9094), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n8718), .CLK(n9133), .Q(
        g6377), .QN(n8426) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n8728), .CLK(n9143), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n8733), .CLK(n9148), .Q(
        g5615) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n8743), .CLK(n9158), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n8677), .CLK(n9092), .Q(
        test_so4), .QN(n8611) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n8683), .CLK(n9098), 
        .Q(g6287) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n8724), .CLK(n9139), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n8649), .CLK(n9064), .Q(
        g2563) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n8730), .CLK(n9145), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n8707), .CLK(n9122), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n8707), .CLK(n9122), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n8711), .CLK(n9126), .Q(
        g2295) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n8647), .CLK(n9062), .Q(
        g1384), .QN(n8055) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n8726), .CLK(n9141), .Q(
        g1339) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n8726), .CLK(n9141), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n8702), .CLK(n9117), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n8656), .CLK(n9071), .Q(
        g1024), .QN(n8157) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n8645), .CLK(n9060), .Q(
        test_so5) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n8677), .CLK(n9092), 
        .Q(g3598), .QN(n8205) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n8700), .CLK(n9115), .Q(
        g4264) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n8675), .CLK(n9090), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n8676), .CLK(n9091), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n8740), .CLK(n9155), .Q(
        g13865) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n8698), .CLK(n9113), .Q(
        g2089) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n8702), .CLK(n9117), .Q(
        g4933) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n8686), .CLK(n9101), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n8686), .CLK(n9101), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n8728), .CLK(n9143), .Q(
        g16656), .QN(n8396) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n8684), .CLK(n9099), .Q(
        g6291) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n8663), .CLK(n9078), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n8747), .CLK(n9162), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n8727), .CLK(n9142), 
        .Q(g9617) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n8660), .CLK(n9075), .Q(
        g9741), .QN(n8084) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n8660), .CLK(n9075), .Q(
        g3813), .QN(n8125) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n8660), .CLK(n9075), .Q(
        g562) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n8661), .CLK(n9076), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n8735), .CLK(n9150), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n8652), .CLK(n9067), .Q(
        g3909), .QN(n8330) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n8683), .CLK(n9098), .Q(
        g6259), .QN(n8427) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n8667), .CLK(n9082), .Q(
        g5905) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n8668), .CLK(n9083), .Q(
        g921), .QN(n8505) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n8641), .CLK(n9056), .Q(
        g2955) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n8713), .CLK(n9128), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n8713), .CLK(n9128), .Q(
        test_so7), .QN(n8588) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n8719), .CLK(n9134), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n8720), .CLK(n9135), .Q(
        g5204) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n8721), .CLK(n9136), .Q(
        g17604), .QN(n8382) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n8722), .CLK(n9137), .Q(
        g3606), .QN(n8395) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n8694), .CLK(n9109), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n8698), .CLK(n9113), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n8730), .CLK(n9145), .Q(
        g3586) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n8663), .CLK(n9078), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n8730), .CLK(n9145), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n8730), .CLK(n9145), .Q(
        g3570) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n8730), .CLK(n9145), .Q(
        g9048), .QN(n8045) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n8730), .CLK(n9145), .Q(
        g17607), .QN(n8270) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n8736), .CLK(n9151), .Q(
        test_so8), .QN(n8586) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n8651), .CLK(n9066), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n8723), .CLK(n9138), .Q(
        g843), .QN(n8148) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n8707), .CLK(n9122), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n8685), .CLK(n9100), .Q(
        g4153), .QN(n8542) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n8685), .CLK(n9100), .Q(
        g17711), .QN(n8287) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n8678), .CLK(n9093), .Q(
        g6336) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n8661), .CLK(n9076), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n8716), .CLK(n9131), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n8716), .CLK(n9131), .Q(
        g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n8716), .CLK(n9131), .Q(
        g17685), .QN(n8401) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n8728), .CLK(n9143), .Q(
        g3111), .QN(n8122) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n8665), .CLK(n9080), .Q(
        g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n8665), .CLK(n9080), .Q(
        test_so9) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n8663), .CLK(n9078), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(n335), .SI(g939), .SE(n8663), .CLK(n9078), .Q(g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n8717), .CLK(n9132), .Q(
        g4492) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n8717), .CLK(n9132), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n8656), .CLK(n9071), .Q(
        g1036), .QN(n8515) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n8710), .CLK(n9125), .Q(
        g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n8710), .CLK(n9125), .Q(
        g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n8741), .CLK(n9156), .Q(
        g3239) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n8741), .CLK(n9156), .Q(
        g718), .QN(n8552) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n8741), .CLK(n9156), .Q(
        g6195) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n8647), .CLK(n9062), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n8739), .CLK(n9154), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n8663), .CLK(n9078), .Q(
        test_so10), .QN(n8613) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n8745), .CLK(n9160), 
        .Q(g554), .QN(n8144) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n8669), .CLK(n9084), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n8669), .CLK(n9084), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n8670), .CLK(n9085), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n8670), .CLK(n9085), .Q(
        g17404), .QN(n8160) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n8744), .CLK(n9159), .Q(
        g8344) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n8745), .CLK(n9160), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n8662), .CLK(n9077), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n8642), .CLK(n9057), .Q(
        n9357), .QN(DFF_150_n1) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n8642), .CLK(n9057), .Q(
        g5555), .QN(n8413) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n8709), .CLK(n9124), .Q(
        g14096) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n8678), .CLK(n9093), .Q(
        g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n8690), .CLK(n9105), .Q(
        test_so11), .QN(n8598) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n8652), .CLK(n9067), 
        .Q(g2941), .QN(n8460) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n8652), .CLK(n9067), .Q(
        g3905), .QN(n8387) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n8675), .CLK(n9090), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n8683), .CLK(n9098), .Q(
        g6255), .QN(n8339) );
  SDFFX1 DFF_159_Q_reg ( .D(n1526), .SI(g6255), .SE(n8659), .CLK(n9074), .Q(
        g4375), .QN(n8560) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n8717), .CLK(n9132), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n8717), .CLK(n9132), .Q(
        g4722), .QN(n5345) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n8661), .CLK(n9076), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n8737), .CLK(n9152), .Q(
        g13099) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n8677), .CLK(n9092), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n8675), .CLK(n9090), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n8650), .CLK(n9065), .Q(
        g3100), .QN(n8522) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n8737), .CLK(n9152), .Q(
        test_so12), .QN(n8632) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n8704), .CLK(n9119), 
        .Q(g1437) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n8679), .CLK(n9094), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n8726), .CLK(n9141), .Q(
        g1579) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n8733), .CLK(n9148), .Q(
        g5567), .QN(n8411) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n8651), .CLK(n9066), .Q(
        g1752) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n8740), .CLK(n9155), .Q(
        g1917), .QN(n8480) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n8675), .CLK(n9090), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n8717), .CLK(n9132), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n8717), .CLK(n9132), .Q(
        g8132), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n8692), .CLK(n9107), .Q(
        g6267) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n8706), .CLK(n9121), .Q(
        g16659), .QN(n8274) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n8706), .CLK(n9121), .Q(
        g1442), .QN(n8440) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n8706), .CLK(n9121), .Q(
        test_so13), .QN(n8626) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n8700), .CLK(n9115), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n8705), .CLK(n9120), .Q(
        g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n8705), .CLK(n9120), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n8655), .CLK(n9070), .Q(
        g5264), .QN(n8371) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n8678), .CLK(n9093), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n8715), .CLK(n9130), .Q(
        g2610), .QN(n8482) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n8715), .CLK(n9130), .Q(
        g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n8737), .CLK(n9152), .Q(
        g5933) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n8648), .CLK(n9063), .Q(
        g1454) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n8681), .CLK(n9096), .Q(
        g753), .QN(n8551) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n8681), .CLK(n9096), .Q(
        g1296) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n8681), .CLK(n9096), .Q(
        g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(n424), .SI(g3151), .SE(n8681), .CLK(n9096), .Q(
        test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n8690), .CLK(n9105), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n8716), .CLK(n9131), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(n8684), .CLK(n9099), .Q(
        g4104), .QN(n8312) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n8700), .CLK(n9115), .Q(
        g1532), .QN(n8307) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n8700), .CLK(n9115), .Q(
        g9251) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n8670), .CLK(n9085), .Q(
        n9352) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n8654), .CLK(n9069), .Q(
        n9351), .QN(DFF_206_n1) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n8654), .CLK(n9069), .Q(
        g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n8710), .CLK(n9125), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n8710), .CLK(n9125), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n8711), .CLK(n9126), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n8648), .CLK(n9063), .Q(
        g1389) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n8703), .CLK(n9118), .Q(
        test_so15), .QN(n8621) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n8667), .CLK(n9082), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n8693), .CLK(n9108), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n8700), .CLK(n9115), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n8744), .CLK(n9159), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n8682), .CLK(n9097), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n8728), .CLK(n9143), .Q(
        g5611) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n8728), .CLK(n9143), .Q(
        g16627), .QN(n8278) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n8644), .CLK(n9059), .Q(
        g4572), .QN(n8120) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n8746), .CLK(n9161), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n8656), .CLK(n9071), .Q(
        g2898) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n8703), .CLK(n9118), .Q(
        g3343), .QN(n8297) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n8703), .CLK(n9118), .Q(
        g3235) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n8743), .CLK(n9158), .Q(
        test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n8716), .CLK(n9131), 
        .Q(g3566) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n8672), .CLK(n9087), .Q(
        n9348), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n8672), .CLK(n9087), .Q(
        g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n8740), .CLK(n9155), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n8670), .CLK(n9085), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n8665), .CLK(n9080), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n8659), .CLK(n9074), .Q(
        g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n8659), .CLK(n9074), .Q(
        g5802), .QN(n8523) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n8702), .CLK(n9117), .Q(
        g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n8723), .CLK(n9138), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n8653), .CLK(n9068), .Q(
        g681), .QN(n8158) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n8657), .CLK(n9072), .Q(
        g437), .QN(n8164) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n8735), .CLK(n9150), .Q(
        test_so17), .QN(n8609) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n8667), .CLK(n9082), 
        .Q(g5901), .QN(n8409) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n8656), .CLK(n9071), .Q(
        g2886), .QN(n8462) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n8645), .CLK(n9060), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n8645), .CLK(n9060), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n8716), .CLK(n9131), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n8716), .CLK(n9131), .Q(
        g1604) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n8641), .CLK(n9056), .Q(
        g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n8706), .CLK(n9121), .Q(
        g4831) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n8706), .CLK(n9121), .Q(
        g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n8678), .CLK(n9093), .Q(
        g6386), .QN(n8299) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n8736), .CLK(n9151), .Q(
        g479), .QN(n8151) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n8648), .CLK(n9063), .Q(
        g3965), .QN(n8218) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n8668), .CLK(n9083), .Q(
        test_so18), .QN(n8635) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n8698), .CLK(n9113), 
        .Q(g2008) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n8710), .CLK(n9125), .Q(
        g736), .QN(n8514) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n8744), .CLK(n9159), .Q(
        g3933) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n8658), .CLK(n9073), .Q(
        g222), .QN(n8470) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n8650), .CLK(n9065), .Q(
        g3050), .QN(n5998) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n8695), .CLK(n9110), .Q(
        g1052), .QN(n8502) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n8695), .CLK(n9110), .Q(
        g17580), .QN(n8272) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n8643), .CLK(n9058), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n8713), .CLK(n9128), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n8713), .CLK(n9128), .Q(
        g5889) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n8713), .CLK(n9128), .Q(
        g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n8713), .CLK(n9128), .Q(
        g8719) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n8731), .CLK(n9146), .Q(
        test_so19), .QN(n8628) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n8694), .CLK(n9109), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n8666), .CLK(n9081), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n8688), .CLK(n9103), .Q(
        g2433) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n8643), .CLK(n9058), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n8731), .CLK(n9146), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n8731), .CLK(n9146), .Q(
        g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n8693), .CLK(n9108), .Q(
        g1070) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n8738), .CLK(n9153), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n8738), .CLK(n9153), .Q(
        g17715), .QN(n8375) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n8662), .CLK(n9077), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n8663), .CLK(n9078), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n8745), .CLK(n9160), .Q(
        g4164), .QN(n8450) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n8657), .CLK(n9072), .Q(
        test_so20), .QN(n8612) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n8664), .CLK(n9079), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n8743), .CLK(n9158), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n8679), .CLK(n9094), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n8679), .CLK(n9094), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n8679), .CLK(n9094), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n8739), .CLK(n9154), .Q(
        g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n8672), .CLK(n9087), .Q(
        g6637) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n8723), .CLK(n9138), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n8647), .CLK(n9062), .Q(
        g1682), .QN(n8135) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n8735), .CLK(n9150), .Q(
        g355), .QN(n8439) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n8735), .CLK(n9150), .Q(
        g1087), .QN(n8446) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n8695), .CLK(n9110), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n8727), .CLK(n9142), .Q(
        test_so21), .QN(n8591) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n8684), .CLK(n9099), 
        .Q(g6307) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n8744), .CLK(n9159), .Q(
        g3802), .QN(n8524) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n8744), .CLK(n9159), .Q(
        g6159), .QN(n8137) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n8670), .CLK(n9085), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n8665), .CLK(n9080), .Q(
        g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n8662), .CLK(n9077), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n8567), .SI(g911), .SE(n8679), .CLK(n9094), .Q(g43), .QN(n8499) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n8706), .CLK(n9121), .Q(
        g16775), .QN(n8288) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n8651), .CLK(n9066), .Q(
        g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n8645), .CLK(n9060), .Q(
        g5551) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n8735), .CLK(n9150), .Q(
        g3558), .QN(n8336) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n8742), .CLK(n9157), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n8745), .CLK(n9160), .Q(
        test_so22) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n8652), .CLK(n9067), 
        .Q(g3901) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n8683), .CLK(n9098), .Q(
        g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n8683), .CLK(n9098), .Q(
        g6251) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n8683), .CLK(n9098), .Q(
        g17649), .QN(n8279) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n8650), .CLK(n9065), .Q(
        g1373), .QN(n8172) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n8650), .CLK(n9065), .Q(
        g8215) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n8658), .CLK(n9073), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n8694), .CLK(n9109), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n8682), .CLK(n9097), .Q(
        g4281), .QN(n8473) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n8731), .CLK(n9146), .Q(
        g3574) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n8745), .CLK(n9160), .Q(
        g2112) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n8654), .CLK(n9069), .Q(
        g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n8657), .CLK(n9072), .Q(
        test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n8722), .CLK(n9137), .Q(g4297), .QN(n8087) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n8722), .CLK(n9137), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n8724), .CLK(n9139), .Q(
        g13272), .QN(n8521) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n8675), .CLK(n9090), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(n411), .SI(g758), .SE(n8705), .CLK(n9120), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n8746), .CLK(n9161), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n8645), .CLK(n9060), .Q(
        g5543) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n8724), .CLK(n9139), .Q(
        g8475), .QN(n8520) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n8729), .CLK(n9144), .Q(
        g5961) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n8692), .CLK(n9107), .Q(
        g6243) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n8662), .CLK(n9077), .Q(
        n9340), .QN(n15227) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n8662), .CLK(n9077), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n8744), .CLK(n9159), .Q(
        test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n8677), .CLK(n9092), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n8677), .CLK(n9092), .Q(
        g1664) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n8677), .CLK(n9092), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n8671), .CLK(n9086), .Q(
        g6629) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n8680), .CLK(n9095), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n8743), .CLK(n9158), .Q(
        g4049), .QN(n8305) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n8701), .CLK(n9116), .Q(
        g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n8701), .CLK(n9116), .Q(
        g2932), .QN(n8537) );
  SDFFX1 DFF_350_Q_reg ( .D(n1680), .SI(g2932), .SE(n8684), .CLK(n9099), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n8684), .CLK(n9099), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n8713), .CLK(n9128), .Q(
        g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n8723), .CLK(n9138), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n8641), .CLK(n9056), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n8669), .CLK(n9084), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n8669), .CLK(n9084), .Q(
        g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n8707), .CLK(n9122), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n8663), .CLK(n9078), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n8663), .CLK(n9078), .Q(
        g17639), .QN(n8370) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n8667), .CLK(n9082), .Q(
        g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n8689), .CLK(n9104), .Q(
        g239), .QN(n8309) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n8689), .CLK(n9104), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n8642), .CLK(n9057), .Q(
        g2848), .QN(n8544) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n8724), .CLK(n9139), .Q(
        g5022), .QN(n8496) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n8724), .CLK(n9139), .Q(
        g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n8656), .CLK(n9071), .Q(
        g1030), .QN(n8174) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n8728), .CLK(n9143), .Q(
        test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n8732), .CLK(n9147), 
        .Q(g3231) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n8734), .CLK(n9149), .Q(
        g9817), .QN(n8088) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n8734), .CLK(n9149), .Q(
        g1430), .QN(n8444) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n8741), .CLK(n9156), .Q(
        n9336), .QN(n15225) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n8697), .CLK(n9112), .Q(
        g2241), .QN(n8134) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n8734), .CLK(n9149), .Q(
        g1564), .QN(n8443) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n8660), .CLK(n9075), .Q(
        g9680), .QN(n8095) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n8660), .CLK(n9075), 
        .Q(g6148), .QN(n8529) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n8672), .CLK(n9087), .Q(
        g6649), .QN(n8390) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n8664), .CLK(n9079), .Q(
        g110) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n8709), .CLK(n9124), .Q(
        g14147) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n8709), .CLK(n9124), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n8709), .CLK(n9124), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n8713), .CLK(n9128), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n8727), .CLK(n9142), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n8727), .CLK(n9142), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n8727), .CLK(n9142), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n8742), .CLK(n9157), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n8655), .CLK(n9070), .Q(
        g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n8655), .CLK(n9070), .Q(
        g5208) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n8725), .CLK(n9140), .Q(
        g5579) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n8725), .CLK(n9140), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n8726), .CLK(n9141), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n8660), .CLK(n9075), .Q(
        g5752), .QN(n5996) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n8691), .CLK(n9106), .Q(
        g6279) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n8737), .CLK(n9152), .Q(
        test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n8646), .CLK(n9061), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n8679), .CLK(n9094), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n8706), .CLK(n9121), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n8687), .CLK(n9102), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n8648), .CLK(n9063), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n8709), .CLK(n9124), .Q(
        g14125) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n8701), .CLK(n9116), .Q(
        g2370) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n8701), .CLK(n9116), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n8724), .CLK(n9139), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n8658), .CLK(n9073), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n8715), .CLK(n9130), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n8715), .CLK(n9130), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n8729), .CLK(n9144), .Q(
        test_so29), .QN(n8595) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n8681), .CLK(n9096), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n8648), .CLK(n9063), .Q(
        g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n8710), .CLK(n9125), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n8654), .CLK(n9069), .Q(
        g101) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n8655), .CLK(n9070), .Q(
        g8918), .QN(n15231) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n8733), .CLK(n9148), .Q(
        g6625) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n8656), .CLK(n9071), .Q(
        n9332), .QN(DFF_420_n1) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n8656), .CLK(n9071), .Q(
        g1018), .QN(n8173) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n8670), .CLK(n9085), .Q(
        g17320), .QN(n8161) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n8743), .CLK(n9158), .Q(
        g4045), .QN(n8306) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n8743), .CLK(n9158), .Q(
        g1467) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n8673), .CLK(n9088), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n8710), .CLK(n9125), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n8739), .CLK(n9154), 
        .Q(g5990) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n8654), .CLK(n9069), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n8680), .CLK(n9095), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n8690), .CLK(n9105), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n8690), .CLK(n9105), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n8666), .CLK(n9081), .Q(
        g1816), .QN(n8070) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n8742), .CLK(n9157), .Q(
        g4369), .QN(n8310) );
  SDFFX1 DFF_439_Q_reg ( .D(n468), .SI(g4369), .SE(n8742), .CLK(n9157), .Q(
        g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n8742), .CLK(n9157), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n8643), .CLK(n9058), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n8688), .CLK(n9103), .Q(
        g2514), .QN(n8103) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n8702), .CLK(n9117), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n8744), .CLK(n9159), .Q(
        test_so31) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n8660), .CLK(n9075), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n8647), .CLK(n9062), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n8715), .CLK(n9130), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n8665), .CLK(n9080), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n8664), .CLK(n9079), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n8712), .CLK(n9127), .Q(
        g2763), .QN(n8052) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n8729), .CLK(n9144), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n8729), .CLK(n9144), .Q(
        g952) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n8654), .CLK(n9069), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n8696), .CLK(n9111), .Q(
        g1950), .QN(n8133) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n8664), .CLK(n9079), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n8664), .CLK(n9079), .Q(
        g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n8679), .CLK(n9094), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n8644), .CLK(n9059), 
        .Q(g8398), .QN(n8091) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n8644), .CLK(n9059), .Q(
        g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n8712), .CLK(n9127), .Q(
        g2223) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n8667), .CLK(n9082), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n8671), .CLK(n9086), .Q(
        g6645) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n8699), .CLK(n9114), .Q(
        g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n8699), .CLK(n9114), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n8732), .CLK(n9147), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n8738), .CLK(n9153), .Q(
        g2315) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n8664), .CLK(n9079), .Q(
        g2811) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n8729), .CLK(n9144), .Q(
        g5957) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n8693), .CLK(n9108), .Q(
        g2047) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n8704), .CLK(n9119), .Q(
        test_so33), .QN(n8594) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n8678), .CLK(n9093), 
        .Q(g17760), .QN(n8294) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n8645), .CLK(n9060), .Q(
        g5575) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n8643), .CLK(n9058), .Q(
        n9327), .QN(DFF_477_n1) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n8644), .CLK(n9059), .Q(
        g3752), .QN(n5994) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n8744), .CLK(n9159), .Q(
        g3917) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n8649), .CLK(n9064), 
        .Q(g8783), .QN(n15233) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n8649), .CLK(n9064), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n8724), .CLK(n9139), .Q(
        g4388) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n8684), .CLK(n9099), .Q(
        g6275) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n8684), .CLK(n9099), .Q(
        g6311), .QN(n8208) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n8684), .CLK(n9099), .Q(
        g8916) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n8656), .CLK(n9071), .Q(
        g1041), .QN(n8054) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n8665), .CLK(n9080), .Q(
        test_so34), .QN(n8636) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n8674), .CLK(n9089), 
        .Q(g2537) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n8659), .CLK(n9074), .Q(
        g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n8659), .CLK(n9074), .Q(
        g4430), .QN(n8121) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n8739), .CLK(n9154), .Q(
        n9325) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n8684), .CLK(n9099), .Q(
        g4826) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n8692), .CLK(n9107), .Q(
        g6239) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n8709), .CLK(n9124), .Q(
        g232), .QN(n8308) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n8709), .CLK(n9124), .Q(
        g5268) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n8709), .CLK(n9124), .Q(
        g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n8666), .CLK(n9081), .Q(
        n9324) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n8666), .CLK(n9081), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n8680), .CLK(n9095), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n8680), .CLK(n9095), .Q(
        test_so35), .QN(n8090) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n8696), .CLK(n9111), 
        .Q(g1890) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n8687), .CLK(n9102), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n8660), .CLK(n9075), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n8660), .CLK(n9075), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n8684), .CLK(n9099), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n8700), .CLK(n9115), .Q(
        g4308) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n8657), .CLK(n9072), .Q(
        g475) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n8692), .CLK(n9107), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n8692), .CLK(n9107), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n8642), .CLK(n9057), .Q(
        n9322), .QN(DFF_514_n1) );
  SDFFX1 DFF_515_Q_reg ( .D(n422), .SI(n9322), .SE(n8642), .CLK(n9057), .Q(
        g12184), .QN(n8627) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n8642), .CLK(n9057), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n8727), .CLK(n9142), .Q(
        test_so36), .QN(n8599) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n8694), .CLK(n9109), 
        .Q(g1992) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n8694), .CLK(n9109), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n8707), .CLK(n9122), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n8708), .CLK(n9123), .Q(
        g832), .QN(n8519) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n8708), .CLK(n9123), .Q(
        g5897) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n8708), .CLK(n9123), .Q(
        g25689) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n8708), .CLK(n9123), .Q(
        g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n8721), .CLK(n9136), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n8721), .CLK(n9136), .Q(
        g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n8652), .CLK(n9067), .Q(
        g2902), .QN(n8546) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n8734), .CLK(n9149), .Q(
        g333), .QN(n8438) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n8735), .CLK(n9150), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n8746), .CLK(n9161), .Q(
        test_so37) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n8687), .CLK(n9102), 
        .Q(g3684) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n8687), .CLK(n9102), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n8718), .CLK(n9133), .Q(
        g14597) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n8703), .CLK(n9118), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n8680), .CLK(n9095), .Q(
        g5406), .QN(n5992) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n8680), .CLK(n9095), .Q(
        g269), .QN(n8189) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n8657), .CLK(n9072), .Q(
        g401), .QN(n8508) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n8689), .CLK(n9104), .Q(
        g6040), .QN(n8300) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n8657), .CLK(n9072), .Q(
        g441), .QN(n8184) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n8680), .CLK(n9095), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n8643), .CLK(n9058), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n8643), .CLK(n9058), .Q(
        g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n8742), .CLK(n9157), .Q(
        test_so38), .QN(n8584) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n8652), .CLK(n9067), 
        .Q(g3957), .QN(n8385) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n8691), .CLK(n9106), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n8678), .CLK(n9093), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n8678), .CLK(n9093), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n8658), .CLK(n9073), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n8671), .CLK(n9086), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n8716), .CLK(n9131), .Q(
        g3498) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n8661), .CLK(n9076), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n8708), .CLK(n9123), .Q(
        g14201) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n8665), .CLK(n9080), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n8693), .CLK(n9108), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n8703), .CLK(n9118), .Q(
        g1608) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n8704), .CLK(n9119), .Q(
        test_so39) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n8718), .CLK(n9133), 
        .Q(g17577), .QN(n8372) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n8736), .CLK(n9151), .Q(
        g1779) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n8649), .CLK(n9064), .Q(
        g2652), .QN(n8231) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n8649), .CLK(n9064), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n8743), .CLK(n9158), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n8744), .CLK(n9159), .Q(
        g661) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n8687), .CLK(n9102), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n8719), .CLK(n9134), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n8650), .CLK(n9065), .Q(
        g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n8650), .CLK(n9065), .Q(
        g1361), .QN(n8171) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n8691), .CLK(n9106), .Q(
        g6235) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n8722), .CLK(n9137), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n8665), .CLK(n9080), .Q(
        test_so40) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n8658), .CLK(n9073), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n8647), .CLK(n9062), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n8719), .CLK(n9134), .Q(
        g6555), .QN(n8495) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n8708), .CLK(n9123), .Q(
        g14189) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n8699), .CLK(n9114), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n8672), .CLK(n9087), .Q(
        g6621) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n8677), .CLK(n9092), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n8697), .CLK(n9112), .Q(
        g3897) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n8658), .CLK(n9073), .Q(
        g538) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n8687), .CLK(n9102), .Q(
        g2606) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n8687), .CLK(n9102), .Q(
        g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n8659), .CLK(n9074), .Q(
        test_so41), .QN(n8634) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n8679), .CLK(n9094), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n8722), .CLK(n9137), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n8722), .CLK(n9137), .Q(
        g13259), .QN(n8527) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n8658), .CLK(n9073), .Q(
        g405), .QN(n8509) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n8726), .CLK(n9141), .Q(
        g5216), .QN(n8321) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n8734), .CLK(n9149), .Q(
        g6494), .QN(n8528) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n8644), .CLK(n9059), .Q(
        g4669) );
  SDFFX1 DFF_606_Q_reg ( .D(n631), .SI(g4669), .SE(n8705), .CLK(n9120), .Q(
        g996) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n8686), .CLK(n9101), .Q(
        g4531), .QN(n15223) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n8702), .CLK(n9117), .Q(
        g2860), .QN(n8452) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n8668), .CLK(n9083), .Q(
        g4743) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n8671), .CLK(n9086), .Q(
        g6593) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n8671), .CLK(n9086), .Q(
        test_so42) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n8659), .CLK(n9074), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n8700), .CLK(n9115), .Q(
        g1413) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n8700), .CLK(n9115), 
        .Q(g26960) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n8718), .CLK(n9133), .Q(
        g13039), .QN(n8351) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n8734), .CLK(n9149), .Q(
        g6641), .QN(n8202) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n8734), .CLK(n9149), .Q(
        g6), .QN(n8117) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n8714), .CLK(n9129), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n8566), .SI(g1936), .SE(n8714), .CLK(n9129), .Q(
        g55) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n8714), .CLK(n9129), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n8714), .CLK(n9129), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n8700), .CLK(n9115), .Q(
        g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n8701), .CLK(n9116), .Q(
        n9314) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n8730), .CLK(n9145), .Q(
        test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n8645), .CLK(n9060), 
        .Q(g5571) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n8686), .CLK(n9101), .Q(
        g3578) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n8719), .CLK(n9134), .Q(
        g9555) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n8677), .CLK(n9092), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n8677), .CLK(n9092), .Q(
        g3582) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n8683), .CLK(n9098), .Q(
        g6271) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n8731), .CLK(n9146), .Q(
        g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n8711), .CLK(n9126), .Q(
        g2380), .QN(n8102) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n8726), .CLK(n9141), .Q(
        g5196) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n8694), .CLK(n9109), .Q(
        g3227) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n8698), .CLK(n9113), .Q(
        n9312) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n8705), .CLK(n9120), .Q(
        g14518) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n8705), .CLK(n9120), .Q(
        test_so44), .QN(n8617) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n8725), .CLK(n9140), 
        .Q(g6541) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n8703), .CLK(n9118), .Q(
        g3203), .QN(n8368) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n8703), .CLK(n9118), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n8689), .CLK(n9104), .Q(
        g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n8689), .CLK(n9104), .Q(
        g262), .QN(n8188) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n8689), .CLK(n9104), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n8653), .CLK(n9068), .Q(
        g5467), .QN(n8124) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n8653), .CLK(n9068), .Q(
        g460) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n8698), .CLK(n9113), .Q(
        g6209), .QN(n8491) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n8735), .CLK(n9150), .Q(
        g29211) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n8675), .CLK(n9090), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n8675), .CLK(n9090), .Q(
        g655), .QN(n8550) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n8675), .CLK(n9090), .Q(
        test_so45), .QN(n8606) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n8720), .CLK(n9135), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n8720), .CLK(n9135), .Q(
        g5256), .QN(n8213) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n8738), .CLK(n9153), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n8676), .CLK(n9091), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n8724), .CLK(n9139), .Q(
        g13906) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n8644), .CLK(n9059), .Q(
        g4423) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n8644), .CLK(n9059), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n8721), .CLK(n9136), .Q(
        g5685), .QN(n8410) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n8707), .CLK(n9122), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n8653), .CLK(n9068), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n8732), .CLK(n9147), .Q(
        g3247), .QN(n8194) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n8693), .CLK(n9108), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n8693), .CLK(n9108), .Q(
        test_so46), .QN(DFF_672_n1) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n8685), .CLK(n9100), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n8685), .CLK(n9100), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n8692), .CLK(n9107), .Q(
        g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n8692), .CLK(n9107), .Q(
        g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n8679), .CLK(n9094), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n8667), .CLK(n9082), .Q(
        g5817), .QN(n8073) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n8664), .CLK(n9079), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n8740), .CLK(n9155), .Q(
        g2648), .QN(n8106) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n8699), .CLK(n9114), .Q(
        g6736), .QN(n8432) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n8687), .CLK(n9102), .Q(
        g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n8691), .CLK(n9106), .Q(
        g4072), .QN(n8543) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n8735), .CLK(n9150), .Q(
        g7540) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n8735), .CLK(n9150), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n8677), .CLK(n9092), 
        .Q(g3466) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n8685), .CLK(n9100), .Q(
        g4116) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n8680), .CLK(n9095), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n8741), .CLK(n9156), .Q(
        g4434), .QN(n8119) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n8743), .CLK(n9158), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n8668), .CLK(n9083), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n8721), .CLK(n9136), .Q(
        g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n8669), .CLK(n9084), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n8695), .CLK(n9110), .Q(
        g3333) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n8695), .CLK(n9110), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n8731), .CLK(n9146), .Q(
        g4681), .QN(n8436) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n8663), .CLK(n9078), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n8687), .CLK(n9102), .Q(
        test_so48), .QN(n8619) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n8704), .CLK(n9119), 
        .Q(g8789), .QN(n8177) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n8740), .CLK(n9155), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n8702), .CLK(n9117), .Q(
        g2988), .QN(n8485) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n8716), .CLK(n9131), .Q(
        g3538) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n8658), .CLK(n9073), .Q(
        g301), .QN(n8545) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n8738), .CLK(n9153), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n8738), .CLK(n9153), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n8689), .CLK(n9104), .Q(
        g17291), .QN(n8150) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n8687), .CLK(n9102), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n8746), .CLK(n9161), .Q(
        g5011) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n8746), .CLK(n9161), .Q(
        g199), .QN(n8469) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n8668), .CLK(n9083), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n8713), .CLK(n9128), .Q(
        test_so49), .QN(n8608) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n8707), .CLK(n9122), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n8707), .CLK(n9122), .Q(
        g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n8740), .CLK(n9155), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n8740), .CLK(n9155), .Q(
        g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n8641), .CLK(n9056), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n8727), .CLK(n9142), .Q(
        g5863), .QN(n8493) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n8690), .CLK(n9105), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n8674), .CLK(n9089), .Q(
        g2518), .QN(n8230) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n8649), .CLK(n9064), .Q(
        g2567) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n8660), .CLK(n9075), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n8695), .CLK(n9110), .Q(
        g3263), .QN(n8193) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n8671), .CLK(n9086), .Q(
        g6613) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n8688), .CLK(n9103), .Q(
        test_so50), .QN(n8610) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n8734), .CLK(n9149), 
        .Q(g6444), .QN(n5990) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n8646), .CLK(n9061), .Q(
        g2965), .QN(n8536) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n8727), .CLK(n9142), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n8689), .CLK(n9104), .Q(
        n9303) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n8653), .CLK(n9068), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n8730), .CLK(n9145), .Q(
        g17646), .QN(n8377) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n8722), .CLK(n9137), .Q(
        g3562) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n8722), .CLK(n9137), .Q(
        g10122_Tj), .QN(n8086) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n8737), .CLK(n9152), 
        .Q(g1404), .QN(n8167) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n8643), .CLK(n9058), .Q(
        g3817), .QN(n8072) );
  SDFFX1 DFF_743_Q_reg ( .D(n8572), .SI(g3817), .SE(n8668), .CLK(n9083), .Q(
        n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n8713), .CLK(n9128), .Q(
        g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n8723), .CLK(n9138), .Q(
        test_so51), .QN(n8631) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n8686), .CLK(n9101), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n8664), .CLK(n9079), .Q(
        g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n8656), .CLK(n9071), .Q(
        g2878), .QN(n8461) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n8726), .CLK(n9141), .Q(
        g5220) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n8661), .CLK(n9076), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n8661), .CLK(n9076), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n8720), .CLK(n9135), .Q(
        g316) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n8654), .CLK(n9069), .Q(
        g1277), .QN(n8467) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n8668), .CLK(n9083), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n8715), .CLK(n9130), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n8656), .CLK(n9071), .Q(
        g2882), .QN(n8547) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n8662), .CLK(n9077), .Q(
        test_so52), .QN(n8471) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n8714), .CLK(n9129), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n8714), .CLK(n9129), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n8648), .CLK(n9063), .Q(g8), .QN(n8533) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n8650), .CLK(n9065), .Q(
        g2799) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n8709), .CLK(n9124), .Q(
        g14167) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n8718), .CLK(n9133), .Q(
        g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n8740), .CLK(n9155), .Q(
        g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n8745), .CLK(n9160), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n8674), .CLK(n9089), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n8720), .CLK(n9135), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n8659), .CLK(n9074), .Q(
        g550), .QN(n8468) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n8709), .CLK(n9124), .Q(
        g255), .QN(n8187) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n8740), .CLK(n9155), .Q(
        test_so53), .QN(n8633) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n8726), .CLK(n9141), 
        .Q(g5240) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n8704), .CLK(n9119), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n8704), .CLK(n9119), .Q(
        g3863), .QN(n8494) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n8740), .CLK(n9155), .Q(
        g1959), .QN(n8229) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n8644), .CLK(n9059), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n8672), .CLK(n9087), .Q(
        g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n8737), .CLK(n9152), .Q(
        g17764), .QN(n8389) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n8655), .CLK(n9070), .Q(
        g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n8683), .CLK(n9098), .Q(
        g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n8721), .CLK(n9136), .Q(
        g17678), .QN(n8380) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n8705), .CLK(n9120), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n8705), .CLK(n9120), .Q(
        g16693), .QN(n8386) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n8736), .CLK(n9151), .Q(
        test_so54) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n8657), .CLK(n9072), 
        .Q(g1002), .QN(n8166) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n8676), .CLK(n9091), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n8676), .CLK(n9091), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n8705), .CLK(n9120), .Q(
        g1236), .QN(n8152) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n8730), .CLK(n9145), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n8674), .CLK(n9089), .Q(
        g2476), .QN(n8481) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n8677), .CLK(n9092), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n8711), .CLK(n9126), .Q(
        g2375), .QN(n8132) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n8644), .CLK(n9059), .Q(
        g63) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n8722), .CLK(n9137), .Q(
        g17739), .QN(n8285) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n8722), .CLK(n9137), .Q(
        g358), .QN(n8190) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n8722), .CLK(n9137), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n8723), .CLK(n9138), .Q(
        test_so55), .QN(n8607) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n8728), .CLK(n9143), 
        .Q(g3161), .QN(n8475) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n8701), .CLK(n9116), .Q(
        g2384), .QN(n8225) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n8699), .CLK(n9114), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n8738), .CLK(n9153), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n8739), .CLK(n9154), .Q(
        g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n8698), .CLK(n9113), .Q(
        g2024) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n8717), .CLK(n9132), .Q(
        g3451), .QN(n8530) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n8693), .CLK(n9108), .Q(
        g2795) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n8661), .CLK(n9076), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n8739), .CLK(n9154), .Q(
        g4527), .QN(n8448) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n8666), .CLK(n9081), .Q(
        g1844) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n8666), .CLK(n9081), .Q(
        g5937) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n8743), .CLK(n9158), .Q(
        test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n8674), .CLK(n9089), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n8721), .CLK(n9136), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n8704), .CLK(n9119), .Q(
        g2643), .QN(n8131) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n8704), .CLK(n9119), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n8658), .CLK(n9073), .Q(
        g8358), .QN(n8169) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n8674), .CLK(n9089), .Q(
        n9295) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n8674), .CLK(n9089), .Q(
        g5156) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n8674), .CLK(n9089), .Q(
        g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n8675), .CLK(n9090), .Q(
        n9294), .QN(DFF_829_n1) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n8717), .CLK(n9132), .Q(
        g8279) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n8682), .CLK(n9097), .Q(
        g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n8696), .CLK(n9111), .Q(
        g1955), .QN(n8099) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n8739), .CLK(n9154), .Q(
        test_so57), .QN(n8597) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n8671), .CLK(n9086), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n8737), .CLK(n9152), .Q(
        g14749) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n8678), .CLK(n9093), .Q(
        g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n8660), .CLK(n9075), .Q(
        g6098), .QN(n5988) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n8728), .CLK(n9143), .Q(
        g3147) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n8741), .CLK(n9156), .Q(
        g3347), .QN(n8296) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n8670), .CLK(n9085), .Q(
        g2269) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n8670), .CLK(n9085), .Q(
        g191), .QN(n8170) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n8671), .CLK(n9086), .Q(
        g2712), .QN(n8083) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n8662), .CLK(n9077), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n8664), .CLK(n9079), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n8682), .CLK(n9097), .Q(
        test_so58), .QN(n8587) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n8688), .CLK(n9103), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n8731), .CLK(n9146), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n8652), .CLK(n9067), .Q(
        g2927), .QN(n8538) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n8706), .CLK(n9121), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n8729), .CLK(n9144), .Q(
        g5929) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n8740), .CLK(n9155), .Q(
        g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n8740), .CLK(n9155), .Q(
        g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n8648), .CLK(n9063), .Q(
        g4035) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n8649), .CLK(n9064), .Q(
        g2946), .QN(n8541) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n8662), .CLK(n9077), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n8691), .CLK(n9106), .Q(
        g4082), .QN(n8163) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n8734), .CLK(n9149), .Q(
        g9743) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n8693), .CLK(n9108), .Q(
        test_so59), .QN(n8637) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n8661), .CLK(n9076), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n8741), .CLK(n9156), .Q(
        g1620) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n8651), .CLK(n9066), .Q(
        g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n8651), .CLK(n9066), .Q(
        g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n8662), .CLK(n9077), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n8697), .CLK(n9112), .Q(
        g3937) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n8707), .CLK(n9122), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n8714), .CLK(n9129), .Q(
        g1249) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n8707), .CLK(n9122), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n8728), .CLK(n9143), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n8661), .CLK(n9076), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n8642), .CLK(n9057), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n8710), .CLK(n9125), .Q(
        test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n8737), .CLK(n9152), 
        .Q(g5949), .QN(n8216) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n8668), .CLK(n9083), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n8668), .CLK(n9083), .Q(
        g904) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n8702), .CLK(n9117), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n8746), .CLK(n9161), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n8641), .CLK(n9056), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n8645), .CLK(n9060), .Q(
        g5603), .QN(n8198) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n8673), .CLK(n9088), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n8673), .CLK(n9088), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n8688), .CLK(n9103), .Q(
        g2437) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n8688), .CLK(n9103), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n8712), .CLK(n9127), .Q(
        g2208), .QN(n8479) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n8649), .CLK(n9064), .Q(
        test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n8691), .CLK(n9106), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n8644), .CLK(n9059), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n8665), .CLK(n9080), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n8730), .CLK(n9145), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n8733), .CLK(n9148), .Q(
        g5583) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n8676), .CLK(n9091), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n8719), .CLK(n9134), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n8718), .CLK(n9133), .Q(
        g17743), .QN(n8399) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n8652), .CLK(n9067), .Q(
        g2917), .QN(n8548) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n8653), .CLK(n9068), .Q(
        g686) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n8654), .CLK(n9069), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n8651), .CLK(n9066), .Q(
        g671), .QN(n8079) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n8720), .CLK(n9135), .Q(
        test_so62), .QN(n8620) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n8692), .CLK(n9107), 
        .Q(g6283) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n8718), .CLK(n9133), .Q(
        g14705) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n8718), .CLK(n9133), .Q(
        g17519), .QN(n8268) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n8718), .CLK(n9133), .Q(
        g8784), .QN(n15234) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n8717), .CLK(n9132), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n8717), .CLK(n9132), .Q(
        g4489) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n8736), .CLK(n9151), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n8654), .CLK(n9069), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n8682), .CLK(n9097), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n8691), .CLK(n9106), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n8653), .CLK(n9068), .Q(
        g3929) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n8653), .CLK(n9068), .Q(
        g5503) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n8655), .CLK(n9070), .Q(
        test_so63), .QN(n8464) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n8727), .CLK(n9142), 
        .Q(g5925) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n8695), .CLK(n9110), .Q(
        g1124) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n8673), .CLK(n9088), .Q(
        g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n8726), .CLK(n9141), .Q(
        g5224) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n8698), .CLK(n9113), .Q(
        g2012) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n8698), .CLK(n9113), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n8675), .CLK(n9090), .Q(
        g5120), .QN(n8123) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n8675), .CLK(n9090), .Q(
        g17674), .QN(n8283) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n8701), .CLK(n9116), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n8701), .CLK(n9116), .Q(
        g4438), .QN(n8442) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n8688), .CLK(n9103), .Q(
        g2429) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n8693), .CLK(n9108), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n8654), .CLK(n9069), .Q(
        test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n8646), .CLK(n9061), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n8685), .CLK(n9100), .Q(
        g18881), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n8719), .CLK(n9134), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n8692), .CLK(n9107), .Q(
        g1199), .QN(n8486) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n8648), .CLK(n9063), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n8645), .CLK(n9060), .Q(
        g5547) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n8660), .CLK(n9075), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n8732), .CLK(n9147), .Q(
        g16744), .QN(n8292) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n8738), .CLK(n9153), .Q(
        g2338) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n8738), .CLK(n9153), .Q(
        g8919), .QN(n15232) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n8683), .CLK(n9098), .Q(
        g6247), .QN(n8429) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n8696), .CLK(n9111), .Q(
        g2791) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n8697), .CLK(n9112), .Q(
        test_so65), .QN(n8618) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n8641), .CLK(n9056), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n8729), .CLK(n9144), .Q(
        g5945) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n8711), .CLK(n9126), .Q(
        g5244) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n8712), .CLK(n9127), .Q(
        g2759), .QN(n8051) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n8683), .CLK(n9098), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n8676), .CLK(n9091), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n8654), .CLK(n9069), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n8645), .CLK(n9060), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n8658), .CLK(n9073), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n8725), .CLK(n9140), .Q(
        g6609) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n8725), .CLK(n9140), .Q(
        g5517), .QN(n8492) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n8745), .CLK(n9160), .Q(
        g2449) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n8745), .CLK(n9160), .Q(
        test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n8685), .CLK(n9100), 
        .Q(n9281) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n8685), .CLK(n9100), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n8662), .CLK(n9077), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n8690), .CLK(n9105), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n8690), .CLK(n9105), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n8661), .CLK(n9076), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n8734), .CLK(n9149), .Q(
        g6589) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n8696), .CLK(n9111), .Q(
        n9280) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n8718), .CLK(n9133), .Q(
        g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n8737), .CLK(n9152), .Q(
        g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n8657), .CLK(n9072), .Q(
        g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n8696), .CLK(n9111), .Q(
        g1870) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n8696), .CLK(n9111), .Q(
        test_so67), .QN(n8624) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n8745), .CLK(n9160), 
        .Q(g1825), .QN(n8223) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n8656), .CLK(n9071), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n8719), .CLK(n9134), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n8719), .CLK(n9134), 
        .Q(g8283) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n8720), .CLK(n9135), .Q(
        g3546) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n8726), .CLK(n9141), .Q(
        g5236) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n8651), .CLK(n9066), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n8736), .CLK(n9151), .Q(
        g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n8652), .CLK(n9067), .Q(
        g3925) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n8668), .CLK(n9083), .Q(
        g6509), .QN(n8111) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n8680), .CLK(n9095), .Q(
        g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n8674), .CLK(n9089), .Q(
        g2504), .QN(n8484) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n8724), .CLK(n9139), .Q(
        test_so68), .QN(n8602) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n8673), .CLK(n9088), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n8673), .CLK(n9088), .Q(
        g8917), .QN(n15230) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n8712), .CLK(n9127), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n8702), .CLK(n9117), .Q(
        g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n8743), .CLK(n9158), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n8693), .CLK(n9108), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n8717), .CLK(n9132), .Q(
        g8235) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n8685), .CLK(n9100), .Q(
        g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n8705), .CLK(n9120), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n8706), .CLK(n9121), .Q(
        g4405), .QN(n8561) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n8709), .CLK(n9124), .Q(
        g872) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n8679), .CLK(n9094), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n8719), .CLK(n9134), .Q(
        test_so69), .QN(n8614) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n8678), .CLK(n9093), 
        .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n8733), .CLK(n9148), .Q(
        g5563), .QN(n8327) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n8714), .CLK(n9129), .Q(
        g1395), .QN(n8501) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n8714), .CLK(n9129), .Q(
        g1913) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n8711), .CLK(n9126), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n8691), .CLK(n9106), .Q(
        g6263) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n8648), .CLK(n9063), .Q(
        n9276), .QN(DFF_1012_n1) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n8648), .CLK(n9063), .Q(
        g3945) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n8735), .CLK(n9150), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n8742), .CLK(n9157), .Q(
        g4473), .QN(n8140) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n8742), .CLK(n9157), .Q(
        g1266), .QN(n8504) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n8742), .CLK(n9157), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n8651), .CLK(n9066), .Q(
        test_so70), .QN(n8603) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n8710), .CLK(n9125), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n8642), .CLK(n9057), .Q(
        g5471), .QN(n8080) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n8690), .CLK(n9105), .Q(
        g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n8690), .CLK(n9105), .Q(
        g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n8672), .CLK(n9087), .Q(
        g6605) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n8673), .CLK(n9088), .Q(
        n9274) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n8670), .CLK(n9085), .Q(
        g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n8682), .CLK(n9097), .Q(
        g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n8682), .CLK(n9097), .Q(
        g2491) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n8682), .CLK(n9097), .Q(
        g4849), .QN(n8557) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n8697), .CLK(n9112), .Q(
        g2169) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n8671), .CLK(n9086), .Q(
        n9273), .QN(n15229) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n8671), .CLK(n9086), .Q(
        test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n8665), .CLK(n9080), 
        .Q(g29219) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n8665), .CLK(n9080), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n8702), .CLK(n9117), .Q(
        g2868), .QN(n8451) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n8677), .CLK(n9092), .Q(
        g2767) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n8678), .CLK(n9093), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n8721), .CLK(n9136), .Q(
        g16718), .QN(n8281) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n8681), .CLK(n9096), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n8682), .CLK(n9097), .Q(
        g5212), .QN(n8373) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n8682), .CLK(n9097), .Q(
        g4245), .QN(n5640) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n8653), .CLK(n9068), .Q(
        g645), .QN(n8182) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n8682), .CLK(n9097), .Q(
        g4291), .QN(n8472) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n8744), .CLK(n9159), .Q(
        g29212) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n8658), .CLK(n9073), 
        .Q(test_so72), .QN(n8593) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n8696), .CLK(n9111), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n8720), .CLK(n9135), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n8704), .CLK(n9119), .Q(
        g8788) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n8697), .CLK(n9112), .Q(
        g2246), .QN(n8105) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n8666), .CLK(n9081), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n8731), .CLK(n9146), .Q(
        g3590) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n8657), .CLK(n9072), .Q(
        g392), .QN(n8510) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n8703), .CLK(n9118), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n8725), .CLK(n9140), .Q(
        g6505), .QN(n8138) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n8735), .CLK(n9150), .Q(
        g1221), .QN(n8445) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n8708), .CLK(n9123), .Q(
        g5921) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n8708), .CLK(n9123), .Q(
        g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n8747), .CLK(n9162), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n8671), .CLK(
        n9086), .Q(g218), .QN(n8441) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n8694), .CLK(n9109), .Q(
        g1932) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n8712), .CLK(n9127), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n8680), .CLK(n9095), .Q(
        g5062), .QN(n8498) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n8642), .CLK(n9057), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n8642), .CLK(n9057), .Q(
        g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n8725), .CLK(n9140), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n8689), .CLK(n9104), .Q(
        g1677) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n8689), .CLK(n9104), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n8646), .CLK(n9061), .Q(
        g2671) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n8726), .CLK(n9141), .Q(
        g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n8706), .CLK(n9121), 
        .Q(g7243), .QN(n8562) );
  SDFFX1 DFF_1074_Q_reg ( .D(n8566), .SI(g7243), .SE(n8714), .CLK(n9129), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n8746), .CLK(n9161), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n8641), .CLK(n9056), .Q(
        g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n8641), .CLK(n9056), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n8710), .CLK(n9125), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n8710), .CLK(n9125), .Q(
        g11678) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n8649), .CLK(n9064), 
        .Q(g2638), .QN(n8512) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n8685), .CLK(n9100), .Q(
        g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n8729), .CLK(n9144), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n8729), .CLK(n9144), .Q(
        g5941) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n8688), .CLK(n9103), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n8688), .CLK(n9103), .Q(
        g13068), .QN(n8408) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n8688), .CLK(n9103), .Q(
        g25) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n8646), .CLK(n9061), .Q(
        test_so75) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n8661), .CLK(n9076), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n8712), .CLK(n9127), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n8648), .CLK(n9063), .Q(
        n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n8712), .CLK(n9127), .Q(
        g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n8722), .CLK(n9137), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n8726), .CLK(n9141), .Q(
        g5252) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n8697), .CLK(n9112), .Q(
        g2165) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n8649), .CLK(n9064), .Q(
        g2571) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n8701), .CLK(n9116), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n8719), .CLK(n9134), .Q(
        g8403) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n8720), .CLK(n9135), .Q(
        g14673) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n8689), .CLK(n9104), 
        .Q(test_so76), .QN(n8604) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n8665), .CLK(n9080), 
        .Q(g2827) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n8708), .CLK(n9123), .Q(
        g14217) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n8736), .CLK(n9151), 
        .Q(g4859), .QN(n8555) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n8657), .CLK(n9072), .Q(
        g424), .QN(n8507) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n8654), .CLK(n9069), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n8670), .CLK(n9085), .Q(
        g17423), .QN(n8159) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n8694), .CLK(n9109), 
        .Q(n9265), .QN(n8630) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n8650), .CLK(n9065), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n8666), .CLK(n9081), .Q(
        g1821), .QN(n8100) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n8688), .CLK(n9103), .Q(
        g2509), .QN(n8130) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n8641), .CLK(n9056), .Q(
        g5073), .QN(n8128) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n8742), .CLK(n9157), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n8717), .CLK(n9132), 
        .Q(g8353) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n8718), .CLK(n9133), .Q(
        g13085), .QN(n8428) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n8672), .CLK(n9087), 
        .Q(g6633) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n8655), .CLK(n9070), .Q(
        g5124), .QN(n8071) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n8705), .CLK(n9120), 
        .Q(g17400), .QN(n8155) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n8683), .CLK(n9098), 
        .Q(g6303) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n8641), .CLK(n9056), .Q(
        g5069), .QN(n8127) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n8701), .CLK(n9116), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n8736), .CLK(n9151), .Q(
        g650), .QN(n8183) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n8736), .CLK(n9151), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n8697), .CLK(n9112), .Q(
        g3921) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n8690), .CLK(n9105), .Q(
        test_so78) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n8699), .CLK(n9114), 
        .Q(g6732), .QN(n8433) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n8699), .CLK(n9114), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n8699), .CLK(n9114), .Q(
        g1061), .QN(n8168) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n8716), .CLK(n9131), .Q(
        g3462), .QN(n8126) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n8698), .CLK(n9113), .Q(
        g2181) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n8698), .CLK(n9113), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n8651), .CLK(n9066), .Q(
        g1756) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n8727), .CLK(n9142), .Q(
        g5849) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n8684), .CLK(n9099), .Q(
        g4112), .QN(n8431) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n8646), .CLK(n9061), .Q(
        n9262), .QN(n15224) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n8646), .CLK(n9061), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n8673), .CLK(n9088), .Q(
        test_so79), .QN(n8585) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n8656), .CLK(n9071), 
        .Q(g1046) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n8723), .CLK(n9138), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n8723), .CLK(n9138), .Q(
        g4401) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n8725), .CLK(n9140), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n8725), .CLK(n9140), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n8725), .CLK(n9140), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n8681), .CLK(n9096), .Q(
        g2950), .QN(n8458) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n8681), .CLK(n9096), .Q(
        g1345), .QN(n8165) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n8669), .CLK(n9084), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n8669), .CLK(n9084), .Q(
        g14421) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n8669), .CLK(n9084), 
        .Q(g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n8699), .CLK(n9114), .Q(
        test_so80), .QN(n8592) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n8700), .CLK(n9115), 
        .Q(g1536) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n8652), .CLK(n9067), .Q(
        g3941) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n8723), .CLK(n9138), .Q(
        g370), .QN(n8539) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n8667), .CLK(n9082), .Q(
        g5694), .QN(n8304) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n8746), .CLK(n9161), .Q(
        g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n8653), .CLK(n9068), .Q(
        g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n8732), .CLK(n9147), .Q(
        g3219) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n8745), .CLK(n9160), .Q(
        g1811) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n8672), .CLK(n9087), .Q(
        g6601), .QN(n8333) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n8673), .CLK(n9088), .Q(
        g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n8696), .CLK(n9111), .Q(
        g1874) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n8707), .CLK(n9122), .Q(
        test_so81), .QN(n8590) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n8725), .CLK(n9140), 
        .Q(g6581) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n8671), .CLK(n9086), .Q(
        g6597), .QN(n8392) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n8719), .CLK(n9134), .Q(
        g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n8686), .CLK(n9101), .Q(
        g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n8702), .CLK(n9117), .Q(
        g2890), .QN(n8465) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n8736), .CLK(n9151), .Q(
        g1978) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n8689), .CLK(n9104), .Q(
        g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n8646), .CLK(n9061), .Q(
        g112), .QN(n8185) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n8643), .CLK(n9058), .Q(
        g2856), .QN(n8549) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n8736), .CLK(n9151), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n8711), .CLK(n9126), .Q(
        g17722), .QN(n8391) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n8711), .CLK(n9126), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n8685), .CLK(n9100), 
        .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n8678), .CLK(n9093), .Q(
        g6390), .QN(n8298) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n8700), .CLK(n9115), .Q(
        g1542), .QN(n8487) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n8700), .CLK(n9115), .Q(
        g4258) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n8718), .CLK(n9133), .Q(
        g4818), .QN(n5636) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n8680), .CLK(n9095), .Q(
        g5033), .QN(n8518) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n8692), .CLK(n9107), .Q(
        g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n8734), .CLK(n9149), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n8699), .CLK(n9114), .Q(
        g3849) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n8699), .CLK(n9114), .Q(
        g17778), .QN(n8290) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n8741), .CLK(n9156), 
        .Q(g3199) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n8746), .CLK(n9161), .Q(
        test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n8683), .CLK(n9098), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n8676), .CLK(n9091), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n8729), .CLK(n9144), .Q(
        g5913), .QN(n8407) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n8696), .CLK(n9111), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n8679), .CLK(n9094), .Q(
        g6163) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n8708), .CLK(n9123), .Q(
        g4125), .QN(n8430) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n8733), .CLK(n9148), .Q(
        g4821) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n8742), .CLK(n9157), .Q(
        g4939), .QN(n5776) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n8695), .CLK(n9110), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n8694), .CLK(n9109), 
        .Q(g3207), .QN(n8318) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n8694), .CLK(n9109), .Q(
        g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n8695), .CLK(n9110), .Q(
        test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n8746), .CLK(n9161), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n8655), .CLK(n9070), .Q(
        g5248) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n8643), .CLK(n9058), .Q(
        g2126) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n8733), .CLK(n9148), .Q(
        g3694), .QN(n8302) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n8642), .CLK(n9057), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n8642), .CLK(n9057), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n8641), .CLK(n9056), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n8732), .CLK(n9147), .Q(
        g3215) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n8732), .CLK(n9147), .Q(
        g16748), .QN(n8384) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n8732), .CLK(n9147), 
        .Q(n9255), .QN(n8629) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n8659), .CLK(n9074), .Q(
        g4427), .QN(n8179) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n8659), .CLK(n9074), .Q(
        test_so85), .QN(n8589) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n8651), .CLK(n9066), 
        .Q(g2779) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n8704), .CLK(n9119), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n8741), .CLK(n9156), .Q(
        g7245), .QN(DFF_1225_n1) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n8647), .CLK(n9062), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n8724), .CLK(n9139), .Q(
        g1367), .QN(n8156) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n8724), .CLK(n9139), .Q(
        g5112), .QN(n8096) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n8724), .CLK(n9139), .Q(
        g19), .QN(n8532) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n8684), .CLK(n9099), .Q(
        g4145), .QN(n8449) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n8697), .CLK(n9112), .Q(
        g2161) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n8723), .CLK(n9138), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n8711), .CLK(n9126), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n8649), .CLK(n9064), .Q(
        test_so86) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n8661), .CLK(n9076), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n8690), .CLK(n9105), .Q(
        g2051), .QN(n8483) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n8693), .CLK(n9108), .Q(
        g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n8664), .CLK(n9079), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n8662), .CLK(n9077), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n8662), .CLK(n9077), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n8666), .CLK(n9081), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n8686), .CLK(n9101), .Q(
        g3594) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n8701), .CLK(n9116), .Q(
        g2999), .QN(n8466) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n8711), .CLK(n9126), .Q(
        g2303) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n8711), .CLK(n9126), .Q(
        g17688), .QN(n8276) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n8653), .CLK(n9068), 
        .Q(test_so87) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n8738), .CLK(n9153), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n8739), .CLK(n9154), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n8659), .CLK(n9074), .Q(
        g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n8737), .CLK(n9152), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n8666), .CLK(n9081), .Q(
        g5953) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n8650), .CLK(n9065), .Q(
        g8277), .QN(n8097) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n8650), .CLK(n9065), .Q(
        g1740) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n8731), .CLK(n9146), .Q(
        g3550) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n8643), .CLK(n9058), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n8643), .CLK(n9058), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n8721), .CLK(n9136), .Q(
        g14635) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n8732), .CLK(n9147), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n8652), .CLK(n9067), 
        .Q(g3913) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n8644), .CLK(n9059), .Q(
        g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n8647), .CLK(n9062), 
        .Q(g1687), .QN(n8104) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n8646), .CLK(n9061), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n8713), .CLK(n9128), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n8715), .CLK(n9130), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n8715), .CLK(n9130), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(n503), .SI(g2697), .SE(n8715), .CLK(n9130), .Q(
        g4417), .QN(n8048) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n8715), .CLK(n9130), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n8713), .CLK(n9128), .Q(
        g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n8714), .CLK(n9129), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n8666), .CLK(n9081), 
        .Q(test_so89), .QN(n8615) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n8647), .CLK(n9062), 
        .Q(g1710) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n8668), .CLK(n9083), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n8741), .CLK(n9156), .Q(
        g3255), .QN(n8366) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n8745), .CLK(n9160), .Q(
        g1691), .QN(n8227) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n8681), .CLK(n9096), .Q(
        g2936), .QN(n8459) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n8668), .CLK(n9083), .Q(
        g5644) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n8747), .CLK(n9162), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n8663), .CLK(n9078), .Q(
        g5352), .QN(n8434) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n8663), .CLK(n9078), .Q(
        g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n8651), .CLK(n9066), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n8681), .CLK(n9096), .Q(
        g2922) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n8695), .CLK(n9110), .Q(
        test_so90) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n8708), .CLK(n9123), 
        .Q(g5893) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n8721), .CLK(n9136), .Q(
        g16603), .QN(n8266) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n8672), .CLK(n9087), 
        .Q(g6617) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n8712), .CLK(n9127), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n8644), .CLK(n9059), .Q(
        g4512) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n8733), .CLK(n9148), .Q(
        g5599) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n8733), .CLK(n9148), .Q(
        g3401), .QN(n5986) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n8739), .CLK(n9154), .Q(
        g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n8739), .CLK(n9154), 
        .Q(g16722), .QN(n8394) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n8739), .CLK(n9154), 
        .Q(g29214), .QN(n5342) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n8669), .CLK(n9084), 
        .Q(g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n8703), .CLK(n9118), .Q(
        test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n8701), .CLK(n9116), 
        .Q(g5170), .QN(n8489) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n8720), .CLK(n9135), .Q(
        g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n8667), .CLK(n9082), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n8692), .CLK(n9107), .Q(
        g6299) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n8692), .CLK(n9107), .Q(
        g8416), .QN(n8526) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n8690), .CLK(n9105), .Q(
        g2079), .QN(n8513) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n8664), .CLK(n9079), .Q(
        g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n8687), .CLK(n9102), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n8687), .CLK(n9102), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n8657), .CLK(n9072), .Q(
        n9247), .QN(n15226) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n8657), .CLK(n9072), .Q(
        g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n8744), .CLK(n9159), .Q(
        test_so92) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n8697), .CLK(n9112), 
        .Q(g3953) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n8697), .CLK(n9112), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n8676), .CLK(n9091), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n8676), .CLK(n9091), .Q(
        n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n8739), .CLK(n9154), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n8691), .CLK(n9106), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n8735), .CLK(n9150), .Q(
        g5200), .QN(n8215) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n8736), .CLK(n9151), .Q(
        g4843), .QN(n8556) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n8680), .CLK(n9095), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n8670), .CLK(n9085), .Q(
        g2250), .QN(n8221) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n8720), .CLK(n9135), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n8743), .CLK(n9158), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n8674), .CLK(n9089), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n8667), .CLK(n9082), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n8667), .CLK(n9082), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n8681), .CLK(n9096), 
        .Q(g2912) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n8664), .CLK(n9079), .Q(
        g2357) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n8738), .CLK(n9153), .Q(
        g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n8658), .CLK(n9073), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n8655), .CLK(n9070), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n8725), .CLK(n9140), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n8669), .CLK(n9084), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n8648), .CLK(n9063), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n8712), .CLK(n9127), .Q(
        test_so94), .QN(n8596) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n8673), .CLK(n9088), 
        .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n8655), .CLK(n9070), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n8741), .CLK(n9156), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n8672), .CLK(n9087), .Q(
        g6657), .QN(n8201) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n8672), .CLK(n9087), .Q(
        g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n8697), .CLK(n9112), .Q(
        g3893), .QN(n8220) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n8694), .CLK(n9109), .Q(
        g3211) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n8721), .CLK(n9136), .Q(
        g13049), .QN(n8412) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n8721), .CLK(n9136), 
        .Q(g16624), .QN(n8367) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n8727), .CLK(n9142), 
        .Q(g5595) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n8686), .CLK(n9101), .Q(
        g3614), .QN(n8204) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n8702), .CLK(n9117), .Q(
        test_so95), .QN(n8625) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n8702), .CLK(n9117), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n8703), .CLK(n9118), .Q(
        g16686), .QN(n8365) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n8643), .CLK(n9058), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n8691), .CLK(n9106), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n8691), .CLK(n9106), .Q(
        g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n8709), .CLK(n9124), .Q(
        g5272), .QN(n8212) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n8710), .CLK(n9125), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n8744), .CLK(n9159), .Q(
        g728), .QN(n8192) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n8691), .CLK(n9106), .Q(
        g6295), .QN(n8209) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n8646), .CLK(n9061), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n8737), .CLK(n9152), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n8737), .CLK(n9152), .Q(
        test_so96), .QN(n8601) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n8734), .CLK(n9149), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n8669), .CLK(n9084), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n8731), .CLK(n9146), .Q(
        g4659), .QN(n8554) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n8731), .CLK(n9146), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n8678), .CLK(n9093), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n8698), .CLK(n9113), .Q(
        g2084), .QN(n8129) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n8728), .CLK(n9143), .Q(
        g3187) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n8729), .CLK(n9144), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n8649), .CLK(n9064), .Q(
        g2583) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n8646), .CLK(n9061), .Q(
        n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n8647), .CLK(n9062), .Q(
        g1094) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n8699), .CLK(n9114), .Q(
        test_so97), .QN(n8623) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n8682), .CLK(n9097), 
        .Q(g4284), .QN(n8511) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n8732), .CLK(n9147), .Q(
        g3191), .QN(n8196) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n8732), .CLK(n9147), .Q(
        g4239), .QN(n8142) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n8704), .CLK(n9119), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n8652), .CLK(n9067), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n8659), .CLK(n9074), .Q(
        g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n8723), .CLK(n9138), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n8698), .CLK(n9113), .Q(
        g2004) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n8674), .CLK(n9089), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n8719), .CLK(n9134), .Q(
        g5456), .QN(n8525) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n8746), .CLK(n9161), .Q(
        n6007), .QN(n8180) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n8746), .CLK(n9161), .Q(
        test_so98), .QN(n8622) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n8742), .CLK(n9157), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n8663), .CLK(n9078), .Q(
        g5348), .QN(n8435) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n8741), .CLK(n9156), .Q(
        g3223) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n8745), .CLK(n9160), .Q(
        g2970), .QN(n8455) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n8667), .CLK(n9082), .Q(
        g5698), .QN(n8303) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n8712), .CLK(n9127), .Q(
        g5260) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n8712), .CLK(n9127), .Q(
        g1521) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n8716), .CLK(n9131), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n8669), .CLK(n9084), .Q(
        g3115) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n8703), .CLK(n9118), .Q(
        g3251) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n8706), .CLK(n9121), .Q(
        g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n8706), .CLK(n9121), 
        .Q(test_so99), .QN(n8600) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n8693), .CLK(n9108), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n8733), .CLK(n9148), .Q(
        g8342), .QN(n8074) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n8686), .CLK(n9101), .Q(
        g4515), .QN(n8437) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n8704), .CLK(n9119), .Q(
        g8787) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n8655), .CLK(n9070), .Q(
        g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n8647), .CLK(n9062), .Q(
        n9236), .QN(n15228) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n8647), .CLK(n9062), .Q(
        g1379), .QN(n8516) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n8732), .CLK(n9147), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n8696), .CLK(n9111), 
        .Q(g1878) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n8733), .CLK(n9148), .Q(
        g5619), .QN(n8197) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n8673), .CLK(n9088), .Q(
        g71) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n8673), .CLK(n9088), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1415), .SI(g4704), .SE(n8714), .CLK(n9129), .Q(
        g22), .QN(n8154) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n8723), .CLK(n9138), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n8686), .CLK(n9101), .Q(
        g2729), .QN(n8186) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n8640), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n8639), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n8640), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n8639), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n8640), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n8639), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n8640), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n8639), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n8640), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n8639), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n8640), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n8639), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n8640), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n8639), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n8640), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n8639), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n8640), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n8639), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n8640), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n8639), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n8640), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n8639), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n58), .QN(
        n87) );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n59), .QN(
        n37) );
  NAND3X0 Trojan_U17 ( .IN1(n2601), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n53), .IN3(n8568), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U8562 ( .INP(n87), .ZN(n8638) );
  INVX0 U8563 ( .INP(n8638), .ZN(n8639) );
  INVX0 U8564 ( .INP(n8638), .ZN(n8640) );
  NBUFFX2 U8565 ( .INP(n8769), .Z(n8642) );
  NBUFFX2 U8566 ( .INP(n8769), .Z(n8641) );
  NBUFFX2 U8567 ( .INP(n8754), .Z(n8714) );
  NBUFFX2 U8568 ( .INP(n8757), .Z(n8699) );
  NBUFFX2 U8569 ( .INP(n8755), .Z(n8712) );
  NBUFFX2 U8570 ( .INP(n8762), .Z(n8673) );
  NBUFFX2 U8571 ( .INP(n8760), .Z(n8687) );
  NBUFFX2 U8572 ( .INP(n8759), .Z(n8691) );
  NBUFFX2 U8573 ( .INP(n8752), .Z(n8725) );
  NBUFFX2 U8574 ( .INP(n8758), .Z(n8697) );
  NBUFFX2 U8575 ( .INP(n8750), .Z(n8734) );
  NBUFFX2 U8576 ( .INP(n8751), .Z(n8732) );
  NBUFFX2 U8577 ( .INP(n8759), .Z(n8689) );
  NBUFFX2 U8578 ( .INP(n8757), .Z(n8701) );
  NBUFFX2 U8579 ( .INP(n8761), .Z(n8680) );
  NBUFFX2 U8580 ( .INP(n8763), .Z(n8671) );
  NBUFFX2 U8581 ( .INP(n8749), .Z(n8742) );
  NBUFFX2 U8582 ( .INP(n8764), .Z(n8664) );
  NBUFFX2 U8583 ( .INP(n8768), .Z(n8643) );
  NBUFFX2 U8584 ( .INP(n8765), .Z(n8658) );
  NBUFFX2 U8585 ( .INP(n8766), .Z(n8657) );
  NBUFFX2 U8586 ( .INP(n8763), .Z(n8672) );
  NBUFFX2 U8587 ( .INP(n8768), .Z(n8644) );
  NBUFFX2 U8588 ( .INP(n8761), .Z(n8682) );
  NBUFFX2 U8589 ( .INP(n8758), .Z(n8693) );
  NBUFFX2 U8590 ( .INP(n8766), .Z(n8654) );
  NBUFFX2 U8591 ( .INP(n8767), .Z(n8648) );
  NBUFFX2 U8592 ( .INP(n8756), .Z(n8706) );
  NBUFFX2 U8593 ( .INP(n8759), .Z(n8692) );
  NBUFFX2 U8594 ( .INP(n8756), .Z(n8704) );
  NBUFFX2 U8595 ( .INP(n8750), .Z(n8737) );
  NBUFFX2 U8596 ( .INP(n8765), .Z(n8659) );
  NBUFFX2 U8597 ( .INP(n8759), .Z(n8690) );
  NBUFFX2 U8598 ( .INP(n8755), .Z(n8709) );
  NBUFFX2 U8599 ( .INP(n8765), .Z(n8662) );
  NBUFFX2 U8600 ( .INP(n8763), .Z(n8669) );
  NBUFFX2 U8601 ( .INP(n8749), .Z(n8739) );
  NBUFFX2 U8602 ( .INP(n8749), .Z(n8741) );
  NBUFFX2 U8603 ( .INP(n8755), .Z(n8710) );
  NBUFFX2 U8604 ( .INP(n8754), .Z(n8717) );
  NBUFFX2 U8605 ( .INP(n8764), .Z(n8665) );
  NBUFFX2 U8606 ( .INP(n8761), .Z(n8678) );
  NBUFFX2 U8607 ( .INP(n8752), .Z(n8723) );
  NBUFFX2 U8608 ( .INP(n8750), .Z(n8736) );
  NBUFFX2 U8609 ( .INP(n8753), .Z(n8722) );
  NBUFFX2 U8610 ( .INP(n8753), .Z(n8721) );
  NBUFFX2 U8611 ( .INP(n8753), .Z(n8719) );
  NBUFFX2 U8612 ( .INP(n8754), .Z(n8713) );
  NBUFFX2 U8613 ( .INP(n8763), .Z(n8668) );
  NBUFFX2 U8614 ( .INP(n8767), .Z(n8652) );
  NBUFFX2 U8615 ( .INP(n8750), .Z(n8735) );
  NBUFFX2 U8616 ( .INP(n8765), .Z(n8661) );
  NBUFFX2 U8617 ( .INP(n8765), .Z(n8660) );
  NBUFFX2 U8618 ( .INP(n8764), .Z(n8663) );
  NBUFFX2 U8619 ( .INP(n8760), .Z(n8684) );
  NBUFFX2 U8620 ( .INP(n8757), .Z(n8698) );
  NBUFFX2 U8621 ( .INP(n8749), .Z(n8740) );
  NBUFFX2 U8622 ( .INP(n8757), .Z(n8700) );
  NBUFFX2 U8623 ( .INP(n8766), .Z(n8656) );
  NBUFFX2 U8624 ( .INP(n8757), .Z(n8702) );
  NBUFFX2 U8625 ( .INP(n8752), .Z(n8726) );
  NBUFFX2 U8626 ( .INP(n8767), .Z(n8649) );
  NBUFFX2 U8627 ( .INP(n8752), .Z(n8724) );
  NBUFFX2 U8628 ( .INP(n8760), .Z(n8683) );
  NBUFFX2 U8629 ( .INP(n8762), .Z(n8677) );
  NBUFFX2 U8630 ( .INP(n8753), .Z(n8718) );
  NBUFFX2 U8631 ( .INP(n8761), .Z(n8679) );
  NBUFFX2 U8632 ( .INP(n8754), .Z(n8715) );
  NBUFFX2 U8633 ( .INP(n8764), .Z(n8667) );
  NBUFFX2 U8634 ( .INP(n8768), .Z(n8646) );
  NBUFFX2 U8635 ( .INP(n8768), .Z(n8645) );
  NBUFFX2 U8636 ( .INP(n8756), .Z(n8705) );
  NBUFFX2 U8637 ( .INP(n8758), .Z(n8694) );
  NBUFFX2 U8638 ( .INP(n8750), .Z(n8733) );
  NBUFFX2 U8639 ( .INP(n8755), .Z(n8708) );
  NBUFFX2 U8640 ( .INP(n8763), .Z(n8670) );
  NBUFFX2 U8641 ( .INP(n8751), .Z(n8728) );
  NBUFFX2 U8642 ( .INP(n8768), .Z(n8647) );
  NBUFFX2 U8643 ( .INP(n8756), .Z(n8703) );
  NBUFFX2 U8644 ( .INP(n8749), .Z(n8738) );
  NBUFFX2 U8645 ( .INP(n8759), .Z(n8688) );
  NBUFFX2 U8646 ( .INP(n8754), .Z(n8716) );
  NBUFFX2 U8647 ( .INP(n8762), .Z(n8675) );
  NBUFFX2 U8648 ( .INP(n8760), .Z(n8686) );
  NBUFFX2 U8649 ( .INP(n8760), .Z(n8685) );
  NBUFFX2 U8650 ( .INP(n8756), .Z(n8707) );
  NBUFFX2 U8651 ( .INP(n8762), .Z(n8676) );
  NBUFFX2 U8652 ( .INP(n8751), .Z(n8731) );
  NBUFFX2 U8653 ( .INP(n8764), .Z(n8666) );
  NBUFFX2 U8654 ( .INP(n8751), .Z(n8729) );
  NBUFFX2 U8655 ( .INP(n8767), .Z(n8650) );
  NBUFFX2 U8656 ( .INP(n8761), .Z(n8681) );
  NBUFFX2 U8657 ( .INP(n8752), .Z(n8727) );
  NBUFFX2 U8658 ( .INP(n8766), .Z(n8655) );
  NBUFFX2 U8659 ( .INP(n8753), .Z(n8720) );
  NBUFFX2 U8660 ( .INP(n8766), .Z(n8653) );
  NBUFFX2 U8661 ( .INP(n8758), .Z(n8695) );
  NBUFFX2 U8662 ( .INP(n8751), .Z(n8730) );
  NBUFFX2 U8663 ( .INP(n8762), .Z(n8674) );
  NBUFFX2 U8664 ( .INP(n8755), .Z(n8711) );
  NBUFFX2 U8665 ( .INP(n8758), .Z(n8696) );
  NBUFFX2 U8666 ( .INP(n8767), .Z(n8651) );
  NBUFFX2 U8667 ( .INP(n9184), .Z(n9057) );
  NBUFFX2 U8668 ( .INP(n9184), .Z(n9056) );
  NBUFFX2 U8669 ( .INP(n9169), .Z(n9129) );
  NBUFFX2 U8670 ( .INP(n9172), .Z(n9114) );
  NBUFFX2 U8671 ( .INP(n9170), .Z(n9127) );
  NBUFFX2 U8672 ( .INP(n9177), .Z(n9088) );
  NBUFFX2 U8673 ( .INP(n9175), .Z(n9102) );
  NBUFFX2 U8674 ( .INP(n9174), .Z(n9106) );
  NBUFFX2 U8675 ( .INP(n9167), .Z(n9140) );
  NBUFFX2 U8676 ( .INP(n9173), .Z(n9112) );
  NBUFFX2 U8677 ( .INP(n9165), .Z(n9149) );
  NBUFFX2 U8678 ( .INP(n9166), .Z(n9147) );
  NBUFFX2 U8679 ( .INP(n9174), .Z(n9104) );
  NBUFFX2 U8680 ( .INP(n9172), .Z(n9116) );
  NBUFFX2 U8681 ( .INP(n9176), .Z(n9095) );
  NBUFFX2 U8682 ( .INP(n9178), .Z(n9086) );
  NBUFFX2 U8683 ( .INP(n9164), .Z(n9157) );
  NBUFFX2 U8684 ( .INP(n9179), .Z(n9079) );
  NBUFFX2 U8685 ( .INP(n9183), .Z(n9058) );
  NBUFFX2 U8686 ( .INP(n9180), .Z(n9073) );
  NBUFFX2 U8687 ( .INP(n9181), .Z(n9072) );
  NBUFFX2 U8688 ( .INP(n9178), .Z(n9087) );
  NBUFFX2 U8689 ( .INP(n9183), .Z(n9059) );
  NBUFFX2 U8690 ( .INP(n9176), .Z(n9097) );
  NBUFFX2 U8691 ( .INP(n9173), .Z(n9108) );
  NBUFFX2 U8692 ( .INP(n9181), .Z(n9069) );
  NBUFFX2 U8693 ( .INP(n9182), .Z(n9063) );
  NBUFFX2 U8694 ( .INP(n9171), .Z(n9121) );
  NBUFFX2 U8695 ( .INP(n9174), .Z(n9107) );
  NBUFFX2 U8696 ( .INP(n9171), .Z(n9119) );
  NBUFFX2 U8697 ( .INP(n9165), .Z(n9152) );
  NBUFFX2 U8698 ( .INP(n9180), .Z(n9074) );
  NBUFFX2 U8699 ( .INP(n9174), .Z(n9105) );
  NBUFFX2 U8700 ( .INP(n9170), .Z(n9124) );
  NBUFFX2 U8701 ( .INP(n9180), .Z(n9077) );
  NBUFFX2 U8702 ( .INP(n9178), .Z(n9084) );
  NBUFFX2 U8703 ( .INP(n9164), .Z(n9154) );
  NBUFFX2 U8704 ( .INP(n9164), .Z(n9156) );
  NBUFFX2 U8705 ( .INP(n9170), .Z(n9125) );
  NBUFFX2 U8706 ( .INP(n9169), .Z(n9132) );
  NBUFFX2 U8707 ( .INP(n9179), .Z(n9080) );
  NBUFFX2 U8708 ( .INP(n9176), .Z(n9093) );
  NBUFFX2 U8709 ( .INP(n9167), .Z(n9138) );
  NBUFFX2 U8710 ( .INP(n9165), .Z(n9151) );
  NBUFFX2 U8711 ( .INP(n9168), .Z(n9137) );
  NBUFFX2 U8712 ( .INP(n9168), .Z(n9136) );
  NBUFFX2 U8713 ( .INP(n9168), .Z(n9134) );
  NBUFFX2 U8714 ( .INP(n9169), .Z(n9128) );
  NBUFFX2 U8715 ( .INP(n9178), .Z(n9083) );
  NBUFFX2 U8716 ( .INP(n9182), .Z(n9067) );
  NBUFFX2 U8717 ( .INP(n9165), .Z(n9150) );
  NBUFFX2 U8718 ( .INP(n9180), .Z(n9076) );
  NBUFFX2 U8719 ( .INP(n9180), .Z(n9075) );
  NBUFFX2 U8720 ( .INP(n9179), .Z(n9078) );
  NBUFFX2 U8721 ( .INP(n9175), .Z(n9099) );
  NBUFFX2 U8722 ( .INP(n9172), .Z(n9113) );
  NBUFFX2 U8723 ( .INP(n9164), .Z(n9155) );
  NBUFFX2 U8724 ( .INP(n9172), .Z(n9115) );
  NBUFFX2 U8725 ( .INP(n9181), .Z(n9071) );
  NBUFFX2 U8726 ( .INP(n9172), .Z(n9117) );
  NBUFFX2 U8727 ( .INP(n9167), .Z(n9141) );
  NBUFFX2 U8728 ( .INP(n9182), .Z(n9064) );
  NBUFFX2 U8729 ( .INP(n9167), .Z(n9139) );
  NBUFFX2 U8730 ( .INP(n9175), .Z(n9098) );
  NBUFFX2 U8731 ( .INP(n9177), .Z(n9092) );
  NBUFFX2 U8732 ( .INP(n9168), .Z(n9133) );
  NBUFFX2 U8733 ( .INP(n9176), .Z(n9094) );
  NBUFFX2 U8734 ( .INP(n9169), .Z(n9130) );
  NBUFFX2 U8735 ( .INP(n9179), .Z(n9082) );
  NBUFFX2 U8736 ( .INP(n9183), .Z(n9061) );
  NBUFFX2 U8737 ( .INP(n9183), .Z(n9060) );
  NBUFFX2 U8738 ( .INP(n9171), .Z(n9120) );
  NBUFFX2 U8739 ( .INP(n9173), .Z(n9109) );
  NBUFFX2 U8740 ( .INP(n9165), .Z(n9148) );
  NBUFFX2 U8741 ( .INP(n9170), .Z(n9123) );
  NBUFFX2 U8742 ( .INP(n9178), .Z(n9085) );
  NBUFFX2 U8743 ( .INP(n9166), .Z(n9143) );
  NBUFFX2 U8744 ( .INP(n9183), .Z(n9062) );
  NBUFFX2 U8745 ( .INP(n9171), .Z(n9118) );
  NBUFFX2 U8746 ( .INP(n9164), .Z(n9153) );
  NBUFFX2 U8747 ( .INP(n9174), .Z(n9103) );
  NBUFFX2 U8748 ( .INP(n9169), .Z(n9131) );
  NBUFFX2 U8749 ( .INP(n9177), .Z(n9090) );
  NBUFFX2 U8750 ( .INP(n9175), .Z(n9101) );
  NBUFFX2 U8751 ( .INP(n9175), .Z(n9100) );
  NBUFFX2 U8752 ( .INP(n9171), .Z(n9122) );
  NBUFFX2 U8753 ( .INP(n9177), .Z(n9091) );
  NBUFFX2 U8754 ( .INP(n9166), .Z(n9146) );
  NBUFFX2 U8755 ( .INP(n9179), .Z(n9081) );
  NBUFFX2 U8756 ( .INP(n9166), .Z(n9144) );
  NBUFFX2 U8757 ( .INP(n9182), .Z(n9065) );
  NBUFFX2 U8758 ( .INP(n9176), .Z(n9096) );
  NBUFFX2 U8759 ( .INP(n9167), .Z(n9142) );
  NBUFFX2 U8760 ( .INP(n9181), .Z(n9070) );
  NBUFFX2 U8761 ( .INP(n9168), .Z(n9135) );
  NBUFFX2 U8762 ( .INP(n9181), .Z(n9068) );
  NBUFFX2 U8763 ( .INP(n9173), .Z(n9110) );
  NBUFFX2 U8764 ( .INP(n9166), .Z(n9145) );
  NBUFFX2 U8765 ( .INP(n9177), .Z(n9089) );
  NBUFFX2 U8766 ( .INP(n9170), .Z(n9126) );
  NBUFFX2 U8767 ( .INP(n9173), .Z(n9111) );
  NBUFFX2 U8768 ( .INP(n9182), .Z(n9066) );
  INVX0 U8769 ( .INP(n8782), .ZN(n8926) );
  INVX0 U8770 ( .INP(n8794), .ZN(n8948) );
  INVX0 U8771 ( .INP(n8797), .ZN(n8955) );
  INVX0 U8772 ( .INP(n8798), .ZN(n8956) );
  INVX0 U8773 ( .INP(n8795), .ZN(n8950) );
  INVX0 U8774 ( .INP(n8797), .ZN(n8954) );
  INVX0 U8775 ( .INP(n8795), .ZN(n8951) );
  INVX0 U8776 ( .INP(n8794), .ZN(n8949) );
  INVX0 U8777 ( .INP(n8796), .ZN(n8953) );
  INVX0 U8778 ( .INP(n8796), .ZN(n8952) );
  INVX0 U8779 ( .INP(n8800), .ZN(n8960) );
  INVX0 U8780 ( .INP(n8801), .ZN(n8962) );
  INVX0 U8781 ( .INP(n8802), .ZN(n8965) );
  INVX0 U8782 ( .INP(n8802), .ZN(n8964) );
  INVX0 U8783 ( .INP(n8801), .ZN(n8963) );
  INVX0 U8784 ( .INP(n8799), .ZN(n8958) );
  INVX0 U8785 ( .INP(n8799), .ZN(n8959) );
  INVX0 U8786 ( .INP(n8800), .ZN(n8961) );
  INVX0 U8787 ( .INP(n8846), .ZN(n9051) );
  INVX0 U8788 ( .INP(n8847), .ZN(n9053) );
  INVX0 U8789 ( .INP(n8847), .ZN(n9054) );
  INVX0 U8790 ( .INP(n8848), .ZN(n9055) );
  INVX0 U8791 ( .INP(n8846), .ZN(n9052) );
  INVX0 U8792 ( .INP(n8803), .ZN(n8966) );
  INVX0 U8793 ( .INP(n8792), .ZN(n8945) );
  INVX0 U8794 ( .INP(n8793), .ZN(n8947) );
  INVX0 U8795 ( .INP(n8793), .ZN(n8946) );
  INVX0 U8796 ( .INP(n8792), .ZN(n8944) );
  INVX0 U8797 ( .INP(n8782), .ZN(n8927) );
  INVX0 U8798 ( .INP(n8798), .ZN(n8957) );
  INVX0 U8799 ( .INP(n8781), .ZN(n8925) );
  INVX0 U8800 ( .INP(n8837), .ZN(n9033) );
  INVX0 U8801 ( .INP(n8818), .ZN(n8996) );
  INVX0 U8802 ( .INP(n8813), .ZN(n8986) );
  INVX0 U8803 ( .INP(n8825), .ZN(n9010) );
  INVX0 U8804 ( .INP(n8831), .ZN(n9021) );
  INVX0 U8805 ( .INP(n8824), .ZN(n9008) );
  INVX0 U8806 ( .INP(n8811), .ZN(n8982) );
  INVX0 U8807 ( .INP(n8816), .ZN(n8992) );
  INVX0 U8808 ( .INP(n8843), .ZN(n9046) );
  INVX0 U8809 ( .INP(n8814), .ZN(n8987) );
  INVX0 U8810 ( .INP(n8815), .ZN(n8990) );
  INVX0 U8811 ( .INP(n8839), .ZN(n9038) );
  INVX0 U8812 ( .INP(n8842), .ZN(n9044) );
  INVX0 U8813 ( .INP(n8806), .ZN(n8973) );
  INVX0 U8814 ( .INP(n8829), .ZN(n9018) );
  INVX0 U8815 ( .INP(n8808), .ZN(n8977) );
  INVX0 U8816 ( .INP(n8840), .ZN(n9039) );
  INVX0 U8817 ( .INP(n8824), .ZN(n9007) );
  INVX0 U8818 ( .INP(n8817), .ZN(n8993) );
  INVX0 U8819 ( .INP(n8815), .ZN(n8989) );
  INVX0 U8820 ( .INP(n8805), .ZN(n8970) );
  INVX0 U8821 ( .INP(n8825), .ZN(n9009) );
  INVX0 U8822 ( .INP(n8813), .ZN(n8985) );
  INVX0 U8823 ( .INP(n8821), .ZN(n9002) );
  INVX0 U8824 ( .INP(n8810), .ZN(n8981) );
  INVX0 U8825 ( .INP(n8827), .ZN(n9014) );
  INVX0 U8826 ( .INP(n8834), .ZN(n9028) );
  INVX0 U8827 ( .INP(n8803), .ZN(n8967) );
  INVX0 U8828 ( .INP(n8829), .ZN(n9017) );
  INVX0 U8829 ( .INP(n8838), .ZN(n9035) );
  INVX0 U8830 ( .INP(n8819), .ZN(n8997) );
  INVX0 U8831 ( .INP(n8841), .ZN(n9042) );
  INVX0 U8832 ( .INP(n8842), .ZN(n9043) );
  INVX0 U8833 ( .INP(n8844), .ZN(n9047) );
  INVX0 U8834 ( .INP(n8816), .ZN(n8991) );
  INVX0 U8835 ( .INP(n8828), .ZN(n9016) );
  INVX0 U8836 ( .INP(n8817), .ZN(n8994) );
  INVX0 U8837 ( .INP(n8828), .ZN(n9015) );
  INVX0 U8838 ( .INP(n8823), .ZN(n9006) );
  INVX0 U8839 ( .INP(n8833), .ZN(n9026) );
  INVX0 U8840 ( .INP(n8805), .ZN(n8971) );
  INVX0 U8841 ( .INP(n8808), .ZN(n8976) );
  INVX0 U8842 ( .INP(n8807), .ZN(n8974) );
  INVX0 U8843 ( .INP(n8835), .ZN(n9029) );
  INVX0 U8844 ( .INP(n8827), .ZN(n9013) );
  INVX0 U8845 ( .INP(n8837), .ZN(n9034) );
  INVX0 U8846 ( .INP(n8839), .ZN(n9037) );
  INVX0 U8847 ( .INP(n8806), .ZN(n8972) );
  INVX0 U8848 ( .INP(n8832), .ZN(n9024) );
  INVX0 U8849 ( .INP(n8814), .ZN(n8988) );
  INVX0 U8850 ( .INP(n8843), .ZN(n9045) );
  INVX0 U8851 ( .INP(n8818), .ZN(n8995) );
  INVX0 U8852 ( .INP(n8807), .ZN(n8975) );
  INVX0 U8853 ( .INP(n8841), .ZN(n9041) );
  INVX0 U8854 ( .INP(n8830), .ZN(n9020) );
  INVX0 U8855 ( .INP(n8812), .ZN(n8984) );
  INVX0 U8856 ( .INP(n8821), .ZN(n9001) );
  INVX0 U8857 ( .INP(n8831), .ZN(n9022) );
  INVX0 U8858 ( .INP(n8820), .ZN(n8999) );
  INVX0 U8859 ( .INP(n8838), .ZN(n9036) );
  INVX0 U8860 ( .INP(n8804), .ZN(n8969) );
  INVX0 U8861 ( .INP(n8836), .ZN(n9031) );
  INVX0 U8862 ( .INP(n8844), .ZN(n9048) );
  INVX0 U8863 ( .INP(n8835), .ZN(n9030) );
  INVX0 U8864 ( .INP(n8833), .ZN(n9025) );
  INVX0 U8865 ( .INP(n8819), .ZN(n8998) );
  INVX0 U8866 ( .INP(n8811), .ZN(n8983) );
  INVX0 U8867 ( .INP(n8809), .ZN(n8979) );
  INVX0 U8868 ( .INP(n8804), .ZN(n8968) );
  INVX0 U8869 ( .INP(n8823), .ZN(n9005) );
  INVX0 U8870 ( .INP(n8840), .ZN(n9040) );
  INVX0 U8871 ( .INP(n8845), .ZN(n9049) );
  INVX0 U8872 ( .INP(n8826), .ZN(n9012) );
  INVX0 U8873 ( .INP(n8826), .ZN(n9011) );
  INVX0 U8874 ( .INP(n8836), .ZN(n9032) );
  INVX0 U8875 ( .INP(n8822), .ZN(n9004) );
  INVX0 U8876 ( .INP(n8830), .ZN(n9019) );
  INVX0 U8877 ( .INP(n8834), .ZN(n9027) );
  INVX0 U8878 ( .INP(n8809), .ZN(n8978) );
  INVX0 U8879 ( .INP(n8810), .ZN(n8980) );
  INVX0 U8880 ( .INP(n8820), .ZN(n9000) );
  INVX0 U8881 ( .INP(n8822), .ZN(n9003) );
  INVX0 U8882 ( .INP(n8832), .ZN(n9023) );
  INVX0 U8883 ( .INP(n8845), .ZN(n9050) );
  INVX0 U8884 ( .INP(n8781), .ZN(n8924) );
  INVX0 U8885 ( .INP(n8788), .ZN(n8936) );
  INVX0 U8886 ( .INP(n8790), .ZN(n8941) );
  INVX0 U8887 ( .INP(n8791), .ZN(n8943) );
  INVX0 U8888 ( .INP(n8786), .ZN(n8932) );
  INVX0 U8889 ( .INP(n8789), .ZN(n8938) );
  INVX0 U8890 ( .INP(n8785), .ZN(n8931) );
  INVX0 U8891 ( .INP(n8786), .ZN(n8933) );
  INVX0 U8892 ( .INP(n8790), .ZN(n8940) );
  INVX0 U8893 ( .INP(n8791), .ZN(n8942) );
  INVX0 U8894 ( .INP(n8787), .ZN(n8935) );
  INVX0 U8895 ( .INP(n8789), .ZN(n8939) );
  INVX0 U8896 ( .INP(n8788), .ZN(n8937) );
  INVX0 U8897 ( .INP(n8787), .ZN(n8934) );
  INVX0 U8898 ( .INP(n8783), .ZN(n8928) );
  INVX0 U8899 ( .INP(n8783), .ZN(n8929) );
  INVX0 U8900 ( .INP(n8784), .ZN(n8930) );
  NBUFFX2 U8901 ( .INP(n8748), .Z(n8746) );
  NBUFFX2 U8902 ( .INP(n8748), .Z(n8744) );
  NBUFFX2 U8903 ( .INP(n8748), .Z(n8745) );
  NBUFFX2 U8904 ( .INP(n8748), .Z(n8743) );
  NBUFFX2 U8905 ( .INP(n9163), .Z(n9161) );
  NBUFFX2 U8906 ( .INP(n9163), .Z(n9159) );
  NBUFFX2 U8907 ( .INP(n9163), .Z(n9160) );
  NBUFFX2 U8908 ( .INP(n9163), .Z(n9158) );
  NBUFFX2 U8909 ( .INP(n8748), .Z(n8747) );
  NBUFFX2 U8910 ( .INP(n8863), .Z(n8783) );
  NBUFFX2 U8911 ( .INP(n8863), .Z(n8781) );
  NBUFFX2 U8912 ( .INP(n8863), .Z(n8782) );
  NBUFFX2 U8913 ( .INP(n8863), .Z(n8784) );
  NBUFFX2 U8914 ( .INP(n8862), .Z(n8788) );
  NBUFFX2 U8915 ( .INP(n8860), .Z(n8794) );
  NBUFFX2 U8916 ( .INP(n8861), .Z(n8790) );
  NBUFFX2 U8917 ( .INP(n8861), .Z(n8791) );
  NBUFFX2 U8918 ( .INP(n8862), .Z(n8786) );
  NBUFFX2 U8919 ( .INP(n8862), .Z(n8785) );
  NBUFFX2 U8920 ( .INP(n8861), .Z(n8792) );
  NBUFFX2 U8921 ( .INP(n8860), .Z(n8797) );
  NBUFFX2 U8922 ( .INP(n8861), .Z(n8789) );
  NBUFFX2 U8923 ( .INP(n8861), .Z(n8793) );
  NBUFFX2 U8924 ( .INP(n8859), .Z(n8800) );
  NBUFFX2 U8925 ( .INP(n8860), .Z(n8798) );
  NBUFFX2 U8926 ( .INP(n8859), .Z(n8801) );
  NBUFFX2 U8927 ( .INP(n8862), .Z(n8787) );
  NBUFFX2 U8928 ( .INP(n8859), .Z(n8802) );
  NBUFFX2 U8929 ( .INP(n8860), .Z(n8795) );
  NBUFFX2 U8930 ( .INP(n8853), .Z(n8824) );
  NBUFFX2 U8931 ( .INP(n8855), .Z(n8815) );
  NBUFFX2 U8932 ( .INP(n8853), .Z(n8825) );
  NBUFFX2 U8933 ( .INP(n8856), .Z(n8813) );
  NBUFFX2 U8934 ( .INP(n8859), .Z(n8799) );
  NBUFFX2 U8935 ( .INP(n8859), .Z(n8803) );
  NBUFFX2 U8936 ( .INP(n8852), .Z(n8829) );
  NBUFFX2 U8937 ( .INP(n8850), .Z(n8842) );
  NBUFFX2 U8938 ( .INP(n8855), .Z(n8816) );
  NBUFFX2 U8939 ( .INP(n8849), .Z(n8847) );
  NBUFFX2 U8940 ( .INP(n8855), .Z(n8817) );
  NBUFFX2 U8941 ( .INP(n8853), .Z(n8828) );
  NBUFFX2 U8942 ( .INP(n8858), .Z(n8805) );
  NBUFFX2 U8943 ( .INP(n8849), .Z(n8848) );
  NBUFFX2 U8944 ( .INP(n8858), .Z(n8808) );
  NBUFFX2 U8945 ( .INP(n8853), .Z(n8827) );
  NBUFFX2 U8946 ( .INP(n8851), .Z(n8837) );
  NBUFFX2 U8947 ( .INP(n8850), .Z(n8839) );
  NBUFFX2 U8948 ( .INP(n8858), .Z(n8806) );
  NBUFFX2 U8949 ( .INP(n8856), .Z(n8814) );
  NBUFFX2 U8950 ( .INP(n8850), .Z(n8843) );
  NBUFFX2 U8951 ( .INP(n8855), .Z(n8818) );
  NBUFFX2 U8952 ( .INP(n8858), .Z(n8807) );
  NBUFFX2 U8953 ( .INP(n8850), .Z(n8841) );
  NBUFFX2 U8954 ( .INP(n8856), .Z(n8812) );
  NBUFFX2 U8955 ( .INP(n8854), .Z(n8821) );
  NBUFFX2 U8956 ( .INP(n8852), .Z(n8831) );
  NBUFFX2 U8957 ( .INP(n8851), .Z(n8838) );
  NBUFFX2 U8958 ( .INP(n8849), .Z(n8844) );
  NBUFFX2 U8959 ( .INP(n8851), .Z(n8835) );
  NBUFFX2 U8960 ( .INP(n8852), .Z(n8833) );
  NBUFFX2 U8961 ( .INP(n8855), .Z(n8819) );
  NBUFFX2 U8962 ( .INP(n8857), .Z(n8811) );
  NBUFFX2 U8963 ( .INP(n8849), .Z(n8846) );
  NBUFFX2 U8964 ( .INP(n8858), .Z(n8804) );
  NBUFFX2 U8965 ( .INP(n8854), .Z(n8823) );
  NBUFFX2 U8966 ( .INP(n8850), .Z(n8840) );
  NBUFFX2 U8967 ( .INP(n8853), .Z(n8826) );
  NBUFFX2 U8968 ( .INP(n8851), .Z(n8836) );
  NBUFFX2 U8969 ( .INP(n8852), .Z(n8830) );
  NBUFFX2 U8970 ( .INP(n8851), .Z(n8834) );
  NBUFFX2 U8971 ( .INP(n8857), .Z(n8809) );
  NBUFFX2 U8972 ( .INP(n8857), .Z(n8810) );
  NBUFFX2 U8973 ( .INP(n8854), .Z(n8820) );
  NBUFFX2 U8976 ( .INP(n8854), .Z(n8822) );
  NBUFFX2 U8977 ( .INP(n8852), .Z(n8832) );
  NBUFFX2 U8978 ( .INP(n8849), .Z(n8845) );
  NBUFFX2 U8979 ( .INP(n8860), .Z(n8796) );
  NBUFFX2 U8980 ( .INP(n9163), .Z(n9162) );
  NBUFFX2 U8981 ( .INP(n8777), .Z(n8748) );
  NBUFFX2 U8982 ( .INP(n8776), .Z(n8749) );
  NBUFFX2 U8983 ( .INP(n8776), .Z(n8750) );
  NBUFFX2 U8984 ( .INP(n8776), .Z(n8751) );
  NBUFFX2 U8985 ( .INP(n8775), .Z(n8752) );
  NBUFFX2 U8986 ( .INP(n8775), .Z(n8753) );
  NBUFFX2 U8987 ( .INP(n8775), .Z(n8754) );
  NBUFFX2 U8988 ( .INP(n8774), .Z(n8755) );
  NBUFFX2 U8989 ( .INP(n8774), .Z(n8756) );
  NBUFFX2 U8990 ( .INP(n8774), .Z(n8757) );
  NBUFFX2 U8991 ( .INP(n8773), .Z(n8758) );
  NBUFFX2 U8992 ( .INP(n8773), .Z(n8759) );
  NBUFFX2 U8993 ( .INP(n8773), .Z(n8760) );
  NBUFFX2 U8994 ( .INP(n8772), .Z(n8761) );
  NBUFFX2 U8995 ( .INP(n8772), .Z(n8762) );
  NBUFFX2 U8996 ( .INP(n8772), .Z(n8763) );
  NBUFFX2 U8997 ( .INP(n8771), .Z(n8764) );
  NBUFFX2 U8998 ( .INP(n8771), .Z(n8765) );
  NBUFFX2 U8999 ( .INP(n8771), .Z(n8766) );
  NBUFFX2 U9000 ( .INP(n8770), .Z(n8767) );
  NBUFFX2 U9001 ( .INP(n8770), .Z(n8768) );
  NBUFFX2 U9002 ( .INP(n8770), .Z(n8769) );
  NBUFFX2 U9003 ( .INP(n8780), .Z(n8770) );
  NBUFFX2 U9004 ( .INP(n8780), .Z(n8771) );
  NBUFFX2 U9005 ( .INP(n8779), .Z(n8772) );
  NBUFFX2 U9006 ( .INP(n8779), .Z(n8773) );
  NBUFFX2 U9007 ( .INP(n8779), .Z(n8774) );
  NBUFFX2 U9008 ( .INP(n8778), .Z(n8775) );
  NBUFFX2 U9009 ( .INP(n8778), .Z(n8776) );
  NBUFFX2 U9010 ( .INP(n8778), .Z(n8777) );
  NBUFFX2 U9011 ( .INP(test_se), .Z(n8778) );
  NBUFFX2 U9012 ( .INP(test_se), .Z(n8779) );
  NBUFFX2 U9013 ( .INP(test_se), .Z(n8780) );
  NBUFFX2 U9014 ( .INP(n8868), .Z(n8849) );
  NBUFFX2 U9015 ( .INP(n8868), .Z(n8850) );
  NBUFFX2 U9016 ( .INP(n8868), .Z(n8851) );
  NBUFFX2 U9017 ( .INP(n8867), .Z(n8852) );
  NBUFFX2 U9018 ( .INP(n8867), .Z(n8853) );
  NBUFFX2 U9019 ( .INP(n8867), .Z(n8854) );
  NBUFFX2 U9020 ( .INP(n8866), .Z(n8855) );
  NBUFFX2 U9021 ( .INP(n8866), .Z(n8856) );
  NBUFFX2 U9022 ( .INP(n8866), .Z(n8857) );
  NBUFFX2 U9023 ( .INP(n8865), .Z(n8858) );
  NBUFFX2 U9024 ( .INP(n8865), .Z(n8859) );
  NBUFFX2 U9025 ( .INP(n8865), .Z(n8860) );
  NBUFFX2 U9026 ( .INP(n8864), .Z(n8861) );
  NBUFFX2 U9027 ( .INP(n8864), .Z(n8862) );
  NBUFFX2 U9028 ( .INP(n8864), .Z(n8863) );
  NBUFFX2 U9029 ( .INP(g35), .Z(n8864) );
  NBUFFX2 U9030 ( .INP(g35), .Z(n8865) );
  NBUFFX2 U9031 ( .INP(g35), .Z(n8866) );
  NBUFFX2 U9032 ( .INP(g35), .Z(n8867) );
  NBUFFX2 U9033 ( .INP(g35), .Z(n8868) );
  INVX0 U9034 ( .INP(n8966), .ZN(n8869) );
  INVX0 U9035 ( .INP(n8966), .ZN(n8870) );
  INVX0 U9036 ( .INP(n8965), .ZN(n8871) );
  INVX0 U9037 ( .INP(n8965), .ZN(n8872) );
  INVX0 U9038 ( .INP(n8963), .ZN(n8873) );
  INVX0 U9039 ( .INP(n8965), .ZN(n8874) );
  INVX0 U9040 ( .INP(n8965), .ZN(n8875) );
  INVX0 U9041 ( .INP(n8962), .ZN(n8876) );
  INVX0 U9042 ( .INP(n8965), .ZN(n8877) );
  INVX0 U9043 ( .INP(n8962), .ZN(n8878) );
  INVX0 U9044 ( .INP(n8965), .ZN(n8879) );
  INVX0 U9045 ( .INP(n8962), .ZN(n8880) );
  INVX0 U9046 ( .INP(n8964), .ZN(n8881) );
  INVX0 U9047 ( .INP(n8964), .ZN(n8882) );
  INVX0 U9048 ( .INP(n8964), .ZN(n8883) );
  INVX0 U9049 ( .INP(n8964), .ZN(n8884) );
  INVX0 U9050 ( .INP(n8961), .ZN(n8885) );
  INVX0 U9051 ( .INP(n8964), .ZN(n8886) );
  INVX0 U9052 ( .INP(n8964), .ZN(n8887) );
  INVX0 U9053 ( .INP(n8961), .ZN(n8888) );
  INVX0 U9054 ( .INP(n8963), .ZN(n8889) );
  INVX0 U9055 ( .INP(n8963), .ZN(n8890) );
  INVX0 U9056 ( .INP(n8963), .ZN(n8891) );
  INVX0 U9057 ( .INP(n8963), .ZN(n8892) );
  INVX0 U9058 ( .INP(n8960), .ZN(n8893) );
  INVX0 U9059 ( .INP(n8963), .ZN(n8894) );
  INVX0 U9060 ( .INP(n8960), .ZN(n8895) );
  INVX0 U9061 ( .INP(n8962), .ZN(n8896) );
  INVX0 U9062 ( .INP(n8962), .ZN(n8897) );
  INVX0 U9063 ( .INP(n8959), .ZN(n8898) );
  INVX0 U9064 ( .INP(n8962), .ZN(n8899) );
  INVX0 U9066 ( .INP(n8959), .ZN(n8900) );
  INVX0 U9067 ( .INP(n8961), .ZN(n8901) );
  INVX0 U9068 ( .INP(n8961), .ZN(n8902) );
  INVX0 U9069 ( .INP(n8958), .ZN(n8903) );
  INVX0 U9071 ( .INP(n8961), .ZN(n8904) );
  INVX0 U9072 ( .INP(n8961), .ZN(n8905) );
  INVX0 U9073 ( .INP(n8958), .ZN(n8906) );
  INVX0 U9074 ( .INP(n8960), .ZN(n8907) );
  INVX0 U9077 ( .INP(n8960), .ZN(n8908) );
  INVX0 U9078 ( .INP(n8960), .ZN(n8909) );
  INVX0 U9079 ( .INP(n8960), .ZN(n8910) );
  INVX0 U9081 ( .INP(n8957), .ZN(n8911) );
  INVX0 U9082 ( .INP(n8959), .ZN(n8912) );
  INVX0 U9083 ( .INP(n8959), .ZN(n8913) );
  INVX0 U9087 ( .INP(n8957), .ZN(n8914) );
  INVX0 U9088 ( .INP(n8959), .ZN(n8915) );
  INVX0 U9089 ( .INP(n8959), .ZN(n8916) );
  INVX0 U9091 ( .INP(n8957), .ZN(n8917) );
  INVX0 U9092 ( .INP(n8958), .ZN(n8918) );
  INVX0 U9093 ( .INP(n8958), .ZN(n8919) );
  INVX0 U9094 ( .INP(n8958), .ZN(n8920) );
  INVX0 U9095 ( .INP(n8958), .ZN(n8921) );
  INVX0 U9096 ( .INP(n8957), .ZN(n8922) );
  INVX0 U9097 ( .INP(n8957), .ZN(n8923) );
  NBUFFX2 U9100 ( .INP(n9192), .Z(n9163) );
  NBUFFX2 U9102 ( .INP(n9191), .Z(n9164) );
  NBUFFX2 U9103 ( .INP(n9191), .Z(n9165) );
  NBUFFX2 U9104 ( .INP(n9191), .Z(n9166) );
  NBUFFX2 U9105 ( .INP(n9190), .Z(n9167) );
  NBUFFX2 U9106 ( .INP(n9190), .Z(n9168) );
  NBUFFX2 U9108 ( .INP(n9190), .Z(n9169) );
  NBUFFX2 U9109 ( .INP(n9189), .Z(n9170) );
  NBUFFX2 U9110 ( .INP(n9189), .Z(n9171) );
  NBUFFX2 U9112 ( .INP(n9189), .Z(n9172) );
  NBUFFX2 U9113 ( .INP(n9188), .Z(n9173) );
  NBUFFX2 U9114 ( .INP(n9188), .Z(n9174) );
  NBUFFX2 U9115 ( .INP(n9188), .Z(n9175) );
  NBUFFX2 U9117 ( .INP(n9187), .Z(n9176) );
  NBUFFX2 U9118 ( .INP(n9187), .Z(n9177) );
  NBUFFX2 U9119 ( .INP(n9187), .Z(n9178) );
  NBUFFX2 U9121 ( .INP(n9186), .Z(n9179) );
  NBUFFX2 U9122 ( .INP(n9186), .Z(n9180) );
  NBUFFX2 U9123 ( .INP(n9186), .Z(n9181) );
  NBUFFX2 U9125 ( .INP(n9185), .Z(n9182) );
  NBUFFX2 U9126 ( .INP(n9185), .Z(n9183) );
  NBUFFX2 U9127 ( .INP(n9185), .Z(n9184) );
  NBUFFX2 U9129 ( .INP(n9195), .Z(n9185) );
  NBUFFX2 U9130 ( .INP(n9195), .Z(n9186) );
  NBUFFX2 U9131 ( .INP(n9194), .Z(n9187) );
  NBUFFX2 U9133 ( .INP(n9194), .Z(n9188) );
  NBUFFX2 U9134 ( .INP(n9194), .Z(n9189) );
  NBUFFX2 U9135 ( .INP(n9193), .Z(n9190) );
  NBUFFX2 U9137 ( .INP(n9193), .Z(n9191) );
  NBUFFX2 U9138 ( .INP(n9193), .Z(n9192) );
  NBUFFX2 U9139 ( .INP(CK), .Z(n9193) );
  NBUFFX2 U9140 ( .INP(CK), .Z(n9194) );
  NBUFFX2 U9141 ( .INP(CK), .Z(n9195) );
  NOR3X0 U9142 ( .IN1(n9196), .IN2(n9197), .IN3(n9198), .QN(n8567) );
  INVX0 U9143 ( .INP(n9199), .ZN(n853) );
  INVX0 U9144 ( .INP(n9200), .ZN(n807) );
  NAND2X0 U9145 ( .IN1(n9201), .IN2(n9202), .QN(n631) );
  NAND2X0 U9146 ( .IN1(n8969), .IN2(g1236), .QN(n9202) );
  NAND4X0 U9147 ( .IN1(n9203), .IN2(n9204), .IN3(n9205), .IN4(n9206), .QN(
        n5961) );
  NAND2X0 U9148 ( .IN1(n9207), .IN2(g5348), .QN(n9206) );
  NAND2X0 U9149 ( .IN1(n8435), .IN2(n9208), .QN(n9205) );
  NAND2X0 U9150 ( .IN1(g31860), .IN2(g5352), .QN(n9204) );
  NAND2X0 U9151 ( .IN1(n8434), .IN2(n9209), .QN(n9203) );
  NAND4X0 U9152 ( .IN1(n9210), .IN2(n9211), .IN3(n9212), .IN4(n9213), .QN(
        n5960) );
  NAND2X0 U9153 ( .IN1(n9214), .IN2(g6732), .QN(n9213) );
  NAND2X0 U9154 ( .IN1(n8433), .IN2(n9215), .QN(n9212) );
  NAND2X0 U9155 ( .IN1(n9216), .IN2(g6736), .QN(n9211) );
  NAND2X0 U9156 ( .IN1(n8432), .IN2(n9217), .QN(n9210) );
  NAND2X0 U9157 ( .IN1(n9218), .IN2(n9219), .QN(n503) );
  NAND2X0 U9158 ( .IN1(n9026), .IN2(g4382), .QN(n9219) );
  INVX0 U9159 ( .INP(n9220), .ZN(n468) );
  NOR2X0 U9160 ( .IN1(n9221), .IN2(g29279), .QN(n9220) );
  NOR2X0 U9161 ( .IN1(n8120), .IN2(n8898), .QN(n9221) );
  NAND2X0 U9162 ( .IN1(n9222), .IN2(g1677), .QN(n4459) );
  NAND2X0 U9163 ( .IN1(n9223), .IN2(g1811), .QN(n4448) );
  NAND2X0 U9164 ( .IN1(test_so53), .IN2(n9224), .QN(n4437) );
  NAND2X0 U9165 ( .IN1(n9225), .IN2(g2236), .QN(n4415) );
  NAND2X0 U9166 ( .IN1(n9226), .IN2(g2370), .QN(n4403) );
  NAND2X0 U9167 ( .IN1(n9227), .IN2(g2504), .QN(n4392) );
  NAND2X0 U9168 ( .IN1(n9228), .IN2(g2638), .QN(n4380) );
  NAND4X0 U9169 ( .IN1(n9229), .IN2(n9230), .IN3(n9231), .IN4(n9232), .QN(
        n4305) );
  NOR2X0 U9170 ( .IN1(n9233), .IN2(n9234), .QN(n9232) );
  NOR2X0 U9171 ( .IN1(n5656), .IN2(g4826), .QN(n9234) );
  NOR2X0 U9172 ( .IN1(n5440), .IN2(g4821), .QN(n9233) );
  NAND2X0 U9173 ( .IN1(g4646), .IN2(g29220), .QN(n9231) );
  NAND4X0 U9174 ( .IN1(n5440), .IN2(n9235), .IN3(n9237), .IN4(n8436), .QN(
        n9230) );
  NOR2X0 U9175 ( .IN1(g4688), .IN2(g4646), .QN(n9237) );
  NAND2X0 U9176 ( .IN1(n9238), .IN2(n9239), .QN(n9235) );
  NAND3X0 U9177 ( .IN1(n9241), .IN2(n9242), .IN3(n9243), .QN(n9238) );
  NAND2X0 U9178 ( .IN1(n9244), .IN2(g4776), .QN(n9243) );
  NAND2X0 U9179 ( .IN1(n5368), .IN2(n9246), .QN(n9244) );
  XOR2X1 U9180 ( .IN1(g34657), .IN2(n9248), .Q(n9246) );
  NAND4X0 U9181 ( .IN1(n9249), .IN2(n9250), .IN3(n9251), .IN4(n9252), .QN(
        n9248) );
  NAND2X0 U9182 ( .IN1(n9253), .IN2(g4732), .QN(n9252) );
  NAND2X0 U9183 ( .IN1(n9254), .IN2(g4717), .QN(n9251) );
  NAND2X0 U9184 ( .IN1(n9256), .IN2(g4727), .QN(n9250) );
  NAND2X0 U9185 ( .IN1(n9257), .IN2(g4722), .QN(n9249) );
  NAND2X0 U9186 ( .IN1(n9258), .IN2(g4793), .QN(n9242) );
  NAND2X0 U9187 ( .IN1(n5368), .IN2(n9259), .QN(n9241) );
  NAND2X0 U9188 ( .IN1(n8595), .IN2(n9260), .QN(n9259) );
  NAND4X0 U9189 ( .IN1(n5707), .IN2(n9261), .IN3(n9263), .IN4(n9264), .QN(
        n9260) );
  NAND2X0 U9190 ( .IN1(n9256), .IN2(n5867), .QN(n9261) );
  NAND2X0 U9191 ( .IN1(g4831), .IN2(g4681), .QN(n9229) );
  NAND4X0 U9192 ( .IN1(n9266), .IN2(n9268), .IN3(n9269), .IN4(n9270), .QN(
        n4283) );
  NOR2X0 U9193 ( .IN1(n9271), .IN2(n9272), .QN(n9270) );
  NOR2X0 U9194 ( .IN1(n5318), .IN2(g3333), .QN(n9272) );
  NOR2X0 U9195 ( .IN1(n5283), .IN2(g4035), .QN(n9271) );
  NAND2X0 U9196 ( .IN1(g4871), .IN2(g3684), .QN(n9269) );
  NAND4X0 U9197 ( .IN1(n5283), .IN2(n9275), .IN3(n9277), .IN4(n5713), .QN(
        n9268) );
  NOR2X0 U9198 ( .IN1(g4864), .IN2(g4871), .QN(n9277) );
  NAND2X0 U9199 ( .IN1(n9278), .IN2(n9279), .QN(n9275) );
  NAND3X0 U9200 ( .IN1(n9282), .IN2(n9283), .IN3(n9284), .QN(n9278) );
  NAND2X0 U9201 ( .IN1(n9285), .IN2(g4966), .QN(n9284) );
  NAND2X0 U9202 ( .IN1(n5367), .IN2(n9286), .QN(n9285) );
  XOR2X1 U9203 ( .IN1(g34649), .IN2(n9287), .Q(n9286) );
  NAND4X0 U9204 ( .IN1(n9288), .IN2(n9289), .IN3(n9290), .IN4(n9291), .QN(
        n9287) );
  NAND2X0 U9205 ( .IN1(n9292), .IN2(g4912), .QN(n9291) );
  NAND2X0 U9206 ( .IN1(n9293), .IN2(g4917), .QN(n9290) );
  NAND2X0 U9207 ( .IN1(n9296), .IN2(g4922), .QN(n9289) );
  NAND2X0 U9208 ( .IN1(n9297), .IN2(g4907), .QN(n9288) );
  NAND2X0 U9209 ( .IN1(n9298), .IN2(g4983), .QN(n9283) );
  NAND2X0 U9210 ( .IN1(n5367), .IN2(n9299), .QN(n9282) );
  NAND2X0 U9211 ( .IN1(n8587), .IN2(n9300), .QN(n9299) );
  NAND4X0 U9212 ( .IN1(n5706), .IN2(n9301), .IN3(n9304), .IN4(n9305), .QN(
        n9300) );
  NAND2X0 U9213 ( .IN1(n9293), .IN2(n5879), .QN(n9301) );
  NAND2X0 U9214 ( .IN1(g4836), .IN2(g5011), .QN(n9266) );
  INVX0 U9215 ( .INP(n9307), .ZN(n424) );
  NOR2X0 U9216 ( .IN1(n9308), .IN2(n9309), .QN(n9307) );
  NOR2X0 U9217 ( .IN1(n8900), .IN2(n8462), .QN(n9309) );
  NOR2X0 U9218 ( .IN1(n9310), .IN2(n8938), .QN(n9308) );
  NOR2X0 U9219 ( .IN1(test_so74), .IN2(test_so14), .QN(n9310) );
  INVX0 U9220 ( .INP(n9311), .ZN(n422) );
  NOR2X0 U9221 ( .IN1(n9313), .IN2(g24212), .QN(n9311) );
  NOR2X0 U9222 ( .IN1(n8551), .IN2(n8898), .QN(n9313) );
  NOR3X0 U9223 ( .IN1(g3161), .IN2(g3155), .IN3(g3167), .QN(n4034) );
  NOR3X0 U9224 ( .IN1(g3512), .IN2(g3506), .IN3(g3518), .QN(n4002) );
  NOR3X0 U9225 ( .IN1(g3863), .IN2(test_so33), .IN3(g3857), .QN(n3969) );
  NOR4X0 U9226 ( .IN1(n8499), .IN2(n1782), .IN3(n9198), .IN4(n9196), .QN(n3933) );
  INVX0 U9227 ( .INP(n9315), .ZN(n9196) );
  INVX0 U9228 ( .INP(n9316), .ZN(n9198) );
  NOR3X0 U9229 ( .IN1(g5176), .IN2(g5164), .IN3(g5170), .QN(n3926) );
  NOR3X0 U9230 ( .IN1(g5523), .IN2(g5511), .IN3(g5517), .QN(n3893) );
  NOR3X0 U9231 ( .IN1(g5863), .IN2(g5857), .IN3(g5869), .QN(n3860) );
  NOR3X0 U9232 ( .IN1(g6209), .IN2(g6203), .IN3(g6215), .QN(n3826) );
  NOR3X0 U9233 ( .IN1(g6561), .IN2(g6549), .IN3(g6555), .QN(n3792) );
  NAND4X0 U9234 ( .IN1(n5358), .IN2(n5520), .IN3(n9317), .IN4(n9318), .QN(
        n3675) );
  NAND2X0 U9235 ( .IN1(n8510), .IN2(n9319), .QN(n9318) );
  NAND2X0 U9236 ( .IN1(n9320), .IN2(n5629), .QN(n9319) );
  XOR2X1 U9237 ( .IN1(g174), .IN2(test_so72), .Q(n9320) );
  NAND2X0 U9238 ( .IN1(n9321), .IN2(g392), .QN(n9317) );
  NAND2X0 U9239 ( .IN1(n9323), .IN2(n8184), .QN(n9321) );
  XOR2X1 U9240 ( .IN1(n8313), .IN2(n8593), .Q(n9323) );
  NAND3X0 U9241 ( .IN1(g2741), .IN2(n5300), .IN3(n5516), .QN(n3635) );
  INVX0 U9242 ( .INP(n9326), .ZN(n335) );
  NAND3X0 U9243 ( .IN1(n9328), .IN2(n8869), .IN3(n9329), .QN(n9326) );
  NOR2X0 U9244 ( .IN1(n9330), .IN2(n9331), .QN(n3174) );
  XOR2X1 U9245 ( .IN1(g482), .IN2(g72), .Q(n9331) );
  XOR2X1 U9246 ( .IN1(g490), .IN2(g73), .Q(n9330) );
  NOR2X0 U9247 ( .IN1(n1782), .IN2(n6010), .QN(n3084) );
  NAND3X0 U9248 ( .IN1(n8897), .IN2(g4104), .IN3(n9333), .QN(n3065) );
  NAND2X0 U9249 ( .IN1(n9334), .IN2(g4108), .QN(n9333) );
  XOR2X1 U9250 ( .IN1(n5323), .IN2(n2607), .Q(n2608) );
  NAND2X0 U9251 ( .IN1(n9335), .IN2(g34979), .QN(n2461) );
  NOR2X0 U9252 ( .IN1(n9337), .IN2(n9338), .QN(n2396) );
  INVX0 U9253 ( .INP(n9339), .ZN(n192) );
  NAND2X0 U9254 ( .IN1(n9341), .IN2(n9342), .QN(n1680) );
  INVX0 U9255 ( .INP(g29277), .ZN(n9342) );
  NAND2X0 U9256 ( .IN1(n9019), .IN2(test_so100), .QN(n9341) );
  INVX0 U9257 ( .INP(n9343), .ZN(n1526) );
  NOR2X0 U9258 ( .IN1(n9344), .IN2(g26953), .QN(n9343) );
  NOR2X0 U9259 ( .IN1(n8179), .IN2(n8898), .QN(n9344) );
  NAND2X0 U9260 ( .IN1(n9345), .IN2(g2079), .QN(n1411) );
  INVX0 U9261 ( .INP(n9346), .ZN(n9345) );
  NAND2X0 U9262 ( .IN1(n9347), .IN2(n9349), .QN(g34980) );
  NAND2X0 U9263 ( .IN1(test_so14), .IN2(n8960), .QN(n9349) );
  NAND2X0 U9264 ( .IN1(n9350), .IN2(n8908), .QN(n9347) );
  NAND2X0 U9265 ( .IN1(n5842), .IN2(n9353), .QN(n9350) );
  NAND4X0 U9266 ( .IN1(n8566), .IN2(n9354), .IN3(n9355), .IN4(n9356), .QN(
        n9353) );
  INVX0 U9267 ( .INP(g54), .ZN(n9355) );
  NAND2X0 U9268 ( .IN1(n9358), .IN2(g22), .QN(g34972) );
  INVX0 U9269 ( .INP(n8566), .ZN(n9358) );
  XOR3X1 U9270 ( .IN1(g34975), .IN2(g34976), .IN3(n9359), .Q(n8566) );
  XOR3X1 U9271 ( .IN1(n9360), .IN2(n9361), .IN3(g34978), .Q(n9359) );
  XOR3X1 U9272 ( .IN1(g34974), .IN2(n9362), .IN3(n9363), .Q(n9361) );
  XOR3X1 U9273 ( .IN1(g34977), .IN2(g34971), .IN3(n9364), .Q(n9360) );
  NAND2X0 U9274 ( .IN1(g55), .IN2(n9365), .QN(n9364) );
  NAND2X0 U9275 ( .IN1(g54), .IN2(n9356), .QN(n9365) );
  NAND2X0 U9276 ( .IN1(n9363), .IN2(g22), .QN(g34927) );
  INVX0 U9277 ( .INP(g34979), .ZN(n9363) );
  NAND4X0 U9278 ( .IN1(n9366), .IN2(n9368), .IN3(n9369), .IN4(n9370), .QN(
        g34979) );
  NOR4X0 U9279 ( .IN1(n9371), .IN2(n9372), .IN3(n9373), .IN4(n9374), .QN(n9370) );
  NOR2X0 U9280 ( .IN1(n5415), .IN2(n9375), .QN(n9374) );
  NOR2X0 U9281 ( .IN1(n5635), .IN2(n9376), .QN(n9373) );
  NOR2X0 U9282 ( .IN1(n5308), .IN2(n9377), .QN(n9372) );
  NOR2X0 U9283 ( .IN1(n9378), .IN2(DFF_420_n1), .QN(n9371) );
  NOR2X0 U9284 ( .IN1(n9379), .IN2(n9380), .QN(n9369) );
  NOR2X0 U9285 ( .IN1(n9381), .IN2(n8624), .QN(n9380) );
  NAND2X0 U9286 ( .IN1(n1415), .IN2(n9382), .QN(n9368) );
  NAND2X0 U9287 ( .IN1(n9383), .IN2(n9384), .QN(n9382) );
  NOR4X0 U9288 ( .IN1(n9385), .IN2(n9386), .IN3(n9387), .IN4(n9388), .QN(n9384) );
  NOR2X0 U9289 ( .IN1(n9389), .IN2(g23612), .QN(n9388) );
  NOR2X0 U9290 ( .IN1(n5293), .IN2(n9390), .QN(n9387) );
  NOR2X0 U9291 ( .IN1(n5470), .IN2(n9391), .QN(n9386) );
  NAND3X0 U9292 ( .IN1(n9392), .IN2(n9393), .IN3(n9394), .QN(n9385) );
  NAND2X0 U9293 ( .IN1(g127), .IN2(n9395), .QN(n9394) );
  NAND2X0 U9294 ( .IN1(test_so14), .IN2(n9335), .QN(n9393) );
  INVX0 U9295 ( .INP(n9338), .ZN(n9335) );
  NAND2X0 U9296 ( .IN1(g92), .IN2(n9396), .QN(n9392) );
  NOR4X0 U9297 ( .IN1(n9397), .IN2(n9398), .IN3(n9399), .IN4(n9400), .QN(n9383) );
  NOR2X0 U9298 ( .IN1(n8455), .IN2(n9401), .QN(n9400) );
  NOR2X0 U9299 ( .IN1(n5981), .IN2(n9402), .QN(n9399) );
  NOR2X0 U9300 ( .IN1(n8462), .IN2(n9403), .QN(n9398) );
  NAND3X0 U9301 ( .IN1(n9404), .IN2(n9405), .IN3(n9406), .QN(n9397) );
  NAND2X0 U9302 ( .IN1(n9407), .IN2(g2975), .QN(n9406) );
  NAND2X0 U9303 ( .IN1(n9408), .IN2(g568), .QN(n9405) );
  NAND2X0 U9304 ( .IN1(n9409), .IN2(g604), .QN(n9404) );
  NAND2X0 U9305 ( .IN1(n9410), .IN2(g2138), .QN(n9366) );
  INVX0 U9306 ( .INP(n9411), .ZN(g34925) );
  NOR2X0 U9307 ( .IN1(g34978), .IN2(n8154), .QN(n9411) );
  NAND4X0 U9308 ( .IN1(n9412), .IN2(n9413), .IN3(n9414), .IN4(n9415), .QN(
        g34978) );
  NOR4X0 U9309 ( .IN1(n9416), .IN2(n9417), .IN3(n9418), .IN4(n9419), .QN(n9415) );
  NOR2X0 U9310 ( .IN1(n9375), .IN2(g952), .QN(n9419) );
  NOR2X0 U9311 ( .IN1(n9376), .IN2(g1296), .QN(n9418) );
  NOR2X0 U9312 ( .IN1(n5347), .IN2(n9377), .QN(n9417) );
  NOR2X0 U9313 ( .IN1(n9378), .IN2(DFF_1012_n1), .QN(n9416) );
  NOR2X0 U9314 ( .IN1(n9379), .IN2(n9420), .QN(n9414) );
  NOR2X0 U9316 ( .IN1(n5484), .IN2(n9381), .QN(n9420) );
  NAND2X0 U9317 ( .IN1(n1415), .IN2(n9421), .QN(n9413) );
  NAND4X0 U9318 ( .IN1(n9422), .IN2(n9423), .IN3(n9424), .IN4(n9425), .QN(
        n9421) );
  NOR4X0 U9319 ( .IN1(n9426), .IN2(n9427), .IN3(n9428), .IN4(n9429), .QN(n9425) );
  NOR2X0 U9320 ( .IN1(n5488), .IN2(n9430), .QN(n9429) );
  NOR2X0 U9321 ( .IN1(n5342), .IN2(n9431), .QN(n9428) );
  NOR2X0 U9322 ( .IN1(n5292), .IN2(n9390), .QN(n9427) );
  NAND3X0 U9323 ( .IN1(n9432), .IN2(n9433), .IN3(n9434), .QN(n9426) );
  NAND2X0 U9324 ( .IN1(n9408), .IN2(g572), .QN(n9434) );
  NAND2X0 U9325 ( .IN1(n8468), .IN2(n9435), .QN(n9433) );
  NAND2X0 U9326 ( .IN1(test_so2), .IN2(n9436), .QN(n9432) );
  NOR3X0 U9327 ( .IN1(n9437), .IN2(n9438), .IN3(n9439), .QN(n9424) );
  NOR2X0 U9328 ( .IN1(n8536), .IN2(n9440), .QN(n9439) );
  NOR2X0 U9329 ( .IN1(n5475), .IN2(n9441), .QN(n9438) );
  NOR2X0 U9330 ( .IN1(n5494), .IN2(n9402), .QN(n9437) );
  NAND2X0 U9331 ( .IN1(test_so22), .IN2(n9442), .QN(n9423) );
  NAND2X0 U9332 ( .IN1(n9443), .IN2(g2878), .QN(n9422) );
  NAND2X0 U9333 ( .IN1(n9410), .IN2(g2130), .QN(n9412) );
  INVX0 U9334 ( .INP(n9444), .ZN(g34923) );
  NOR2X0 U9335 ( .IN1(g34977), .IN2(n8154), .QN(n9444) );
  NAND4X0 U9336 ( .IN1(n9445), .IN2(n9446), .IN3(n9447), .IN4(n9448), .QN(
        g34977) );
  NOR4X0 U9337 ( .IN1(n9449), .IN2(n9450), .IN3(n9451), .IN4(n9452), .QN(n9448) );
  NOR2X0 U9338 ( .IN1(n5286), .IN2(n9375), .QN(n9452) );
  NOR2X0 U9339 ( .IN1(n2549), .IN2(n9376), .QN(n9451) );
  NOR2X0 U9340 ( .IN1(n9453), .IN2(g4927), .QN(n9450) );
  NOR2X0 U9341 ( .IN1(n9454), .IN2(g4737), .QN(n9449) );
  NOR2X0 U9342 ( .IN1(n9379), .IN2(n9455), .QN(n9447) );
  NOR2X0 U9343 ( .IN1(n5639), .IN2(n9381), .QN(n9455) );
  NAND2X0 U9344 ( .IN1(n1415), .IN2(n9456), .QN(n9446) );
  NAND2X0 U9345 ( .IN1(n9457), .IN2(n9458), .QN(n9456) );
  NOR4X0 U9346 ( .IN1(n9459), .IN2(n9460), .IN3(n9461), .IN4(n9462), .QN(n9458) );
  NOR2X0 U9347 ( .IN1(n9431), .IN2(g30327), .QN(n9462) );
  NOR2X0 U9348 ( .IN1(n8451), .IN2(n9430), .QN(n9460) );
  NAND3X0 U9349 ( .IN1(n9463), .IN2(n9464), .IN3(n9465), .QN(n9459) );
  NAND2X0 U9350 ( .IN1(n9436), .IN2(g758), .QN(n9465) );
  NAND2X0 U9351 ( .IN1(n9466), .IN2(g794), .QN(n9464) );
  NAND2X0 U9352 ( .IN1(n9435), .IN2(g534), .QN(n9463) );
  NOR4X0 U9353 ( .IN1(n9467), .IN2(n9468), .IN3(n9469), .IN4(n9470), .QN(n9457) );
  NOR2X0 U9354 ( .IN1(n8458), .IN2(n9401), .QN(n9470) );
  NOR2X0 U9355 ( .IN1(n5493), .IN2(n9402), .QN(n9469) );
  NOR2X0 U9356 ( .IN1(n8547), .IN2(n9403), .QN(n9468) );
  NAND3X0 U9357 ( .IN1(n9471), .IN2(n9472), .IN3(n9473), .QN(n9467) );
  NAND2X0 U9358 ( .IN1(n9407), .IN2(g2955), .QN(n9473) );
  NAND2X0 U9359 ( .IN1(n9408), .IN2(g586), .QN(n9472) );
  NAND2X0 U9360 ( .IN1(n9409), .IN2(g613), .QN(n9471) );
  INVX0 U9361 ( .INP(n9441), .ZN(n9409) );
  NAND2X0 U9362 ( .IN1(n9245), .IN2(n9474), .QN(n9445) );
  INVX0 U9363 ( .INP(n9378), .ZN(n9474) );
  NAND2X0 U9364 ( .IN1(n9475), .IN2(g22), .QN(g34921) );
  INVX0 U9365 ( .INP(g34976), .ZN(n9475) );
  NAND4X0 U9366 ( .IN1(n9476), .IN2(n9477), .IN3(n9478), .IN4(n9479), .QN(
        g34976) );
  NOR4X0 U9367 ( .IN1(n9480), .IN2(n9481), .IN3(n9482), .IN4(n9483), .QN(n9479) );
  NOR2X0 U9368 ( .IN1(n5297), .IN2(n9453), .QN(n9483) );
  NOR2X0 U9369 ( .IN1(n5345), .IN2(n9454), .QN(n9482) );
  NOR2X0 U9370 ( .IN1(n5497), .IN2(n9377), .QN(n9481) );
  NOR2X0 U9371 ( .IN1(n9378), .IN2(DFF_150_n1), .QN(n9480) );
  NOR3X0 U9372 ( .IN1(n9484), .IN2(n9379), .IN3(n9485), .QN(n9478) );
  NOR2X0 U9373 ( .IN1(n9376), .IN2(n9486), .QN(n9485) );
  NOR2X0 U9374 ( .IN1(n9375), .IN2(n9487), .QN(n9484) );
  NAND2X0 U9375 ( .IN1(n1415), .IN2(n9488), .QN(n9477) );
  NAND4X0 U9376 ( .IN1(n9489), .IN2(n9490), .IN3(n9491), .IN4(n9492), .QN(
        n9488) );
  NOR4X0 U9377 ( .IN1(n9493), .IN2(n9494), .IN3(n9461), .IN4(n9495), .QN(n9492) );
  NOR2X0 U9378 ( .IN1(n8485), .IN2(n9430), .QN(n9495) );
  NOR2X0 U9379 ( .IN1(n5479), .IN2(n9390), .QN(n9494) );
  NAND3X0 U9380 ( .IN1(n9496), .IN2(n9497), .IN3(n9498), .QN(n9493) );
  NAND2X0 U9381 ( .IN1(n9408), .IN2(g577), .QN(n9498) );
  NAND2X0 U9382 ( .IN1(test_so41), .IN2(n9435), .QN(n9497) );
  NAND2X0 U9383 ( .IN1(n9436), .IN2(g763), .QN(n9496) );
  NOR3X0 U9384 ( .IN1(n9499), .IN2(n9500), .IN3(n9501), .QN(n9491) );
  NOR2X0 U9385 ( .IN1(n8460), .IN2(n9440), .QN(n9501) );
  NOR2X0 U9386 ( .IN1(n5339), .IN2(n9441), .QN(n9500) );
  NOR2X0 U9387 ( .IN1(n9402), .IN2(n8625), .QN(n9499) );
  NAND2X0 U9388 ( .IN1(n9442), .IN2(g2936), .QN(n9490) );
  NAND2X0 U9389 ( .IN1(n9443), .IN2(g2898), .QN(n9489) );
  NAND2X0 U9390 ( .IN1(n9410), .IN2(g5160), .QN(n9476) );
  INVX0 U9391 ( .INP(n9502), .ZN(g34919) );
  NOR2X0 U9392 ( .IN1(g34975), .IN2(n8154), .QN(n9502) );
  NAND4X0 U9393 ( .IN1(n9503), .IN2(n9504), .IN3(n9505), .IN4(n9506), .QN(
        g34975) );
  NOR4X0 U9394 ( .IN1(n9507), .IN2(n9508), .IN3(n9509), .IN4(n9510), .QN(n9506) );
  NOR2X0 U9395 ( .IN1(n5295), .IN2(n9453), .QN(n9510) );
  NOR2X0 U9396 ( .IN1(n5344), .IN2(n9454), .QN(n9509) );
  NOR2X0 U9397 ( .IN1(n5495), .IN2(n9377), .QN(n9508) );
  NOR2X0 U9398 ( .IN1(n9378), .IN2(DFF_829_n1), .QN(n9507) );
  NOR3X0 U9399 ( .IN1(n9511), .IN2(n9379), .IN3(n9512), .QN(n9505) );
  NOR2X0 U9400 ( .IN1(n9376), .IN2(n9513), .QN(n9512) );
  NOR2X0 U9401 ( .IN1(n9375), .IN2(n9514), .QN(n9511) );
  NAND2X0 U9402 ( .IN1(n1415), .IN2(n9515), .QN(n9504) );
  NAND4X0 U9403 ( .IN1(n9516), .IN2(n9517), .IN3(n9518), .IN4(n9519), .QN(
        n9515) );
  NOR4X0 U9404 ( .IN1(n9520), .IN2(n9521), .IN3(n9522), .IN4(n9523), .QN(n9519) );
  NOR2X0 U9405 ( .IN1(n8144), .IN2(n9390), .QN(n9523) );
  NOR2X0 U9406 ( .IN1(n9430), .IN2(g2994), .QN(n9522) );
  NOR2X0 U9407 ( .IN1(n5492), .IN2(n9389), .QN(n9521) );
  NAND2X0 U9408 ( .IN1(n9524), .IN2(n9525), .QN(n9520) );
  NAND2X0 U9409 ( .IN1(n9436), .IN2(g767), .QN(n9525) );
  NAND2X0 U9410 ( .IN1(n9408), .IN2(g582), .QN(n9524) );
  NOR3X0 U9411 ( .IN1(n9526), .IN2(n9527), .IN3(n9528), .QN(n9518) );
  NOR2X0 U9412 ( .IN1(n8538), .IN2(n9440), .QN(n9528) );
  NOR2X0 U9413 ( .IN1(n5672), .IN2(n9441), .QN(n9527) );
  NOR2X0 U9414 ( .IN1(n8452), .IN2(n9402), .QN(n9526) );
  NAND2X0 U9415 ( .IN1(n9442), .IN2(g2922), .QN(n9517) );
  NAND2X0 U9416 ( .IN1(n9443), .IN2(g2864), .QN(n9516) );
  NAND2X0 U9417 ( .IN1(n9410), .IN2(g5507), .QN(n9503) );
  NAND2X0 U9418 ( .IN1(n9529), .IN2(g22), .QN(g34917) );
  INVX0 U9419 ( .INP(g34974), .ZN(n9529) );
  NAND4X0 U9420 ( .IN1(n9530), .IN2(n9531), .IN3(n9532), .IN4(n9533), .QN(
        g34974) );
  NOR4X0 U9421 ( .IN1(n9534), .IN2(n9535), .IN3(n9536), .IN4(n9537), .QN(n9533) );
  NOR2X0 U9422 ( .IN1(n5346), .IN2(n9453), .QN(n9537) );
  NOR2X0 U9423 ( .IN1(n5296), .IN2(n9454), .QN(n9536) );
  NOR2X0 U9424 ( .IN1(n9377), .IN2(n8606), .QN(n9535) );
  NOR2X0 U9425 ( .IN1(n9378), .IN2(DFF_477_n1), .QN(n9534) );
  NOR2X0 U9426 ( .IN1(n9538), .IN2(n9539), .QN(n9532) );
  NOR2X0 U9427 ( .IN1(n5499), .IN2(n9540), .QN(n9539) );
  NOR2X0 U9428 ( .IN1(n9541), .IN2(n9542), .QN(n9538) );
  NOR4X0 U9429 ( .IN1(n9543), .IN2(n9544), .IN3(n9545), .IN4(n9546), .QN(n9541) );
  NOR2X0 U9430 ( .IN1(n5288), .IN2(n9441), .QN(n9546) );
  NOR2X0 U9431 ( .IN1(n5472), .IN2(n9547), .QN(n9545) );
  NAND3X0 U9432 ( .IN1(n9548), .IN2(n9549), .IN3(n9550), .QN(n9544) );
  NAND2X0 U9433 ( .IN1(n9436), .IN2(g772), .QN(n9550) );
  NAND2X0 U9434 ( .IN1(n9395), .IN2(g2999), .QN(n9548) );
  NAND4X0 U9435 ( .IN1(n9551), .IN2(n9552), .IN3(n9553), .IN4(n9554), .QN(
        n9543) );
  NAND2X0 U9436 ( .IN1(n9407), .IN2(g2917), .QN(n9554) );
  NAND2X0 U9437 ( .IN1(n9555), .IN2(g2852), .QN(n9553) );
  NAND2X0 U9438 ( .IN1(n9442), .IN2(g2912), .QN(n9552) );
  NAND2X0 U9439 ( .IN1(n9443), .IN2(g2856), .QN(n9551) );
  INVX0 U9440 ( .INP(n9556), .ZN(n9531) );
  NOR2X0 U9441 ( .IN1(n9557), .IN2(n9376), .QN(n9556) );
  INVX0 U9442 ( .INP(n9558), .ZN(n9530) );
  NOR2X0 U9443 ( .IN1(n9559), .IN2(n9375), .QN(n9558) );
  NAND2X0 U9444 ( .IN1(n9337), .IN2(g22), .QN(g34915) );
  INVX0 U9445 ( .INP(g34971), .ZN(n9337) );
  NAND4X0 U9446 ( .IN1(n9560), .IN2(n9561), .IN3(n9562), .IN4(n9563), .QN(
        g34971) );
  NOR4X0 U9447 ( .IN1(n9379), .IN2(n9564), .IN3(n9565), .IN4(n9566), .QN(n9563) );
  NOR2X0 U9448 ( .IN1(n5307), .IN2(n9540), .QN(n9566) );
  NOR2X0 U9449 ( .IN1(n9567), .IN2(n9542), .QN(n9565) );
  NOR4X0 U9450 ( .IN1(n9568), .IN2(n9569), .IN3(n9570), .IN4(n9571), .QN(n9567) );
  NOR2X0 U9451 ( .IN1(n5983), .IN2(n9402), .QN(n9571) );
  NOR2X0 U9452 ( .IN1(n5550), .IN2(n9441), .QN(n9570) );
  NAND3X0 U9454 ( .IN1(n9572), .IN2(n9573), .IN3(n9574), .QN(n9569) );
  NAND2X0 U9455 ( .IN1(n9408), .IN2(g562), .QN(n9574) );
  INVX0 U9456 ( .INP(n9547), .ZN(n9408) );
  NAND2X0 U9457 ( .IN1(n9435), .IN2(g199), .QN(n9573) );
  NAND2X0 U9458 ( .IN1(test_so60), .IN2(n9436), .QN(n9572) );
  NAND4X0 U9459 ( .IN1(n9575), .IN2(n9576), .IN3(n9577), .IN4(n9578), .QN(
        n9568) );
  NAND2X0 U9460 ( .IN1(g100), .IN2(n9396), .QN(n9578) );
  INVX0 U9461 ( .INP(n9431), .ZN(n9396) );
  NAND3X0 U9462 ( .IN1(n9579), .IN2(g28), .IN3(n9580), .QN(n9431) );
  NOR2X0 U9463 ( .IN1(n9461), .IN2(n9581), .QN(n9577) );
  NOR2X0 U9464 ( .IN1(n5842), .IN2(n9338), .QN(n9581) );
  NAND4X0 U9465 ( .IN1(n9582), .IN2(test_so25), .IN3(n5324), .IN4(n8532), .QN(
        n9338) );
  INVX0 U9466 ( .INP(n9583), .ZN(n9461) );
  NAND4X0 U9467 ( .IN1(n9582), .IN2(g28), .IN3(g19), .IN4(n5477), .QN(n9583)
         );
  NAND2X0 U9468 ( .IN1(n9395), .IN2(g2890), .QN(n9576) );
  INVX0 U9469 ( .INP(n9430), .ZN(n9395) );
  NAND2X0 U9470 ( .IN1(n9580), .IN2(n9584), .QN(n9430) );
  NAND2X0 U9471 ( .IN1(n9466), .IN2(g781), .QN(n9575) );
  NOR2X0 U9472 ( .IN1(n5640), .IN2(n9381), .QN(n9564) );
  NAND2X0 U9473 ( .IN1(n9585), .IN2(n9584), .QN(n9381) );
  INVX0 U9474 ( .INP(n9586), .ZN(n9379) );
  NAND2X0 U9475 ( .IN1(n1415), .IN2(n9587), .QN(n9586) );
  NAND2X0 U9476 ( .IN1(n9549), .IN2(n9588), .QN(n9587) );
  NAND2X0 U9477 ( .IN1(n9466), .IN2(n8948), .QN(n9588) );
  INVX0 U9478 ( .INP(n9390), .ZN(n9466) );
  NAND2X0 U9479 ( .IN1(n9584), .IN2(n9589), .QN(n9390) );
  NOR2X0 U9480 ( .IN1(n9590), .IN2(n9591), .QN(n9562) );
  NOR2X0 U9481 ( .IN1(n5377), .IN2(n9377), .QN(n9591) );
  NOR2X0 U9482 ( .IN1(n9378), .IN2(DFF_206_n1), .QN(n9590) );
  NAND2X0 U9483 ( .IN1(test_so64), .IN2(n9592), .QN(n9561) );
  INVX0 U9484 ( .INP(n9376), .ZN(n9592) );
  INVX0 U9485 ( .INP(n9593), .ZN(n9560) );
  NOR2X0 U9486 ( .IN1(n9375), .IN2(n15226), .QN(n9593) );
  NAND2X0 U9487 ( .IN1(n9362), .IN2(g22), .QN(g34913) );
  INVX0 U9488 ( .INP(g34970), .ZN(n9362) );
  NAND4X0 U9489 ( .IN1(n9594), .IN2(n9595), .IN3(n9596), .IN4(n9597), .QN(
        g34970) );
  NOR4X0 U9490 ( .IN1(n9598), .IN2(n9599), .IN3(n9600), .IN4(n9601), .QN(n9597) );
  NOR2X0 U9491 ( .IN1(n5408), .IN2(n9453), .QN(n9601) );
  NAND3X0 U9492 ( .IN1(n1415), .IN2(n9584), .IN3(n2527), .QN(n9453) );
  NOR2X0 U9493 ( .IN1(n5312), .IN2(n9454), .QN(n9600) );
  NAND3X0 U9494 ( .IN1(n1415), .IN2(n9602), .IN3(n2527), .QN(n9454) );
  NOR2X0 U9495 ( .IN1(n5641), .IN2(n9377), .QN(n9599) );
  NAND3X0 U9496 ( .IN1(n9579), .IN2(n5324), .IN3(n9585), .QN(n9377) );
  NOR2X0 U9497 ( .IN1(n9378), .IN2(DFF_514_n1), .QN(n9598) );
  NAND2X0 U9498 ( .IN1(n9354), .IN2(n9542), .QN(n9378) );
  NOR2X0 U9499 ( .IN1(n9603), .IN2(n9604), .QN(n9596) );
  NOR2X0 U9500 ( .IN1(n9605), .IN2(n9542), .QN(n9604) );
  NOR4X0 U9501 ( .IN1(n9606), .IN2(n9607), .IN3(n9608), .IN4(n9609), .QN(n9605) );
  NOR2X0 U9502 ( .IN1(n15227), .IN2(n9441), .QN(n9609) );
  NOR2X0 U9503 ( .IN1(n5476), .IN2(n9547), .QN(n9608) );
  NAND3X0 U9504 ( .IN1(n9610), .IN2(n9549), .IN3(n9611), .QN(n9607) );
  NAND2X0 U9505 ( .IN1(n9436), .IN2(g776), .QN(n9611) );
  INVX0 U9506 ( .INP(n9391), .ZN(n9436) );
  NAND2X0 U9507 ( .IN1(n9012), .IN2(n9612), .QN(n9549) );
  NAND3X0 U9508 ( .IN1(n9547), .IN2(n9441), .IN3(n9391), .QN(n9612) );
  NAND3X0 U9509 ( .IN1(n9589), .IN2(g28), .IN3(n9579), .QN(n9391) );
  NAND2X0 U9510 ( .IN1(n2552), .IN2(n9602), .QN(n9441) );
  NAND3X0 U9511 ( .IN1(n2552), .IN2(n5324), .IN3(n9579), .QN(n9547) );
  INVX0 U9512 ( .INP(n9613), .ZN(n9579) );
  NAND4X0 U9513 ( .IN1(n8533), .IN2(n8117), .IN3(g31), .IN4(n8589), .QN(n9613)
         );
  NAND2X0 U9514 ( .IN1(n9435), .IN2(g538), .QN(n9610) );
  INVX0 U9515 ( .INP(n9389), .ZN(n9435) );
  NAND2X0 U9516 ( .IN1(n9602), .IN2(n9589), .QN(n9389) );
  NOR2X0 U9517 ( .IN1(g9), .IN2(n9614), .QN(n9589) );
  NAND4X0 U9518 ( .IN1(n9615), .IN2(n9616), .IN3(n9617), .IN4(n9618), .QN(
        n9606) );
  NAND2X0 U9519 ( .IN1(n9407), .IN2(g2902), .QN(n9618) );
  INVX0 U9520 ( .INP(n9440), .ZN(n9407) );
  NAND3X0 U9521 ( .IN1(n5324), .IN2(n9619), .IN3(n9582), .QN(n9440) );
  NAND2X0 U9522 ( .IN1(n9555), .IN2(g2844), .QN(n9617) );
  INVX0 U9523 ( .INP(n9402), .ZN(n9555) );
  NAND3X0 U9524 ( .IN1(n9619), .IN2(g9), .IN3(n9602), .QN(n9402) );
  NAND2X0 U9525 ( .IN1(test_so1), .IN2(n9442), .QN(n9616) );
  INVX0 U9526 ( .INP(n9401), .ZN(n9442) );
  NAND3X0 U9527 ( .IN1(n9619), .IN2(g28), .IN3(n9582), .QN(n9401) );
  NOR4X0 U9528 ( .IN1(n8589), .IN2(n9620), .IN3(n5468), .IN4(n8533), .QN(n9582) );
  INVX0 U9529 ( .INP(n3395), .ZN(n9620) );
  NAND2X0 U9530 ( .IN1(n9443), .IN2(g2848), .QN(n9615) );
  INVX0 U9531 ( .INP(n9403), .ZN(n9443) );
  NAND3X0 U9532 ( .IN1(n9619), .IN2(g9), .IN3(n9584), .QN(n9403) );
  INVX0 U9533 ( .INP(n9614), .ZN(n9619) );
  NAND2X0 U9534 ( .IN1(n8532), .IN2(n5477), .QN(n9614) );
  NOR2X0 U9535 ( .IN1(n9376), .IN2(n9621), .QN(n9603) );
  NAND3X0 U9536 ( .IN1(n1415), .IN2(n9602), .IN3(n9580), .QN(n9376) );
  NOR3X0 U9537 ( .IN1(g9), .IN2(g19), .IN3(n5477), .QN(n9580) );
  INVX0 U9538 ( .INP(n9622), .ZN(n9595) );
  NOR2X0 U9539 ( .IN1(n9623), .IN2(n9375), .QN(n9622) );
  NAND3X0 U9540 ( .IN1(n2552), .IN2(n9584), .IN3(n1415), .QN(n9375) );
  INVX0 U9541 ( .INP(n9542), .ZN(n1415) );
  NOR2X0 U9542 ( .IN1(n9624), .IN2(n5324), .QN(n9584) );
  NAND2X0 U9543 ( .IN1(n9410), .IN2(g6199), .QN(n9594) );
  INVX0 U9544 ( .INP(n9540), .ZN(n9410) );
  NAND2X0 U9545 ( .IN1(n9585), .IN2(n9602), .QN(n9540) );
  NOR2X0 U9546 ( .IN1(g28), .IN2(n9624), .QN(n9602) );
  NAND4X0 U9547 ( .IN1(n8533), .IN2(n8117), .IN3(n5469), .IN4(n8589), .QN(
        n9624) );
  NOR4X0 U9548 ( .IN1(n9542), .IN2(n5468), .IN3(n8532), .IN4(test_so25), .QN(
        n9585) );
  NAND4X0 U9549 ( .IN1(g54), .IN2(n9354), .IN3(n9625), .IN4(n9356), .QN(n9542)
         );
  INVX0 U9550 ( .INP(g56), .ZN(n9356) );
  NOR2X0 U9551 ( .IN1(test_so74), .IN2(g57), .QN(n9625) );
  INVX0 U9552 ( .INP(g53), .ZN(n9354) );
  NAND2X0 U9553 ( .IN1(n9626), .IN2(n9627), .QN(g34911) );
  NAND2X0 U9554 ( .IN1(n9628), .IN2(g807), .QN(n9627) );
  NAND2X0 U9555 ( .IN1(n8906), .IN2(n9629), .QN(n9628) );
  NAND2X0 U9556 ( .IN1(n2404), .IN2(g554), .QN(n9626) );
  NAND2X0 U9557 ( .IN1(n9630), .IN2(n9631), .QN(g34882) );
  NAND2X0 U9558 ( .IN1(n9012), .IN2(g4366), .QN(n9631) );
  NAND2X0 U9559 ( .IN1(n9632), .IN2(n8909), .QN(n9630) );
  NAND3X0 U9560 ( .IN1(n9633), .IN2(n9634), .IN3(n9635), .QN(n9632) );
  NAND3X0 U9561 ( .IN1(n5653), .IN2(n9636), .IN3(n9637), .QN(n9635) );
  NAND2X0 U9562 ( .IN1(n9638), .IN2(n5348), .QN(n9636) );
  INVX0 U9563 ( .INP(n9639), .ZN(n9638) );
  NAND3X0 U9564 ( .IN1(test_so81), .IN2(g4340), .IN3(g4358), .QN(n9634) );
  NAND3X0 U9565 ( .IN1(n9639), .IN2(n8590), .IN3(n5348), .QN(n9633) );
  NAND4X0 U9566 ( .IN1(n5653), .IN2(n8590), .IN3(n9640), .IN4(n9641), .QN(
        n9639) );
  NAND2X0 U9567 ( .IN1(n5540), .IN2(n9642), .QN(n9641) );
  NAND3X0 U9568 ( .IN1(n9643), .IN2(n9644), .IN3(n9645), .QN(n9642) );
  NAND2X0 U9569 ( .IN1(n8437), .IN2(g4322), .QN(n9644) );
  NAND3X0 U9570 ( .IN1(g90), .IN2(n5634), .IN3(n5506), .QN(n9643) );
  NAND3X0 U9571 ( .IN1(n5506), .IN2(g4311), .IN3(g4332), .QN(n9640) );
  NAND3X0 U9572 ( .IN1(n9646), .IN2(n9647), .IN3(n9648), .QN(g34881) );
  NAND2X0 U9573 ( .IN1(n9012), .IN2(g794), .QN(n9648) );
  NAND3X0 U9574 ( .IN1(n2404), .IN2(n9629), .IN3(g807), .QN(n9647) );
  INVX0 U9575 ( .INP(n2405), .ZN(n9629) );
  NAND2X0 U9576 ( .IN1(n2405), .IN2(n5479), .QN(n9646) );
  NAND3X0 U9577 ( .IN1(n9649), .IN2(n9650), .IN3(n9651), .QN(g34880) );
  NAND2X0 U9578 ( .IN1(n9012), .IN2(g626), .QN(n9651) );
  NAND3X0 U9579 ( .IN1(n2421), .IN2(n9652), .IN3(n9340), .QN(n9650) );
  INVX0 U9580 ( .INP(n2422), .ZN(n9652) );
  NAND2X0 U9581 ( .IN1(n2422), .IN2(n15227), .QN(n9649) );
  NAND3X0 U9582 ( .IN1(n9653), .IN2(n9654), .IN3(n9655), .QN(g34850) );
  NAND2X0 U9583 ( .IN1(n9012), .IN2(g790), .QN(n9655) );
  NAND3X0 U9584 ( .IN1(n2404), .IN2(n9656), .IN3(g794), .QN(n9654) );
  INVX0 U9585 ( .INP(n2419), .ZN(n9656) );
  NAND2X0 U9586 ( .IN1(n2419), .IN2(n5291), .QN(n9653) );
  NAND3X0 U9587 ( .IN1(n9657), .IN2(n9658), .IN3(n9659), .QN(g34849) );
  NAND2X0 U9588 ( .IN1(n9013), .IN2(g622), .QN(n9659) );
  NAND3X0 U9589 ( .IN1(n2421), .IN2(n9660), .IN3(g626), .QN(n9658) );
  INVX0 U9590 ( .INP(n2423), .ZN(n9660) );
  NAND2X0 U9591 ( .IN1(n2423), .IN2(n5288), .QN(n9657) );
  NOR2X0 U9592 ( .IN1(n8310), .IN2(n9661), .QN(g34839) );
  NOR3X0 U9593 ( .IN1(g4366), .IN2(n9662), .IN3(n9663), .QN(n9661) );
  NOR2X0 U9594 ( .IN1(n9664), .IN2(g4332), .QN(n9663) );
  NOR3X0 U9595 ( .IN1(g4311), .IN2(g73), .IN3(n9665), .QN(n9664) );
  NOR2X0 U9596 ( .IN1(n5540), .IN2(n9666), .QN(n9662) );
  NOR3X0 U9597 ( .IN1(n9667), .IN2(n9665), .IN3(g4311), .QN(n9666) );
  NAND2X0 U9598 ( .IN1(n9668), .IN2(n9669), .QN(g34808) );
  NAND2X0 U9599 ( .IN1(n9013), .IN2(g2955), .QN(n9669) );
  NAND2X0 U9600 ( .IN1(n9670), .IN2(n8909), .QN(n9668) );
  NAND3X0 U9601 ( .IN1(g91), .IN2(n9671), .IN3(n8536), .QN(n9670) );
  NAND2X0 U9602 ( .IN1(n9672), .IN2(n9673), .QN(g34807) );
  NAND2X0 U9603 ( .IN1(n9013), .IN2(g2941), .QN(n9673) );
  NAND2X0 U9604 ( .IN1(n9674), .IN2(n8909), .QN(n9672) );
  NAND4X0 U9605 ( .IN1(n9675), .IN2(n9676), .IN3(n9677), .IN4(n9678), .QN(
        n9674) );
  NOR4X0 U9606 ( .IN1(n9679), .IN2(n9680), .IN3(g2955), .IN4(g2946), .QN(n9678) );
  NOR2X0 U9607 ( .IN1(n9681), .IN2(n9682), .QN(n9677) );
  NAND2X0 U9608 ( .IN1(n9683), .IN2(n9684), .QN(g34806) );
  NAND2X0 U9609 ( .IN1(n9013), .IN2(g2927), .QN(n9684) );
  NAND2X0 U9610 ( .IN1(n9685), .IN2(n8910), .QN(n9683) );
  NAND3X0 U9611 ( .IN1(n8542), .IN2(n8460), .IN3(n8543), .QN(n9685) );
  NOR2X0 U9612 ( .IN1(n8949), .IN2(n9686), .QN(g34805) );
  INVX0 U9613 ( .INP(n9687), .ZN(n9686) );
  NAND2X0 U9614 ( .IN1(n8466), .IN2(n8537), .QN(n9687) );
  NAND2X0 U9615 ( .IN1(n9688), .IN2(n9689), .QN(g34804) );
  NAND2X0 U9616 ( .IN1(n9013), .IN2(g2965), .QN(n9689) );
  NAND2X0 U9617 ( .IN1(n9690), .IN2(n8910), .QN(n9688) );
  NAND3X0 U9618 ( .IN1(g962), .IN2(g1306), .IN3(n5750), .QN(n9690) );
  NAND2X0 U9619 ( .IN1(n9691), .IN2(n9692), .QN(g34803) );
  NAND2X0 U9620 ( .IN1(n9013), .IN2(g2917), .QN(n9692) );
  NAND2X0 U9621 ( .IN1(n9693), .IN2(n8910), .QN(n9691) );
  NAND3X0 U9622 ( .IN1(g44), .IN2(n8537), .IN3(n8538), .QN(n9693) );
  NAND2X0 U9623 ( .IN1(n9694), .IN2(n9695), .QN(g34802) );
  NAND2X0 U9624 ( .IN1(n9013), .IN2(g2902), .QN(n9695) );
  NAND2X0 U9625 ( .IN1(n9696), .IN2(n8910), .QN(n9694) );
  NAND3X0 U9626 ( .IN1(n9697), .IN2(n9698), .IN3(n8548), .QN(n9696) );
  NAND2X0 U9627 ( .IN1(n9699), .IN2(n9700), .QN(g34801) );
  NAND2X0 U9628 ( .IN1(n9014), .IN2(g2970), .QN(n9700) );
  NAND2X0 U9629 ( .IN1(n9701), .IN2(n8910), .QN(n9699) );
  NAND4X0 U9630 ( .IN1(n8546), .IN2(n8545), .IN3(n5595), .IN4(g691), .QN(n9701) );
  NAND2X0 U9631 ( .IN1(n9702), .IN2(n9703), .QN(g34799) );
  NAND2X0 U9632 ( .IN1(n9014), .IN2(g2873), .QN(n9703) );
  NAND2X0 U9633 ( .IN1(n9704), .IN2(n8911), .QN(n9702) );
  NAND2X0 U9634 ( .IN1(n8465), .IN2(g44), .QN(n9704) );
  NAND2X0 U9635 ( .IN1(n9705), .IN2(n9706), .QN(g34798) );
  NAND2X0 U9636 ( .IN1(n9014), .IN2(g2878), .QN(n9706) );
  NAND2X0 U9637 ( .IN1(n9707), .IN2(n8911), .QN(n9705) );
  NAND2X0 U9638 ( .IN1(n8462), .IN2(n8541), .QN(n9707) );
  NAND2X0 U9639 ( .IN1(n9708), .IN2(n9709), .QN(g34797) );
  NAND2X0 U9640 ( .IN1(n9014), .IN2(g2882), .QN(n9709) );
  NAND2X0 U9641 ( .IN1(n9710), .IN2(n8911), .QN(n9708) );
  NAND2X0 U9642 ( .IN1(n8461), .IN2(g91), .QN(n9710) );
  NAND2X0 U9643 ( .IN1(n9711), .IN2(n9712), .QN(g34796) );
  NAND2X0 U9644 ( .IN1(n9014), .IN2(g2898), .QN(n9712) );
  NAND2X0 U9645 ( .IN1(n9713), .IN2(n8912), .QN(n9711) );
  NAND2X0 U9646 ( .IN1(n8547), .IN2(n9671), .QN(n9713) );
  NOR2X0 U9647 ( .IN1(n9714), .IN2(n9715), .QN(n9671) );
  NAND2X0 U9648 ( .IN1(n9716), .IN2(n9717), .QN(g34795) );
  NAND2X0 U9649 ( .IN1(n9014), .IN2(g2864), .QN(n9717) );
  NAND2X0 U9650 ( .IN1(n9718), .IN2(n8912), .QN(n9716) );
  INVX0 U9651 ( .INP(n9719), .ZN(n9718) );
  NOR2X0 U9652 ( .IN1(g2898), .IN2(n9681), .QN(n9719) );
  NAND4X0 U9653 ( .IN1(n5882), .IN2(n5861), .IN3(n9720), .IN4(n9721), .QN(
        n9681) );
  NAND2X0 U9654 ( .IN1(n9722), .IN2(n9723), .QN(g34794) );
  NAND2X0 U9655 ( .IN1(n9014), .IN2(g2856), .QN(n9723) );
  NAND2X0 U9656 ( .IN1(n9724), .IN2(n8913), .QN(n9722) );
  INVX0 U9657 ( .INP(n9725), .ZN(n9724) );
  NOR2X0 U9658 ( .IN1(g2864), .IN2(n9682), .QN(n9725) );
  NAND3X0 U9659 ( .IN1(n9726), .IN2(n9727), .IN3(n9728), .QN(n9682) );
  NAND2X0 U9660 ( .IN1(n9729), .IN2(n9730), .QN(g34793) );
  NAND2X0 U9661 ( .IN1(n9015), .IN2(g2848), .QN(n9730) );
  NAND2X0 U9662 ( .IN1(n9731), .IN2(n8913), .QN(n9729) );
  NAND3X0 U9663 ( .IN1(n9732), .IN2(n9675), .IN3(n8549), .QN(n9731) );
  INVX0 U9664 ( .INP(n9679), .ZN(n9732) );
  NAND2X0 U9665 ( .IN1(n9733), .IN2(n9734), .QN(g34792) );
  NAND2X0 U9666 ( .IN1(n9015), .IN2(g29214), .QN(n9734) );
  NAND2X0 U9667 ( .IN1(n9735), .IN2(n8913), .QN(n9733) );
  NAND3X0 U9668 ( .IN1(n9736), .IN2(n9676), .IN3(n8544), .QN(n9735) );
  INVX0 U9669 ( .INP(n9680), .ZN(n9736) );
  NAND3X0 U9670 ( .IN1(n9737), .IN2(n9738), .IN3(n9739), .QN(g34791) );
  NAND2X0 U9671 ( .IN1(n9015), .IN2(g785), .QN(n9739) );
  NAND3X0 U9672 ( .IN1(n2404), .IN2(n9740), .IN3(g790), .QN(n9738) );
  INVX0 U9673 ( .INP(n2425), .ZN(n9740) );
  NAND2X0 U9674 ( .IN1(n2425), .IN2(n5292), .QN(n9737) );
  NAND3X0 U9675 ( .IN1(n9741), .IN2(n9742), .IN3(n9743), .QN(g34790) );
  NAND2X0 U9676 ( .IN1(n9015), .IN2(g617), .QN(n9743) );
  NAND3X0 U9677 ( .IN1(n2421), .IN2(n9744), .IN3(g622), .QN(n9742) );
  INVX0 U9678 ( .INP(n2427), .ZN(n9744) );
  NAND2X0 U9679 ( .IN1(n2427), .IN2(n5672), .QN(n9741) );
  NOR2X0 U9680 ( .IN1(n5305), .IN2(n9745), .QN(g34788) );
  NOR2X0 U9681 ( .IN1(n8151), .IN2(n9746), .QN(n9745) );
  INVX0 U9682 ( .INP(n3195), .ZN(n9746) );
  NAND2X0 U9683 ( .IN1(n9747), .IN2(n9748), .QN(g34783) );
  NAND3X0 U9684 ( .IN1(n9749), .IN2(n9750), .IN3(n9751), .QN(n9748) );
  NAND3X0 U9685 ( .IN1(n9752), .IN2(n9753), .IN3(n9754), .QN(n9747) );
  NAND2X0 U9686 ( .IN1(n9755), .IN2(n9756), .QN(g34735) );
  NAND2X0 U9687 ( .IN1(n9015), .IN2(g4297), .QN(n9756) );
  NAND2X0 U9688 ( .IN1(n9757), .IN2(n8913), .QN(n9755) );
  NAND2X0 U9689 ( .IN1(n5639), .IN2(n8464), .QN(n9757) );
  NAND2X0 U9690 ( .IN1(n9758), .IN2(n9759), .QN(g34734) );
  NAND2X0 U9691 ( .IN1(n9015), .IN2(g4172), .QN(n9759) );
  NAND2X0 U9692 ( .IN1(n9760), .IN2(n8913), .QN(n9758) );
  NAND2X0 U9693 ( .IN1(n5494), .IN2(n8543), .QN(n9760) );
  NOR2X0 U9694 ( .IN1(n8950), .IN2(n9761), .QN(g34733) );
  NOR2X0 U9695 ( .IN1(g4153), .IN2(g4172), .QN(n9761) );
  NAND2X0 U9696 ( .IN1(n9762), .IN2(n9763), .QN(g34732) );
  NAND2X0 U9697 ( .IN1(n8902), .IN2(g2994), .QN(n9763) );
  NAND2X0 U9698 ( .IN1(n9015), .IN2(g2999), .QN(n9762) );
  INVX0 U9699 ( .INP(n9764), .ZN(g34731) );
  NOR2X0 U9700 ( .IN1(n9765), .IN2(n9766), .QN(n9764) );
  NOR2X0 U9701 ( .IN1(n8900), .IN2(n5635), .QN(n9766) );
  NOR2X0 U9702 ( .IN1(n9767), .IN2(n8927), .QN(n9765) );
  NOR2X0 U9703 ( .IN1(n9768), .IN2(test_so64), .QN(n9767) );
  NAND2X0 U9704 ( .IN1(n9769), .IN2(n9770), .QN(g34730) );
  NAND2X0 U9705 ( .IN1(n9016), .IN2(g1296), .QN(n9770) );
  NAND2X0 U9706 ( .IN1(n9771), .IN2(n8913), .QN(n9769) );
  NAND2X0 U9707 ( .IN1(n8467), .IN2(n5635), .QN(n9771) );
  NAND3X0 U9708 ( .IN1(n9772), .IN2(n9773), .IN3(n9774), .QN(g34729) );
  INVX0 U9709 ( .INP(n2499), .ZN(n9774) );
  NAND2X0 U9710 ( .IN1(n5796), .IN2(n8912), .QN(n9773) );
  INVX0 U9711 ( .INP(n9775), .ZN(n9772) );
  NOR2X0 U9712 ( .IN1(n8900), .IN2(n2549), .QN(n9775) );
  NAND2X0 U9713 ( .IN1(n9776), .IN2(n9777), .QN(g34728) );
  NAND2X0 U9714 ( .IN1(n9016), .IN2(g939), .QN(n9777) );
  NAND2X0 U9715 ( .IN1(n9778), .IN2(n8912), .QN(n9776) );
  NAND2X0 U9716 ( .IN1(n15226), .IN2(n9697), .QN(n9778) );
  NAND2X0 U9717 ( .IN1(n9779), .IN2(n9780), .QN(g34727) );
  NAND2X0 U9718 ( .IN1(n9016), .IN2(g952), .QN(n9780) );
  NAND2X0 U9719 ( .IN1(n9781), .IN2(n8911), .QN(n9779) );
  NAND2X0 U9720 ( .IN1(n5415), .IN2(n8471), .QN(n9781) );
  NAND3X0 U9721 ( .IN1(n9782), .IN2(n9783), .IN3(n9784), .QN(g34726) );
  INVX0 U9722 ( .INP(n2505), .ZN(n9784) );
  NAND2X0 U9723 ( .IN1(n5630), .IN2(n8911), .QN(n9783) );
  INVX0 U9724 ( .INP(n9785), .ZN(n9782) );
  NOR2X0 U9725 ( .IN1(n8900), .IN2(n5286), .QN(n9785) );
  NAND3X0 U9726 ( .IN1(n9786), .IN2(n9787), .IN3(n9788), .QN(g34725) );
  NAND2X0 U9727 ( .IN1(n9016), .IN2(g781), .QN(n9788) );
  NAND3X0 U9728 ( .IN1(n2404), .IN2(n9789), .IN3(g785), .QN(n9787) );
  INVX0 U9729 ( .INP(n2485), .ZN(n9789) );
  NAND2X0 U9730 ( .IN1(n2485), .IN2(n5293), .QN(n9786) );
  NAND3X0 U9731 ( .IN1(n9790), .IN2(n9791), .IN3(n9792), .QN(g34724) );
  NAND2X0 U9732 ( .IN1(n9016), .IN2(g613), .QN(n9792) );
  NAND3X0 U9733 ( .IN1(n2421), .IN2(n9793), .IN3(g617), .QN(n9791) );
  INVX0 U9734 ( .INP(n2487), .ZN(n9793) );
  NAND2X0 U9735 ( .IN1(n2487), .IN2(n5339), .QN(n9790) );
  NAND2X0 U9736 ( .IN1(n9794), .IN2(n9795), .QN(g34723) );
  NAND2X0 U9737 ( .IN1(test_so41), .IN2(n8965), .QN(n9795) );
  NAND2X0 U9738 ( .IN1(n9796), .IN2(n8910), .QN(n9794) );
  NAND2X0 U9739 ( .IN1(n5490), .IN2(n8545), .QN(n9796) );
  NAND2X0 U9740 ( .IN1(n9797), .IN2(n9798), .QN(g34722) );
  NAND2X0 U9741 ( .IN1(n9016), .IN2(g538), .QN(n9798) );
  NAND2X0 U9742 ( .IN1(n9799), .IN2(n8910), .QN(n9797) );
  NAND2X0 U9743 ( .IN1(n5492), .IN2(g691), .QN(n9799) );
  NAND2X0 U9744 ( .IN1(n9800), .IN2(n9801), .QN(g34721) );
  NAND2X0 U9745 ( .IN1(g29221), .IN2(n9051), .QN(n9801) );
  NAND2X0 U9746 ( .IN1(n9802), .IN2(n8910), .QN(n9800) );
  NAND2X0 U9747 ( .IN1(n8470), .IN2(n8469), .QN(n9802) );
  NAND2X0 U9748 ( .IN1(n9803), .IN2(n9804), .QN(g34720) );
  NAND2X0 U9749 ( .IN1(n9016), .IN2(g534), .QN(n9804) );
  NAND2X0 U9750 ( .IN1(n9805), .IN2(n8910), .QN(n9803) );
  NAND2X0 U9751 ( .IN1(n8468), .IN2(g29212), .QN(n9805) );
  NOR2X0 U9752 ( .IN1(n8950), .IN2(n9806), .QN(g34719) );
  NOR2X0 U9753 ( .IN1(g209), .IN2(g538), .QN(n9806) );
  NOR2X0 U9754 ( .IN1(n5497), .IN2(n8927), .QN(g34647) );
  NOR2X0 U9755 ( .IN1(n5644), .IN2(n8937), .QN(g34646) );
  NOR2X0 U9756 ( .IN1(n5499), .IN2(n8927), .QN(g34645) );
  NOR2X0 U9757 ( .IN1(n5643), .IN2(n8936), .QN(g34644) );
  NOR2X0 U9758 ( .IN1(n5498), .IN2(n8930), .QN(g34643) );
  NAND2X0 U9759 ( .IN1(n9807), .IN2(n9808), .QN(g34642) );
  NAND2X0 U9760 ( .IN1(n8903), .IN2(g4927), .QN(n9808) );
  NAND2X0 U9761 ( .IN1(n9017), .IN2(g4912), .QN(n9807) );
  NAND2X0 U9762 ( .IN1(n9809), .IN2(n9810), .QN(g34641) );
  NAND2X0 U9763 ( .IN1(n8903), .IN2(g4912), .QN(n9810) );
  NAND2X0 U9764 ( .IN1(n9017), .IN2(g4907), .QN(n9809) );
  NAND2X0 U9765 ( .IN1(n9811), .IN2(n9812), .QN(g34640) );
  NAND2X0 U9766 ( .IN1(n8903), .IN2(g4907), .QN(n9812) );
  NAND2X0 U9767 ( .IN1(n9017), .IN2(g4922), .QN(n9811) );
  NAND2X0 U9768 ( .IN1(n9813), .IN2(n9814), .QN(g34639) );
  NAND2X0 U9769 ( .IN1(n8903), .IN2(g4922), .QN(n9814) );
  NAND2X0 U9770 ( .IN1(n9017), .IN2(g4917), .QN(n9813) );
  NOR2X0 U9771 ( .IN1(n5408), .IN2(n8940), .QN(g34638) );
  NAND2X0 U9772 ( .IN1(n9815), .IN2(n9816), .QN(g34637) );
  NAND2X0 U9773 ( .IN1(n8903), .IN2(g4737), .QN(n9816) );
  NAND2X0 U9774 ( .IN1(n9017), .IN2(g4722), .QN(n9815) );
  NAND2X0 U9775 ( .IN1(n9817), .IN2(n9818), .QN(g34636) );
  NAND2X0 U9776 ( .IN1(n8903), .IN2(g4722), .QN(n9818) );
  NAND2X0 U9777 ( .IN1(n9017), .IN2(g4717), .QN(n9817) );
  NAND2X0 U9778 ( .IN1(n9819), .IN2(n9820), .QN(g34635) );
  NAND2X0 U9779 ( .IN1(n8903), .IN2(g4717), .QN(n9820) );
  NAND2X0 U9780 ( .IN1(n9017), .IN2(g4732), .QN(n9819) );
  NAND2X0 U9781 ( .IN1(n9821), .IN2(n9822), .QN(g34634) );
  NAND2X0 U9782 ( .IN1(n8903), .IN2(g4732), .QN(n9822) );
  NAND2X0 U9783 ( .IN1(n9018), .IN2(g4727), .QN(n9821) );
  NOR2X0 U9784 ( .IN1(n5312), .IN2(n8934), .QN(g34633) );
  NAND2X0 U9785 ( .IN1(n9823), .IN2(n9824), .QN(g34632) );
  NAND2X0 U9786 ( .IN1(n8903), .IN2(g4245), .QN(n9824) );
  NAND2X0 U9787 ( .IN1(test_so67), .IN2(n9052), .QN(n9823) );
  NAND2X0 U9788 ( .IN1(n9825), .IN2(n9826), .QN(g34631) );
  NAND2X0 U9789 ( .IN1(test_so67), .IN2(n8909), .QN(n9826) );
  NAND2X0 U9790 ( .IN1(n9018), .IN2(g4253), .QN(n9825) );
  NAND2X0 U9791 ( .IN1(n9827), .IN2(n9828), .QN(g34630) );
  NAND2X0 U9792 ( .IN1(n8903), .IN2(g4253), .QN(n9828) );
  NAND2X0 U9793 ( .IN1(n9018), .IN2(g4300), .QN(n9827) );
  NAND2X0 U9794 ( .IN1(n9829), .IN2(n9830), .QN(g34629) );
  NAND2X0 U9795 ( .IN1(n8903), .IN2(g4157), .QN(n9830) );
  NAND2X0 U9796 ( .IN1(n9018), .IN2(g4146), .QN(n9829) );
  NAND2X0 U9797 ( .IN1(n9831), .IN2(n9832), .QN(g34628) );
  NAND2X0 U9798 ( .IN1(n8903), .IN2(g4146), .QN(n9832) );
  NAND2X0 U9799 ( .IN1(n9018), .IN2(g4176), .QN(n9831) );
  NOR2X0 U9800 ( .IN1(n5641), .IN2(n8935), .QN(g34627) );
  NOR2X0 U9801 ( .IN1(n8952), .IN2(n8606), .QN(g34626) );
  NOR2X0 U9802 ( .IN1(n5495), .IN2(n8931), .QN(g34625) );
  NAND2X0 U9803 ( .IN1(n9833), .IN2(n9834), .QN(g34624) );
  NAND2X0 U9804 ( .IN1(n8904), .IN2(g2988), .QN(n9834) );
  NAND2X0 U9805 ( .IN1(n9018), .IN2(g2994), .QN(n9833) );
  NAND2X0 U9806 ( .IN1(n9835), .IN2(n9836), .QN(g34623) );
  NAND2X0 U9807 ( .IN1(n8904), .IN2(g2970), .QN(n9836) );
  NAND2X0 U9808 ( .IN1(test_so22), .IN2(n9052), .QN(n9835) );
  NAND2X0 U9809 ( .IN1(n9837), .IN2(n9838), .QN(g34622) );
  NAND2X0 U9810 ( .IN1(test_so22), .IN2(n8908), .QN(n9838) );
  NAND2X0 U9811 ( .IN1(n9018), .IN2(g2950), .QN(n9837) );
  NAND2X0 U9812 ( .IN1(n9839), .IN2(n9840), .QN(g34621) );
  NAND2X0 U9813 ( .IN1(n8904), .IN2(g2950), .QN(n9840) );
  NAND2X0 U9814 ( .IN1(n9019), .IN2(g2936), .QN(n9839) );
  NAND2X0 U9815 ( .IN1(n9841), .IN2(n9842), .QN(g34620) );
  NAND2X0 U9816 ( .IN1(n8904), .IN2(g2936), .QN(n9842) );
  NAND2X0 U9817 ( .IN1(n9019), .IN2(g2922), .QN(n9841) );
  NAND2X0 U9818 ( .IN1(n9843), .IN2(n9844), .QN(g34619) );
  NAND2X0 U9819 ( .IN1(n8904), .IN2(g2922), .QN(n9844) );
  NAND2X0 U9820 ( .IN1(n9019), .IN2(g2912), .QN(n9843) );
  NAND2X0 U9821 ( .IN1(n9845), .IN2(n9846), .QN(g34618) );
  NAND2X0 U9822 ( .IN1(n8904), .IN2(g2912), .QN(n9846) );
  NAND2X0 U9823 ( .IN1(test_so1), .IN2(n9053), .QN(n9845) );
  NAND2X0 U9824 ( .IN1(n9847), .IN2(n9848), .QN(g34617) );
  NAND2X0 U9826 ( .IN1(test_so1), .IN2(n8908), .QN(n9848) );
  NAND2X0 U9827 ( .IN1(n9019), .IN2(g2984), .QN(n9847) );
  NAND2X0 U9828 ( .IN1(n9849), .IN2(n9850), .QN(g34616) );
  NAND2X0 U9829 ( .IN1(n8904), .IN2(g2868), .QN(n9850) );
  NAND2X0 U9830 ( .IN1(n9019), .IN2(g2988), .QN(n9849) );
  NAND2X0 U9831 ( .IN1(n9851), .IN2(n9852), .QN(g34615) );
  NAND2X0 U9832 ( .IN1(n8904), .IN2(g2873), .QN(n9852) );
  NAND2X0 U9833 ( .IN1(n9019), .IN2(g2868), .QN(n9851) );
  NAND2X0 U9834 ( .IN1(n9853), .IN2(n9854), .QN(g34614) );
  NAND2X0 U9835 ( .IN1(n8904), .IN2(g29214), .QN(n9854) );
  NAND2X0 U9836 ( .IN1(g37), .IN2(n9053), .QN(n9853) );
  NAND2X0 U9837 ( .IN1(n9855), .IN2(n9856), .QN(g34613) );
  NAND2X0 U9838 ( .IN1(test_so95), .IN2(n9053), .QN(n9856) );
  NAND2X0 U9839 ( .IN1(g37), .IN2(n8907), .QN(n9855) );
  NAND2X0 U9840 ( .IN1(n9857), .IN2(n9858), .QN(g34612) );
  NAND2X0 U9841 ( .IN1(test_so95), .IN2(n8907), .QN(n9858) );
  NAND2X0 U9842 ( .IN1(n9020), .IN2(g2860), .QN(n9857) );
  NAND2X0 U9843 ( .IN1(n9859), .IN2(n9860), .QN(g34611) );
  NAND2X0 U9844 ( .IN1(n8904), .IN2(g2860), .QN(n9860) );
  NAND2X0 U9845 ( .IN1(n9020), .IN2(g2852), .QN(n9859) );
  NAND2X0 U9846 ( .IN1(n9861), .IN2(n9862), .QN(g34610) );
  NAND2X0 U9847 ( .IN1(n8904), .IN2(g2852), .QN(n9862) );
  NAND2X0 U9848 ( .IN1(n9020), .IN2(g2844), .QN(n9861) );
  NAND2X0 U9849 ( .IN1(n9863), .IN2(n9864), .QN(g34609) );
  NAND2X0 U9850 ( .IN1(n8904), .IN2(g2844), .QN(n9864) );
  NAND2X0 U9851 ( .IN1(n9020), .IN2(g2890), .QN(n9863) );
  NAND2X0 U9852 ( .IN1(n9865), .IN2(n9866), .QN(g34608) );
  NAND2X0 U9853 ( .IN1(n8904), .IN2(g2704), .QN(n9866) );
  NAND2X0 U9854 ( .IN1(n9020), .IN2(g2697), .QN(n9865) );
  NAND2X0 U9855 ( .IN1(n9867), .IN2(n9868), .QN(g34607) );
  NAND2X0 U9856 ( .IN1(n8905), .IN2(g2697), .QN(n9868) );
  NAND2X0 U9857 ( .IN1(n9020), .IN2(g2689), .QN(n9867) );
  NOR2X0 U9858 ( .IN1(n5347), .IN2(n8933), .QN(g34606) );
  NAND2X0 U9859 ( .IN1(n9869), .IN2(n9870), .QN(g34605) );
  NAND2X0 U9860 ( .IN1(n8902), .IN2(g2145), .QN(n9870) );
  NAND2X0 U9861 ( .IN1(n9020), .IN2(g2138), .QN(n9869) );
  NAND2X0 U9862 ( .IN1(n9871), .IN2(n9872), .QN(g34604) );
  NAND2X0 U9863 ( .IN1(n8905), .IN2(g2138), .QN(n9872) );
  NAND2X0 U9864 ( .IN1(n9021), .IN2(g2130), .QN(n9871) );
  NOR2X0 U9865 ( .IN1(n5487), .IN2(n8933), .QN(g34603) );
  NOR2X0 U9866 ( .IN1(n2549), .IN2(n8934), .QN(g34602) );
  NOR2X0 U9867 ( .IN1(n5286), .IN2(n8934), .QN(g34601) );
  NAND3X0 U9868 ( .IN1(n9873), .IN2(n9874), .IN3(n9875), .QN(g34600) );
  NAND2X0 U9869 ( .IN1(n9021), .IN2(g776), .QN(n9875) );
  NAND3X0 U9870 ( .IN1(n2404), .IN2(n9876), .IN3(g781), .QN(n9874) );
  INVX0 U9871 ( .INP(n2507), .ZN(n9876) );
  NAND2X0 U9872 ( .IN1(n2507), .IN2(n5551), .QN(n9873) );
  NAND3X0 U9873 ( .IN1(n9877), .IN2(n9878), .IN3(n9879), .QN(g34599) );
  NAND2X0 U9874 ( .IN1(n9021), .IN2(g608), .QN(n9879) );
  NAND3X0 U9875 ( .IN1(n2421), .IN2(n9880), .IN3(g613), .QN(n9878) );
  INVX0 U9876 ( .INP(n2509), .ZN(n9880) );
  NAND2X0 U9877 ( .IN1(n2509), .IN2(n5474), .QN(n9877) );
  NAND2X0 U9878 ( .IN1(n9881), .IN2(n9882), .QN(g34598) );
  NAND2X0 U9879 ( .IN1(n9021), .IN2(g550), .QN(n9882) );
  NAND2X0 U9880 ( .IN1(g29221), .IN2(n8918), .QN(n9881) );
  NAND2X0 U9881 ( .IN1(n9883), .IN2(n9884), .QN(g34468) );
  NAND2X0 U9882 ( .IN1(n9885), .IN2(g4854), .QN(n9884) );
  NAND2X0 U9883 ( .IN1(n9886), .IN2(n8919), .QN(n9885) );
  NAND2X0 U9884 ( .IN1(n9887), .IN2(n9888), .QN(n9886) );
  NAND2X0 U9885 ( .IN1(n9889), .IN2(g4859), .QN(n9883) );
  NAND2X0 U9887 ( .IN1(n9890), .IN2(n9891), .QN(g34467) );
  NAND2X0 U9888 ( .IN1(n9892), .IN2(n9889), .QN(n9891) );
  XOR2X1 U9889 ( .IN1(g4854), .IN2(n9888), .Q(n9892) );
  NOR2X0 U9890 ( .IN1(n9893), .IN2(n8557), .QN(n9888) );
  INVX0 U9891 ( .INP(n2563), .ZN(n9893) );
  NAND2X0 U9892 ( .IN1(n9021), .IN2(g4849), .QN(n9890) );
  NAND2X0 U9893 ( .IN1(n9894), .IN2(n9895), .QN(g34466) );
  NAND2X0 U9894 ( .IN1(n9896), .IN2(g4878), .QN(n9895) );
  NAND2X0 U9895 ( .IN1(n9897), .IN2(n8919), .QN(n9896) );
  NAND2X0 U9896 ( .IN1(n8556), .IN2(n9887), .QN(n9897) );
  NAND3X0 U9897 ( .IN1(n9889), .IN2(g4843), .IN3(n5283), .QN(n9894) );
  NAND3X0 U9898 ( .IN1(n9898), .IN2(n9899), .IN3(n9900), .QN(g34465) );
  NAND2X0 U9899 ( .IN1(n9021), .IN2(g4843), .QN(n9900) );
  NAND3X0 U9900 ( .IN1(n9887), .IN2(n2563), .IN3(n8557), .QN(n9899) );
  NAND2X0 U9901 ( .IN1(n2567), .IN2(n9889), .QN(n9898) );
  INVX0 U9902 ( .INP(n9901), .ZN(n9889) );
  NAND2X0 U9903 ( .IN1(n9902), .IN2(n9903), .QN(g34464) );
  NAND2X0 U9904 ( .IN1(n9904), .IN2(g4664), .QN(n9903) );
  NAND2X0 U9905 ( .IN1(n9905), .IN2(n8919), .QN(n9904) );
  NAND2X0 U9906 ( .IN1(n9906), .IN2(n9907), .QN(n9905) );
  NAND2X0 U9907 ( .IN1(n9908), .IN2(g4669), .QN(n9902) );
  NAND2X0 U9908 ( .IN1(n9909), .IN2(n9910), .QN(g34463) );
  NAND2X0 U9909 ( .IN1(n9911), .IN2(n9908), .QN(n9910) );
  XOR2X1 U9910 ( .IN1(g4664), .IN2(n9907), .Q(n9911) );
  NOR2X0 U9911 ( .IN1(n9912), .IN2(n8554), .QN(n9907) );
  INVX0 U9912 ( .INP(n2573), .ZN(n9912) );
  NAND2X0 U9913 ( .IN1(n9021), .IN2(g4659), .QN(n9909) );
  NAND2X0 U9914 ( .IN1(n9913), .IN2(n9914), .QN(g34462) );
  NAND2X0 U9915 ( .IN1(n9915), .IN2(g4688), .QN(n9914) );
  NAND2X0 U9916 ( .IN1(n9916), .IN2(n8919), .QN(n9915) );
  NAND2X0 U9917 ( .IN1(n9906), .IN2(n8628), .QN(n9916) );
  NAND3X0 U9918 ( .IN1(n9908), .IN2(test_so19), .IN3(n5656), .QN(n9913) );
  NAND3X0 U9919 ( .IN1(n9917), .IN2(n9918), .IN3(n9919), .QN(g34461) );
  NAND2X0 U9920 ( .IN1(test_so19), .IN2(n9054), .QN(n9919) );
  NAND3X0 U9921 ( .IN1(n9906), .IN2(n2573), .IN3(n8554), .QN(n9918) );
  NAND2X0 U9922 ( .IN1(n2577), .IN2(n9908), .QN(n9917) );
  INVX0 U9923 ( .INP(n9920), .ZN(n9908) );
  NAND2X0 U9924 ( .IN1(n9921), .IN2(n9922), .QN(g34460) );
  NAND2X0 U9925 ( .IN1(n9923), .IN2(g4639), .QN(n9922) );
  NAND2X0 U9926 ( .IN1(n9924), .IN2(n8919), .QN(n9923) );
  NAND2X0 U9928 ( .IN1(n9925), .IN2(n8605), .QN(n9924) );
  NAND2X0 U9929 ( .IN1(n411), .IN2(test_so3), .QN(n9921) );
  INVX0 U9930 ( .INP(n9926), .ZN(n411) );
  NAND2X0 U9931 ( .IN1(n9927), .IN2(n9928), .QN(g34459) );
  NAND2X0 U9932 ( .IN1(n9022), .IN2(g4643), .QN(n9928) );
  NAND2X0 U9933 ( .IN1(n9929), .IN2(n8919), .QN(n9927) );
  NAND2X0 U9934 ( .IN1(n9930), .IN2(n9931), .QN(n9929) );
  NAND2X0 U9935 ( .IN1(n9932), .IN2(n9933), .QN(n9931) );
  NAND2X0 U9936 ( .IN1(n5653), .IN2(n9934), .QN(n9932) );
  NAND2X0 U9937 ( .IN1(test_so99), .IN2(n9935), .QN(n9934) );
  NAND2X0 U9938 ( .IN1(n9936), .IN2(n9937), .QN(g34458) );
  NAND2X0 U9939 ( .IN1(n9938), .IN2(g4633), .QN(n9937) );
  NAND2X0 U9940 ( .IN1(n9939), .IN2(n9940), .QN(n9938) );
  NAND3X0 U9941 ( .IN1(n8894), .IN2(n8600), .IN3(n9925), .QN(n9940) );
  INVX0 U9942 ( .INP(n9941), .ZN(n9939) );
  NAND2X0 U9943 ( .IN1(test_so99), .IN2(n9942), .QN(n9936) );
  NAND2X0 U9944 ( .IN1(n9943), .IN2(n8919), .QN(n9942) );
  NAND4X0 U9945 ( .IN1(n5844), .IN2(n9925), .IN3(test_so3), .IN4(g4639), .QN(
        n9943) );
  NAND2X0 U9946 ( .IN1(n9944), .IN2(n9945), .QN(g34457) );
  NAND2X0 U9947 ( .IN1(test_so3), .IN2(n9946), .QN(n9945) );
  NAND2X0 U9948 ( .IN1(n9947), .IN2(n8919), .QN(n9946) );
  NAND3X0 U9949 ( .IN1(g4639), .IN2(n8600), .IN3(n9925), .QN(n9947) );
  NAND2X0 U9950 ( .IN1(test_so99), .IN2(n9941), .QN(n9944) );
  NAND2X0 U9951 ( .IN1(n9926), .IN2(n9948), .QN(n9941) );
  NAND3X0 U9952 ( .IN1(n8894), .IN2(n8605), .IN3(n9925), .QN(n9948) );
  INVX0 U9954 ( .INP(n9949), .ZN(n9925) );
  NAND3X0 U9955 ( .IN1(n5382), .IN2(n9950), .IN3(n5727), .QN(n9926) );
  NAND2X0 U9956 ( .IN1(n9951), .IN2(n9952), .QN(g34456) );
  NAND2X0 U9959 ( .IN1(n9953), .IN2(g4608), .QN(n9952) );
  NAND2X0 U9960 ( .IN1(n9954), .IN2(n8919), .QN(n9953) );
  NAND2X0 U9961 ( .IN1(n2590), .IN2(n9955), .QN(n9954) );
  NAND2X0 U9962 ( .IN1(n9956), .IN2(g4616), .QN(n9951) );
  NAND2X0 U9963 ( .IN1(n9957), .IN2(n9958), .QN(g34455) );
  NAND2X0 U9964 ( .IN1(n9959), .IN2(g4322), .QN(n9958) );
  NAND2X0 U9965 ( .IN1(n9960), .IN2(n8919), .QN(n9959) );
  NAND3X0 U9966 ( .IN1(n9961), .IN2(n9930), .IN3(n2594), .QN(n9960) );
  NAND2X0 U9967 ( .IN1(n2595), .IN2(g4332), .QN(n9957) );
  NAND2X0 U9969 ( .IN1(n9962), .IN2(n9963), .QN(g34454) );
  NAND2X0 U9970 ( .IN1(n9964), .IN2(n9956), .QN(n9963) );
  XOR2X1 U9971 ( .IN1(n2590), .IN2(g4608), .Q(n9964) );
  NAND2X0 U9973 ( .IN1(n9022), .IN2(g4601), .QN(n9962) );
  NAND3X0 U9974 ( .IN1(n9965), .IN2(n9966), .IN3(n9967), .QN(g34453) );
  NAND2X0 U9975 ( .IN1(n9022), .IN2(g4593), .QN(n9967) );
  NAND3X0 U9976 ( .IN1(n9956), .IN2(n9968), .IN3(g4601), .QN(n9966) );
  INVX0 U9977 ( .INP(n2598), .ZN(n9968) );
  NAND3X0 U9978 ( .IN1(n2598), .IN2(n9955), .IN3(n5365), .QN(n9965) );
  INVX0 U9979 ( .INP(n9969), .ZN(n9955) );
  NAND2X0 U9980 ( .IN1(n9970), .IN2(n9971), .QN(g34452) );
  NAND2X0 U9981 ( .IN1(n9972), .IN2(n9956), .QN(n9971) );
  XOR2X1 U9982 ( .IN1(g4593), .IN2(n2601), .Q(n9972) );
  NAND2X0 U9983 ( .IN1(n9022), .IN2(g4584), .QN(n9970) );
  NAND2X0 U9984 ( .IN1(n9973), .IN2(n9974), .QN(g34451) );
  NAND2X0 U9985 ( .IN1(n9975), .IN2(n9956), .QN(n9974) );
  NOR2X0 U9986 ( .IN1(n9969), .IN2(n8942), .QN(n9956) );
  NAND2X0 U9987 ( .IN1(n9930), .IN2(n9976), .QN(n9969) );
  NAND2X0 U9988 ( .IN1(n2601), .IN2(g4616), .QN(n9976) );
  NOR2X0 U9989 ( .IN1(n9961), .IN2(n5539), .QN(n2601) );
  XOR2X1 U9990 ( .IN1(n9961), .IN2(n5539), .Q(n9975) );
  NAND2X0 U9991 ( .IN1(n9022), .IN2(g4332), .QN(n9973) );
  NAND3X0 U9993 ( .IN1(n9977), .IN2(n9978), .IN3(n9979), .QN(g34450) );
  NAND2X0 U9994 ( .IN1(n9022), .IN2(g4311), .QN(n9979) );
  NAND3X0 U9995 ( .IN1(n2595), .IN2(n9980), .IN3(g4322), .QN(n9978) );
  INVX0 U9996 ( .INP(n2594), .ZN(n9980) );
  INVX0 U9997 ( .INP(n9981), .ZN(n2595) );
  NAND2X0 U9998 ( .IN1(n9950), .IN2(n9961), .QN(n9981) );
  NAND3X0 U9999 ( .IN1(g4322), .IN2(g4332), .IN3(n2607), .QN(n9961) );
  NOR2X0 U10000 ( .IN1(n9982), .IN2(n5348), .QN(n2607) );
  NAND3X0 U10001 ( .IN1(n2594), .IN2(n9930), .IN3(n5506), .QN(n9977) );
  NAND3X0 U10002 ( .IN1(n9983), .IN2(n9984), .IN3(n9985), .QN(g34448) );
  NAND2X0 U10003 ( .IN1(n9022), .IN2(g2827), .QN(n9985) );
  NAND3X0 U10004 ( .IN1(n8894), .IN2(g2819), .IN3(n9986), .QN(n9984) );
  NAND3X0 U10005 ( .IN1(n9987), .IN2(n9988), .IN3(n9989), .QN(n9983) );
  NAND2X0 U10006 ( .IN1(n9218), .IN2(g2827), .QN(n9988) );
  NAND3X0 U10007 ( .IN1(n9990), .IN2(n9991), .IN3(n9992), .QN(g34447) );
  NAND2X0 U10008 ( .IN1(n9023), .IN2(g2815), .QN(n9992) );
  NAND3X0 U10009 ( .IN1(n8895), .IN2(g2807), .IN3(n9993), .QN(n9991) );
  NAND3X0 U10010 ( .IN1(n9987), .IN2(n9994), .IN3(n9995), .QN(n9990) );
  NAND2X0 U10011 ( .IN1(n9218), .IN2(g2811), .QN(n9994) );
  NAND3X0 U10012 ( .IN1(n9996), .IN2(n9997), .IN3(n9998), .QN(g34446) );
  NAND2X0 U10013 ( .IN1(n9023), .IN2(g2819), .QN(n9998) );
  NAND3X0 U10014 ( .IN1(n8894), .IN2(g2815), .IN3(n9999), .QN(n9997) );
  NAND3X0 U10015 ( .IN1(n9987), .IN2(n10000), .IN3(n10001), .QN(n9996) );
  NAND2X0 U10016 ( .IN1(test_so37), .IN2(n9218), .QN(n10000) );
  NAND3X0 U10017 ( .IN1(n10002), .IN2(n10003), .IN3(n10004), .QN(g34445) );
  NAND2X0 U10018 ( .IN1(n9023), .IN2(g2807), .QN(n10004) );
  NAND3X0 U10019 ( .IN1(n8895), .IN2(g2803), .IN3(n10005), .QN(n10003) );
  NAND3X0 U10020 ( .IN1(n9987), .IN2(n10006), .IN3(n10007), .QN(n10002) );
  NAND2X0 U10021 ( .IN1(n9218), .IN2(g2799), .QN(n10006) );
  NOR2X0 U10022 ( .IN1(n10008), .IN2(n8942), .QN(n9987) );
  NOR2X0 U10023 ( .IN1(n1782), .IN2(n8629), .QN(n10008) );
  NAND3X0 U10024 ( .IN1(n10009), .IN2(n10010), .IN3(n10011), .QN(g34444) );
  NAND2X0 U10025 ( .IN1(n9023), .IN2(g2795), .QN(n10011) );
  NAND3X0 U10026 ( .IN1(n8896), .IN2(g2787), .IN3(n9986), .QN(n10010) );
  INVX0 U10027 ( .INP(n9989), .ZN(n9986) );
  NAND3X0 U10028 ( .IN1(n10012), .IN2(n10013), .IN3(n9989), .QN(n10009) );
  NOR2X0 U10029 ( .IN1(n10014), .IN2(n10015), .QN(n9989) );
  NAND2X0 U10030 ( .IN1(n9218), .IN2(g2795), .QN(n10013) );
  NAND3X0 U10031 ( .IN1(n10016), .IN2(n10017), .IN3(n10018), .QN(g34443) );
  NAND2X0 U10032 ( .IN1(n9023), .IN2(g2783), .QN(n10018) );
  NAND3X0 U10033 ( .IN1(n8895), .IN2(g2775), .IN3(n9993), .QN(n10017) );
  INVX0 U10034 ( .INP(n9995), .ZN(n9993) );
  NAND3X0 U10035 ( .IN1(n10012), .IN2(n10019), .IN3(n9995), .QN(n10016) );
  NOR2X0 U10036 ( .IN1(n10020), .IN2(n10015), .QN(n9995) );
  NAND2X0 U10037 ( .IN1(n9218), .IN2(g2779), .QN(n10019) );
  NAND3X0 U10038 ( .IN1(n10021), .IN2(n10022), .IN3(n10023), .QN(g34442) );
  NAND2X0 U10039 ( .IN1(n9023), .IN2(g2787), .QN(n10023) );
  NAND3X0 U10040 ( .IN1(n8896), .IN2(g2783), .IN3(n9999), .QN(n10022) );
  INVX0 U10041 ( .INP(n10001), .ZN(n9999) );
  NAND3X0 U10042 ( .IN1(n10012), .IN2(n10024), .IN3(n10001), .QN(n10021) );
  NOR2X0 U10043 ( .IN1(n10025), .IN2(n10015), .QN(n10001) );
  NAND2X0 U10044 ( .IN1(n9218), .IN2(g2791), .QN(n10024) );
  NAND3X0 U10045 ( .IN1(n10026), .IN2(n10027), .IN3(n10028), .QN(g34441) );
  NAND2X0 U10046 ( .IN1(n9023), .IN2(g2775), .QN(n10028) );
  NAND3X0 U10047 ( .IN1(n8896), .IN2(g2771), .IN3(n10005), .QN(n10027) );
  INVX0 U10048 ( .INP(n10007), .ZN(n10005) );
  NAND3X0 U10049 ( .IN1(n10012), .IN2(n10029), .IN3(n10007), .QN(n10026) );
  NOR2X0 U10050 ( .IN1(n10015), .IN2(n10030), .QN(n10007) );
  NAND2X0 U10051 ( .IN1(n9218), .IN2(g2767), .QN(n10029) );
  NOR2X0 U10052 ( .IN1(n10031), .IN2(n8934), .QN(n10012) );
  NOR2X0 U10053 ( .IN1(n1782), .IN2(n8630), .QN(n10031) );
  NAND2X0 U10054 ( .IN1(n10032), .IN2(n10033), .QN(g34440) );
  NAND2X0 U10055 ( .IN1(n9024), .IN2(g446), .QN(n10033) );
  NAND2X0 U10056 ( .IN1(n10034), .IN2(n8919), .QN(n10032) );
  NAND2X0 U10057 ( .IN1(n10035), .IN2(n10036), .QN(n10034) );
  NAND2X0 U10058 ( .IN1(n10037), .IN2(g862), .QN(n10036) );
  NAND2X0 U10059 ( .IN1(g896), .IN2(n10038), .QN(n10037) );
  NAND2X0 U10060 ( .IN1(n10039), .IN2(n10040), .QN(n10038) );
  NAND3X0 U10061 ( .IN1(n10041), .IN2(n10042), .IN3(n5821), .QN(n10039) );
  NAND2X0 U10062 ( .IN1(g890), .IN2(g896), .QN(n10035) );
  NAND3X0 U10063 ( .IN1(n10043), .IN2(n10044), .IN3(n10045), .QN(g34439) );
  NAND2X0 U10064 ( .IN1(n9024), .IN2(g772), .QN(n10045) );
  NAND3X0 U10065 ( .IN1(n2404), .IN2(n10046), .IN3(g776), .QN(n10044) );
  INVX0 U10066 ( .INP(n2554), .ZN(n10046) );
  NAND2X0 U10067 ( .IN1(n2554), .IN2(n5330), .QN(n10043) );
  NAND3X0 U10068 ( .IN1(n10047), .IN2(n10048), .IN3(n10049), .QN(g34438) );
  NAND2X0 U10069 ( .IN1(n9024), .IN2(g604), .QN(n10049) );
  NAND3X0 U10070 ( .IN1(n2421), .IN2(n10050), .IN3(g608), .QN(n10048) );
  INVX0 U10071 ( .INP(n2556), .ZN(n10050) );
  NAND2X0 U10072 ( .IN1(n2556), .IN2(n5475), .QN(n10047) );
  NOR4X0 U10073 ( .IN1(n10051), .IN2(g4064), .IN3(g4057), .IN4(g4125), .QN(
        g34435) );
  NOR3X0 U10074 ( .IN1(g4082), .IN2(n10052), .IN3(g4141), .QN(n10051) );
  NOR4X0 U10075 ( .IN1(n8431), .IN2(n10053), .IN3(g4098), .IN4(n8598), .QN(
        n10052) );
  NAND2X0 U10076 ( .IN1(n2730), .IN2(n10054), .QN(g34425) );
  INVX0 U10077 ( .INP(n8572), .ZN(n10054) );
  NAND2X0 U10078 ( .IN1(n10055), .IN2(n10056), .QN(n8572) );
  NAND2X0 U10079 ( .IN1(n10057), .IN2(g4358), .QN(n10056) );
  NAND2X0 U10080 ( .IN1(n10058), .IN2(n10059), .QN(n10057) );
  NAND2X0 U10081 ( .IN1(test_so81), .IN2(n10060), .QN(n10059) );
  NAND2X0 U10082 ( .IN1(n10061), .IN2(n10062), .QN(n10060) );
  NAND2X0 U10083 ( .IN1(n10063), .IN2(n9753), .QN(n10062) );
  NAND2X0 U10084 ( .IN1(n10064), .IN2(n9750), .QN(n10061) );
  NAND2X0 U10085 ( .IN1(n10065), .IN2(n8590), .QN(n10058) );
  NAND2X0 U10086 ( .IN1(n10066), .IN2(n10067), .QN(n10065) );
  NAND2X0 U10087 ( .IN1(n10068), .IN2(n9753), .QN(n10067) );
  NAND2X0 U10088 ( .IN1(n10069), .IN2(n9750), .QN(n10066) );
  NAND2X0 U10089 ( .IN1(n10070), .IN2(n5348), .QN(n10055) );
  NAND2X0 U10090 ( .IN1(n10071), .IN2(n10072), .QN(n10070) );
  NAND2X0 U10091 ( .IN1(test_so81), .IN2(n10073), .QN(n10072) );
  NAND2X0 U10092 ( .IN1(n10074), .IN2(n10075), .QN(n10073) );
  NAND2X0 U10093 ( .IN1(n10076), .IN2(n9753), .QN(n10075) );
  NAND2X0 U10094 ( .IN1(n10077), .IN2(n9750), .QN(n10074) );
  NAND2X0 U10095 ( .IN1(n10078), .IN2(n8590), .QN(n10071) );
  NAND2X0 U10096 ( .IN1(n10079), .IN2(n10080), .QN(n10078) );
  NAND2X0 U10097 ( .IN1(g31860), .IN2(n9753), .QN(n10080) );
  NAND2X0 U10098 ( .IN1(n9216), .IN2(n9750), .QN(n10079) );
  NOR2X0 U10099 ( .IN1(n10081), .IN2(n10082), .QN(n2730) );
  NOR2X0 U10100 ( .IN1(n9750), .IN2(n9753), .QN(n10082) );
  NAND3X0 U10101 ( .IN1(n10083), .IN2(n10084), .IN3(n10085), .QN(g34383) );
  INVX0 U10102 ( .INP(g34843), .ZN(n10084) );
  NAND4X0 U10103 ( .IN1(n10086), .IN2(n10087), .IN3(n10088), .IN4(n10089), 
        .QN(g34843) );
  NOR4X0 U10104 ( .IN1(n10090), .IN2(n10091), .IN3(n10092), .IN4(n10093), .QN(
        n10089) );
  NOR2X0 U10105 ( .IN1(n10094), .IN2(n10095), .QN(n10093) );
  INVX0 U10106 ( .INP(g25259), .ZN(n10095) );
  NOR2X0 U10107 ( .IN1(n2727), .IN2(n10096), .QN(n10092) );
  NOR2X0 U10108 ( .IN1(n10097), .IN2(n10098), .QN(n10091) );
  NOR2X0 U10109 ( .IN1(n3146), .IN2(n10099), .QN(n10090) );
  INVX0 U10110 ( .INP(n10100), .ZN(n10099) );
  NOR2X0 U10111 ( .IN1(n10101), .IN2(n10102), .QN(n10088) );
  NOR3X0 U10112 ( .IN1(g2040), .IN2(n5535), .IN3(n10103), .QN(n10102) );
  NAND3X0 U10113 ( .IN1(n10104), .IN2(g1802), .IN3(n5504), .QN(n10087) );
  NAND2X0 U10114 ( .IN1(n10105), .IN2(n10106), .QN(n10086) );
  NAND4X0 U10115 ( .IN1(n10107), .IN2(n10094), .IN3(n10098), .IN4(n10108), 
        .QN(n10083) );
  NOR4X0 U10116 ( .IN1(n10109), .IN2(n10110), .IN3(n10106), .IN4(n10111), .QN(
        n10108) );
  NAND2X0 U10117 ( .IN1(n10112), .IN2(n10113), .QN(g34269) );
  NAND2X0 U10118 ( .IN1(n9024), .IN2(g4961), .QN(n10113) );
  NAND3X0 U10119 ( .IN1(n10114), .IN2(n10115), .IN3(n10116), .QN(n10112) );
  NAND3X0 U10120 ( .IN1(n5614), .IN2(n10117), .IN3(n10118), .QN(n10115) );
  NAND3X0 U10121 ( .IN1(n5770), .IN2(n10119), .IN3(n10120), .QN(n10114) );
  NAND2X0 U10122 ( .IN1(n10121), .IN2(n10122), .QN(g34268) );
  NAND2X0 U10123 ( .IN1(n9024), .IN2(g4950), .QN(n10122) );
  NAND3X0 U10124 ( .IN1(n10123), .IN2(n10124), .IN3(n10116), .QN(n10121) );
  NAND3X0 U10125 ( .IN1(n5875), .IN2(n10117), .IN3(n10125), .QN(n10124) );
  NAND3X0 U10126 ( .IN1(n5772), .IN2(n10119), .IN3(n10126), .QN(n10123) );
  NAND2X0 U10127 ( .IN1(n10127), .IN2(n10128), .QN(g34267) );
  NAND2X0 U10128 ( .IN1(n10129), .IN2(n8919), .QN(n10128) );
  NAND2X0 U10129 ( .IN1(n10119), .IN2(n10130), .QN(n10129) );
  NAND3X0 U10130 ( .IN1(n10117), .IN2(g4933), .IN3(n10131), .QN(n10130) );
  NAND2X0 U10131 ( .IN1(n10132), .IN2(g4939), .QN(n10127) );
  NAND2X0 U10132 ( .IN1(n10133), .IN2(n8920), .QN(n10132) );
  NAND2X0 U10133 ( .IN1(n10134), .IN2(n10117), .QN(n10133) );
  NAND2X0 U10134 ( .IN1(n10135), .IN2(n10136), .QN(g34266) );
  NAND2X0 U10135 ( .IN1(n9024), .IN2(g4894), .QN(n10136) );
  NAND3X0 U10136 ( .IN1(n10137), .IN2(n10138), .IN3(n10116), .QN(n10135) );
  INVX0 U10137 ( .INP(n10139), .ZN(n10116) );
  NAND2X0 U10138 ( .IN1(n10140), .IN2(n8920), .QN(n10139) );
  NAND2X0 U10139 ( .IN1(n10141), .IN2(n10119), .QN(n10140) );
  NAND3X0 U10140 ( .IN1(n5863), .IN2(n10117), .IN3(n10142), .QN(n10138) );
  NAND3X0 U10141 ( .IN1(n5774), .IN2(n10119), .IN3(n9749), .QN(n10137) );
  NAND2X0 U10142 ( .IN1(n10141), .IN2(g71), .QN(n10119) );
  INVX0 U10143 ( .INP(n10117), .ZN(n10141) );
  NAND3X0 U10144 ( .IN1(n2668), .IN2(DFF_672_n1), .IN3(n5637), .QN(n10117) );
  NOR4X0 U10145 ( .IN1(g4864), .IN2(g4871), .IN3(g4836), .IN4(n9901), .QN(
        g34265) );
  NAND2X0 U10146 ( .IN1(n9887), .IN2(n8920), .QN(n9901) );
  NOR2X0 U10147 ( .IN1(n10143), .IN2(n9751), .QN(n9887) );
  NAND2X0 U10148 ( .IN1(n10144), .IN2(n10145), .QN(g34264) );
  NAND2X0 U10149 ( .IN1(n9024), .IN2(g4771), .QN(n10145) );
  NAND3X0 U10150 ( .IN1(n10146), .IN2(n10147), .IN3(n10148), .QN(n10144) );
  NAND3X0 U10151 ( .IN1(n5613), .IN2(n10149), .IN3(n10150), .QN(n10147) );
  NAND3X0 U10152 ( .IN1(n5769), .IN2(n10151), .IN3(n10152), .QN(n10146) );
  NAND2X0 U10153 ( .IN1(n10153), .IN2(n10154), .QN(g34263) );
  NAND2X0 U10154 ( .IN1(n9025), .IN2(g4760), .QN(n10154) );
  NAND3X0 U10155 ( .IN1(n10155), .IN2(n10156), .IN3(n10148), .QN(n10153) );
  NAND3X0 U10156 ( .IN1(n5877), .IN2(n10149), .IN3(n10157), .QN(n10156) );
  NAND3X0 U10157 ( .IN1(n5775), .IN2(n10151), .IN3(n10158), .QN(n10155) );
  NAND2X0 U10158 ( .IN1(n10159), .IN2(n10160), .QN(g34262) );
  NAND2X0 U10159 ( .IN1(n10161), .IN2(n8920), .QN(n10160) );
  NAND2X0 U10160 ( .IN1(n10151), .IN2(n10162), .QN(n10161) );
  NAND3X0 U10161 ( .IN1(n10149), .IN2(g4743), .IN3(n10163), .QN(n10162) );
  NAND2X0 U10162 ( .IN1(test_so18), .IN2(n10164), .QN(n10159) );
  NAND2X0 U10163 ( .IN1(n10165), .IN2(n8920), .QN(n10164) );
  NAND2X0 U10164 ( .IN1(n10166), .IN2(n10149), .QN(n10165) );
  NAND2X0 U10165 ( .IN1(n10167), .IN2(n10168), .QN(g34261) );
  NAND2X0 U10166 ( .IN1(n9025), .IN2(g4704), .QN(n10168) );
  NAND3X0 U10167 ( .IN1(n10169), .IN2(n10170), .IN3(n10148), .QN(n10167) );
  INVX0 U10168 ( .INP(n10171), .ZN(n10148) );
  NAND2X0 U10169 ( .IN1(n10172), .IN2(n8920), .QN(n10171) );
  NAND2X0 U10170 ( .IN1(n10173), .IN2(n10151), .QN(n10172) );
  NAND3X0 U10171 ( .IN1(n5862), .IN2(n10149), .IN3(n10174), .QN(n10170) );
  NAND3X0 U10172 ( .IN1(n5771), .IN2(n10151), .IN3(n9752), .QN(n10169) );
  NAND2X0 U10173 ( .IN1(n10173), .IN2(g101), .QN(n10151) );
  INVX0 U10174 ( .INP(n10149), .ZN(n10173) );
  NAND3X0 U10175 ( .IN1(n2668), .IN2(DFF_178_n1), .IN3(n5636), .QN(n10149) );
  NOR4X0 U10176 ( .IN1(g4674), .IN2(g4646), .IN3(g4681), .IN4(n9920), .QN(
        g34260) );
  NAND2X0 U10177 ( .IN1(n9906), .IN2(n8920), .QN(n9920) );
  NOR2X0 U10178 ( .IN1(n10175), .IN2(n9754), .QN(n9906) );
  NOR2X0 U10179 ( .IN1(n5844), .IN2(n10176), .QN(g34259) );
  NOR2X0 U10180 ( .IN1(n8953), .IN2(n10177), .QN(n10176) );
  NOR2X0 U10181 ( .IN1(n10178), .IN2(n9949), .QN(n10177) );
  NAND2X0 U10182 ( .IN1(n5382), .IN2(n9930), .QN(n9949) );
  NAND3X0 U10183 ( .IN1(n10179), .IN2(n10180), .IN3(n10181), .QN(g34258) );
  NAND2X0 U10184 ( .IN1(test_so81), .IN2(n9055), .QN(n10181) );
  NAND3X0 U10185 ( .IN1(n9950), .IN2(n9982), .IN3(g4358), .QN(n10180) );
  NAND3X0 U10186 ( .IN1(n10182), .IN2(n9930), .IN3(n5348), .QN(n10179) );
  INVX0 U10187 ( .INP(n9982), .ZN(n10182) );
  NAND2X0 U10188 ( .IN1(n10183), .IN2(test_so81), .QN(n9982) );
  NAND3X0 U10189 ( .IN1(n10184), .IN2(n10185), .IN3(n10186), .QN(g34257) );
  NAND2X0 U10190 ( .IN1(n9025), .IN2(g4340), .QN(n10186) );
  NAND3X0 U10191 ( .IN1(n9950), .IN2(test_so81), .IN3(n9933), .QN(n10185) );
  INVX0 U10192 ( .INP(n10187), .ZN(n9950) );
  NAND2X0 U10193 ( .IN1(n9930), .IN2(n8920), .QN(n10187) );
  NAND3X0 U10194 ( .IN1(n9930), .IN2(n8590), .IN3(n10183), .QN(n10184) );
  INVX0 U10195 ( .INP(n9933), .ZN(n10183) );
  NAND3X0 U10196 ( .IN1(n9935), .IN2(g4340), .IN3(test_so99), .QN(n9933) );
  INVX0 U10197 ( .INP(n10178), .ZN(n9935) );
  NAND2X0 U10198 ( .IN1(n9281), .IN2(n10188), .QN(n9930) );
  NAND2X0 U10199 ( .IN1(n9645), .IN2(n1782), .QN(n10188) );
  NAND2X0 U10200 ( .IN1(n10189), .IN2(n10190), .QN(g34256) );
  NAND2X0 U10201 ( .IN1(n9025), .IN2(g4369), .QN(n10190) );
  NAND2X0 U10202 ( .IN1(n10191), .IN2(n8920), .QN(n10189) );
  NAND3X0 U10203 ( .IN1(n10192), .IN2(n10193), .IN3(n5765), .QN(n10191) );
  NAND2X0 U10204 ( .IN1(n5671), .IN2(g4473), .QN(n10192) );
  NAND4X0 U10205 ( .IN1(n5671), .IN2(n10194), .IN3(n10193), .IN4(n8901), .QN(
        g34255) );
  NAND2X0 U10206 ( .IN1(test_so38), .IN2(g4473), .QN(n10194) );
  NAND2X0 U10207 ( .IN1(n10195), .IN2(n10196), .QN(g34254) );
  NAND2X0 U10208 ( .IN1(n10197), .IN2(g4473), .QN(n10196) );
  NAND4X0 U10209 ( .IN1(n8902), .IN2(g4643), .IN3(g4462), .IN4(n8584), .QN(
        n10197) );
  NAND2X0 U10210 ( .IN1(n10198), .IN2(n8920), .QN(n10195) );
  NOR2X0 U10211 ( .IN1(n8952), .IN2(n10199), .QN(g34253) );
  NOR3X0 U10212 ( .IN1(n8584), .IN2(n5671), .IN3(n10198), .QN(n10199) );
  INVX0 U10213 ( .INP(n10193), .ZN(n10198) );
  NAND3X0 U10214 ( .IN1(n10200), .IN2(g26960), .IN3(n5849), .QN(n10193) );
  NAND2X0 U10215 ( .IN1(n9645), .IN2(n10201), .QN(n10200) );
  NAND2X0 U10216 ( .IN1(n5846), .IN2(n2668), .QN(n10201) );
  NAND3X0 U10217 ( .IN1(n10202), .IN2(n10203), .IN3(n10204), .QN(g34252) );
  NAND2X0 U10218 ( .IN1(n9025), .IN2(g767), .QN(n10204) );
  NAND3X0 U10219 ( .IN1(n2404), .IN2(n10205), .IN3(g772), .QN(n10203) );
  INVX0 U10220 ( .INP(n2647), .ZN(n10205) );
  NAND2X0 U10221 ( .IN1(n2647), .IN2(n5334), .QN(n10202) );
  NAND3X0 U10222 ( .IN1(n10206), .IN2(n10207), .IN3(n10208), .QN(g34251) );
  NAND2X0 U10223 ( .IN1(n9025), .IN2(g599), .QN(n10208) );
  NAND3X0 U10224 ( .IN1(n2421), .IN2(n10209), .IN3(g604), .QN(n10207) );
  INVX0 U10225 ( .INP(n2649), .ZN(n10209) );
  NAND2X0 U10226 ( .IN1(n2649), .IN2(n5473), .QN(n10206) );
  NAND3X0 U10227 ( .IN1(n10210), .IN2(n10211), .IN3(n10212), .QN(g34250) );
  NAND2X0 U10228 ( .IN1(n9025), .IN2(g298), .QN(n10212) );
  NAND3X0 U10229 ( .IN1(n8568), .IN2(n10213), .IN3(g142), .QN(n10211) );
  INVX0 U10230 ( .INP(n2707), .ZN(n10213) );
  NAND2X0 U10231 ( .IN1(n5724), .IN2(n2707), .QN(n10210) );
  NAND3X0 U10232 ( .IN1(n10214), .IN2(n10215), .IN3(n10216), .QN(g34249) );
  NAND2X0 U10233 ( .IN1(n9026), .IN2(g157), .QN(n10216) );
  NAND3X0 U10234 ( .IN1(n10217), .IN2(n10218), .IN3(g160), .QN(n10215) );
  INVX0 U10235 ( .INP(n2710), .ZN(n10218) );
  NAND2X0 U10236 ( .IN1(n2710), .IN2(n5843), .QN(n10214) );
  NAND3X0 U10237 ( .IN1(n10219), .IN2(n10220), .IN3(n10085), .QN(g34201) );
  INVX0 U10238 ( .INP(g34781), .ZN(n10220) );
  NAND4X0 U10239 ( .IN1(n10221), .IN2(n10222), .IN3(n10223), .IN4(n10224), 
        .QN(g34781) );
  NOR4X0 U10240 ( .IN1(n10225), .IN2(n10226), .IN3(n10227), .IN4(n10228), .QN(
        n10224) );
  NOR3X0 U10241 ( .IN1(g2217), .IN2(n8479), .IN3(n3569), .QN(n10228) );
  NOR3X0 U10242 ( .IN1(g2351), .IN2(n3550), .IN3(n8591), .QN(n10227) );
  NOR3X0 U10243 ( .IN1(g2485), .IN2(n8481), .IN3(n3007), .QN(n10226) );
  NOR3X0 U10244 ( .IN1(g2619), .IN2(n8482), .IN3(n3006), .QN(n10225) );
  NOR2X0 U10245 ( .IN1(n10229), .IN2(n10230), .QN(n10223) );
  NOR2X0 U10246 ( .IN1(n3003), .IN2(n10231), .QN(n10230) );
  NOR3X0 U10247 ( .IN1(g1792), .IN2(n5596), .IN3(n1721), .QN(n10229) );
  NAND3X0 U10248 ( .IN1(n10232), .IN2(g2051), .IN3(n5507), .QN(n10222) );
  NAND3X0 U10249 ( .IN1(n10233), .IN2(g1917), .IN3(n5510), .QN(n10221) );
  NAND4X0 U10250 ( .IN1(n3588), .IN2(n3606), .IN3(n10234), .IN4(n10235), .QN(
        n10219) );
  NOR4X0 U10251 ( .IN1(n10236), .IN2(n10237), .IN3(n10238), .IN4(n10239), .QN(
        n10235) );
  NOR2X0 U10252 ( .IN1(n3005), .IN2(n10240), .QN(n10234) );
  NAND2X0 U10253 ( .IN1(n10241), .IN2(n10242), .QN(g34041) );
  NAND2X0 U10254 ( .IN1(n10243), .IN2(n10244), .QN(n10242) );
  XOR2X1 U10255 ( .IN1(n10245), .IN2(n5367), .Q(n10243) );
  NAND2X0 U10256 ( .IN1(n9026), .IN2(g5008), .QN(n10241) );
  NAND3X0 U10257 ( .IN1(n10246), .IN2(n10247), .IN3(n10248), .QN(g34040) );
  NAND2X0 U10258 ( .IN1(n9026), .IN2(g4975), .QN(n10248) );
  NAND2X0 U10259 ( .IN1(n10249), .IN2(n10250), .QN(n10247) );
  NAND2X0 U10260 ( .IN1(n10251), .IN2(n10252), .QN(n10249) );
  NAND2X0 U10261 ( .IN1(n10253), .IN2(n9297), .QN(n10252) );
  NAND2X0 U10262 ( .IN1(n9296), .IN2(n8920), .QN(n10251) );
  NAND2X0 U10263 ( .IN1(n10244), .IN2(g4899), .QN(n10246) );
  NAND2X0 U10264 ( .IN1(n10254), .IN2(n10255), .QN(g34039) );
  NAND2X0 U10265 ( .IN1(test_so58), .IN2(n10256), .QN(n10255) );
  NAND2X0 U10266 ( .IN1(n10257), .IN2(n8920), .QN(n10256) );
  NAND2X0 U10267 ( .IN1(n10258), .IN2(n10259), .QN(n10257) );
  NAND2X0 U10268 ( .IN1(n10244), .IN2(g4966), .QN(n10254) );
  NAND3X0 U10269 ( .IN1(n10260), .IN2(n10261), .IN3(n10262), .QN(g34038) );
  NAND2X0 U10270 ( .IN1(n9026), .IN2(g4983), .QN(n10262) );
  NAND3X0 U10271 ( .IN1(n10258), .IN2(n10259), .IN3(n8587), .QN(n10261) );
  INVX0 U10272 ( .INP(n10263), .ZN(n10259) );
  NAND3X0 U10273 ( .IN1(n10244), .IN2(n10263), .IN3(test_so58), .QN(n10260) );
  NAND3X0 U10274 ( .IN1(n10264), .IN2(n10265), .IN3(n10266), .QN(g34037) );
  NAND2X0 U10275 ( .IN1(n9004), .IN2(g4966), .QN(n10266) );
  NAND2X0 U10276 ( .IN1(n10244), .IN2(g4975), .QN(n10265) );
  INVX0 U10277 ( .INP(n10267), .ZN(n10244) );
  NAND2X0 U10278 ( .IN1(n10258), .IN2(n8920), .QN(n10267) );
  NOR2X0 U10279 ( .IN1(n10143), .IN2(n10253), .QN(n10258) );
  INVX0 U10280 ( .INP(n10250), .ZN(n10143) );
  NAND3X0 U10281 ( .IN1(n10253), .IN2(n10250), .IN3(n5360), .QN(n10264) );
  NOR2X0 U10282 ( .IN1(n10263), .IN2(n5706), .QN(n10253) );
  NAND2X0 U10283 ( .IN1(n9751), .IN2(g4983), .QN(n10263) );
  INVX0 U10284 ( .INP(n10245), .ZN(n9751) );
  NAND2X0 U10285 ( .IN1(n10268), .IN2(g4878), .QN(n10245) );
  NOR2X0 U10286 ( .IN1(n5443), .IN2(n10269), .QN(g34036) );
  NOR2X0 U10287 ( .IN1(n5318), .IN2(n10269), .QN(g34035) );
  NOR2X0 U10288 ( .IN1(n5713), .IN2(n10269), .QN(g34034) );
  NOR2X0 U10289 ( .IN1(n10250), .IN2(n8931), .QN(n10269) );
  NAND3X0 U10290 ( .IN1(n2760), .IN2(g63), .IN3(n9750), .QN(n10250) );
  NAND2X0 U10291 ( .IN1(n10270), .IN2(n10271), .QN(g34033) );
  NAND2X0 U10292 ( .IN1(n10272), .IN2(n10273), .QN(n10271) );
  XOR2X1 U10293 ( .IN1(g4793), .IN2(n9754), .Q(n10272) );
  NAND2X0 U10294 ( .IN1(n9049), .IN2(g4818), .QN(n10270) );
  NAND3X0 U10295 ( .IN1(n10274), .IN2(n10275), .IN3(n10276), .QN(g34032) );
  NAND2X0 U10296 ( .IN1(n9034), .IN2(g4785), .QN(n10276) );
  NAND2X0 U10297 ( .IN1(n10277), .IN2(n10278), .QN(n10275) );
  NAND2X0 U10298 ( .IN1(n10279), .IN2(n10280), .QN(n10277) );
  NAND2X0 U10299 ( .IN1(n10281), .IN2(n9254), .QN(n10280) );
  NAND2X0 U10300 ( .IN1(n9253), .IN2(n8920), .QN(n10279) );
  NAND2X0 U10301 ( .IN1(n10273), .IN2(g4709), .QN(n10274) );
  NAND2X0 U10302 ( .IN1(n10282), .IN2(n10283), .QN(g34031) );
  NAND2X0 U10303 ( .IN1(test_so29), .IN2(n10284), .QN(n10283) );
  NAND2X0 U10304 ( .IN1(n10285), .IN2(n8921), .QN(n10284) );
  NAND2X0 U10305 ( .IN1(n10286), .IN2(n10287), .QN(n10285) );
  NAND2X0 U10306 ( .IN1(n10273), .IN2(g4776), .QN(n10282) );
  NAND3X0 U10307 ( .IN1(n10288), .IN2(n10289), .IN3(n10290), .QN(g34030) );
  NAND2X0 U10308 ( .IN1(n9033), .IN2(g4793), .QN(n10290) );
  NAND3X0 U10309 ( .IN1(n10286), .IN2(n10287), .IN3(n8595), .QN(n10289) );
  INVX0 U10310 ( .INP(n10291), .ZN(n10287) );
  NAND3X0 U10311 ( .IN1(n10273), .IN2(n10291), .IN3(test_so29), .QN(n10288) );
  NAND3X0 U10312 ( .IN1(n10292), .IN2(n10293), .IN3(n10294), .QN(g34029) );
  NAND2X0 U10313 ( .IN1(n9040), .IN2(g4776), .QN(n10294) );
  NAND2X0 U10315 ( .IN1(n10273), .IN2(g4785), .QN(n10293) );
  INVX0 U10316 ( .INP(n10295), .ZN(n10273) );
  NAND2X0 U10317 ( .IN1(n10286), .IN2(n8921), .QN(n10295) );
  NOR2X0 U10319 ( .IN1(n10175), .IN2(n10281), .QN(n10286) );
  INVX0 U10320 ( .INP(n10278), .ZN(n10175) );
  NAND3X0 U10321 ( .IN1(n10281), .IN2(n10278), .IN3(n5361), .QN(n10292) );
  NOR2X0 U10322 ( .IN1(n10291), .IN2(n5707), .QN(n10281) );
  NAND2X0 U10323 ( .IN1(n9754), .IN2(g4793), .QN(n10291) );
  NOR2X0 U10324 ( .IN1(n10296), .IN2(n5656), .QN(n9754) );
  NOR2X0 U10325 ( .IN1(n5440), .IN2(n2774), .QN(g34027) );
  NOR2X0 U10326 ( .IN1(n5712), .IN2(n2774), .QN(g34026) );
  NOR2X0 U10327 ( .IN1(n10278), .IN2(n8957), .QN(n2774) );
  NAND3X0 U10328 ( .IN1(n2760), .IN2(g63), .IN3(n9753), .QN(n10278) );
  NAND4X0 U10329 ( .IN1(n10297), .IN2(n10298), .IN3(n10299), .IN4(n10300), 
        .QN(g34024) );
  NAND2X0 U10330 ( .IN1(n9039), .IN2(g4492), .QN(n10300) );
  NAND2X0 U10331 ( .IN1(n10301), .IN2(n8921), .QN(n10299) );
  NAND2X0 U10332 ( .IN1(n10302), .IN2(n10303), .QN(n10301) );
  NAND2X0 U10333 ( .IN1(n10304), .IN2(g4512), .QN(n10303) );
  NAND2X0 U10334 ( .IN1(n10305), .IN2(n9645), .QN(n10302) );
  NAND4X0 U10335 ( .IN1(n10306), .IN2(n10307), .IN3(n10297), .IN4(n10298), 
        .QN(g34023) );
  NAND3X0 U10336 ( .IN1(n8897), .IN2(g2988), .IN3(n9645), .QN(n10297) );
  NAND3X0 U10337 ( .IN1(n8898), .IN2(g4552), .IN3(n10304), .QN(n10307) );
  NAND2X0 U10338 ( .IN1(n10308), .IN2(n9325), .QN(n10306) );
  NAND2X0 U10339 ( .IN1(n10309), .IN2(n8922), .QN(n10308) );
  NAND4X0 U10340 ( .IN1(n9645), .IN2(g4555), .IN3(g4558), .IN4(g4561), .QN(
        n10309) );
  INVX0 U10341 ( .INP(n10304), .ZN(n9645) );
  NAND4X0 U10342 ( .IN1(n10310), .IN2(n9200), .IN3(n10311), .IN4(n10312), .QN(
        g34022) );
  NAND3X0 U10343 ( .IN1(n10313), .IN2(g2763), .IN3(n8889), .QN(n10312) );
  NAND2X0 U10344 ( .IN1(n9041), .IN2(g2759), .QN(n10311) );
  NAND2X0 U10345 ( .IN1(n10314), .IN2(n8052), .QN(n10310) );
  INVX0 U10346 ( .INP(n10313), .ZN(n10314) );
  NAND2X0 U10347 ( .IN1(n10315), .IN2(g2759), .QN(n10313) );
  NAND3X0 U10348 ( .IN1(n10316), .IN2(n10317), .IN3(n10318), .QN(g34021) );
  NAND2X0 U10349 ( .IN1(n9042), .IN2(g2648), .QN(n10318) );
  NAND2X0 U10350 ( .IN1(n10319), .IN2(n10320), .QN(n10317) );
  NAND2X0 U10351 ( .IN1(n10321), .IN2(g2567), .QN(n10316) );
  NAND2X0 U10352 ( .IN1(n10322), .IN2(n10323), .QN(g34020) );
  NAND2X0 U10353 ( .IN1(n10324), .IN2(g2629), .QN(n10323) );
  NAND2X0 U10354 ( .IN1(n10325), .IN2(n8923), .QN(n10324) );
  NAND2X0 U10355 ( .IN1(n10326), .IN2(g2643), .QN(n10325) );
  NAND2X0 U10356 ( .IN1(n10327), .IN2(n8913), .QN(n10322) );
  NAND2X0 U10357 ( .IN1(n10328), .IN2(n10329), .QN(n10327) );
  NAND2X0 U10358 ( .IN1(n10330), .IN2(n10331), .QN(n10329) );
  NAND2X0 U10359 ( .IN1(n10332), .IN2(n10333), .QN(n10331) );
  NAND2X0 U10360 ( .IN1(n8131), .IN2(n10334), .QN(n10333) );
  NAND2X0 U10361 ( .IN1(n10335), .IN2(g2643), .QN(n10328) );
  NAND2X0 U10362 ( .IN1(n10334), .IN2(n10336), .QN(n10335) );
  NAND2X0 U10363 ( .IN1(n10326), .IN2(g2555), .QN(n10336) );
  INVX0 U10364 ( .INP(n10330), .ZN(n10326) );
  NAND2X0 U10365 ( .IN1(n10337), .IN2(n10338), .QN(n10330) );
  NAND2X0 U10366 ( .IN1(n5755), .IN2(n10339), .QN(n10338) );
  NAND2X0 U10367 ( .IN1(n10340), .IN2(n10341), .QN(n10337) );
  NAND2X0 U10368 ( .IN1(n10342), .IN2(n9621), .QN(n10340) );
  NAND3X0 U10369 ( .IN1(n10343), .IN2(n10344), .IN3(n10345), .QN(g34019) );
  NAND2X0 U10370 ( .IN1(n10346), .IN2(n10320), .QN(n10345) );
  NAND3X0 U10371 ( .IN1(n10347), .IN2(g2583), .IN3(n8893), .QN(n10344) );
  INVX0 U10372 ( .INP(n10346), .ZN(n10347) );
  NOR2X0 U10373 ( .IN1(n10348), .IN2(n5521), .QN(n10346) );
  NAND2X0 U10374 ( .IN1(n9045), .IN2(g2571), .QN(n10343) );
  NAND3X0 U10375 ( .IN1(n10349), .IN2(n10350), .IN3(n10351), .QN(g34018) );
  NAND2X0 U10376 ( .IN1(n8999), .IN2(g2583), .QN(n10351) );
  NAND3X0 U10377 ( .IN1(n10320), .IN2(n5351), .IN3(n10352), .QN(n10350) );
  NAND2X0 U10378 ( .IN1(test_so61), .IN2(n10353), .QN(n10349) );
  INVX0 U10379 ( .INP(n10354), .ZN(n10353) );
  NOR2X0 U10380 ( .IN1(n10355), .IN2(n10356), .QN(n10354) );
  NOR2X0 U10381 ( .IN1(n10352), .IN2(n8932), .QN(n10356) );
  NAND3X0 U10382 ( .IN1(n10357), .IN2(n10358), .IN3(n10359), .QN(g34017) );
  NAND2X0 U10383 ( .IN1(n10360), .IN2(n10320), .QN(n10359) );
  INVX0 U10384 ( .INP(n10361), .ZN(n10360) );
  NAND3X0 U10385 ( .IN1(test_so66), .IN2(n10361), .IN3(n8893), .QN(n10358) );
  NAND3X0 U10386 ( .IN1(g2555), .IN2(g2629), .IN3(n10334), .QN(n10361) );
  NAND2X0 U10387 ( .IN1(test_so61), .IN2(n8945), .QN(n10357) );
  NAND3X0 U10388 ( .IN1(n10362), .IN2(n10363), .IN3(n10364), .QN(g34016) );
  NAND2X0 U10389 ( .IN1(n10365), .IN2(n10320), .QN(n10364) );
  INVX0 U10390 ( .INP(n10366), .ZN(n10365) );
  NAND3X0 U10391 ( .IN1(n10366), .IN2(g2571), .IN3(n8893), .QN(n10363) );
  NAND2X0 U10392 ( .IN1(n10352), .IN2(n5521), .QN(n10366) );
  NAND2X0 U10393 ( .IN1(n8999), .IN2(g2563), .QN(n10362) );
  NAND3X0 U10394 ( .IN1(n10367), .IN2(n10368), .IN3(n10369), .QN(g34015) );
  NAND2X0 U10395 ( .IN1(n10370), .IN2(n10320), .QN(n10369) );
  INVX0 U10396 ( .INP(n10371), .ZN(n10320) );
  NAND3X0 U10397 ( .IN1(n10372), .IN2(n10373), .IN3(n8893), .QN(n10371) );
  NAND2X0 U10398 ( .IN1(n10339), .IN2(g1585), .QN(n10373) );
  INVX0 U10399 ( .INP(n10341), .ZN(n10339) );
  NAND3X0 U10400 ( .IN1(n10342), .IN2(n9621), .IN3(n10341), .QN(n10372) );
  NAND3X0 U10401 ( .IN1(n10374), .IN2(g2563), .IN3(n8893), .QN(n10368) );
  INVX0 U10402 ( .INP(n10370), .ZN(n10374) );
  NOR2X0 U10403 ( .IN1(n10348), .IN2(n5351), .QN(n10370) );
  NAND2X0 U10404 ( .IN1(n8999), .IN2(g2567), .QN(n10367) );
  NAND3X0 U10405 ( .IN1(n10375), .IN2(n10376), .IN3(n10377), .QN(g34014) );
  NAND2X0 U10406 ( .IN1(n8999), .IN2(g2514), .QN(n10377) );
  NAND2X0 U10407 ( .IN1(n10378), .IN2(n10379), .QN(n10376) );
  NAND2X0 U10408 ( .IN1(n10380), .IN2(g2433), .QN(n10375) );
  NAND2X0 U10409 ( .IN1(n10381), .IN2(n10382), .QN(g34013) );
  NAND2X0 U10410 ( .IN1(n10383), .IN2(g2495), .QN(n10382) );
  NAND2X0 U10411 ( .IN1(n10384), .IN2(n8913), .QN(n10383) );
  NAND2X0 U10412 ( .IN1(n10385), .IN2(g2509), .QN(n10384) );
  NAND2X0 U10413 ( .IN1(n10386), .IN2(n8913), .QN(n10381) );
  NAND2X0 U10414 ( .IN1(n10387), .IN2(n10388), .QN(n10386) );
  NAND2X0 U10415 ( .IN1(n10389), .IN2(n10390), .QN(n10388) );
  NAND2X0 U10416 ( .IN1(n10391), .IN2(n10392), .QN(n10390) );
  NAND2X0 U10417 ( .IN1(n8130), .IN2(n10393), .QN(n10392) );
  NAND2X0 U10418 ( .IN1(n10394), .IN2(g2509), .QN(n10387) );
  NAND2X0 U10419 ( .IN1(n10393), .IN2(n10395), .QN(n10394) );
  NAND2X0 U10420 ( .IN1(test_so79), .IN2(n10385), .QN(n10395) );
  INVX0 U10421 ( .INP(n10389), .ZN(n10385) );
  NAND2X0 U10422 ( .IN1(n10396), .IN2(n10397), .QN(n10389) );
  NAND2X0 U10423 ( .IN1(n10398), .IN2(g1589), .QN(n10397) );
  NAND2X0 U10424 ( .IN1(n10399), .IN2(n10400), .QN(n10396) );
  NAND3X0 U10425 ( .IN1(n10401), .IN2(n10402), .IN3(n10403), .QN(g34012) );
  NAND2X0 U10426 ( .IN1(n8999), .IN2(g2437), .QN(n10403) );
  NAND3X0 U10427 ( .IN1(n10404), .IN2(n10393), .IN3(n10378), .QN(n10402) );
  NAND2X0 U10428 ( .IN1(n10405), .IN2(g2449), .QN(n10401) );
  NAND2X0 U10429 ( .IN1(n10406), .IN2(n10407), .QN(n10405) );
  NAND2X0 U10430 ( .IN1(n10096), .IN2(n8913), .QN(n10407) );
  NAND3X0 U10431 ( .IN1(n10408), .IN2(n10409), .IN3(n10410), .QN(g34011) );
  NAND2X0 U10432 ( .IN1(n10411), .IN2(n10378), .QN(n10410) );
  INVX0 U10433 ( .INP(n10412), .ZN(n10411) );
  NAND3X0 U10434 ( .IN1(n10412), .IN2(n9274), .IN3(n8893), .QN(n10409) );
  NAND2X0 U10435 ( .IN1(n10413), .IN2(n8585), .QN(n10412) );
  NAND2X0 U10436 ( .IN1(n8999), .IN2(g2449), .QN(n10408) );
  NAND3X0 U10437 ( .IN1(n10414), .IN2(n10415), .IN3(n10416), .QN(g34010) );
  NAND2X0 U10438 ( .IN1(n10417), .IN2(n10378), .QN(n10416) );
  INVX0 U10439 ( .INP(n10418), .ZN(n10417) );
  NAND3X0 U10440 ( .IN1(n10418), .IN2(g2441), .IN3(n8893), .QN(n10415) );
  NAND2X0 U10441 ( .IN1(n10419), .IN2(g2495), .QN(n10418) );
  NAND2X0 U10442 ( .IN1(n8999), .IN2(n9274), .QN(n10414) );
  NAND3X0 U10443 ( .IN1(n10420), .IN2(n10421), .IN3(n10422), .QN(g34009) );
  NAND2X0 U10444 ( .IN1(n10423), .IN2(n10378), .QN(n10422) );
  INVX0 U10445 ( .INP(n10424), .ZN(n10423) );
  NAND3X0 U10446 ( .IN1(n10424), .IN2(g2437), .IN3(n8893), .QN(n10421) );
  NAND2X0 U10447 ( .IN1(n10413), .IN2(n5522), .QN(n10424) );
  NAND2X0 U10448 ( .IN1(n9000), .IN2(g2429), .QN(n10420) );
  NAND3X0 U10449 ( .IN1(n10425), .IN2(n10426), .IN3(n10427), .QN(g34008) );
  NAND2X0 U10450 ( .IN1(n10428), .IN2(n10378), .QN(n10427) );
  NOR3X0 U10451 ( .IN1(n10429), .IN2(n10430), .IN3(n8924), .QN(n10378) );
  NOR2X0 U10452 ( .IN1(n10399), .IN2(n10398), .QN(n10430) );
  INVX0 U10453 ( .INP(n10400), .ZN(n10398) );
  NAND2X0 U10454 ( .IN1(n10342), .IN2(n9557), .QN(n10399) );
  NOR2X0 U10455 ( .IN1(g1585), .IN2(n10400), .QN(n10429) );
  INVX0 U10456 ( .INP(n10431), .ZN(n10428) );
  NAND3X0 U10457 ( .IN1(n10431), .IN2(g2429), .IN3(n8892), .QN(n10426) );
  NAND2X0 U10458 ( .IN1(n10419), .IN2(n5523), .QN(n10431) );
  NAND2X0 U10459 ( .IN1(n9000), .IN2(g2433), .QN(n10425) );
  NAND3X0 U10460 ( .IN1(n10432), .IN2(n10433), .IN3(n10434), .QN(g34007) );
  NAND2X0 U10461 ( .IN1(n9000), .IN2(g2380), .QN(n10434) );
  NAND2X0 U10462 ( .IN1(n10435), .IN2(n10436), .QN(n10433) );
  NAND2X0 U10463 ( .IN1(n10437), .IN2(g2299), .QN(n10432) );
  NAND2X0 U10464 ( .IN1(n10438), .IN2(n10439), .QN(g34006) );
  NAND2X0 U10465 ( .IN1(n10440), .IN2(g2361), .QN(n10439) );
  NAND2X0 U10466 ( .IN1(n10441), .IN2(n8914), .QN(n10440) );
  NAND2X0 U10467 ( .IN1(n10442), .IN2(g2375), .QN(n10441) );
  NAND2X0 U10468 ( .IN1(n10443), .IN2(n8913), .QN(n10438) );
  NAND2X0 U10469 ( .IN1(n10444), .IN2(n10445), .QN(n10443) );
  NAND2X0 U10470 ( .IN1(n10446), .IN2(n10447), .QN(n10445) );
  NAND2X0 U10471 ( .IN1(n10448), .IN2(n10449), .QN(n10447) );
  NAND2X0 U10472 ( .IN1(n8132), .IN2(n10450), .QN(n10449) );
  NAND2X0 U10473 ( .IN1(n10451), .IN2(g2375), .QN(n10444) );
  NAND2X0 U10474 ( .IN1(n10450), .IN2(n10452), .QN(n10451) );
  NAND2X0 U10475 ( .IN1(n10442), .IN2(g2287), .QN(n10452) );
  INVX0 U10476 ( .INP(n10446), .ZN(n10442) );
  NAND2X0 U10477 ( .IN1(n10453), .IN2(n10454), .QN(n10446) );
  NAND2X0 U10478 ( .IN1(n10455), .IN2(n5755), .QN(n10454) );
  NAND2X0 U10479 ( .IN1(n10456), .IN2(n10457), .QN(n10453) );
  NAND3X0 U10480 ( .IN1(n10458), .IN2(n10459), .IN3(n10460), .QN(g34005) );
  NAND2X0 U10481 ( .IN1(n10461), .IN2(n10435), .QN(n10460) );
  NAND3X0 U10482 ( .IN1(n10462), .IN2(g2315), .IN3(n8892), .QN(n10459) );
  INVX0 U10483 ( .INP(n10461), .ZN(n10462) );
  NOR2X0 U10484 ( .IN1(n10463), .IN2(n5537), .QN(n10461) );
  NAND2X0 U10485 ( .IN1(n9000), .IN2(g2303), .QN(n10458) );
  NAND3X0 U10486 ( .IN1(n10464), .IN2(n10465), .IN3(n10466), .QN(g34004) );
  NAND2X0 U10487 ( .IN1(n9000), .IN2(g2315), .QN(n10466) );
  NAND3X0 U10488 ( .IN1(n10435), .IN2(n5353), .IN3(n10467), .QN(n10465) );
  NAND2X0 U10489 ( .IN1(n10468), .IN2(n9314), .QN(n10464) );
  INVX0 U10490 ( .INP(n10469), .ZN(n10468) );
  NOR2X0 U10491 ( .IN1(n10470), .IN2(n10471), .QN(n10469) );
  NOR2X0 U10492 ( .IN1(n10467), .IN2(n8928), .QN(n10471) );
  NAND3X0 U10493 ( .IN1(n10472), .IN2(n10473), .IN3(n10474), .QN(g34003) );
  NAND2X0 U10494 ( .IN1(n10475), .IN2(n10435), .QN(n10474) );
  INVX0 U10495 ( .INP(n10476), .ZN(n10475) );
  NAND3X0 U10496 ( .IN1(n10476), .IN2(g2307), .IN3(n8892), .QN(n10473) );
  NAND3X0 U10497 ( .IN1(g2287), .IN2(g2361), .IN3(n10450), .QN(n10476) );
  NAND2X0 U10498 ( .IN1(n9000), .IN2(n9314), .QN(n10472) );
  NAND3X0 U10499 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .QN(g34002) );
  NAND2X0 U10500 ( .IN1(n10480), .IN2(n10435), .QN(n10479) );
  INVX0 U10501 ( .INP(n10481), .ZN(n10480) );
  NAND3X0 U10502 ( .IN1(n10481), .IN2(g2303), .IN3(n8892), .QN(n10478) );
  NAND2X0 U10503 ( .IN1(n10467), .IN2(n5537), .QN(n10481) );
  NAND2X0 U10504 ( .IN1(n9000), .IN2(g2295), .QN(n10477) );
  NAND3X0 U10505 ( .IN1(n10482), .IN2(n10483), .IN3(n10484), .QN(g34001) );
  NAND2X0 U10506 ( .IN1(n10485), .IN2(n10435), .QN(n10484) );
  NOR3X0 U10507 ( .IN1(n10486), .IN2(n10487), .IN3(n8924), .QN(n10435) );
  NOR2X0 U10508 ( .IN1(n10457), .IN2(n5757), .QN(n10487) );
  NOR2X0 U10509 ( .IN1(n10456), .IN2(n10455), .QN(n10486) );
  INVX0 U10510 ( .INP(n10457), .ZN(n10455) );
  NAND2X0 U10511 ( .IN1(n10342), .IN2(n9513), .QN(n10456) );
  NAND3X0 U10512 ( .IN1(n10488), .IN2(g2295), .IN3(n8892), .QN(n10483) );
  INVX0 U10513 ( .INP(n10485), .ZN(n10488) );
  NOR2X0 U10514 ( .IN1(n10463), .IN2(n5353), .QN(n10485) );
  NAND2X0 U10515 ( .IN1(n9001), .IN2(g2299), .QN(n10482) );
  NAND3X0 U10516 ( .IN1(n10489), .IN2(n10490), .IN3(n10491), .QN(g34000) );
  NAND2X0 U10517 ( .IN1(n9001), .IN2(g2246), .QN(n10491) );
  NAND2X0 U10518 ( .IN1(n10492), .IN2(n10493), .QN(n10490) );
  NAND2X0 U10519 ( .IN1(n10494), .IN2(g2165), .QN(n10489) );
  NAND2X0 U10520 ( .IN1(n10495), .IN2(n10496), .QN(g33999) );
  NAND2X0 U10521 ( .IN1(n10497), .IN2(g2227), .QN(n10496) );
  NAND2X0 U10522 ( .IN1(n10498), .IN2(n8914), .QN(n10497) );
  NAND2X0 U10523 ( .IN1(n10499), .IN2(g2241), .QN(n10498) );
  NAND2X0 U10524 ( .IN1(n10500), .IN2(n8914), .QN(n10495) );
  NAND2X0 U10525 ( .IN1(n10501), .IN2(n10502), .QN(n10500) );
  NAND2X0 U10526 ( .IN1(n10503), .IN2(n10504), .QN(n10502) );
  NAND2X0 U10527 ( .IN1(n10505), .IN2(n10506), .QN(n10504) );
  NAND2X0 U10528 ( .IN1(n8134), .IN2(n10507), .QN(n10506) );
  NAND2X0 U10529 ( .IN1(n10508), .IN2(g2241), .QN(n10501) );
  NAND2X0 U10530 ( .IN1(n10507), .IN2(n10509), .QN(n10508) );
  NAND2X0 U10531 ( .IN1(n10499), .IN2(g2153), .QN(n10509) );
  INVX0 U10532 ( .INP(n10503), .ZN(n10499) );
  NAND2X0 U10533 ( .IN1(n10510), .IN2(n10511), .QN(n10503) );
  NAND2X0 U10534 ( .IN1(n10512), .IN2(g1589), .QN(n10511) );
  NAND2X0 U10535 ( .IN1(n10513), .IN2(n10514), .QN(n10510) );
  NAND3X0 U10536 ( .IN1(n10515), .IN2(n10516), .IN3(n10517), .QN(g33998) );
  NAND2X0 U10537 ( .IN1(n10518), .IN2(n10492), .QN(n10517) );
  NAND3X0 U10538 ( .IN1(n10519), .IN2(g2181), .IN3(n8892), .QN(n10516) );
  INVX0 U10539 ( .INP(n10518), .ZN(n10519) );
  NOR2X0 U10540 ( .IN1(n10520), .IN2(n5538), .QN(n10518) );
  NAND2X0 U10541 ( .IN1(n9001), .IN2(g2169), .QN(n10515) );
  NAND3X0 U10542 ( .IN1(n10521), .IN2(n10522), .IN3(n10523), .QN(g33997) );
  NAND2X0 U10543 ( .IN1(n9001), .IN2(g2181), .QN(n10523) );
  NAND3X0 U10544 ( .IN1(n10492), .IN2(n5356), .IN3(n10524), .QN(n10522) );
  NAND2X0 U10545 ( .IN1(n10525), .IN2(n9352), .QN(n10521) );
  INVX0 U10546 ( .INP(n10526), .ZN(n10525) );
  NOR2X0 U10547 ( .IN1(n10527), .IN2(n10528), .QN(n10526) );
  NOR2X0 U10548 ( .IN1(n10524), .IN2(n8929), .QN(n10528) );
  NAND3X0 U10549 ( .IN1(n10529), .IN2(n10530), .IN3(n10531), .QN(g33996) );
  NAND2X0 U10550 ( .IN1(n10532), .IN2(n10492), .QN(n10531) );
  INVX0 U10551 ( .INP(n10533), .ZN(n10532) );
  NAND3X0 U10552 ( .IN1(n10533), .IN2(g2173), .IN3(n8892), .QN(n10530) );
  NAND3X0 U10553 ( .IN1(g2153), .IN2(g2227), .IN3(n10507), .QN(n10533) );
  NAND2X0 U10554 ( .IN1(n9001), .IN2(n9352), .QN(n10529) );
  NAND3X0 U10555 ( .IN1(n10534), .IN2(n10535), .IN3(n10536), .QN(g33995) );
  NAND2X0 U10556 ( .IN1(n10537), .IN2(n10492), .QN(n10536) );
  INVX0 U10557 ( .INP(n10538), .ZN(n10537) );
  NAND3X0 U10558 ( .IN1(n10538), .IN2(g2169), .IN3(n8892), .QN(n10535) );
  NAND2X0 U10559 ( .IN1(n10524), .IN2(n5538), .QN(n10538) );
  NAND2X0 U10560 ( .IN1(n9001), .IN2(g2161), .QN(n10534) );
  NAND3X0 U10561 ( .IN1(n10539), .IN2(n10540), .IN3(n10541), .QN(g33994) );
  NAND2X0 U10562 ( .IN1(n10542), .IN2(n10492), .QN(n10541) );
  NOR3X0 U10563 ( .IN1(n10543), .IN2(n10544), .IN3(n8925), .QN(n10492) );
  NOR2X0 U10564 ( .IN1(n10513), .IN2(n10512), .QN(n10544) );
  INVX0 U10565 ( .INP(n10514), .ZN(n10512) );
  NAND2X0 U10566 ( .IN1(n10342), .IN2(n9486), .QN(n10513) );
  INVX0 U10567 ( .INP(n10545), .ZN(n10342) );
  NAND2X0 U10568 ( .IN1(n10546), .IN2(g4180), .QN(n10545) );
  NOR2X0 U10569 ( .IN1(n10514), .IN2(g1585), .QN(n10543) );
  NAND3X0 U10570 ( .IN1(n10547), .IN2(g2161), .IN3(n8892), .QN(n10540) );
  INVX0 U10571 ( .INP(n10542), .ZN(n10547) );
  NOR2X0 U10572 ( .IN1(n10520), .IN2(n5356), .QN(n10542) );
  NAND2X0 U10573 ( .IN1(n9001), .IN2(g2165), .QN(n10539) );
  NAND3X0 U10574 ( .IN1(n10548), .IN2(n10549), .IN3(n10550), .QN(g33993) );
  NAND2X0 U10575 ( .IN1(n9002), .IN2(g2089), .QN(n10550) );
  NAND2X0 U10576 ( .IN1(n10551), .IN2(n10552), .QN(n10549) );
  NAND2X0 U10577 ( .IN1(n10553), .IN2(g2008), .QN(n10548) );
  NAND2X0 U10578 ( .IN1(n10554), .IN2(n10555), .QN(g33992) );
  NAND2X0 U10579 ( .IN1(n10556), .IN2(g2070), .QN(n10555) );
  NAND2X0 U10580 ( .IN1(n10557), .IN2(n8914), .QN(n10556) );
  NAND2X0 U10581 ( .IN1(n10558), .IN2(g2084), .QN(n10557) );
  NAND2X0 U10582 ( .IN1(n10559), .IN2(n8914), .QN(n10554) );
  NAND2X0 U10583 ( .IN1(n10560), .IN2(n10561), .QN(n10559) );
  NAND2X0 U10584 ( .IN1(n10562), .IN2(n10563), .QN(n10561) );
  NAND2X0 U10585 ( .IN1(n10564), .IN2(n10565), .QN(n10563) );
  NAND2X0 U10586 ( .IN1(n8129), .IN2(n10566), .QN(n10565) );
  NAND2X0 U10587 ( .IN1(n10567), .IN2(g2084), .QN(n10560) );
  NAND2X0 U10588 ( .IN1(n10566), .IN2(n10568), .QN(n10567) );
  NAND2X0 U10589 ( .IN1(n10558), .IN2(g1996), .QN(n10568) );
  INVX0 U10590 ( .INP(n10562), .ZN(n10558) );
  NAND2X0 U10591 ( .IN1(n10569), .IN2(n10570), .QN(n10562) );
  NAND2X0 U10592 ( .IN1(n5756), .IN2(n10571), .QN(n10570) );
  NAND2X0 U10593 ( .IN1(n10572), .IN2(n10573), .QN(n10569) );
  NAND2X0 U10594 ( .IN1(n10574), .IN2(n9623), .QN(n10572) );
  NAND3X0 U10595 ( .IN1(n10575), .IN2(n10576), .IN3(n10577), .QN(g33991) );
  NAND2X0 U10596 ( .IN1(n10578), .IN2(n10552), .QN(n10577) );
  NAND3X0 U10597 ( .IN1(n10579), .IN2(g2024), .IN3(n8891), .QN(n10576) );
  INVX0 U10598 ( .INP(n10578), .ZN(n10579) );
  NOR2X0 U10599 ( .IN1(n10580), .IN2(n5535), .QN(n10578) );
  NAND2X0 U10600 ( .IN1(n9002), .IN2(g2012), .QN(n10575) );
  NAND3X0 U10601 ( .IN1(n10581), .IN2(n10582), .IN3(n10583), .QN(g33990) );
  NAND2X0 U10602 ( .IN1(n9002), .IN2(g2024), .QN(n10583) );
  NAND3X0 U10603 ( .IN1(n10552), .IN2(n5355), .IN3(n10584), .QN(n10582) );
  NAND2X0 U10604 ( .IN1(n10585), .IN2(n9312), .QN(n10581) );
  INVX0 U10605 ( .INP(n10586), .ZN(n10585) );
  NOR2X0 U10606 ( .IN1(n10587), .IN2(n10588), .QN(n10586) );
  NOR2X0 U10607 ( .IN1(n10584), .IN2(n8928), .QN(n10588) );
  NAND3X0 U10608 ( .IN1(n10589), .IN2(n10590), .IN3(n10591), .QN(g33989) );
  NAND2X0 U10609 ( .IN1(n10592), .IN2(n10552), .QN(n10591) );
  INVX0 U10610 ( .INP(n10593), .ZN(n10592) );
  NAND3X0 U10611 ( .IN1(n10593), .IN2(g2016), .IN3(n8891), .QN(n10590) );
  NAND3X0 U10612 ( .IN1(g1996), .IN2(g2070), .IN3(n10566), .QN(n10593) );
  NAND2X0 U10613 ( .IN1(n9002), .IN2(n9312), .QN(n10589) );
  NAND3X0 U10614 ( .IN1(n10594), .IN2(n10595), .IN3(n10596), .QN(g33988) );
  NAND2X0 U10615 ( .IN1(n10597), .IN2(n10552), .QN(n10596) );
  INVX0 U10616 ( .INP(n10598), .ZN(n10597) );
  NAND3X0 U10617 ( .IN1(n10598), .IN2(g2012), .IN3(n8891), .QN(n10595) );
  NAND2X0 U10618 ( .IN1(n10584), .IN2(n5535), .QN(n10598) );
  NAND2X0 U10619 ( .IN1(n9002), .IN2(g2004), .QN(n10594) );
  NAND3X0 U10620 ( .IN1(n10599), .IN2(n10600), .IN3(n10601), .QN(g33987) );
  NAND2X0 U10621 ( .IN1(n10602), .IN2(n10552), .QN(n10601) );
  INVX0 U10622 ( .INP(n10603), .ZN(n10552) );
  NAND3X0 U10623 ( .IN1(n10604), .IN2(n10605), .IN3(n8891), .QN(n10603) );
  NAND2X0 U10624 ( .IN1(n10571), .IN2(g30332), .QN(n10605) );
  INVX0 U10625 ( .INP(n10573), .ZN(n10571) );
  NAND3X0 U10626 ( .IN1(n10574), .IN2(n9623), .IN3(n10573), .QN(n10604) );
  NAND3X0 U10627 ( .IN1(n10606), .IN2(g2004), .IN3(n8891), .QN(n10600) );
  INVX0 U10628 ( .INP(n10602), .ZN(n10606) );
  NOR2X0 U10629 ( .IN1(n10580), .IN2(n5355), .QN(n10602) );
  NAND2X0 U10630 ( .IN1(n9002), .IN2(g2008), .QN(n10599) );
  NAND3X0 U10631 ( .IN1(n10607), .IN2(n10608), .IN3(n10609), .QN(g33986) );
  NAND2X0 U10632 ( .IN1(n9002), .IN2(g1955), .QN(n10609) );
  NAND2X0 U10633 ( .IN1(n10610), .IN2(n10611), .QN(n10608) );
  NAND2X0 U10634 ( .IN1(n10612), .IN2(g1874), .QN(n10607) );
  NAND2X0 U10635 ( .IN1(n10613), .IN2(n10614), .QN(g33985) );
  NAND2X0 U10636 ( .IN1(n10615), .IN2(g1936), .QN(n10614) );
  NAND2X0 U10637 ( .IN1(n10616), .IN2(n8914), .QN(n10615) );
  NAND2X0 U10638 ( .IN1(n10617), .IN2(g1950), .QN(n10616) );
  NAND2X0 U10639 ( .IN1(n10618), .IN2(n8914), .QN(n10613) );
  NAND2X0 U10640 ( .IN1(n10619), .IN2(n10620), .QN(n10618) );
  NAND2X0 U10641 ( .IN1(n10621), .IN2(n10622), .QN(n10620) );
  NAND2X0 U10642 ( .IN1(n10623), .IN2(n10624), .QN(n10622) );
  NAND2X0 U10643 ( .IN1(n8133), .IN2(n10625), .QN(n10624) );
  NAND2X0 U10644 ( .IN1(n10626), .IN2(g1950), .QN(n10619) );
  NAND2X0 U10645 ( .IN1(n10625), .IN2(n10627), .QN(n10626) );
  NAND2X0 U10646 ( .IN1(test_so8), .IN2(n10617), .QN(n10627) );
  INVX0 U10647 ( .INP(n10621), .ZN(n10617) );
  NAND2X0 U10648 ( .IN1(n10628), .IN2(n10629), .QN(n10621) );
  NAND2X0 U10649 ( .IN1(n10630), .IN2(g1246), .QN(n10629) );
  NAND2X0 U10650 ( .IN1(n10631), .IN2(n10632), .QN(n10628) );
  NAND3X0 U10651 ( .IN1(n10633), .IN2(n10634), .IN3(n10635), .QN(g33984) );
  NAND2X0 U10652 ( .IN1(n10636), .IN2(n10610), .QN(n10635) );
  INVX0 U10653 ( .INP(n10637), .ZN(n10636) );
  NAND3X0 U10654 ( .IN1(n10637), .IN2(g1890), .IN3(n8891), .QN(n10634) );
  NAND2X0 U10655 ( .IN1(n10638), .IN2(n10625), .QN(n10637) );
  NAND2X0 U10656 ( .IN1(n9003), .IN2(g1878), .QN(n10633) );
  NAND3X0 U10657 ( .IN1(n10639), .IN2(n10640), .IN3(n10641), .QN(g33983) );
  NAND2X0 U10658 ( .IN1(n10642), .IN2(n10610), .QN(n10641) );
  INVX0 U10659 ( .INP(n10643), .ZN(n10642) );
  NAND3X0 U10660 ( .IN1(n10643), .IN2(n9280), .IN3(n8891), .QN(n10640) );
  NAND2X0 U10661 ( .IN1(n10644), .IN2(n8586), .QN(n10643) );
  NAND2X0 U10662 ( .IN1(n9003), .IN2(g1890), .QN(n10639) );
  NAND3X0 U10663 ( .IN1(n10645), .IN2(n10646), .IN3(n10647), .QN(g33982) );
  NAND2X0 U10664 ( .IN1(n10648), .IN2(n10610), .QN(n10647) );
  INVX0 U10665 ( .INP(n10649), .ZN(n10648) );
  NAND3X0 U10666 ( .IN1(n10649), .IN2(g1882), .IN3(n8891), .QN(n10646) );
  NAND2X0 U10667 ( .IN1(n10650), .IN2(g1936), .QN(n10649) );
  NAND2X0 U10668 ( .IN1(n9003), .IN2(n9280), .QN(n10645) );
  NAND3X0 U10669 ( .IN1(n10651), .IN2(n10652), .IN3(n10653), .QN(g33981) );
  NAND2X0 U10670 ( .IN1(n10654), .IN2(n10610), .QN(n10653) );
  INVX0 U10671 ( .INP(n10655), .ZN(n10654) );
  NAND3X0 U10672 ( .IN1(n10655), .IN2(g1878), .IN3(n8890), .QN(n10652) );
  NAND2X0 U10673 ( .IN1(n10644), .IN2(n5534), .QN(n10655) );
  NAND2X0 U10674 ( .IN1(n9003), .IN2(g1870), .QN(n10651) );
  NAND3X0 U10675 ( .IN1(n10656), .IN2(n10657), .IN3(n10658), .QN(g33980) );
  NAND2X0 U10676 ( .IN1(n10659), .IN2(n10610), .QN(n10658) );
  NOR3X0 U10677 ( .IN1(n10660), .IN2(n10661), .IN3(n8924), .QN(n10610) );
  NOR2X0 U10678 ( .IN1(n10631), .IN2(n10630), .QN(n10661) );
  INVX0 U10679 ( .INP(n10632), .ZN(n10630) );
  NAND2X0 U10680 ( .IN1(n10574), .IN2(n9559), .QN(n10631) );
  NOR2X0 U10681 ( .IN1(g30332), .IN2(n10632), .QN(n10660) );
  INVX0 U10682 ( .INP(n10662), .ZN(n10659) );
  NAND3X0 U10683 ( .IN1(n10662), .IN2(g1870), .IN3(n8890), .QN(n10657) );
  NAND2X0 U10684 ( .IN1(n10650), .IN2(n5503), .QN(n10662) );
  NAND2X0 U10685 ( .IN1(n9003), .IN2(g1874), .QN(n10656) );
  NAND3X0 U10686 ( .IN1(n10663), .IN2(n10664), .IN3(n10665), .QN(g33979) );
  NAND2X0 U10687 ( .IN1(n9003), .IN2(g1821), .QN(n10665) );
  NAND2X0 U10688 ( .IN1(n10666), .IN2(n10667), .QN(n10664) );
  NAND2X0 U10689 ( .IN1(n10668), .IN2(g1740), .QN(n10663) );
  NAND2X0 U10690 ( .IN1(n10669), .IN2(n10670), .QN(g33978) );
  NAND2X0 U10691 ( .IN1(n10671), .IN2(g1802), .QN(n10670) );
  NAND2X0 U10692 ( .IN1(n10672), .IN2(n8915), .QN(n10671) );
  NAND2X0 U10693 ( .IN1(n10673), .IN2(g1816), .QN(n10672) );
  NAND2X0 U10694 ( .IN1(n10674), .IN2(n8915), .QN(n10669) );
  NAND2X0 U10695 ( .IN1(n10675), .IN2(n10676), .QN(n10674) );
  NAND2X0 U10696 ( .IN1(n10677), .IN2(n10678), .QN(n10676) );
  NAND2X0 U10697 ( .IN1(n10679), .IN2(n10680), .QN(n10678) );
  NAND2X0 U10698 ( .IN1(n8070), .IN2(n10681), .QN(n10680) );
  NAND2X0 U10699 ( .IN1(n10682), .IN2(g1816), .QN(n10675) );
  NAND2X0 U10700 ( .IN1(n10681), .IN2(n10683), .QN(n10682) );
  NAND2X0 U10701 ( .IN1(n10673), .IN2(g1728), .QN(n10683) );
  INVX0 U10702 ( .INP(n10677), .ZN(n10673) );
  NAND2X0 U10703 ( .IN1(n10684), .IN2(n10685), .QN(n10677) );
  NAND2X0 U10704 ( .IN1(n10686), .IN2(n5756), .QN(n10685) );
  NAND2X0 U10705 ( .IN1(n10687), .IN2(n10688), .QN(n10684) );
  NAND3X0 U10706 ( .IN1(n10689), .IN2(n10690), .IN3(n10691), .QN(g33977) );
  NAND2X0 U10707 ( .IN1(n10692), .IN2(n10666), .QN(n10691) );
  NAND3X0 U10708 ( .IN1(n10693), .IN2(g1756), .IN3(n8890), .QN(n10690) );
  INVX0 U10709 ( .INP(n10692), .ZN(n10693) );
  NOR2X0 U10710 ( .IN1(n10694), .IN2(n5536), .QN(n10692) );
  NAND2X0 U10711 ( .IN1(n9003), .IN2(g1744), .QN(n10689) );
  NAND3X0 U10712 ( .IN1(n10695), .IN2(n10696), .IN3(n10697), .QN(g33976) );
  NAND2X0 U10713 ( .IN1(n9004), .IN2(g1756), .QN(n10697) );
  NAND3X0 U10714 ( .IN1(n10666), .IN2(n5352), .IN3(n10698), .QN(n10696) );
  NAND2X0 U10715 ( .IN1(n10699), .IN2(g1752), .QN(n10695) );
  INVX0 U10716 ( .INP(n10700), .ZN(n10699) );
  NOR2X0 U10717 ( .IN1(n10701), .IN2(n10702), .QN(n10700) );
  NOR2X0 U10718 ( .IN1(n10698), .IN2(n8930), .QN(n10702) );
  NAND3X0 U10719 ( .IN1(n10703), .IN2(n10704), .IN3(n10705), .QN(g33975) );
  NAND2X0 U10720 ( .IN1(n10706), .IN2(n10666), .QN(n10705) );
  INVX0 U10721 ( .INP(n10707), .ZN(n10706) );
  NAND3X0 U10722 ( .IN1(n10707), .IN2(g1748), .IN3(n8890), .QN(n10704) );
  NAND3X0 U10723 ( .IN1(g1728), .IN2(g1802), .IN3(n10681), .QN(n10707) );
  NAND2X0 U10724 ( .IN1(n9004), .IN2(g1752), .QN(n10703) );
  NAND3X0 U10725 ( .IN1(n10708), .IN2(n10709), .IN3(n10710), .QN(g33974) );
  NAND2X0 U10726 ( .IN1(n10711), .IN2(n10666), .QN(n10710) );
  INVX0 U10727 ( .INP(n10712), .ZN(n10711) );
  NAND3X0 U10728 ( .IN1(n10712), .IN2(g1744), .IN3(n8890), .QN(n10709) );
  NAND2X0 U10729 ( .IN1(n10698), .IN2(n5536), .QN(n10712) );
  NAND2X0 U10730 ( .IN1(n9004), .IN2(g1736), .QN(n10708) );
  NAND3X0 U10731 ( .IN1(n10713), .IN2(n10714), .IN3(n10715), .QN(g33973) );
  NAND2X0 U10732 ( .IN1(n10716), .IN2(n10666), .QN(n10715) );
  NOR3X0 U10733 ( .IN1(n10717), .IN2(n10718), .IN3(n8924), .QN(n10666) );
  NOR2X0 U10734 ( .IN1(n10688), .IN2(n5526), .QN(n10718) );
  NOR2X0 U10735 ( .IN1(n10687), .IN2(n10686), .QN(n10717) );
  INVX0 U10736 ( .INP(n10688), .ZN(n10686) );
  NAND2X0 U10737 ( .IN1(n10574), .IN2(n9514), .QN(n10687) );
  NAND3X0 U10738 ( .IN1(n10719), .IN2(g1736), .IN3(n8890), .QN(n10714) );
  INVX0 U10739 ( .INP(n10716), .ZN(n10719) );
  NOR2X0 U10740 ( .IN1(n10694), .IN2(n5352), .QN(n10716) );
  NAND2X0 U10741 ( .IN1(n9004), .IN2(g1740), .QN(n10713) );
  NAND3X0 U10742 ( .IN1(n10720), .IN2(n10721), .IN3(n10722), .QN(g33972) );
  NAND2X0 U10743 ( .IN1(n9004), .IN2(g1687), .QN(n10722) );
  INVX0 U10744 ( .INP(n10723), .ZN(n10721) );
  NOR2X0 U10745 ( .IN1(n10724), .IN2(n10725), .QN(n10723) );
  NAND2X0 U10746 ( .IN1(n10726), .IN2(g1604), .QN(n10720) );
  NAND2X0 U10747 ( .IN1(n10727), .IN2(n10728), .QN(g33971) );
  NAND2X0 U10748 ( .IN1(n10729), .IN2(g1668), .QN(n10728) );
  NAND2X0 U10749 ( .IN1(n10730), .IN2(n8915), .QN(n10729) );
  NAND2X0 U10750 ( .IN1(n10731), .IN2(g1682), .QN(n10730) );
  NAND2X0 U10751 ( .IN1(n10732), .IN2(n8915), .QN(n10727) );
  NAND2X0 U10752 ( .IN1(n10733), .IN2(n10734), .QN(n10732) );
  NAND2X0 U10753 ( .IN1(n10735), .IN2(n10736), .QN(n10734) );
  NAND2X0 U10754 ( .IN1(n10724), .IN2(n10737), .QN(n10736) );
  NAND2X0 U10755 ( .IN1(n8135), .IN2(n10738), .QN(n10737) );
  NAND2X0 U10756 ( .IN1(n10739), .IN2(g1682), .QN(n10733) );
  NAND2X0 U10757 ( .IN1(n10738), .IN2(n10740), .QN(n10739) );
  NAND2X0 U10758 ( .IN1(n10731), .IN2(g1592), .QN(n10740) );
  INVX0 U10759 ( .INP(n10735), .ZN(n10731) );
  NAND2X0 U10760 ( .IN1(n10741), .IN2(n10742), .QN(n10735) );
  NAND2X0 U10761 ( .IN1(n10743), .IN2(g1246), .QN(n10742) );
  NAND2X0 U10762 ( .IN1(n10744), .IN2(n10745), .QN(n10741) );
  NAND2X0 U10763 ( .IN1(n10574), .IN2(n9487), .QN(n10744) );
  NAND3X0 U10764 ( .IN1(n10746), .IN2(n10747), .IN3(n10748), .QN(g33970) );
  INVX0 U10765 ( .INP(n10749), .ZN(n10748) );
  NOR2X0 U10766 ( .IN1(n10750), .IN2(n10725), .QN(n10749) );
  NAND3X0 U10767 ( .IN1(n10750), .IN2(g1620), .IN3(n8890), .QN(n10747) );
  NAND2X0 U10768 ( .IN1(g25259), .IN2(n10738), .QN(n10750) );
  NAND2X0 U10769 ( .IN1(n9004), .IN2(g1608), .QN(n10746) );
  NAND3X0 U10770 ( .IN1(n10751), .IN2(n10752), .IN3(n10753), .QN(g33969) );
  INVX0 U10771 ( .INP(n10754), .ZN(n10753) );
  NOR2X0 U10772 ( .IN1(n10755), .IN2(n10725), .QN(n10754) );
  NAND3X0 U10773 ( .IN1(n10755), .IN2(n9303), .IN3(n8890), .QN(n10752) );
  NAND2X0 U10774 ( .IN1(n10756), .IN2(n5362), .QN(n10755) );
  NAND2X0 U10775 ( .IN1(n9005), .IN2(g1620), .QN(n10751) );
  NAND3X0 U10776 ( .IN1(n10757), .IN2(n10758), .IN3(n10759), .QN(g33968) );
  INVX0 U10777 ( .INP(n10760), .ZN(n10759) );
  NOR2X0 U10778 ( .IN1(n10761), .IN2(n10725), .QN(n10760) );
  NAND3X0 U10779 ( .IN1(n10761), .IN2(g1612), .IN3(n8889), .QN(n10758) );
  NAND2X0 U10780 ( .IN1(n10762), .IN2(g1668), .QN(n10761) );
  NAND2X0 U10781 ( .IN1(n9005), .IN2(n9303), .QN(n10757) );
  NAND3X0 U10782 ( .IN1(n10763), .IN2(n10764), .IN3(n10765), .QN(g33967) );
  INVX0 U10783 ( .INP(n10766), .ZN(n10765) );
  NOR2X0 U10784 ( .IN1(n10767), .IN2(n10725), .QN(n10766) );
  NAND3X0 U10785 ( .IN1(n10767), .IN2(g1608), .IN3(n8889), .QN(n10764) );
  NAND2X0 U10786 ( .IN1(n10756), .IN2(n5598), .QN(n10767) );
  NAND2X0 U10787 ( .IN1(n9005), .IN2(g1600), .QN(n10763) );
  NAND3X0 U10788 ( .IN1(n10768), .IN2(n10769), .IN3(n10770), .QN(g33966) );
  INVX0 U10789 ( .INP(n10771), .ZN(n10770) );
  NOR2X0 U10790 ( .IN1(n10772), .IN2(n10725), .QN(n10771) );
  NAND3X0 U10791 ( .IN1(n10773), .IN2(n10774), .IN3(n8889), .QN(n10725) );
  NAND3X0 U10792 ( .IN1(n10574), .IN2(n9487), .IN3(n10745), .QN(n10774) );
  INVX0 U10793 ( .INP(n10775), .ZN(n10574) );
  NAND2X0 U10794 ( .IN1(n10776), .IN2(g4180), .QN(n10775) );
  NAND2X0 U10795 ( .IN1(n10743), .IN2(n5526), .QN(n10773) );
  INVX0 U10796 ( .INP(n10745), .ZN(n10743) );
  NAND3X0 U10797 ( .IN1(n10772), .IN2(g1600), .IN3(n8889), .QN(n10769) );
  NAND2X0 U10798 ( .IN1(n10762), .IN2(n5549), .QN(n10772) );
  NAND2X0 U10799 ( .IN1(n9005), .IN2(g1604), .QN(n10768) );
  NAND3X0 U10800 ( .IN1(n10777), .IN2(n10778), .IN3(n10779), .QN(g33965) );
  NAND2X0 U10801 ( .IN1(n9005), .IN2(g763), .QN(n10779) );
  NAND3X0 U10802 ( .IN1(n2404), .IN2(n10780), .IN3(g767), .QN(n10778) );
  INVX0 U10803 ( .INP(n2704), .ZN(n10780) );
  NAND2X0 U10804 ( .IN1(n2704), .IN2(n5333), .QN(n10777) );
  NAND3X0 U10805 ( .IN1(n10781), .IN2(n10782), .IN3(n10783), .QN(g33964) );
  NAND2X0 U10806 ( .IN1(n9005), .IN2(g595), .QN(n10783) );
  NAND3X0 U10807 ( .IN1(n2421), .IN2(n10784), .IN3(g599), .QN(n10782) );
  INVX0 U10808 ( .INP(n2706), .ZN(n10784) );
  NAND2X0 U10809 ( .IN1(n2706), .IN2(n5550), .QN(n10781) );
  NAND2X0 U10810 ( .IN1(n10785), .IN2(n10786), .QN(g33963) );
  NAND2X0 U10811 ( .IN1(n9005), .IN2(g29215), .QN(n10786) );
  NAND3X0 U10812 ( .IN1(n10787), .IN2(n10788), .IN3(n8889), .QN(n10785) );
  NAND3X0 U10813 ( .IN1(n10789), .IN2(n10790), .IN3(n10791), .QN(n10788) );
  NAND2X0 U10814 ( .IN1(g72), .IN2(g262), .QN(n10791) );
  NAND2X0 U10815 ( .IN1(n10792), .IN2(g269), .QN(n10789) );
  NAND2X0 U10816 ( .IN1(g73), .IN2(n10793), .QN(n10787) );
  NAND2X0 U10817 ( .IN1(n10792), .IN2(g255), .QN(n10793) );
  NAND2X0 U10818 ( .IN1(n10794), .IN2(n10795), .QN(g33962) );
  NAND2X0 U10819 ( .IN1(n9006), .IN2(g479), .QN(n10795) );
  NAND3X0 U10820 ( .IN1(n10796), .IN2(n10797), .IN3(n8889), .QN(n10794) );
  NAND3X0 U10821 ( .IN1(n10798), .IN2(n10790), .IN3(n10799), .QN(n10797) );
  NAND2X0 U10822 ( .IN1(g72), .IN2(g239), .QN(n10799) );
  INVX0 U10823 ( .INP(g73), .ZN(n10790) );
  NAND2X0 U10824 ( .IN1(n10792), .IN2(g246), .QN(n10798) );
  NAND2X0 U10825 ( .IN1(g73), .IN2(n10800), .QN(n10796) );
  NAND2X0 U10826 ( .IN1(n10801), .IN2(n10802), .QN(n10800) );
  NAND2X0 U10827 ( .IN1(n5597), .IN2(g72), .QN(n10802) );
  INVX0 U10828 ( .INP(n10803), .ZN(n10801) );
  NOR2X0 U10829 ( .IN1(g232), .IN2(g72), .QN(n10803) );
  NAND3X0 U10830 ( .IN1(n10804), .IN2(n10805), .IN3(n10806), .QN(g33961) );
  NAND2X0 U10831 ( .IN1(n9006), .IN2(g294), .QN(n10806) );
  NAND3X0 U10832 ( .IN1(n8568), .IN2(n10807), .IN3(g298), .QN(n10805) );
  INVX0 U10833 ( .INP(n2989), .ZN(n10807) );
  NAND2X0 U10834 ( .IN1(n2989), .IN2(n5675), .QN(n10804) );
  NAND3X0 U10835 ( .IN1(n10808), .IN2(n10809), .IN3(n10810), .QN(g33960) );
  NAND2X0 U10836 ( .IN1(n9006), .IN2(g153), .QN(n10810) );
  NAND3X0 U10837 ( .IN1(n10217), .IN2(n10811), .IN3(g157), .QN(n10809) );
  INVX0 U10838 ( .INP(n2991), .ZN(n10811) );
  NAND2X0 U10839 ( .IN1(n2991), .IN2(n5678), .QN(n10808) );
  NAND4X0 U10840 ( .IN1(n2668), .IN2(n9298), .IN3(g8403), .IN4(g8283), .QN(
        g33935) );
  INVX0 U10841 ( .INP(g34649), .ZN(n9298) );
  NAND4X0 U10842 ( .IN1(n10812), .IN2(n10813), .IN3(n10814), .IN4(n10815), 
        .QN(g34649) );
  NAND2X0 U10843 ( .IN1(n9292), .IN2(g4888), .QN(n10815) );
  NAND2X0 U10844 ( .IN1(n9293), .IN2(g4955), .QN(n10814) );
  NAND2X0 U10845 ( .IN1(n9296), .IN2(g4944), .QN(n10813) );
  NAND2X0 U10846 ( .IN1(n9297), .IN2(g4933), .QN(n10812) );
  NAND3X0 U10847 ( .IN1(n2668), .IN2(g4507), .IN3(n5541), .QN(g33874) );
  NAND4X0 U10848 ( .IN1(n9197), .IN2(n10085), .IN3(n9315), .IN4(n9316), .QN(
        g33659) );
  XNOR2X1 U10849 ( .IN1(g4104), .IN2(g73), .Q(n9316) );
  XNOR2X1 U10850 ( .IN1(g4108), .IN2(g72), .Q(n9315) );
  INVX0 U10851 ( .INP(n10081), .ZN(n10085) );
  NAND2X0 U10852 ( .IN1(g113), .IN2(n2668), .QN(n10081) );
  INVX0 U10853 ( .INP(n10816), .ZN(n9197) );
  NAND2X0 U10854 ( .IN1(n10817), .IN2(n10818), .QN(n10816) );
  NAND2X0 U10855 ( .IN1(n5350), .IN2(n10819), .QN(n10818) );
  NAND3X0 U10856 ( .IN1(n10820), .IN2(n10821), .IN3(n10822), .QN(n10819) );
  NAND2X0 U10857 ( .IN1(n10823), .IN2(n10824), .QN(n10822) );
  NAND3X0 U10858 ( .IN1(n10825), .IN2(n10826), .IN3(g4093), .QN(n10821) );
  NAND2X0 U10859 ( .IN1(n5480), .IN2(n10827), .QN(n10826) );
  NAND2X0 U10860 ( .IN1(n10828), .IN2(g4087), .QN(n10825) );
  NAND2X0 U10861 ( .IN1(g32975), .IN2(n10829), .QN(n10820) );
  NAND2X0 U10862 ( .IN1(n10830), .IN2(g4098), .QN(n10817) );
  NAND3X0 U10863 ( .IN1(n10831), .IN2(n10832), .IN3(n10833), .QN(n10830) );
  NAND2X0 U10864 ( .IN1(n10834), .IN2(n10824), .QN(n10833) );
  NAND3X0 U10865 ( .IN1(n10835), .IN2(n10836), .IN3(g4093), .QN(n10832) );
  NAND2X0 U10866 ( .IN1(n5480), .IN2(n10837), .QN(n10836) );
  NAND2X0 U10867 ( .IN1(n10838), .IN2(g4087), .QN(n10835) );
  NAND2X0 U10868 ( .IN1(n10839), .IN2(n10829), .QN(n10831) );
  NAND4X0 U10869 ( .IN1(n2668), .IN2(n9258), .IN3(g8353), .IN4(g8235), .QN(
        g33636) );
  INVX0 U10870 ( .INP(g34657), .ZN(n9258) );
  NAND4X0 U10871 ( .IN1(n10840), .IN2(n10841), .IN3(n10842), .IN4(n10843), 
        .QN(g34657) );
  NAND2X0 U10872 ( .IN1(n9253), .IN2(g4754), .QN(n10843) );
  NAND2X0 U10873 ( .IN1(n9254), .IN2(g4743), .QN(n10842) );
  NAND2X0 U10874 ( .IN1(n9256), .IN2(g4765), .QN(n10841) );
  NAND2X0 U10875 ( .IN1(n9257), .IN2(g4698), .QN(n10840) );
  NAND2X0 U10876 ( .IN1(n10844), .IN2(n10845), .QN(n2668) );
  NAND2X0 U10877 ( .IN1(g99), .IN2(g37), .QN(n10845) );
  NAND3X0 U10878 ( .IN1(n10846), .IN2(n10847), .IN3(n10848), .QN(g33627) );
  NAND3X0 U10879 ( .IN1(n10849), .IN2(n10850), .IN3(n9217), .QN(n10848) );
  NAND2X0 U10880 ( .IN1(n9006), .IN2(g6741), .QN(n10847) );
  NAND2X0 U10881 ( .IN1(n10851), .IN2(n8915), .QN(n10846) );
  NAND2X0 U10882 ( .IN1(n10852), .IN2(n10853), .QN(n10851) );
  NAND2X0 U10883 ( .IN1(n8575), .IN2(g6682), .QN(n10853) );
  NAND2X0 U10884 ( .IN1(n9214), .IN2(n10849), .QN(n10852) );
  NAND3X0 U10885 ( .IN1(n10854), .IN2(n10855), .IN3(n10856), .QN(g33626) );
  NAND2X0 U10886 ( .IN1(n10857), .IN2(g6741), .QN(n10856) );
  NAND4X0 U10887 ( .IN1(n10849), .IN2(n10850), .IN3(n5398), .IN4(n8901), .QN(
        n10855) );
  NAND2X0 U10888 ( .IN1(n10858), .IN2(n9750), .QN(n10849) );
  NAND2X0 U10889 ( .IN1(n9006), .IN2(g6736), .QN(n10854) );
  NAND3X0 U10890 ( .IN1(n10859), .IN2(n10860), .IN3(n10861), .QN(g33625) );
  NAND3X0 U10891 ( .IN1(n10862), .IN2(n10863), .IN3(n10864), .QN(n10861) );
  NAND2X0 U10892 ( .IN1(n9006), .IN2(g6395), .QN(n10860) );
  NAND2X0 U10893 ( .IN1(n10865), .IN2(n8915), .QN(n10859) );
  NAND2X0 U10894 ( .IN1(n10866), .IN2(n10867), .QN(n10865) );
  NAND2X0 U10895 ( .IN1(n10868), .IN2(g6336), .QN(n10867) );
  NAND2X0 U10896 ( .IN1(n10869), .IN2(n10863), .QN(n10866) );
  NAND3X0 U10897 ( .IN1(n10870), .IN2(n10871), .IN3(n10872), .QN(g33624) );
  NAND2X0 U10898 ( .IN1(n10873), .IN2(g6395), .QN(n10872) );
  NAND4X0 U10899 ( .IN1(n10862), .IN2(n10863), .IN3(n5396), .IN4(n8902), .QN(
        n10871) );
  NAND2X0 U10900 ( .IN1(n10874), .IN2(n9753), .QN(n10863) );
  NAND2X0 U10901 ( .IN1(n9006), .IN2(g6390), .QN(n10870) );
  NAND3X0 U10902 ( .IN1(n10875), .IN2(n10876), .IN3(n10877), .QN(g33623) );
  NAND3X0 U10903 ( .IN1(n10878), .IN2(n10879), .IN3(n10880), .QN(n10877) );
  NAND2X0 U10904 ( .IN1(test_so57), .IN2(n9053), .QN(n10876) );
  NAND2X0 U10905 ( .IN1(n10881), .IN2(n8915), .QN(n10875) );
  NAND2X0 U10906 ( .IN1(n10882), .IN2(n10883), .QN(n10881) );
  NAND2X0 U10907 ( .IN1(n10884), .IN2(g5990), .QN(n10883) );
  NAND2X0 U10908 ( .IN1(n10885), .IN2(n10879), .QN(n10882) );
  NAND3X0 U10909 ( .IN1(n10886), .IN2(n10887), .IN3(n10888), .QN(g33622) );
  NAND2X0 U10910 ( .IN1(n10889), .IN2(test_so57), .QN(n10888) );
  NAND4X0 U10911 ( .IN1(n10879), .IN2(n8597), .IN3(n10878), .IN4(n8900), .QN(
        n10887) );
  NAND2X0 U10912 ( .IN1(n10890), .IN2(n9753), .QN(n10879) );
  NAND2X0 U10913 ( .IN1(test_so50), .IN2(n9053), .QN(n10886) );
  NAND3X0 U10914 ( .IN1(n10891), .IN2(n10892), .IN3(n10893), .QN(g33621) );
  NAND3X0 U10915 ( .IN1(n10894), .IN2(n10895), .IN3(n10896), .QN(n10893) );
  NAND2X0 U10916 ( .IN1(n9007), .IN2(g5703), .QN(n10892) );
  NAND2X0 U10917 ( .IN1(n10897), .IN2(n8915), .QN(n10891) );
  NAND2X0 U10918 ( .IN1(n10898), .IN2(n10899), .QN(n10897) );
  NAND2X0 U10919 ( .IN1(n10900), .IN2(g5644), .QN(n10899) );
  NAND2X0 U10920 ( .IN1(n10901), .IN2(n10895), .QN(n10898) );
  NAND3X0 U10921 ( .IN1(n10902), .IN2(n10903), .IN3(n10904), .QN(g33620) );
  NAND2X0 U10922 ( .IN1(n10905), .IN2(g5703), .QN(n10904) );
  NAND4X0 U10923 ( .IN1(n10894), .IN2(n10895), .IN3(n5397), .IN4(n8900), .QN(
        n10903) );
  NAND2X0 U10924 ( .IN1(n10906), .IN2(n9753), .QN(n10895) );
  NAND2X0 U10925 ( .IN1(n9007), .IN2(g5698), .QN(n10902) );
  NAND3X0 U10926 ( .IN1(n10907), .IN2(n10908), .IN3(n10909), .QN(g33619) );
  NAND3X0 U10927 ( .IN1(n10910), .IN2(g33959), .IN3(n9209), .QN(n10909) );
  NAND2X0 U10928 ( .IN1(n9007), .IN2(g5357), .QN(n10908) );
  NAND2X0 U10929 ( .IN1(n10911), .IN2(n8915), .QN(n10907) );
  NAND2X0 U10930 ( .IN1(n10912), .IN2(n10913), .QN(n10911) );
  NAND2X0 U10931 ( .IN1(n8570), .IN2(g5297), .QN(n10913) );
  NAND2X0 U10932 ( .IN1(n9207), .IN2(n10910), .QN(n10912) );
  NAND3X0 U10933 ( .IN1(n10914), .IN2(n10915), .IN3(n10916), .QN(g33618) );
  NAND2X0 U10934 ( .IN1(n10917), .IN2(g5357), .QN(n10916) );
  NAND4X0 U10935 ( .IN1(n10910), .IN2(g33959), .IN3(n5393), .IN4(n8901), .QN(
        n10915) );
  NAND2X0 U10936 ( .IN1(n10858), .IN2(n9753), .QN(n10910) );
  NOR2X0 U10937 ( .IN1(g4311), .IN2(n10918), .QN(n9753) );
  NOR2X0 U10938 ( .IN1(n10919), .IN2(test_so81), .QN(n10858) );
  NAND2X0 U10939 ( .IN1(n9007), .IN2(g5352), .QN(n10914) );
  NAND3X0 U10940 ( .IN1(n10920), .IN2(n10298), .IN3(n10921), .QN(g33617) );
  NAND2X0 U10941 ( .IN1(n10922), .IN2(g4552), .QN(n10921) );
  NAND4X0 U10942 ( .IN1(n10923), .IN2(n10924), .IN3(n10925), .IN4(n10298), 
        .QN(g33616) );
  NAND2X0 U10943 ( .IN1(n10926), .IN2(g4512), .QN(n10924) );
  NAND2X0 U10944 ( .IN1(n9007), .IN2(g4515), .QN(n10923) );
  NAND2X0 U10945 ( .IN1(n3064), .IN2(n10927), .QN(g33615) );
  NAND2X0 U10946 ( .IN1(n10928), .IN2(g4108), .QN(n10927) );
  NAND2X0 U10947 ( .IN1(n10929), .IN2(n8915), .QN(n10928) );
  NAND2X0 U10948 ( .IN1(n9334), .IN2(n8312), .QN(n10929) );
  NAND3X0 U10949 ( .IN1(n10930), .IN2(n10931), .IN3(n10932), .QN(g33614) );
  NAND3X0 U10950 ( .IN1(n10933), .IN2(n10934), .IN3(n10935), .QN(n10932) );
  NAND2X0 U10951 ( .IN1(n9007), .IN2(g4054), .QN(n10931) );
  NAND2X0 U10952 ( .IN1(n10936), .IN2(n8915), .QN(n10930) );
  NAND2X0 U10953 ( .IN1(n10937), .IN2(n10938), .QN(n10936) );
  NAND2X0 U10954 ( .IN1(n10939), .IN2(g3990), .QN(n10938) );
  NAND2X0 U10955 ( .IN1(n10940), .IN2(n10934), .QN(n10937) );
  NAND3X0 U10956 ( .IN1(n10941), .IN2(n10942), .IN3(n10943), .QN(g33613) );
  NAND2X0 U10957 ( .IN1(n10944), .IN2(g4054), .QN(n10943) );
  NAND4X0 U10958 ( .IN1(n10933), .IN2(n10934), .IN3(n5395), .IN4(n8901), .QN(
        n10942) );
  NAND2X0 U10959 ( .IN1(n10874), .IN2(n9750), .QN(n10934) );
  NOR2X0 U10960 ( .IN1(n10945), .IN2(n8590), .QN(n10874) );
  NAND2X0 U10961 ( .IN1(n9007), .IN2(g4049), .QN(n10941) );
  NAND3X0 U10962 ( .IN1(n10946), .IN2(n10947), .IN3(n10948), .QN(g33612) );
  NAND3X0 U10963 ( .IN1(n10949), .IN2(n10950), .IN3(n10951), .QN(n10948) );
  NAND2X0 U10964 ( .IN1(n9008), .IN2(g3703), .QN(n10947) );
  NAND2X0 U10965 ( .IN1(n10952), .IN2(n8915), .QN(n10946) );
  NAND2X0 U10966 ( .IN1(n10953), .IN2(n10954), .QN(n10952) );
  NAND2X0 U10967 ( .IN1(n10955), .IN2(g3639), .QN(n10954) );
  NAND2X0 U10968 ( .IN1(n10956), .IN2(n10950), .QN(n10953) );
  NAND3X0 U10969 ( .IN1(n10957), .IN2(n10958), .IN3(n10959), .QN(g33611) );
  NAND2X0 U10970 ( .IN1(n10960), .IN2(g3703), .QN(n10959) );
  NAND4X0 U10971 ( .IN1(n10949), .IN2(n10950), .IN3(n5399), .IN4(n8901), .QN(
        n10958) );
  NAND2X0 U10972 ( .IN1(n10890), .IN2(n9750), .QN(n10950) );
  NOR2X0 U10973 ( .IN1(n10945), .IN2(test_so81), .QN(n10890) );
  INVX0 U10974 ( .INP(n3033), .ZN(n10945) );
  NAND2X0 U10975 ( .IN1(n9008), .IN2(g3698), .QN(n10957) );
  NAND2X0 U10976 ( .IN1(n10961), .IN2(n10962), .QN(g33610) );
  NAND2X0 U10977 ( .IN1(n9008), .IN2(g3352), .QN(n10962) );
  NAND2X0 U10978 ( .IN1(n10963), .IN2(n8915), .QN(n10961) );
  NAND2X0 U10979 ( .IN1(n10964), .IN2(n10965), .QN(n10963) );
  NAND2X0 U10980 ( .IN1(n10966), .IN2(g3288), .QN(n10965) );
  NAND3X0 U10981 ( .IN1(n10967), .IN2(n10968), .IN3(n10969), .QN(n10964) );
  NAND2X0 U10982 ( .IN1(n10970), .IN2(n10971), .QN(n10967) );
  NAND3X0 U10983 ( .IN1(n10972), .IN2(n10973), .IN3(n10974), .QN(g33609) );
  NAND2X0 U10984 ( .IN1(n10975), .IN2(g3352), .QN(n10974) );
  NAND4X0 U10985 ( .IN1(n5604), .IN2(n10968), .IN3(n10969), .IN4(n8901), .QN(
        n10973) );
  NAND2X0 U10986 ( .IN1(n10906), .IN2(n9750), .QN(n10968) );
  NOR2X0 U10987 ( .IN1(n10918), .IN2(n5323), .QN(n9750) );
  INVX0 U10988 ( .INP(n10976), .ZN(n10918) );
  NOR2X0 U10989 ( .IN1(n10977), .IN2(n9665), .QN(n10976) );
  XOR2X1 U10990 ( .IN1(g72), .IN2(g4322), .Q(n9665) );
  XOR2X1 U10991 ( .IN1(g4332), .IN2(g73), .Q(n10977) );
  NOR2X0 U10992 ( .IN1(n10919), .IN2(n8590), .QN(n10906) );
  INVX0 U10993 ( .INP(n3023), .ZN(n10919) );
  NAND2X0 U10994 ( .IN1(n9008), .IN2(g3347), .QN(n10972) );
  NAND4X0 U10995 ( .IN1(n10978), .IN2(n9200), .IN3(n10979), .IN4(n10980), .QN(
        g33608) );
  NAND3X0 U10996 ( .IN1(n10981), .IN2(g2759), .IN3(n8876), .QN(n10980) );
  NAND2X0 U10997 ( .IN1(test_so30), .IN2(n9051), .QN(n10979) );
  NAND2X0 U10998 ( .IN1(n10315), .IN2(n8051), .QN(n10978) );
  INVX0 U10999 ( .INP(n10981), .ZN(n10315) );
  NAND2X0 U11000 ( .IN1(n2790), .IN2(test_so30), .QN(n10981) );
  NAND3X0 U11001 ( .IN1(n10982), .IN2(n10983), .IN3(n10984), .QN(g33607) );
  NAND2X0 U11002 ( .IN1(n9008), .IN2(g2555), .QN(n10984) );
  NAND3X0 U11003 ( .IN1(n10985), .IN2(n10986), .IN3(n686), .QN(n10983) );
  NAND3X0 U11004 ( .IN1(g2629), .IN2(g112), .IN3(n5524), .QN(n10986) );
  NAND2X0 U11005 ( .IN1(n10987), .IN2(n10988), .QN(n10985) );
  NAND2X0 U11006 ( .IN1(n10101), .IN2(n10989), .QN(n10988) );
  NOR3X0 U11007 ( .IN1(n2726), .IN2(n5521), .IN3(g2599), .QN(n10101) );
  NAND2X0 U11008 ( .IN1(n10110), .IN2(n5519), .QN(n2726) );
  NAND2X0 U11009 ( .IN1(n3111), .IN2(n8915), .QN(n10987) );
  NAND2X0 U11010 ( .IN1(n10990), .IN2(g2606), .QN(n10982) );
  NAND2X0 U11011 ( .IN1(n10991), .IN2(n10992), .QN(n10990) );
  NAND2X0 U11012 ( .IN1(n8905), .IN2(n10993), .QN(n10992) );
  INVX0 U11013 ( .INP(n3105), .ZN(n10993) );
  NAND3X0 U11014 ( .IN1(n10994), .IN2(n10995), .IN3(n10996), .QN(g33606) );
  NAND2X0 U11015 ( .IN1(n10321), .IN2(g2675), .QN(n10996) );
  NAND3X0 U11016 ( .IN1(n5457), .IN2(n10319), .IN3(n8876), .QN(n10995) );
  NAND2X0 U11017 ( .IN1(n9008), .IN2(g2671), .QN(n10994) );
  NAND3X0 U11018 ( .IN1(n10997), .IN2(n10998), .IN3(n10999), .QN(g33605) );
  NAND2X0 U11019 ( .IN1(n10321), .IN2(g2671), .QN(n10999) );
  NAND2X0 U11020 ( .IN1(test_so48), .IN2(n11000), .QN(n10998) );
  NAND2X0 U11021 ( .IN1(n11001), .IN2(n8915), .QN(n11000) );
  NAND2X0 U11022 ( .IN1(n10319), .IN2(g2661), .QN(n11001) );
  NAND4X0 U11023 ( .IN1(n10319), .IN2(n8899), .IN3(n5418), .IN4(n8619), .QN(
        n10997) );
  INVX0 U11024 ( .INP(n10332), .ZN(n10319) );
  NAND2X0 U11025 ( .IN1(n11002), .IN2(n11003), .QN(g33604) );
  NAND2X0 U11026 ( .IN1(test_so48), .IN2(n10321), .QN(n11003) );
  NAND2X0 U11027 ( .IN1(n11004), .IN2(g2661), .QN(n11002) );
  NAND2X0 U11028 ( .IN1(n11005), .IN2(n11006), .QN(g33603) );
  NAND2X0 U11029 ( .IN1(n10321), .IN2(g2648), .QN(n11006) );
  INVX0 U11030 ( .INP(n11004), .ZN(n10321) );
  NAND2X0 U11031 ( .IN1(n11004), .IN2(g2643), .QN(n11005) );
  NAND2X0 U11032 ( .IN1(n10332), .IN2(n8915), .QN(n11004) );
  NAND3X0 U11033 ( .IN1(n5351), .IN2(n10334), .IN3(n5521), .QN(n10332) );
  NAND3X0 U11034 ( .IN1(n11007), .IN2(n11008), .IN3(n11009), .QN(g33602) );
  NAND2X0 U11035 ( .IN1(n10352), .IN2(n11010), .QN(n11009) );
  NOR2X0 U11036 ( .IN1(n5524), .IN2(n11011), .QN(n10352) );
  NAND2X0 U11037 ( .IN1(n9008), .IN2(g2599), .QN(n11008) );
  NAND3X0 U11038 ( .IN1(n11011), .IN2(g2629), .IN3(n8876), .QN(n11007) );
  NAND3X0 U11039 ( .IN1(n11012), .IN2(n11013), .IN3(n11014), .QN(g33601) );
  NAND3X0 U11040 ( .IN1(n10334), .IN2(n11010), .IN3(n10355), .QN(n11014) );
  NAND3X0 U11041 ( .IN1(n11011), .IN2(g2599), .IN3(n8875), .QN(n11013) );
  NAND2X0 U11042 ( .IN1(n9009), .IN2(g2606), .QN(n11012) );
  NAND2X0 U11043 ( .IN1(n11015), .IN2(n11016), .QN(g33600) );
  NAND4X0 U11044 ( .IN1(n5521), .IN2(n11017), .IN3(n8898), .IN4(n11010), .QN(
        n11016) );
  INVX0 U11045 ( .INP(n3111), .ZN(n11010) );
  NAND2X0 U11046 ( .IN1(n5351), .IN2(n10348), .QN(n11017) );
  NAND2X0 U11047 ( .IN1(n5524), .IN2(n10334), .QN(n10348) );
  INVX0 U11048 ( .INP(n11011), .ZN(n10334) );
  NAND2X0 U11049 ( .IN1(n10355), .IN2(n11011), .QN(n11015) );
  NOR2X0 U11050 ( .IN1(n10341), .IN2(n686), .QN(n11011) );
  NOR2X0 U11051 ( .IN1(n8444), .IN2(n11018), .QN(n686) );
  NOR3X0 U11052 ( .IN1(n11019), .IN2(test_so49), .IN3(g1514), .QN(n11018) );
  NAND3X0 U11053 ( .IN1(n10546), .IN2(n9621), .IN3(n11020), .QN(n10341) );
  NAND3X0 U11054 ( .IN1(g2689), .IN2(g2704), .IN3(g2697), .QN(n11020) );
  NAND2X0 U11055 ( .IN1(n2549), .IN2(g1300), .QN(n9621) );
  NOR2X0 U11056 ( .IN1(n8955), .IN2(n5351), .QN(n10355) );
  NAND3X0 U11057 ( .IN1(n11021), .IN2(n11022), .IN3(n11023), .QN(g33599) );
  NOR2X0 U11058 ( .IN1(n11024), .IN2(n11025), .QN(n11023) );
  NOR2X0 U11059 ( .IN1(n5619), .IN2(n11026), .QN(n11025) );
  NOR2X0 U11060 ( .IN1(n11027), .IN2(n11028), .QN(n11026) );
  NOR2X0 U11061 ( .IN1(n3125), .IN2(n8937), .QN(n11027) );
  INVX0 U11062 ( .INP(n3121), .ZN(n11024) );
  NAND4X0 U11063 ( .IN1(n3122), .IN2(n10404), .IN3(n11029), .IN4(n8185), .QN(
        n3121) );
  NOR2X0 U11064 ( .IN1(n2727), .IN2(n9218), .QN(n11029) );
  NAND2X0 U11065 ( .IN1(n10110), .IN2(g504), .QN(n2727) );
  INVX0 U11066 ( .INP(n11030), .ZN(n10110) );
  NAND2X0 U11067 ( .IN1(n3116), .IN2(g518), .QN(n11030) );
  NAND2X0 U11068 ( .IN1(test_so79), .IN2(n8963), .QN(n11022) );
  NAND4X0 U11069 ( .IN1(n3122), .IN2(n11031), .IN3(n3131), .IN4(n8901), .QN(
        n11021) );
  NAND2X0 U11070 ( .IN1(n10404), .IN2(g112), .QN(n11031) );
  INVX0 U11071 ( .INP(n10096), .ZN(n10404) );
  NAND2X0 U11072 ( .IN1(n5523), .IN2(g2495), .QN(n10096) );
  NAND3X0 U11073 ( .IN1(n11032), .IN2(n11033), .IN3(n11034), .QN(g33598) );
  NAND2X0 U11074 ( .IN1(n10380), .IN2(g2541), .QN(n11034) );
  NAND3X0 U11075 ( .IN1(n5461), .IN2(n10379), .IN3(n8875), .QN(n11033) );
  NAND2X0 U11076 ( .IN1(n9009), .IN2(g2537), .QN(n11032) );
  NAND3X0 U11077 ( .IN1(n11035), .IN2(n11036), .IN3(n11037), .QN(g33597) );
  NAND2X0 U11078 ( .IN1(n10380), .IN2(g2537), .QN(n11037) );
  NAND2X0 U11079 ( .IN1(n11038), .IN2(g2533), .QN(n11036) );
  NAND2X0 U11080 ( .IN1(n11039), .IN2(n8915), .QN(n11038) );
  NAND2X0 U11081 ( .IN1(n10379), .IN2(g2527), .QN(n11039) );
  NAND4X0 U11082 ( .IN1(n10379), .IN2(n8898), .IN3(n5420), .IN4(n5761), .QN(
        n11035) );
  INVX0 U11083 ( .INP(n10391), .ZN(n10379) );
  NAND2X0 U11084 ( .IN1(n11040), .IN2(n11041), .QN(g33596) );
  NAND2X0 U11085 ( .IN1(n10380), .IN2(g2533), .QN(n11041) );
  NAND2X0 U11086 ( .IN1(n11042), .IN2(g2527), .QN(n11040) );
  NAND2X0 U11087 ( .IN1(n11043), .IN2(n11044), .QN(g33595) );
  NAND2X0 U11088 ( .IN1(n10380), .IN2(g2514), .QN(n11044) );
  INVX0 U11089 ( .INP(n11042), .ZN(n10380) );
  NAND2X0 U11090 ( .IN1(n11042), .IN2(g2509), .QN(n11043) );
  NAND2X0 U11091 ( .IN1(n10391), .IN2(n8915), .QN(n11042) );
  NAND3X0 U11092 ( .IN1(n10393), .IN2(n8585), .IN3(n5522), .QN(n10391) );
  NAND3X0 U11093 ( .IN1(n11045), .IN2(n11046), .IN3(n11047), .QN(g33594) );
  NAND2X0 U11094 ( .IN1(n9009), .IN2(g2465), .QN(n11047) );
  NAND2X0 U11095 ( .IN1(n11048), .IN2(g2495), .QN(n11046) );
  NAND2X0 U11096 ( .IN1(n10413), .IN2(n11049), .QN(n11045) );
  NOR2X0 U11097 ( .IN1(n5523), .IN2(n11050), .QN(n10413) );
  NAND3X0 U11098 ( .IN1(n11051), .IN2(n11052), .IN3(n11053), .QN(g33593) );
  NAND2X0 U11099 ( .IN1(n11048), .IN2(g2465), .QN(n11053) );
  NAND2X0 U11100 ( .IN1(n9009), .IN2(g2472), .QN(n11052) );
  NAND3X0 U11101 ( .IN1(n10419), .IN2(n11049), .IN3(n8875), .QN(n11051) );
  NOR2X0 U11102 ( .IN1(n8585), .IN2(n11050), .QN(n10419) );
  NAND2X0 U11103 ( .IN1(n11054), .IN2(n11055), .QN(g33592) );
  NAND4X0 U11104 ( .IN1(n5522), .IN2(n11056), .IN3(n8898), .IN4(n11049), .QN(
        n11055) );
  INVX0 U11105 ( .INP(n3131), .ZN(n11049) );
  NAND2X0 U11106 ( .IN1(n8585), .IN2(n11057), .QN(n11056) );
  NAND2X0 U11107 ( .IN1(n5523), .IN2(n10393), .QN(n11057) );
  INVX0 U11108 ( .INP(n11050), .ZN(n10393) );
  NAND2X0 U11109 ( .IN1(n11048), .IN2(test_so79), .QN(n11054) );
  INVX0 U11110 ( .INP(n10406), .ZN(n11048) );
  NAND2X0 U11111 ( .IN1(n11050), .IN2(n8915), .QN(n10406) );
  NOR2X0 U11112 ( .IN1(n10400), .IN2(n3122), .QN(n11050) );
  NOR2X0 U11113 ( .IN1(n11058), .IN2(n8159), .QN(n3122) );
  NOR2X0 U11114 ( .IN1(n11059), .IN2(n11019), .QN(n11058) );
  NAND3X0 U11115 ( .IN1(n10546), .IN2(n9557), .IN3(n11060), .QN(n10400) );
  NAND3X0 U11116 ( .IN1(g2697), .IN2(g2689), .IN3(n5377), .QN(n11060) );
  NAND2X0 U11117 ( .IN1(n2549), .IN2(g1472), .QN(n9557) );
  NAND3X0 U11118 ( .IN1(n11061), .IN2(n11062), .IN3(n11063), .QN(g33591) );
  NAND2X0 U11119 ( .IN1(n9009), .IN2(g2287), .QN(n11063) );
  NAND3X0 U11120 ( .IN1(n11064), .IN2(n11065), .IN3(n3141), .QN(n11062) );
  NAND2X0 U11121 ( .IN1(n11066), .IN2(n11067), .QN(n11065) );
  NAND2X0 U11122 ( .IN1(n11068), .IN2(n8916), .QN(n11067) );
  INVX0 U11123 ( .INP(n11069), .ZN(n11068) );
  NAND3X0 U11124 ( .IN1(n10989), .IN2(n10111), .IN3(n10100), .QN(n11066) );
  NAND2X0 U11125 ( .IN1(n10100), .IN2(g112), .QN(n11064) );
  NOR2X0 U11126 ( .IN1(g2331), .IN2(n5537), .QN(n10100) );
  NAND2X0 U11127 ( .IN1(n11070), .IN2(g2338), .QN(n11061) );
  NAND2X0 U11128 ( .IN1(n10991), .IN2(n11071), .QN(n11070) );
  NAND2X0 U11129 ( .IN1(n8905), .IN2(n11072), .QN(n11071) );
  INVX0 U11130 ( .INP(n3145), .ZN(n11072) );
  NAND3X0 U11131 ( .IN1(n11073), .IN2(n11074), .IN3(n11075), .QN(g33590) );
  NAND2X0 U11132 ( .IN1(n10437), .IN2(g2407), .QN(n11075) );
  NAND3X0 U11133 ( .IN1(n5459), .IN2(n10436), .IN3(n8875), .QN(n11074) );
  NAND2X0 U11134 ( .IN1(test_so31), .IN2(n8958), .QN(n11073) );
  NAND3X0 U11135 ( .IN1(n11076), .IN2(n11077), .IN3(n11078), .QN(g33589) );
  NAND2X0 U11136 ( .IN1(test_so31), .IN2(n10437), .QN(n11078) );
  NAND2X0 U11137 ( .IN1(n11079), .IN2(g2399), .QN(n11077) );
  NAND2X0 U11138 ( .IN1(n11080), .IN2(n8916), .QN(n11079) );
  NAND2X0 U11139 ( .IN1(n10436), .IN2(g2393), .QN(n11080) );
  NAND4X0 U11140 ( .IN1(n10436), .IN2(n8899), .IN3(n5421), .IN4(n5762), .QN(
        n11076) );
  INVX0 U11141 ( .INP(n10448), .ZN(n10436) );
  NAND2X0 U11142 ( .IN1(n11081), .IN2(n11082), .QN(g33588) );
  NAND2X0 U11143 ( .IN1(n10437), .IN2(g2399), .QN(n11082) );
  NAND2X0 U11144 ( .IN1(n11083), .IN2(g2393), .QN(n11081) );
  NAND2X0 U11145 ( .IN1(n11084), .IN2(n11085), .QN(g33587) );
  NAND2X0 U11146 ( .IN1(n10437), .IN2(g2380), .QN(n11085) );
  INVX0 U11147 ( .INP(n11083), .ZN(n10437) );
  NAND2X0 U11148 ( .IN1(n11083), .IN2(g2375), .QN(n11084) );
  NAND2X0 U11149 ( .IN1(n10448), .IN2(n8916), .QN(n11083) );
  NAND3X0 U11150 ( .IN1(n5353), .IN2(n10450), .IN3(n5537), .QN(n10448) );
  NAND3X0 U11151 ( .IN1(n11086), .IN2(n11087), .IN3(n11088), .QN(g33586) );
  NAND2X0 U11152 ( .IN1(n10467), .IN2(n11069), .QN(n11088) );
  NOR2X0 U11153 ( .IN1(n5513), .IN2(n11089), .QN(n10467) );
  NAND2X0 U11154 ( .IN1(n9009), .IN2(g2331), .QN(n11087) );
  NAND3X0 U11155 ( .IN1(n11089), .IN2(g2361), .IN3(n8875), .QN(n11086) );
  NAND3X0 U11156 ( .IN1(n11090), .IN2(n11091), .IN3(n11092), .QN(g33585) );
  NAND3X0 U11157 ( .IN1(n11069), .IN2(n10450), .IN3(n10470), .QN(n11092) );
  NAND3X0 U11158 ( .IN1(n11089), .IN2(g2331), .IN3(n8874), .QN(n11091) );
  NAND2X0 U11159 ( .IN1(n9009), .IN2(g2338), .QN(n11090) );
  NAND2X0 U11160 ( .IN1(n11093), .IN2(n11094), .QN(g33584) );
  NAND2X0 U11161 ( .IN1(n10470), .IN2(n11089), .QN(n11094) );
  NOR2X0 U11162 ( .IN1(n8955), .IN2(n5353), .QN(n10470) );
  NAND4X0 U11163 ( .IN1(n5537), .IN2(n11095), .IN3(n11069), .IN4(n8901), .QN(
        n11093) );
  NAND2X0 U11164 ( .IN1(n3115), .IN2(n10111), .QN(n11069) );
  INVX0 U11165 ( .INP(n3146), .ZN(n10111) );
  NAND3X0 U11166 ( .IN1(n5287), .IN2(g504), .IN3(n3116), .QN(n3146) );
  NAND2X0 U11167 ( .IN1(n5353), .IN2(n10463), .QN(n11095) );
  NAND2X0 U11168 ( .IN1(n5513), .IN2(n10450), .QN(n10463) );
  INVX0 U11169 ( .INP(n11089), .ZN(n10450) );
  NOR2X0 U11170 ( .IN1(n10457), .IN2(n3141), .QN(n11089) );
  NOR2X0 U11171 ( .IN1(n11096), .IN2(n8160), .QN(n3141) );
  NOR2X0 U11172 ( .IN1(n11097), .IN2(n11019), .QN(n11096) );
  NAND3X0 U11173 ( .IN1(n10546), .IN2(n9513), .IN3(n11098), .QN(n10457) );
  NAND3X0 U11174 ( .IN1(g2689), .IN2(g2704), .IN3(n5308), .QN(n11098) );
  NAND2X0 U11175 ( .IN1(n2549), .IN2(g1448), .QN(n9513) );
  NAND3X0 U11176 ( .IN1(n11099), .IN2(n11100), .IN3(n11101), .QN(g33583) );
  NAND2X0 U11177 ( .IN1(n9010), .IN2(g2153), .QN(n11101) );
  NAND3X0 U11178 ( .IN1(n11102), .IN2(n11103), .IN3(n700), .QN(n11100) );
  NAND2X0 U11179 ( .IN1(n11104), .IN2(n11105), .QN(n11103) );
  NAND2X0 U11180 ( .IN1(n11106), .IN2(n8916), .QN(n11105) );
  INVX0 U11181 ( .INP(n11107), .ZN(n11106) );
  NAND3X0 U11182 ( .IN1(n10989), .IN2(n10106), .IN3(n10105), .QN(n11104) );
  NAND2X0 U11183 ( .IN1(n10105), .IN2(g112), .QN(n11102) );
  NOR2X0 U11184 ( .IN1(g2197), .IN2(n5538), .QN(n10105) );
  NAND2X0 U11185 ( .IN1(n11108), .IN2(g2204), .QN(n11099) );
  INVX0 U11186 ( .INP(n11109), .ZN(n11108) );
  NOR2X0 U11187 ( .IN1(n11028), .IN2(n11110), .QN(n11109) );
  NOR2X0 U11188 ( .IN1(n8956), .IN2(n3164), .QN(n11110) );
  INVX0 U11189 ( .INP(n10991), .ZN(n11028) );
  NAND3X0 U11190 ( .IN1(n11111), .IN2(n11112), .IN3(n11113), .QN(g33582) );
  NAND2X0 U11191 ( .IN1(n10494), .IN2(g2273), .QN(n11113) );
  NAND3X0 U11192 ( .IN1(n5458), .IN2(n10493), .IN3(n8874), .QN(n11112) );
  NAND2X0 U11193 ( .IN1(n9010), .IN2(g2269), .QN(n11111) );
  NAND3X0 U11194 ( .IN1(n11114), .IN2(n11115), .IN3(n11116), .QN(g33581) );
  NAND2X0 U11195 ( .IN1(n10494), .IN2(g2269), .QN(n11116) );
  NAND2X0 U11196 ( .IN1(test_so62), .IN2(n11117), .QN(n11115) );
  NAND2X0 U11197 ( .IN1(n11118), .IN2(n8916), .QN(n11117) );
  NAND2X0 U11198 ( .IN1(n10493), .IN2(g2259), .QN(n11118) );
  NAND4X0 U11199 ( .IN1(n10493), .IN2(n8900), .IN3(n5419), .IN4(n8620), .QN(
        n11114) );
  INVX0 U11200 ( .INP(n10505), .ZN(n10493) );
  NAND2X0 U11201 ( .IN1(n11119), .IN2(n11120), .QN(g33580) );
  NAND2X0 U11202 ( .IN1(test_so62), .IN2(n10494), .QN(n11120) );
  NAND2X0 U11203 ( .IN1(n11121), .IN2(g2259), .QN(n11119) );
  NAND2X0 U11204 ( .IN1(n11122), .IN2(n11123), .QN(g33579) );
  NAND2X0 U11205 ( .IN1(n10494), .IN2(g2246), .QN(n11123) );
  INVX0 U11206 ( .INP(n11121), .ZN(n10494) );
  NAND2X0 U11207 ( .IN1(n11121), .IN2(g2241), .QN(n11122) );
  NAND2X0 U11208 ( .IN1(n10505), .IN2(n8916), .QN(n11121) );
  NAND3X0 U11209 ( .IN1(n5356), .IN2(n10507), .IN3(n5538), .QN(n10505) );
  NAND3X0 U11210 ( .IN1(n11124), .IN2(n11125), .IN3(n11126), .QN(g33578) );
  NAND2X0 U11211 ( .IN1(n10524), .IN2(n11107), .QN(n11126) );
  NOR2X0 U11212 ( .IN1(n5514), .IN2(n11127), .QN(n10524) );
  NAND2X0 U11213 ( .IN1(n9010), .IN2(g2197), .QN(n11125) );
  NAND3X0 U11214 ( .IN1(n11127), .IN2(g2227), .IN3(n8874), .QN(n11124) );
  NAND3X0 U11215 ( .IN1(n11128), .IN2(n11129), .IN3(n11130), .QN(g33577) );
  NAND3X0 U11216 ( .IN1(n11107), .IN2(n10507), .IN3(n10527), .QN(n11130) );
  NAND3X0 U11217 ( .IN1(n11127), .IN2(g2197), .IN3(n8874), .QN(n11129) );
  NAND2X0 U11218 ( .IN1(n9010), .IN2(g2204), .QN(n11128) );
  NAND2X0 U11219 ( .IN1(n11131), .IN2(n11132), .QN(g33576) );
  NAND2X0 U11220 ( .IN1(n10527), .IN2(n11127), .QN(n11132) );
  NOR2X0 U11221 ( .IN1(n8956), .IN2(n5356), .QN(n10527) );
  NAND4X0 U11222 ( .IN1(n5538), .IN2(n11133), .IN3(n11107), .IN4(n8901), .QN(
        n11131) );
  NAND2X0 U11223 ( .IN1(n3115), .IN2(n10106), .QN(n11107) );
  INVX0 U11224 ( .INP(n3165), .ZN(n10106) );
  NAND3X0 U11225 ( .IN1(n5287), .IN2(n5519), .IN3(n3116), .QN(n3165) );
  NAND2X0 U11226 ( .IN1(n5356), .IN2(n10520), .QN(n11133) );
  NAND2X0 U11227 ( .IN1(n5514), .IN2(n10507), .QN(n10520) );
  INVX0 U11228 ( .INP(n11127), .ZN(n10507) );
  NOR2X0 U11229 ( .IN1(n10514), .IN2(n700), .QN(n11127) );
  NOR2X0 U11230 ( .IN1(n8161), .IN2(n11134), .QN(n700) );
  NOR3X0 U11231 ( .IN1(n5364), .IN2(test_so49), .IN3(n11019), .QN(n11134) );
  NAND4X0 U11232 ( .IN1(n8443), .IN2(n5768), .IN3(test_so68), .IN4(n11135), 
        .QN(n11019) );
  NOR3X0 U11233 ( .IN1(g1548), .IN2(n8167), .IN3(g1559), .QN(n11135) );
  NAND3X0 U11234 ( .IN1(n10546), .IN2(n9486), .IN3(n11136), .QN(n10514) );
  NAND3X0 U11235 ( .IN1(n5377), .IN2(g2689), .IN3(n5308), .QN(n11136) );
  NAND2X0 U11236 ( .IN1(n2549), .IN2(g1478), .QN(n9486) );
  NAND2X0 U11237 ( .IN1(n10844), .IN2(n11137), .QN(n10546) );
  NAND3X0 U11238 ( .IN1(n9698), .IN2(g691), .IN3(n5595), .QN(n11137) );
  NAND4X0 U11239 ( .IN1(n11138), .IN2(n3180), .IN3(n11139), .IN4(n11140), .QN(
        g33575) );
  NAND2X0 U11240 ( .IN1(n9010), .IN2(g1996), .QN(n11140) );
  NAND4X0 U11241 ( .IN1(n11141), .IN2(n11142), .IN3(n11143), .IN4(n8901), .QN(
        n11139) );
  INVX0 U11242 ( .INP(n11144), .ZN(n11143) );
  NAND3X0 U11243 ( .IN1(g2070), .IN2(g112), .IN3(n5505), .QN(n11142) );
  NAND4X0 U11244 ( .IN1(n11145), .IN2(g2070), .IN3(n10989), .IN4(n11146), .QN(
        n3180) );
  NOR2X0 U11245 ( .IN1(g2040), .IN2(g112), .QN(n11146) );
  INVX0 U11246 ( .INP(n11147), .ZN(n11145) );
  NAND2X0 U11247 ( .IN1(n11148), .IN2(g2047), .QN(n11138) );
  NAND2X0 U11248 ( .IN1(n10991), .IN2(n11149), .QN(n11148) );
  NAND2X0 U11249 ( .IN1(n11147), .IN2(n8916), .QN(n11149) );
  NAND2X0 U11250 ( .IN1(n11141), .IN2(n10109), .QN(n11147) );
  NAND3X0 U11251 ( .IN1(n11150), .IN2(n11151), .IN3(n11152), .QN(g33574) );
  NAND2X0 U11252 ( .IN1(n10553), .IN2(g2116), .QN(n11152) );
  NAND3X0 U11253 ( .IN1(n5463), .IN2(n10551), .IN3(n8873), .QN(n11151) );
  NAND2X0 U11254 ( .IN1(n9010), .IN2(g2112), .QN(n11150) );
  NAND3X0 U11255 ( .IN1(n11153), .IN2(n11154), .IN3(n11155), .QN(g33573) );
  NAND2X0 U11256 ( .IN1(n10553), .IN2(g2112), .QN(n11155) );
  NAND2X0 U11257 ( .IN1(n11156), .IN2(g2108), .QN(n11154) );
  NAND2X0 U11258 ( .IN1(n11157), .IN2(n8916), .QN(n11156) );
  NAND2X0 U11259 ( .IN1(n10551), .IN2(g2102), .QN(n11157) );
  NAND4X0 U11260 ( .IN1(n10551), .IN2(n8900), .IN3(n5666), .IN4(n5452), .QN(
        n11153) );
  INVX0 U11261 ( .INP(n10564), .ZN(n10551) );
  NAND2X0 U11262 ( .IN1(n11158), .IN2(n11159), .QN(g33572) );
  NAND2X0 U11263 ( .IN1(n10553), .IN2(g2108), .QN(n11159) );
  NAND2X0 U11264 ( .IN1(n11160), .IN2(g2102), .QN(n11158) );
  NAND2X0 U11265 ( .IN1(n11161), .IN2(n11162), .QN(g33571) );
  NAND2X0 U11266 ( .IN1(n10553), .IN2(g2089), .QN(n11162) );
  INVX0 U11267 ( .INP(n11160), .ZN(n10553) );
  NAND2X0 U11268 ( .IN1(n11160), .IN2(g2084), .QN(n11161) );
  NAND2X0 U11269 ( .IN1(n10564), .IN2(n8916), .QN(n11160) );
  NAND3X0 U11270 ( .IN1(n5355), .IN2(n10566), .IN3(n5535), .QN(n10564) );
  NAND3X0 U11271 ( .IN1(n11163), .IN2(n11164), .IN3(n11165), .QN(g33570) );
  NAND2X0 U11272 ( .IN1(n10584), .IN2(n11144), .QN(n11165) );
  NOR2X0 U11273 ( .IN1(n5505), .IN2(n11166), .QN(n10584) );
  NAND2X0 U11274 ( .IN1(n9010), .IN2(g2040), .QN(n11164) );
  NAND3X0 U11275 ( .IN1(n11166), .IN2(g2070), .IN3(n8873), .QN(n11163) );
  NAND3X0 U11276 ( .IN1(n11167), .IN2(n11168), .IN3(n11169), .QN(g33569) );
  NAND3X0 U11277 ( .IN1(n11144), .IN2(n10566), .IN3(n10587), .QN(n11169) );
  NAND3X0 U11278 ( .IN1(n11166), .IN2(g2040), .IN3(n8873), .QN(n11168) );
  NAND2X0 U11279 ( .IN1(n9011), .IN2(g2047), .QN(n11167) );
  NAND2X0 U11280 ( .IN1(n11170), .IN2(n11171), .QN(g33568) );
  NAND2X0 U11281 ( .IN1(n10587), .IN2(n11166), .QN(n11171) );
  NOR2X0 U11282 ( .IN1(n8956), .IN2(n5355), .QN(n10587) );
  NAND4X0 U11283 ( .IN1(n5535), .IN2(n11172), .IN3(n11144), .IN4(n8902), .QN(
        n11170) );
  NAND2X0 U11284 ( .IN1(n3115), .IN2(n10109), .QN(n11144) );
  INVX0 U11285 ( .INP(n10103), .ZN(n10109) );
  NAND3X0 U11286 ( .IN1(n5519), .IN2(g518), .IN3(n3195), .QN(n10103) );
  NAND2X0 U11287 ( .IN1(n5355), .IN2(n10580), .QN(n11172) );
  NAND2X0 U11288 ( .IN1(n5505), .IN2(n10566), .QN(n10580) );
  INVX0 U11289 ( .INP(n11166), .ZN(n10566) );
  NOR2X0 U11290 ( .IN1(n10573), .IN2(n11141), .QN(n11166) );
  NOR2X0 U11291 ( .IN1(n11173), .IN2(n8446), .QN(n11141) );
  NOR3X0 U11292 ( .IN1(g1171), .IN2(n11174), .IN3(g1183), .QN(n11173) );
  NAND3X0 U11293 ( .IN1(n10776), .IN2(n9623), .IN3(n11175), .QN(n10573) );
  NAND3X0 U11294 ( .IN1(g2145), .IN2(g2130), .IN3(g2138), .QN(n11175) );
  NAND2X0 U11295 ( .IN1(n5286), .IN2(g956), .QN(n9623) );
  NAND3X0 U11296 ( .IN1(n11176), .IN2(n11177), .IN3(n11178), .QN(g33567) );
  NAND2X0 U11297 ( .IN1(test_so8), .IN2(n8950), .QN(n11178) );
  NAND2X0 U11298 ( .IN1(n11179), .IN2(n11180), .QN(n11177) );
  NAND2X0 U11299 ( .IN1(n11181), .IN2(n11182), .QN(n11180) );
  NAND3X0 U11300 ( .IN1(n10097), .IN2(n8871), .IN3(n11183), .QN(n11182) );
  NAND2X0 U11301 ( .IN1(n8185), .IN2(n11184), .QN(n11181) );
  NAND2X0 U11302 ( .IN1(n11185), .IN2(n11186), .QN(n11184) );
  NAND3X0 U11303 ( .IN1(n10638), .IN2(n10989), .IN3(n11187), .QN(n11186) );
  INVX0 U11304 ( .INP(n10097), .ZN(n10638) );
  NAND2X0 U11305 ( .IN1(n5503), .IN2(g1936), .QN(n10097) );
  NAND2X0 U11306 ( .IN1(n11183), .IN2(n8916), .QN(n11185) );
  INVX0 U11307 ( .INP(n11188), .ZN(n11183) );
  NAND2X0 U11308 ( .IN1(n11189), .IN2(g1913), .QN(n11176) );
  NAND2X0 U11309 ( .IN1(n10991), .IN2(n11190), .QN(n11189) );
  NAND2X0 U11310 ( .IN1(n11191), .IN2(n8916), .QN(n11190) );
  NAND2X0 U11311 ( .IN1(n11179), .IN2(n11187), .QN(n11191) );
  NAND3X0 U11312 ( .IN1(n11192), .IN2(n11193), .IN3(n11194), .QN(g33566) );
  NAND2X0 U11313 ( .IN1(n10612), .IN2(g1982), .QN(n11194) );
  NAND3X0 U11314 ( .IN1(n5462), .IN2(n10611), .IN3(n8872), .QN(n11193) );
  NAND2X0 U11315 ( .IN1(n9011), .IN2(g1978), .QN(n11192) );
  NAND3X0 U11316 ( .IN1(n11195), .IN2(n11196), .IN3(n11197), .QN(g33565) );
  NAND2X0 U11317 ( .IN1(n10612), .IN2(g1978), .QN(n11197) );
  NAND2X0 U11318 ( .IN1(n11198), .IN2(g1974), .QN(n11196) );
  NAND2X0 U11319 ( .IN1(n11199), .IN2(n8916), .QN(n11198) );
  NAND2X0 U11320 ( .IN1(n10611), .IN2(g1968), .QN(n11199) );
  NAND4X0 U11321 ( .IN1(n10611), .IN2(n8899), .IN3(n5664), .IN4(n5450), .QN(
        n11195) );
  INVX0 U11322 ( .INP(n10623), .ZN(n10611) );
  NAND2X0 U11323 ( .IN1(n11200), .IN2(n11201), .QN(g33564) );
  NAND2X0 U11324 ( .IN1(n10612), .IN2(g1974), .QN(n11201) );
  NAND2X0 U11325 ( .IN1(n11202), .IN2(g1968), .QN(n11200) );
  NAND2X0 U11326 ( .IN1(n11203), .IN2(n11204), .QN(g33563) );
  NAND2X0 U11327 ( .IN1(n10612), .IN2(g1955), .QN(n11204) );
  INVX0 U11328 ( .INP(n11202), .ZN(n10612) );
  NAND2X0 U11329 ( .IN1(n11202), .IN2(g1950), .QN(n11203) );
  NAND2X0 U11330 ( .IN1(n10623), .IN2(n8916), .QN(n11202) );
  NAND3X0 U11331 ( .IN1(n10625), .IN2(n8586), .IN3(n5534), .QN(n10623) );
  NAND3X0 U11332 ( .IN1(n11205), .IN2(n11206), .IN3(n11207), .QN(g33562) );
  NAND2X0 U11333 ( .IN1(n9011), .IN2(g1906), .QN(n11207) );
  NAND2X0 U11334 ( .IN1(n11208), .IN2(g1936), .QN(n11206) );
  NAND2X0 U11335 ( .IN1(n10644), .IN2(n11188), .QN(n11205) );
  NOR2X0 U11336 ( .IN1(n5503), .IN2(n11209), .QN(n10644) );
  NAND3X0 U11337 ( .IN1(n11210), .IN2(n11211), .IN3(n11212), .QN(g33561) );
  NAND2X0 U11338 ( .IN1(n11208), .IN2(g1906), .QN(n11212) );
  NAND2X0 U11339 ( .IN1(n9011), .IN2(g1913), .QN(n11211) );
  NAND3X0 U11340 ( .IN1(n10650), .IN2(n11188), .IN3(n8873), .QN(n11210) );
  NOR2X0 U11341 ( .IN1(n8586), .IN2(n11209), .QN(n10650) );
  NAND2X0 U11342 ( .IN1(n11213), .IN2(n11214), .QN(g33560) );
  NAND4X0 U11343 ( .IN1(n5534), .IN2(n11215), .IN3(n11188), .IN4(n8901), .QN(
        n11214) );
  NAND2X0 U11344 ( .IN1(n3115), .IN2(n11187), .QN(n11188) );
  INVX0 U11345 ( .INP(n10098), .ZN(n11187) );
  NAND3X0 U11346 ( .IN1(g518), .IN2(g504), .IN3(n3195), .QN(n10098) );
  NAND2X0 U11347 ( .IN1(n8586), .IN2(n11216), .QN(n11215) );
  NAND2X0 U11348 ( .IN1(n5503), .IN2(n10625), .QN(n11216) );
  NAND2X0 U11349 ( .IN1(n11208), .IN2(test_so8), .QN(n11213) );
  NOR2X0 U11350 ( .IN1(n10625), .IN2(n8941), .QN(n11208) );
  INVX0 U11351 ( .INP(n11209), .ZN(n10625) );
  NOR2X0 U11352 ( .IN1(n10632), .IN2(n11179), .QN(n11209) );
  NOR2X0 U11353 ( .IN1(n11217), .IN2(n8155), .QN(n11179) );
  NOR2X0 U11354 ( .IN1(n11218), .IN2(n11174), .QN(n11217) );
  INVX0 U11355 ( .INP(n11219), .ZN(n11218) );
  NAND3X0 U11356 ( .IN1(n10776), .IN2(n9559), .IN3(n11220), .QN(n10632) );
  NAND3X0 U11357 ( .IN1(g2138), .IN2(g2130), .IN3(n5307), .QN(n11220) );
  NAND2X0 U11358 ( .IN1(n5286), .IN2(g1129), .QN(n9559) );
  NAND3X0 U11359 ( .IN1(n11221), .IN2(n11222), .IN3(n11223), .QN(g33559) );
  NAND2X0 U11360 ( .IN1(n9011), .IN2(g1728), .QN(n11223) );
  NAND4X0 U11361 ( .IN1(n11224), .IN2(n10104), .IN3(n11225), .IN4(n11226), 
        .QN(n11222) );
  NAND3X0 U11362 ( .IN1(g1802), .IN2(g112), .IN3(n5504), .QN(n11226) );
  NAND2X0 U11363 ( .IN1(n11227), .IN2(n11228), .QN(n11225) );
  NAND3X0 U11364 ( .IN1(n10989), .IN2(g1802), .IN3(n5504), .QN(n11228) );
  NAND2X0 U11365 ( .IN1(n3115), .IN2(n8916), .QN(n11227) );
  NAND2X0 U11366 ( .IN1(n11229), .IN2(g1779), .QN(n11221) );
  NAND2X0 U11367 ( .IN1(n10991), .IN2(n11230), .QN(n11229) );
  NAND2X0 U11368 ( .IN1(n11231), .IN2(n8916), .QN(n11230) );
  NAND2X0 U11369 ( .IN1(n11224), .IN2(n10104), .QN(n11231) );
  NAND3X0 U11370 ( .IN1(n11232), .IN2(n11233), .IN3(n11234), .QN(g33558) );
  NAND2X0 U11371 ( .IN1(n10668), .IN2(g1848), .QN(n11234) );
  NAND3X0 U11372 ( .IN1(n5464), .IN2(n10667), .IN3(n8872), .QN(n11233) );
  NAND2X0 U11373 ( .IN1(n9011), .IN2(g1844), .QN(n11232) );
  NAND3X0 U11374 ( .IN1(n11235), .IN2(n11236), .IN3(n11237), .QN(g33557) );
  NAND2X0 U11375 ( .IN1(n10668), .IN2(g1844), .QN(n11237) );
  NAND2X0 U11376 ( .IN1(n11238), .IN2(g1840), .QN(n11236) );
  NAND2X0 U11377 ( .IN1(n11239), .IN2(n8916), .QN(n11238) );
  NAND2X0 U11378 ( .IN1(n10667), .IN2(g1834), .QN(n11239) );
  NAND4X0 U11379 ( .IN1(n10667), .IN2(n8899), .IN3(n5665), .IN4(n5451), .QN(
        n11235) );
  INVX0 U11380 ( .INP(n10679), .ZN(n10667) );
  NAND2X0 U11381 ( .IN1(n11240), .IN2(n11241), .QN(g33556) );
  NAND2X0 U11382 ( .IN1(n10668), .IN2(g1840), .QN(n11241) );
  NAND2X0 U11383 ( .IN1(n11242), .IN2(g1834), .QN(n11240) );
  NAND2X0 U11384 ( .IN1(n11243), .IN2(n11244), .QN(g33555) );
  NAND2X0 U11385 ( .IN1(n10668), .IN2(g1821), .QN(n11244) );
  INVX0 U11386 ( .INP(n11242), .ZN(n10668) );
  NAND2X0 U11387 ( .IN1(n11242), .IN2(g1816), .QN(n11243) );
  NAND2X0 U11388 ( .IN1(n10679), .IN2(n8916), .QN(n11242) );
  NAND3X0 U11389 ( .IN1(n5352), .IN2(n10681), .IN3(n5536), .QN(n10679) );
  NAND3X0 U11390 ( .IN1(n11245), .IN2(n11246), .IN3(n11247), .QN(g33554) );
  NAND2X0 U11391 ( .IN1(n10698), .IN2(n11248), .QN(n11247) );
  NOR2X0 U11392 ( .IN1(n5504), .IN2(n11249), .QN(n10698) );
  NAND2X0 U11393 ( .IN1(n9011), .IN2(g1772), .QN(n11246) );
  NAND3X0 U11394 ( .IN1(n11249), .IN2(g1802), .IN3(n8872), .QN(n11245) );
  NAND3X0 U11395 ( .IN1(n11250), .IN2(n11251), .IN3(n11252), .QN(g33553) );
  NAND3X0 U11396 ( .IN1(n11248), .IN2(n10681), .IN3(n10701), .QN(n11252) );
  NAND3X0 U11397 ( .IN1(n11249), .IN2(g1772), .IN3(n8872), .QN(n11251) );
  NAND2X0 U11398 ( .IN1(n9012), .IN2(g1779), .QN(n11250) );
  NAND2X0 U11399 ( .IN1(n11253), .IN2(n11254), .QN(g33552) );
  NAND2X0 U11400 ( .IN1(n10701), .IN2(n11249), .QN(n11254) );
  NOR2X0 U11401 ( .IN1(n8956), .IN2(n5352), .QN(n10701) );
  NAND4X0 U11402 ( .IN1(n5536), .IN2(n11255), .IN3(n11248), .IN4(n8901), .QN(
        n11253) );
  NAND2X0 U11403 ( .IN1(n3115), .IN2(n10104), .QN(n11248) );
  INVX0 U11404 ( .INP(n10107), .ZN(n10104) );
  NAND3X0 U11405 ( .IN1(n5287), .IN2(g504), .IN3(n3195), .QN(n10107) );
  NAND2X0 U11406 ( .IN1(n5352), .IN2(n10694), .QN(n11255) );
  NAND2X0 U11407 ( .IN1(n5504), .IN2(n10681), .QN(n10694) );
  INVX0 U11408 ( .INP(n11249), .ZN(n10681) );
  NOR2X0 U11409 ( .IN1(n10688), .IN2(n11224), .QN(n11249) );
  NOR2X0 U11410 ( .IN1(n8617), .IN2(n11256), .QN(n11224) );
  NOR2X0 U11411 ( .IN1(n11257), .IN2(n11174), .QN(n11256) );
  NAND3X0 U11412 ( .IN1(n10776), .IN2(n9514), .IN3(n11258), .QN(n10688) );
  NAND3X0 U11413 ( .IN1(g2145), .IN2(g2130), .IN3(n5275), .QN(n11258) );
  NAND2X0 U11414 ( .IN1(n5286), .IN2(g1105), .QN(n9514) );
  NAND3X0 U11415 ( .IN1(n11259), .IN2(n11260), .IN3(n11261), .QN(g33551) );
  NAND2X0 U11416 ( .IN1(n9012), .IN2(g1592), .QN(n11261) );
  NAND3X0 U11417 ( .IN1(n11262), .IN2(n11263), .IN3(g33533), .QN(n11260) );
  NAND2X0 U11418 ( .IN1(n11264), .IN2(n11265), .QN(n11263) );
  NAND3X0 U11419 ( .IN1(n11266), .IN2(n8871), .IN3(n3115), .QN(n11265) );
  NAND2X0 U11420 ( .IN1(g25259), .IN2(g112), .QN(n11266) );
  NAND3X0 U11421 ( .IN1(n8185), .IN2(n10989), .IN3(g25259), .QN(n11264) );
  NAND2X0 U11422 ( .IN1(test_so75), .IN2(n11267), .QN(n11259) );
  NAND2X0 U11423 ( .IN1(n10991), .IN2(n11268), .QN(n11267) );
  NAND2X0 U11424 ( .IN1(n11269), .IN2(n8916), .QN(n11268) );
  NAND2X0 U11425 ( .IN1(g33533), .IN2(n11262), .QN(n11269) );
  NAND3X0 U11426 ( .IN1(n11270), .IN2(n11271), .IN3(n11272), .QN(g33550) );
  NAND2X0 U11427 ( .IN1(n10726), .IN2(g1714), .QN(n11272) );
  NAND3X0 U11428 ( .IN1(n5460), .IN2(n11273), .IN3(n8872), .QN(n11271) );
  NAND2X0 U11429 ( .IN1(n9049), .IN2(g1710), .QN(n11270) );
  NAND3X0 U11430 ( .IN1(n11274), .IN2(n11275), .IN3(n11276), .QN(g33549) );
  NAND2X0 U11431 ( .IN1(n10726), .IN2(g1710), .QN(n11276) );
  NAND2X0 U11432 ( .IN1(test_so15), .IN2(n11277), .QN(n11275) );
  NAND2X0 U11433 ( .IN1(n11278), .IN2(n8916), .QN(n11277) );
  NAND2X0 U11434 ( .IN1(n11273), .IN2(g1700), .QN(n11278) );
  NAND4X0 U11435 ( .IN1(n11273), .IN2(n8899), .IN3(n5417), .IN4(n8621), .QN(
        n11274) );
  INVX0 U11436 ( .INP(n10724), .ZN(n11273) );
  NAND2X0 U11437 ( .IN1(n11279), .IN2(n11280), .QN(g33548) );
  NAND2X0 U11438 ( .IN1(test_so15), .IN2(n10726), .QN(n11280) );
  NAND2X0 U11439 ( .IN1(n11281), .IN2(g1700), .QN(n11279) );
  NAND2X0 U11440 ( .IN1(n11282), .IN2(n11283), .QN(g33547) );
  NAND2X0 U11441 ( .IN1(n10726), .IN2(g1687), .QN(n11283) );
  INVX0 U11442 ( .INP(n11281), .ZN(n10726) );
  NAND2X0 U11443 ( .IN1(n11281), .IN2(g1682), .QN(n11282) );
  NAND2X0 U11444 ( .IN1(n10724), .IN2(n8917), .QN(n11281) );
  NAND3X0 U11445 ( .IN1(n5362), .IN2(n10738), .IN3(n5598), .QN(n10724) );
  NAND3X0 U11446 ( .IN1(n11284), .IN2(n11285), .IN3(n11286), .QN(g33546) );
  NAND2X0 U11447 ( .IN1(n9041), .IN2(g1636), .QN(n11286) );
  NAND2X0 U11448 ( .IN1(n11287), .IN2(g1668), .QN(n11285) );
  NAND2X0 U11449 ( .IN1(n10756), .IN2(n11288), .QN(n11284) );
  NOR2X0 U11450 ( .IN1(n5549), .IN2(n11289), .QN(n10756) );
  NAND3X0 U11451 ( .IN1(n11290), .IN2(n11291), .IN3(n11292), .QN(g33545) );
  NAND2X0 U11452 ( .IN1(n11287), .IN2(g1636), .QN(n11292) );
  NAND2X0 U11453 ( .IN1(test_so75), .IN2(n8949), .QN(n11291) );
  NAND3X0 U11454 ( .IN1(n10762), .IN2(n11288), .IN3(n8874), .QN(n11290) );
  NOR2X0 U11455 ( .IN1(n5362), .IN2(n11289), .QN(n10762) );
  NAND2X0 U11456 ( .IN1(n11293), .IN2(n11294), .QN(g33544) );
  NAND2X0 U11457 ( .IN1(n11287), .IN2(g1592), .QN(n11294) );
  NOR2X0 U11458 ( .IN1(n10738), .IN2(n8943), .QN(n11287) );
  NAND4X0 U11459 ( .IN1(n10738), .IN2(n8899), .IN3(n11288), .IN4(n11295), .QN(
        n11293) );
  INVX0 U11460 ( .INP(n11296), .ZN(n11295) );
  NAND2X0 U11461 ( .IN1(n11297), .IN2(n5598), .QN(n11296) );
  NAND2X0 U11462 ( .IN1(n3115), .IN2(n11262), .QN(n11288) );
  INVX0 U11463 ( .INP(n10094), .ZN(n11262) );
  NAND3X0 U11464 ( .IN1(n5287), .IN2(n5519), .IN3(n3195), .QN(n10094) );
  INVX0 U11465 ( .INP(n11289), .ZN(n10738) );
  NOR2X0 U11466 ( .IN1(n10745), .IN2(g33533), .QN(n11289) );
  NAND3X0 U11467 ( .IN1(n10776), .IN2(n9487), .IN3(n11298), .QN(n10745) );
  NAND3X0 U11468 ( .IN1(n5307), .IN2(g2130), .IN3(n5275), .QN(n11298) );
  NAND2X0 U11469 ( .IN1(n5286), .IN2(g1135), .QN(n9487) );
  NAND2X0 U11470 ( .IN1(n10844), .IN2(n11299), .QN(n10776) );
  NAND3X0 U11471 ( .IN1(n9697), .IN2(g691), .IN3(n5595), .QN(n11299) );
  INVX0 U11472 ( .INP(g134), .ZN(n10844) );
  NAND2X0 U11473 ( .IN1(n11300), .IN2(n11301), .QN(g33543) );
  NAND3X0 U11474 ( .IN1(n8896), .IN2(g1379), .IN3(n11302), .QN(n11301) );
  NAND2X0 U11475 ( .IN1(n11303), .IN2(n11304), .QN(n11302) );
  NAND2X0 U11476 ( .IN1(n8172), .IN2(n11305), .QN(n11304) );
  NAND2X0 U11477 ( .IN1(n11306), .IN2(g1373), .QN(n11300) );
  NAND2X0 U11478 ( .IN1(n11307), .IN2(n8917), .QN(n11306) );
  NAND3X0 U11479 ( .IN1(n11303), .IN2(n11305), .IN3(n8516), .QN(n11307) );
  NAND3X0 U11480 ( .IN1(n11308), .IN2(n11309), .IN3(n11310), .QN(g33542) );
  NAND2X0 U11481 ( .IN1(n9043), .IN2(g1270), .QN(n11310) );
  NAND3X0 U11482 ( .IN1(n11311), .IN2(n11312), .IN3(g1274), .QN(n11309) );
  INVX0 U11483 ( .INP(n11313), .ZN(n11308) );
  NOR2X0 U11484 ( .IN1(g1274), .IN2(n11312), .QN(n11313) );
  NAND2X0 U11485 ( .IN1(n11314), .IN2(n11315), .QN(g33541) );
  NAND3X0 U11486 ( .IN1(n8898), .IN2(g1036), .IN3(n11316), .QN(n11315) );
  NAND2X0 U11487 ( .IN1(n11317), .IN2(n11318), .QN(n11316) );
  NAND2X0 U11488 ( .IN1(n8174), .IN2(n11319), .QN(n11318) );
  NAND2X0 U11489 ( .IN1(n11320), .IN2(g1030), .QN(n11314) );
  NAND2X0 U11490 ( .IN1(n11321), .IN2(n8917), .QN(n11320) );
  NAND3X0 U11491 ( .IN1(n11317), .IN2(n11319), .IN3(n8515), .QN(n11321) );
  NAND3X0 U11492 ( .IN1(n11322), .IN2(n11323), .IN3(n11324), .QN(g33540) );
  NAND2X0 U11493 ( .IN1(n9043), .IN2(g925), .QN(n11324) );
  NAND3X0 U11494 ( .IN1(n11325), .IN2(n11326), .IN3(g930), .QN(n11323) );
  INVX0 U11495 ( .INP(n11327), .ZN(n11322) );
  NOR2X0 U11496 ( .IN1(g930), .IN2(n11326), .QN(n11327) );
  NAND3X0 U11497 ( .IN1(n11328), .IN2(n11329), .IN3(n11330), .QN(g33539) );
  NAND2X0 U11498 ( .IN1(n9043), .IN2(g758), .QN(n11330) );
  NAND3X0 U11499 ( .IN1(n2404), .IN2(n11331), .IN3(g763), .QN(n11329) );
  INVX0 U11500 ( .INP(n2980), .ZN(n11331) );
  NAND2X0 U11501 ( .IN1(n2980), .IN2(n5332), .QN(n11328) );
  NAND3X0 U11502 ( .IN1(n11332), .IN2(n11333), .IN3(n11334), .QN(g33538) );
  NAND2X0 U11503 ( .IN1(n9044), .IN2(g590), .QN(n11334) );
  NAND3X0 U11504 ( .IN1(n2421), .IN2(n11335), .IN3(g595), .QN(n11333) );
  INVX0 U11505 ( .INP(n2982), .ZN(n11335) );
  NAND2X0 U11506 ( .IN1(n2982), .IN2(n5476), .QN(n11332) );
  NAND2X0 U11507 ( .IN1(n11336), .IN2(n11337), .QN(g33537) );
  NAND2X0 U11508 ( .IN1(n9045), .IN2(g301), .QN(n11337) );
  NAND3X0 U11509 ( .IN1(n2707), .IN2(g142), .IN3(n8877), .QN(n11336) );
  NOR2X0 U11510 ( .IN1(n5843), .IN2(n11338), .QN(g33536) );
  NOR2X0 U11511 ( .IN1(n2710), .IN2(n8927), .QN(n11338) );
  NAND3X0 U11512 ( .IN1(n11339), .IN2(n11340), .IN3(n11341), .QN(g33535) );
  NAND2X0 U11513 ( .IN1(n9045), .IN2(g291), .QN(n11341) );
  NAND3X0 U11514 ( .IN1(n8568), .IN2(n11342), .IN3(g294), .QN(n11340) );
  INVX0 U11515 ( .INP(n3276), .ZN(n11342) );
  NAND2X0 U11516 ( .IN1(n3276), .IN2(n5680), .QN(n11339) );
  NAND3X0 U11517 ( .IN1(n11343), .IN2(n11344), .IN3(n11345), .QN(g33534) );
  NAND2X0 U11518 ( .IN1(n9046), .IN2(g150), .QN(n11345) );
  NAND3X0 U11519 ( .IN1(n10217), .IN2(n11346), .IN3(g153), .QN(n11344) );
  INVX0 U11520 ( .INP(n3277), .ZN(n11346) );
  NAND2X0 U11521 ( .IN1(n3277), .IN2(n5677), .QN(n11343) );
  NOR2X0 U11522 ( .IN1(n11347), .IN2(n8150), .QN(g33533) );
  NOR2X0 U11523 ( .IN1(n11348), .IN2(n11174), .QN(n11347) );
  NAND4X0 U11524 ( .IN1(n5547), .IN2(n5442), .IN3(n8445), .IN4(n11349), .QN(
        n11174) );
  NOR3X0 U11525 ( .IN1(n5320), .IN2(test_so76), .IN3(n8168), .QN(n11349) );
  INVX0 U11526 ( .INP(n11350), .ZN(n11348) );
  NOR4X0 U11527 ( .IN1(n11351), .IN2(n11352), .IN3(n11353), .IN4(n11354), .QN(
        g33435) );
  NOR2X0 U11528 ( .IN1(n5403), .IN2(n10025), .QN(n11354) );
  NOR2X0 U11529 ( .IN1(n5544), .IN2(n10030), .QN(n11353) );
  NOR2X0 U11530 ( .IN1(n5378), .IN2(n10020), .QN(n11352) );
  NOR2X0 U11531 ( .IN1(n5610), .IN2(n10014), .QN(n11351) );
  NOR4X0 U11532 ( .IN1(n11355), .IN2(n11356), .IN3(n11357), .IN4(n11358), .QN(
        g33079) );
  NOR2X0 U11533 ( .IN1(n5404), .IN2(n10025), .QN(n11358) );
  NAND2X0 U11534 ( .IN1(n5301), .IN2(g2729), .QN(n10025) );
  NOR2X0 U11535 ( .IN1(n5545), .IN2(n10030), .QN(n11357) );
  NOR2X0 U11536 ( .IN1(n5379), .IN2(n10020), .QN(n11356) );
  NAND2X0 U11537 ( .IN1(n8186), .IN2(g2724), .QN(n10020) );
  NOR2X0 U11538 ( .IN1(n5609), .IN2(n10014), .QN(n11355) );
  NAND2X0 U11539 ( .IN1(g2724), .IN2(g2729), .QN(n10014) );
  NAND2X0 U11540 ( .IN1(n11359), .IN2(n11360), .QN(g33070) );
  NAND2X0 U11541 ( .IN1(n11361), .IN2(n11362), .QN(n11360) );
  NAND3X0 U11542 ( .IN1(n11363), .IN2(n11364), .IN3(n11365), .QN(n11361) );
  NAND2X0 U11543 ( .IN1(g25756), .IN2(n5646), .QN(n11365) );
  NAND2X0 U11544 ( .IN1(n11366), .IN2(n8917), .QN(n11363) );
  NAND2X0 U11545 ( .IN1(n9047), .IN2(g6565), .QN(n11359) );
  NAND2X0 U11546 ( .IN1(n11367), .IN2(n11368), .QN(g33069) );
  NAND2X0 U11547 ( .IN1(n11369), .IN2(g6561), .QN(n11368) );
  NAND2X0 U11548 ( .IN1(n11370), .IN2(n8917), .QN(n11369) );
  NAND2X0 U11549 ( .IN1(n5386), .IN2(n11362), .QN(n11370) );
  NAND2X0 U11550 ( .IN1(n11371), .IN2(g6565), .QN(n11367) );
  INVX0 U11551 ( .INP(n11372), .ZN(n11371) );
  NAND2X0 U11552 ( .IN1(n11373), .IN2(n11374), .QN(g33068) );
  NAND3X0 U11553 ( .IN1(n11362), .IN2(n11375), .IN3(n5646), .QN(n11374) );
  NAND2X0 U11554 ( .IN1(n9047), .IN2(g6555), .QN(n11373) );
  NAND2X0 U11555 ( .IN1(n11376), .IN2(n11377), .QN(g33067) );
  NAND2X0 U11556 ( .IN1(n11378), .IN2(n11362), .QN(n11377) );
  NAND2X0 U11557 ( .IN1(n751), .IN2(n11379), .QN(n11378) );
  NAND2X0 U11558 ( .IN1(n8905), .IN2(n11380), .QN(n11379) );
  NAND2X0 U11559 ( .IN1(n9048), .IN2(g6549), .QN(n11376) );
  NAND2X0 U11560 ( .IN1(n11381), .IN2(n11382), .QN(g33065) );
  NAND2X0 U11561 ( .IN1(n11383), .IN2(n11384), .QN(n11382) );
  NAND3X0 U11562 ( .IN1(n11385), .IN2(n11386), .IN3(n11387), .QN(n11383) );
  NAND2X0 U11563 ( .IN1(g25742), .IN2(n5651), .QN(n11387) );
  NAND2X0 U11564 ( .IN1(n8905), .IN2(n11388), .QN(n11385) );
  NAND2X0 U11565 ( .IN1(n9048), .IN2(g6219), .QN(n11381) );
  NAND2X0 U11566 ( .IN1(n11389), .IN2(n11390), .QN(g33064) );
  NAND2X0 U11567 ( .IN1(n11391), .IN2(g6215), .QN(n11390) );
  NAND2X0 U11568 ( .IN1(n11392), .IN2(n8917), .QN(n11391) );
  NAND2X0 U11569 ( .IN1(n5385), .IN2(n11384), .QN(n11392) );
  NAND2X0 U11570 ( .IN1(n11393), .IN2(g6219), .QN(n11389) );
  INVX0 U11571 ( .INP(n11394), .ZN(n11393) );
  NAND2X0 U11572 ( .IN1(n11395), .IN2(n11396), .QN(g33063) );
  NAND3X0 U11573 ( .IN1(n11384), .IN2(n11397), .IN3(n5651), .QN(n11396) );
  NAND2X0 U11574 ( .IN1(n9048), .IN2(g6209), .QN(n11395) );
  NAND2X0 U11575 ( .IN1(n11398), .IN2(n11399), .QN(g33062) );
  NAND2X0 U11576 ( .IN1(n11400), .IN2(n11384), .QN(n11399) );
  NAND2X0 U11577 ( .IN1(n1011), .IN2(n11401), .QN(n11400) );
  NAND2X0 U11578 ( .IN1(n11402), .IN2(n8917), .QN(n11401) );
  NAND2X0 U11579 ( .IN1(n9048), .IN2(g6203), .QN(n11398) );
  NAND2X0 U11580 ( .IN1(n11403), .IN2(n11404), .QN(g33060) );
  NAND2X0 U11581 ( .IN1(n11405), .IN2(n11406), .QN(n11404) );
  NAND3X0 U11582 ( .IN1(n11407), .IN2(n11408), .IN3(n11409), .QN(n11405) );
  NAND2X0 U11583 ( .IN1(g25728), .IN2(n5649), .QN(n11409) );
  NAND2X0 U11584 ( .IN1(n8906), .IN2(n11410), .QN(n11407) );
  NAND2X0 U11585 ( .IN1(n9049), .IN2(g5873), .QN(n11403) );
  NAND2X0 U11586 ( .IN1(n11411), .IN2(n11412), .QN(g33059) );
  NAND2X0 U11587 ( .IN1(n11413), .IN2(g5869), .QN(n11412) );
  NAND2X0 U11588 ( .IN1(n11414), .IN2(n8917), .QN(n11413) );
  NAND2X0 U11589 ( .IN1(n5388), .IN2(n11406), .QN(n11414) );
  NAND2X0 U11590 ( .IN1(n11415), .IN2(g5873), .QN(n11411) );
  INVX0 U11591 ( .INP(n11416), .ZN(n11415) );
  NAND2X0 U11592 ( .IN1(n11417), .IN2(n11418), .QN(g33058) );
  NAND3X0 U11593 ( .IN1(n11406), .IN2(n11419), .IN3(n5649), .QN(n11418) );
  NAND2X0 U11594 ( .IN1(n9049), .IN2(g5863), .QN(n11417) );
  NAND2X0 U11595 ( .IN1(n11420), .IN2(n11421), .QN(g33057) );
  NAND2X0 U11596 ( .IN1(n11422), .IN2(n11406), .QN(n11421) );
  NAND2X0 U11597 ( .IN1(n1075), .IN2(n11423), .QN(n11422) );
  NAND2X0 U11598 ( .IN1(n11424), .IN2(n8917), .QN(n11423) );
  NAND2X0 U11599 ( .IN1(n9050), .IN2(g5857), .QN(n11420) );
  NAND2X0 U11600 ( .IN1(n11425), .IN2(n11426), .QN(g33055) );
  NAND2X0 U11601 ( .IN1(n11427), .IN2(n11428), .QN(n11426) );
  NAND3X0 U11602 ( .IN1(n11429), .IN2(n11430), .IN3(n11431), .QN(n11427) );
  NAND2X0 U11603 ( .IN1(g25714), .IN2(n5647), .QN(n11431) );
  NAND2X0 U11604 ( .IN1(n8906), .IN2(n11432), .QN(n11429) );
  NAND2X0 U11605 ( .IN1(n9050), .IN2(g5527), .QN(n11425) );
  NAND2X0 U11606 ( .IN1(n11433), .IN2(n11434), .QN(g33054) );
  NAND2X0 U11607 ( .IN1(n11435), .IN2(g5523), .QN(n11434) );
  NAND2X0 U11608 ( .IN1(n11436), .IN2(n8917), .QN(n11435) );
  NAND2X0 U11609 ( .IN1(n5389), .IN2(n11428), .QN(n11436) );
  NAND2X0 U11610 ( .IN1(n11437), .IN2(g5527), .QN(n11433) );
  INVX0 U11611 ( .INP(n11438), .ZN(n11437) );
  NAND2X0 U11612 ( .IN1(n11439), .IN2(n11440), .QN(g33053) );
  NAND3X0 U11613 ( .IN1(n11428), .IN2(n11441), .IN3(n5647), .QN(n11440) );
  NAND2X0 U11614 ( .IN1(n9051), .IN2(g5517), .QN(n11439) );
  NAND2X0 U11615 ( .IN1(n11442), .IN2(n11443), .QN(g33052) );
  NAND2X0 U11616 ( .IN1(n11444), .IN2(n11428), .QN(n11443) );
  NAND2X0 U11617 ( .IN1(n495), .IN2(n11445), .QN(n11444) );
  NAND2X0 U11618 ( .IN1(n8905), .IN2(n11446), .QN(n11445) );
  NAND2X0 U11619 ( .IN1(n9041), .IN2(g5511), .QN(n11442) );
  NAND2X0 U11620 ( .IN1(n11447), .IN2(n11448), .QN(g33050) );
  NAND2X0 U11621 ( .IN1(n11449), .IN2(n11450), .QN(n11448) );
  NAND3X0 U11622 ( .IN1(n11451), .IN2(n11452), .IN3(n11453), .QN(n11449) );
  NAND2X0 U11623 ( .IN1(g25700), .IN2(n5650), .QN(n11453) );
  NAND2X0 U11624 ( .IN1(n8905), .IN2(n11454), .QN(n11451) );
  NAND2X0 U11625 ( .IN1(n9051), .IN2(g5180), .QN(n11447) );
  NAND2X0 U11626 ( .IN1(n11455), .IN2(n11456), .QN(g33049) );
  NAND2X0 U11627 ( .IN1(n11457), .IN2(g5176), .QN(n11456) );
  NAND2X0 U11628 ( .IN1(n11458), .IN2(n8917), .QN(n11457) );
  NAND2X0 U11629 ( .IN1(n5384), .IN2(n11450), .QN(n11458) );
  NAND2X0 U11630 ( .IN1(n11459), .IN2(g5180), .QN(n11455) );
  INVX0 U11631 ( .INP(n11460), .ZN(n11459) );
  NAND2X0 U11632 ( .IN1(n11461), .IN2(n11462), .QN(g33048) );
  NAND3X0 U11633 ( .IN1(n11450), .IN2(n11463), .IN3(n5650), .QN(n11462) );
  NAND2X0 U11634 ( .IN1(n9050), .IN2(g5170), .QN(n11461) );
  NAND2X0 U11635 ( .IN1(n11464), .IN2(n11465), .QN(g33047) );
  NAND2X0 U11636 ( .IN1(n11466), .IN2(n11450), .QN(n11465) );
  NAND2X0 U11637 ( .IN1(n745), .IN2(n11467), .QN(n11466) );
  NAND2X0 U11638 ( .IN1(n8906), .IN2(n11468), .QN(n11467) );
  NAND2X0 U11639 ( .IN1(n9051), .IN2(g5164), .QN(n11464) );
  NAND3X0 U11640 ( .IN1(n11469), .IN2(n11470), .IN3(n11471), .QN(g33046) );
  NAND2X0 U11641 ( .IN1(n9050), .IN2(g5052), .QN(n11471) );
  NAND2X0 U11642 ( .IN1(n5615), .IN2(n11472), .QN(n11470) );
  NAND2X0 U11643 ( .IN1(n11473), .IN2(n11474), .QN(n11472) );
  NAND3X0 U11644 ( .IN1(n11475), .IN2(n11474), .IN3(g5057), .QN(n11469) );
  NAND2X0 U11645 ( .IN1(n11476), .IN2(g5052), .QN(n11474) );
  NAND3X0 U11646 ( .IN1(n11477), .IN2(n11478), .IN3(n11479), .QN(g33045) );
  NAND2X0 U11647 ( .IN1(n10922), .IN2(g4567), .QN(n11479) );
  NAND3X0 U11648 ( .IN1(n11478), .IN2(n10298), .IN3(n11480), .QN(g33044) );
  NAND2X0 U11649 ( .IN1(test_so93), .IN2(n10922), .QN(n11480) );
  NAND3X0 U11650 ( .IN1(n11481), .IN2(n10920), .IN3(n11482), .QN(g33043) );
  NAND2X0 U11651 ( .IN1(test_so16), .IN2(n10922), .QN(n11482) );
  NAND3X0 U11652 ( .IN1(n11481), .IN2(n11478), .IN3(n11483), .QN(g33042) );
  NAND2X0 U11653 ( .IN1(n10922), .IN2(g4540), .QN(n11483) );
  NAND2X0 U11654 ( .IN1(n11484), .IN2(g4578), .QN(n11478) );
  NAND3X0 U11655 ( .IN1(n11477), .IN2(n10920), .IN3(n11485), .QN(g33041) );
  NAND2X0 U11656 ( .IN1(test_so56), .IN2(n10922), .QN(n11485) );
  NAND3X0 U11657 ( .IN1(n11486), .IN2(n10298), .IN3(n11487), .QN(g33040) );
  NAND2X0 U11658 ( .IN1(n10922), .IN2(g4504), .QN(n11487) );
  NAND2X0 U11659 ( .IN1(n11484), .IN2(n10304), .QN(n10298) );
  NAND2X0 U11660 ( .IN1(n9667), .IN2(n10792), .QN(n10304) );
  NAND3X0 U11661 ( .IN1(n11477), .IN2(n10925), .IN3(n11488), .QN(g33039) );
  NAND2X0 U11662 ( .IN1(n10922), .IN2(g4501), .QN(n11488) );
  NAND3X0 U11663 ( .IN1(n11477), .IN2(n11486), .IN3(n11489), .QN(g33038) );
  NAND2X0 U11664 ( .IN1(n10922), .IN2(g4498), .QN(n11489) );
  NAND2X0 U11665 ( .IN1(n11484), .IN2(n11490), .QN(n11477) );
  NAND2X0 U11666 ( .IN1(g72), .IN2(n9667), .QN(n11490) );
  INVX0 U11667 ( .INP(g73), .ZN(n9667) );
  NAND3X0 U11668 ( .IN1(n11481), .IN2(n10925), .IN3(n11491), .QN(g33037) );
  NAND2X0 U11669 ( .IN1(n10922), .IN2(g4495), .QN(n11491) );
  NAND3X0 U11670 ( .IN1(n11481), .IN2(n11486), .IN3(n11492), .QN(g33036) );
  NAND2X0 U11671 ( .IN1(n10922), .IN2(g4480), .QN(n11492) );
  INVX0 U11672 ( .INP(n11484), .ZN(n10922) );
  NAND2X0 U11673 ( .IN1(n11484), .IN2(g4572), .QN(n11486) );
  NAND2X0 U11674 ( .IN1(n11484), .IN2(n11493), .QN(n11481) );
  NAND2X0 U11675 ( .IN1(g73), .IN2(n10792), .QN(n11493) );
  INVX0 U11676 ( .INP(g72), .ZN(n10792) );
  NAND4X0 U11677 ( .IN1(n11494), .IN2(n11495), .IN3(n11496), .IN4(n11497), 
        .QN(g33035) );
  NAND3X0 U11678 ( .IN1(n11498), .IN2(g4108), .IN3(n8878), .QN(n11497) );
  NAND2X0 U11679 ( .IN1(n9050), .IN2(g4098), .QN(n11496) );
  NAND2X0 U11680 ( .IN1(n9334), .IN2(n5715), .QN(n11494) );
  INVX0 U11681 ( .INP(n11498), .ZN(n9334) );
  NAND2X0 U11682 ( .IN1(n11499), .IN2(g4098), .QN(n11498) );
  NAND2X0 U11683 ( .IN1(n11500), .IN2(n11501), .QN(g33034) );
  NAND2X0 U11684 ( .IN1(n11502), .IN2(n11503), .QN(n11501) );
  NAND3X0 U11685 ( .IN1(n11504), .IN2(n11505), .IN3(n11506), .QN(n11502) );
  NAND2X0 U11686 ( .IN1(g25676), .IN2(n8594), .QN(n11506) );
  NAND2X0 U11687 ( .IN1(n8905), .IN2(n11507), .QN(n11504) );
  NAND2X0 U11688 ( .IN1(n9050), .IN2(g3873), .QN(n11500) );
  NAND2X0 U11689 ( .IN1(n11508), .IN2(n11509), .QN(g33033) );
  NAND2X0 U11690 ( .IN1(test_so33), .IN2(n11510), .QN(n11509) );
  NAND2X0 U11691 ( .IN1(n11511), .IN2(n8917), .QN(n11510) );
  NAND2X0 U11692 ( .IN1(n5387), .IN2(n11503), .QN(n11511) );
  NAND2X0 U11693 ( .IN1(n11512), .IN2(g3873), .QN(n11508) );
  INVX0 U11694 ( .INP(n11513), .ZN(n11512) );
  NAND2X0 U11695 ( .IN1(n11514), .IN2(n11515), .QN(g33032) );
  NAND3X0 U11696 ( .IN1(n11516), .IN2(n8594), .IN3(n11503), .QN(n11515) );
  NAND2X0 U11697 ( .IN1(n9050), .IN2(g3863), .QN(n11514) );
  NAND2X0 U11698 ( .IN1(n11517), .IN2(n11518), .QN(g33031) );
  NAND2X0 U11699 ( .IN1(n11519), .IN2(n11503), .QN(n11518) );
  NAND2X0 U11700 ( .IN1(n1137), .IN2(n11520), .QN(n11519) );
  NAND2X0 U11701 ( .IN1(n11521), .IN2(n8917), .QN(n11520) );
  NAND2X0 U11702 ( .IN1(n9049), .IN2(g3857), .QN(n11517) );
  NAND2X0 U11703 ( .IN1(n11522), .IN2(n11523), .QN(g33029) );
  NAND2X0 U11704 ( .IN1(n11524), .IN2(n11525), .QN(n11523) );
  NAND3X0 U11705 ( .IN1(n11526), .IN2(n11527), .IN3(n11528), .QN(n11524) );
  NAND2X0 U11706 ( .IN1(g25662), .IN2(n5645), .QN(n11528) );
  NAND2X0 U11707 ( .IN1(n8906), .IN2(n11529), .QN(n11526) );
  NAND2X0 U11708 ( .IN1(n9045), .IN2(g3522), .QN(n11522) );
  NAND2X0 U11709 ( .IN1(n11530), .IN2(n11531), .QN(g33028) );
  NAND2X0 U11710 ( .IN1(n11532), .IN2(g3518), .QN(n11531) );
  NAND2X0 U11711 ( .IN1(n11533), .IN2(n8917), .QN(n11532) );
  NAND2X0 U11712 ( .IN1(n5383), .IN2(n11525), .QN(n11533) );
  NAND2X0 U11713 ( .IN1(n11534), .IN2(g3522), .QN(n11530) );
  INVX0 U11714 ( .INP(n11535), .ZN(n11534) );
  NAND2X0 U11715 ( .IN1(n11536), .IN2(n11537), .QN(g33027) );
  NAND3X0 U11716 ( .IN1(n11525), .IN2(n11538), .IN3(n5645), .QN(n11537) );
  NAND2X0 U11717 ( .IN1(n9049), .IN2(g3512), .QN(n11536) );
  NAND2X0 U11718 ( .IN1(n11539), .IN2(n11540), .QN(g33026) );
  NAND2X0 U11719 ( .IN1(n11541), .IN2(n11525), .QN(n11540) );
  NAND2X0 U11720 ( .IN1(n101), .IN2(n11542), .QN(n11541) );
  NAND2X0 U11721 ( .IN1(n11543), .IN2(n8917), .QN(n11542) );
  NAND2X0 U11722 ( .IN1(n9049), .IN2(g3506), .QN(n11539) );
  NAND3X0 U11723 ( .IN1(n11544), .IN2(n11545), .IN3(n11546), .QN(g33024) );
  NAND2X0 U11724 ( .IN1(g25648), .IN2(n11547), .QN(n11546) );
  NAND2X0 U11725 ( .IN1(n9049), .IN2(g3171), .QN(n11545) );
  NAND3X0 U11726 ( .IN1(n11548), .IN2(n11549), .IN3(n8879), .QN(n11544) );
  NAND2X0 U11727 ( .IN1(n11550), .IN2(n526), .QN(n11548) );
  NAND2X0 U11728 ( .IN1(n11551), .IN2(n11552), .QN(g33023) );
  NAND3X0 U11729 ( .IN1(n8893), .IN2(g3171), .IN3(n11547), .QN(n11552) );
  NAND2X0 U11730 ( .IN1(n11553), .IN2(g3167), .QN(n11551) );
  NAND2X0 U11731 ( .IN1(n11554), .IN2(n8917), .QN(n11553) );
  NAND2X0 U11732 ( .IN1(n5603), .IN2(n11549), .QN(n11554) );
  NAND2X0 U11733 ( .IN1(n11555), .IN2(n11556), .QN(g33022) );
  NAND2X0 U11734 ( .IN1(n11547), .IN2(n11557), .QN(n11556) );
  INVX0 U11735 ( .INP(n11558), .ZN(n11547) );
  NAND2X0 U11736 ( .IN1(n9048), .IN2(g3161), .QN(n11555) );
  NAND2X0 U11737 ( .IN1(n11559), .IN2(n11560), .QN(g33021) );
  NAND2X0 U11738 ( .IN1(n11561), .IN2(n11549), .QN(n11560) );
  NAND2X0 U11739 ( .IN1(n113), .IN2(n11562), .QN(n11561) );
  NAND2X0 U11740 ( .IN1(n11563), .IN2(n8917), .QN(n11562) );
  NAND2X0 U11741 ( .IN1(n9048), .IN2(g3155), .QN(n11559) );
  NAND3X0 U11742 ( .IN1(n11564), .IN2(n11565), .IN3(n9200), .QN(g33019) );
  NAND2X0 U11743 ( .IN1(n9047), .IN2(g2748), .QN(n11565) );
  NAND2X0 U11744 ( .IN1(n11566), .IN2(n8917), .QN(n11564) );
  XOR2X1 U11745 ( .IN1(test_so30), .IN2(n2790), .Q(n11566) );
  NAND4X0 U11746 ( .IN1(n11567), .IN2(n11568), .IN3(n11569), .IN4(n11570), 
        .QN(g33018) );
  NAND2X0 U11747 ( .IN1(n9048), .IN2(g2610), .QN(n11570) );
  NAND4X0 U11748 ( .IN1(n3511), .IN2(n10989), .IN3(n11571), .IN4(n8482), .QN(
        n11569) );
  NOR2X0 U11749 ( .IN1(n5508), .IN2(n11572), .QN(n11571) );
  NAND3X0 U11750 ( .IN1(n3512), .IN2(n11573), .IN3(n3517), .QN(n11568) );
  INVX0 U11751 ( .INP(n3513), .ZN(n11573) );
  NAND2X0 U11752 ( .IN1(n3524), .IN2(n10239), .QN(n3513) );
  INVX0 U11753 ( .INP(n3006), .ZN(n10239) );
  NAND3X0 U11754 ( .IN1(g2619), .IN2(g110), .IN3(n8482), .QN(n3512) );
  NAND2X0 U11755 ( .IN1(test_so40), .IN2(n11574), .QN(n11567) );
  NAND3X0 U11756 ( .IN1(n11575), .IN2(n10991), .IN3(n11576), .QN(n11574) );
  NAND2X0 U11757 ( .IN1(n3006), .IN2(n8917), .QN(n11576) );
  NAND2X0 U11758 ( .IN1(n3525), .IN2(n3505), .QN(n3006) );
  NAND4X0 U11759 ( .IN1(n11577), .IN2(n11578), .IN3(n11579), .IN4(n11580), 
        .QN(g33017) );
  NAND2X0 U11760 ( .IN1(n11581), .IN2(g2619), .QN(n11579) );
  NAND2X0 U11761 ( .IN1(n3517), .IN2(g2610), .QN(n11578) );
  NAND2X0 U11762 ( .IN1(test_so40), .IN2(n9054), .QN(n11577) );
  NAND3X0 U11763 ( .IN1(n11582), .IN2(n11583), .IN3(n11580), .QN(g33016) );
  NAND2X0 U11764 ( .IN1(n11581), .IN2(g2610), .QN(n11583) );
  NAND2X0 U11765 ( .IN1(n11575), .IN2(g2587), .QN(n11582) );
  NAND4X0 U11766 ( .IN1(n11584), .IN2(n11585), .IN3(n11586), .IN4(n11580), 
        .QN(g33015) );
  INVX0 U11767 ( .INP(n3519), .ZN(n11580) );
  NAND3X0 U11768 ( .IN1(n5508), .IN2(n11587), .IN3(n3517), .QN(n11586) );
  NAND2X0 U11769 ( .IN1(n11581), .IN2(g2587), .QN(n11585) );
  NAND2X0 U11770 ( .IN1(test_so34), .IN2(n9054), .QN(n11584) );
  NAND4X0 U11771 ( .IN1(n11588), .IN2(n11589), .IN3(n11590), .IN4(n11591), 
        .QN(g33014) );
  NAND2X0 U11772 ( .IN1(n9047), .IN2(g2476), .QN(n11591) );
  NAND4X0 U11773 ( .IN1(n3530), .IN2(n10989), .IN3(n11592), .IN4(n8481), .QN(
        n11590) );
  NOR2X0 U11774 ( .IN1(n5509), .IN2(n11593), .QN(n11592) );
  NAND3X0 U11775 ( .IN1(n3531), .IN2(n11594), .IN3(n3536), .QN(n11589) );
  INVX0 U11776 ( .INP(n3532), .ZN(n11594) );
  NAND2X0 U11777 ( .IN1(n3524), .IN2(n10238), .QN(n3532) );
  INVX0 U11778 ( .INP(n3007), .ZN(n10238) );
  NAND3X0 U11779 ( .IN1(g2485), .IN2(g110), .IN3(n8481), .QN(n3531) );
  NAND2X0 U11780 ( .IN1(n11595), .IN2(g2491), .QN(n11588) );
  NAND3X0 U11781 ( .IN1(n11596), .IN2(n10991), .IN3(n11597), .QN(n11595) );
  NAND2X0 U11782 ( .IN1(n3007), .IN2(n8917), .QN(n11597) );
  NAND3X0 U11783 ( .IN1(n5349), .IN2(g2748), .IN3(n3525), .QN(n3007) );
  NAND4X0 U11784 ( .IN1(n11598), .IN2(n11599), .IN3(n11600), .IN4(n11601), 
        .QN(g33013) );
  NAND2X0 U11785 ( .IN1(n11602), .IN2(g2485), .QN(n11600) );
  NAND2X0 U11786 ( .IN1(n3536), .IN2(g2476), .QN(n11599) );
  NAND2X0 U11787 ( .IN1(n9047), .IN2(g2491), .QN(n11598) );
  NAND3X0 U11788 ( .IN1(n11603), .IN2(n11604), .IN3(n11601), .QN(g33012) );
  NAND2X0 U11789 ( .IN1(n11602), .IN2(g2476), .QN(n11604) );
  NAND2X0 U11790 ( .IN1(n11596), .IN2(g2453), .QN(n11603) );
  NAND4X0 U11791 ( .IN1(n11605), .IN2(n11606), .IN3(n11607), .IN4(n11601), 
        .QN(g33011) );
  INVX0 U11792 ( .INP(n3538), .ZN(n11601) );
  NAND3X0 U11793 ( .IN1(n5509), .IN2(n11608), .IN3(n3536), .QN(n11607) );
  NAND2X0 U11794 ( .IN1(n11602), .IN2(g2453), .QN(n11606) );
  NAND2X0 U11795 ( .IN1(n9047), .IN2(g2461), .QN(n11605) );
  NAND4X0 U11796 ( .IN1(n11609), .IN2(n11610), .IN3(n11611), .IN4(n11612), 
        .QN(g33010) );
  NAND2X0 U11797 ( .IN1(test_so21), .IN2(n9054), .QN(n11612) );
  NAND4X0 U11798 ( .IN1(n3548), .IN2(n10989), .IN3(n11613), .IN4(n8591), .QN(
        n11611) );
  NOR2X0 U11799 ( .IN1(n5511), .IN2(n11614), .QN(n11613) );
  NAND3X0 U11800 ( .IN1(n3549), .IN2(n11615), .IN3(n3555), .QN(n11610) );
  INVX0 U11801 ( .INP(n3551), .ZN(n11615) );
  NAND2X0 U11802 ( .IN1(n3524), .IN2(n10237), .QN(n3551) );
  INVX0 U11803 ( .INP(n3550), .ZN(n10237) );
  NAND3X0 U11804 ( .IN1(g110), .IN2(n8591), .IN3(g2351), .QN(n3549) );
  NAND2X0 U11805 ( .IN1(n11616), .IN2(g2357), .QN(n11609) );
  NAND3X0 U11806 ( .IN1(n11617), .IN2(n10991), .IN3(n11618), .QN(n11616) );
  NAND2X0 U11807 ( .IN1(n3550), .IN2(n8918), .QN(n11618) );
  NAND3X0 U11808 ( .IN1(n5516), .IN2(g2741), .IN3(n3525), .QN(n3550) );
  NAND4X0 U11809 ( .IN1(n11619), .IN2(n11620), .IN3(n11621), .IN4(n11622), 
        .QN(g33009) );
  NAND2X0 U11810 ( .IN1(n11623), .IN2(g2351), .QN(n11621) );
  NAND2X0 U11811 ( .IN1(n3555), .IN2(test_so21), .QN(n11620) );
  NAND2X0 U11812 ( .IN1(n9047), .IN2(g2357), .QN(n11619) );
  NAND3X0 U11813 ( .IN1(n11624), .IN2(n11625), .IN3(n11622), .QN(g33008) );
  NAND2X0 U11814 ( .IN1(n11623), .IN2(test_so21), .QN(n11625) );
  NAND2X0 U11815 ( .IN1(n11617), .IN2(g2319), .QN(n11624) );
  NAND4X0 U11816 ( .IN1(n11626), .IN2(n11627), .IN3(n11628), .IN4(n11622), 
        .QN(g33007) );
  INVX0 U11817 ( .INP(n3557), .ZN(n11622) );
  NAND3X0 U11818 ( .IN1(n5511), .IN2(n11629), .IN3(n3555), .QN(n11628) );
  NAND2X0 U11819 ( .IN1(n11623), .IN2(g2319), .QN(n11627) );
  NAND2X0 U11820 ( .IN1(n9046), .IN2(g2327), .QN(n11626) );
  NAND4X0 U11821 ( .IN1(n11630), .IN2(n11631), .IN3(n11632), .IN4(n11633), 
        .QN(g33006) );
  NAND2X0 U11822 ( .IN1(n9046), .IN2(g2208), .QN(n11633) );
  NAND4X0 U11823 ( .IN1(n3567), .IN2(n10989), .IN3(n11634), .IN4(n8479), .QN(
        n11632) );
  NOR2X0 U11824 ( .IN1(n5512), .IN2(n11635), .QN(n11634) );
  NAND3X0 U11825 ( .IN1(n3568), .IN2(n11636), .IN3(n3574), .QN(n11631) );
  INVX0 U11826 ( .INP(n3570), .ZN(n11636) );
  NAND2X0 U11827 ( .IN1(n3524), .IN2(n10236), .QN(n3570) );
  INVX0 U11828 ( .INP(n3569), .ZN(n10236) );
  NAND3X0 U11829 ( .IN1(g2217), .IN2(g110), .IN3(n8479), .QN(n3568) );
  NAND2X0 U11830 ( .IN1(n11637), .IN2(g2223), .QN(n11630) );
  NAND3X0 U11831 ( .IN1(n11638), .IN2(n10991), .IN3(n11639), .QN(n11637) );
  NAND2X0 U11832 ( .IN1(n3569), .IN2(n8918), .QN(n11639) );
  NAND3X0 U11833 ( .IN1(n5516), .IN2(n5349), .IN3(n3525), .QN(n3569) );
  NAND4X0 U11834 ( .IN1(n11640), .IN2(n11641), .IN3(n11642), .IN4(n11643), 
        .QN(g33005) );
  NAND2X0 U11835 ( .IN1(n11644), .IN2(g2217), .QN(n11642) );
  NAND2X0 U11836 ( .IN1(n3574), .IN2(g2208), .QN(n11641) );
  NAND2X0 U11837 ( .IN1(n9046), .IN2(g2223), .QN(n11640) );
  NAND3X0 U11838 ( .IN1(n11645), .IN2(n11646), .IN3(n11643), .QN(g33004) );
  NAND2X0 U11839 ( .IN1(n11644), .IN2(g2208), .QN(n11646) );
  NAND2X0 U11840 ( .IN1(n11638), .IN2(g2185), .QN(n11645) );
  NAND4X0 U11841 ( .IN1(n11647), .IN2(n11648), .IN3(n11649), .IN4(n11643), 
        .QN(g33003) );
  INVX0 U11842 ( .INP(n3576), .ZN(n11643) );
  NAND3X0 U11843 ( .IN1(n5512), .IN2(n11650), .IN3(n3574), .QN(n11649) );
  NAND2X0 U11844 ( .IN1(n11644), .IN2(g2185), .QN(n11648) );
  NAND2X0 U11845 ( .IN1(n9046), .IN2(g2193), .QN(n11647) );
  NAND4X0 U11846 ( .IN1(n11651), .IN2(n11652), .IN3(n11653), .IN4(n11654), 
        .QN(g33002) );
  NAND2X0 U11847 ( .IN1(n9046), .IN2(g2051), .QN(n11654) );
  NAND4X0 U11848 ( .IN1(n3586), .IN2(n10989), .IN3(n11655), .IN4(n8483), .QN(
        n11653) );
  NOR2X0 U11849 ( .IN1(n5507), .IN2(n11656), .QN(n11655) );
  NAND3X0 U11850 ( .IN1(n3587), .IN2(n11657), .IN3(n3593), .QN(n11652) );
  INVX0 U11851 ( .INP(n3589), .ZN(n11657) );
  NAND2X0 U11852 ( .IN1(n3524), .IN2(n10232), .QN(n3589) );
  INVX0 U11853 ( .INP(n3588), .ZN(n10232) );
  NAND3X0 U11854 ( .IN1(g2060), .IN2(g110), .IN3(n8483), .QN(n3587) );
  NAND2X0 U11855 ( .IN1(n11658), .IN2(g2066), .QN(n11651) );
  NAND3X0 U11856 ( .IN1(n11659), .IN2(n10991), .IN3(n11660), .QN(n11658) );
  NAND2X0 U11857 ( .IN1(n3588), .IN2(n8918), .QN(n11660) );
  NAND3X0 U11858 ( .IN1(n811), .IN2(n5300), .IN3(n3505), .QN(n3588) );
  NAND4X0 U11859 ( .IN1(n11661), .IN2(n11662), .IN3(n11663), .IN4(n11664), 
        .QN(g33001) );
  NAND2X0 U11860 ( .IN1(n11665), .IN2(g2060), .QN(n11663) );
  NAND2X0 U11861 ( .IN1(n3593), .IN2(g2051), .QN(n11662) );
  NAND2X0 U11862 ( .IN1(n9046), .IN2(g2066), .QN(n11661) );
  NAND3X0 U11863 ( .IN1(n11666), .IN2(n11667), .IN3(n11664), .QN(g33000) );
  NAND2X0 U11864 ( .IN1(n11665), .IN2(g2051), .QN(n11667) );
  NAND2X0 U11865 ( .IN1(n11659), .IN2(g2028), .QN(n11666) );
  NAND4X0 U11866 ( .IN1(n11668), .IN2(n11669), .IN3(n11670), .IN4(n11664), 
        .QN(g32999) );
  INVX0 U11867 ( .INP(n3595), .ZN(n11664) );
  NAND3X0 U11868 ( .IN1(n5507), .IN2(n11671), .IN3(n3593), .QN(n11670) );
  NAND2X0 U11869 ( .IN1(n11665), .IN2(g2028), .QN(n11669) );
  NAND2X0 U11870 ( .IN1(test_so59), .IN2(n9055), .QN(n11668) );
  NAND4X0 U11871 ( .IN1(n11672), .IN2(n11673), .IN3(n11674), .IN4(n11675), 
        .QN(g32998) );
  NAND2X0 U11872 ( .IN1(n9045), .IN2(g1917), .QN(n11675) );
  NAND4X0 U11873 ( .IN1(n3604), .IN2(n10989), .IN3(n11676), .IN4(n8480), .QN(
        n11674) );
  NOR2X0 U11874 ( .IN1(n5510), .IN2(n11677), .QN(n11676) );
  NAND3X0 U11875 ( .IN1(n3605), .IN2(n11678), .IN3(n3611), .QN(n11673) );
  INVX0 U11876 ( .INP(n3607), .ZN(n11678) );
  NAND2X0 U11877 ( .IN1(n3524), .IN2(n10233), .QN(n3607) );
  INVX0 U11878 ( .INP(n3606), .ZN(n10233) );
  NAND3X0 U11879 ( .IN1(g1926), .IN2(g110), .IN3(n8480), .QN(n3605) );
  NAND2X0 U11880 ( .IN1(n11679), .IN2(g1932), .QN(n11672) );
  NAND3X0 U11881 ( .IN1(n11680), .IN2(n10991), .IN3(n11681), .QN(n11679) );
  NAND2X0 U11882 ( .IN1(n3606), .IN2(n8918), .QN(n11681) );
  NAND4X0 U11883 ( .IN1(n811), .IN2(n5349), .IN3(g2748), .IN4(n5300), .QN(
        n3606) );
  NAND4X0 U11884 ( .IN1(n11682), .IN2(n11683), .IN3(n11684), .IN4(n11685), 
        .QN(g32997) );
  NAND2X0 U11885 ( .IN1(n11686), .IN2(g1926), .QN(n11684) );
  NAND2X0 U11886 ( .IN1(n3611), .IN2(g1917), .QN(n11683) );
  NAND2X0 U11887 ( .IN1(n9045), .IN2(g1932), .QN(n11682) );
  NAND3X0 U11888 ( .IN1(n11687), .IN2(n11688), .IN3(n11685), .QN(g32996) );
  NAND2X0 U11889 ( .IN1(n11686), .IN2(g1917), .QN(n11688) );
  NAND2X0 U11890 ( .IN1(n11680), .IN2(g1894), .QN(n11687) );
  NAND4X0 U11891 ( .IN1(n11689), .IN2(n11690), .IN3(n11691), .IN4(n11685), 
        .QN(g32995) );
  INVX0 U11892 ( .INP(n3613), .ZN(n11685) );
  NAND3X0 U11893 ( .IN1(n5510), .IN2(n11692), .IN3(n3611), .QN(n11691) );
  NAND2X0 U11894 ( .IN1(n11686), .IN2(g1894), .QN(n11690) );
  NAND2X0 U11895 ( .IN1(n9045), .IN2(g1902), .QN(n11689) );
  NAND4X0 U11896 ( .IN1(n11693), .IN2(n11694), .IN3(n11695), .IN4(n11696), 
        .QN(g32994) );
  NAND2X0 U11897 ( .IN1(n9042), .IN2(g1783), .QN(n11696) );
  NAND4X0 U11898 ( .IN1(n3622), .IN2(n10989), .IN3(n11697), .IN4(n5596), .QN(
        n11695) );
  NOR2X0 U11899 ( .IN1(n5359), .IN2(n11698), .QN(n11697) );
  NAND3X0 U11900 ( .IN1(n3623), .IN2(n11699), .IN3(n3628), .QN(n11694) );
  INVX0 U11901 ( .INP(n3624), .ZN(n11699) );
  NAND2X0 U11902 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  NAND3X0 U11903 ( .IN1(g1792), .IN2(g110), .IN3(n5596), .QN(n3623) );
  NAND2X0 U11904 ( .IN1(n11700), .IN2(g1798), .QN(n11693) );
  NAND3X0 U11905 ( .IN1(n11701), .IN2(n10991), .IN3(n11702), .QN(n11700) );
  NAND2X0 U11906 ( .IN1(n8905), .IN2(n1721), .QN(n11702) );
  INVX0 U11907 ( .INP(n3005), .ZN(n1721) );
  NAND4X0 U11908 ( .IN1(n11703), .IN2(n11704), .IN3(n11705), .IN4(n11706), 
        .QN(g32993) );
  NAND2X0 U11909 ( .IN1(n11707), .IN2(g1792), .QN(n11705) );
  NAND2X0 U11910 ( .IN1(n3628), .IN2(g1783), .QN(n11704) );
  NAND2X0 U11911 ( .IN1(n9045), .IN2(g1798), .QN(n11703) );
  NAND3X0 U11912 ( .IN1(n11708), .IN2(n11709), .IN3(n11706), .QN(g32992) );
  NAND2X0 U11913 ( .IN1(n11707), .IN2(g1783), .QN(n11709) );
  NAND2X0 U11914 ( .IN1(n11701), .IN2(g1760), .QN(n11708) );
  NAND4X0 U11915 ( .IN1(n11710), .IN2(n11711), .IN3(n11712), .IN4(n11706), 
        .QN(g32991) );
  INVX0 U11916 ( .INP(n3630), .ZN(n11706) );
  NAND3X0 U11917 ( .IN1(n5359), .IN2(n11713), .IN3(n3628), .QN(n11712) );
  NAND2X0 U11918 ( .IN1(n11707), .IN2(g1760), .QN(n11711) );
  NAND2X0 U11919 ( .IN1(n9044), .IN2(g1768), .QN(n11710) );
  NAND4X0 U11920 ( .IN1(n11714), .IN2(n11715), .IN3(n11716), .IN4(n11717), 
        .QN(g32990) );
  NAND2X0 U11921 ( .IN1(test_so94), .IN2(n9055), .QN(n11717) );
  NAND4X0 U11922 ( .IN1(n3640), .IN2(n10989), .IN3(n11718), .IN4(n8596), .QN(
        n11716) );
  NOR2X0 U11923 ( .IN1(n5525), .IN2(n11719), .QN(n11718) );
  INVX0 U11924 ( .INP(n9218), .ZN(n10989) );
  NAND2X0 U11925 ( .IN1(n2760), .IN2(n8918), .QN(n9218) );
  NAND3X0 U11926 ( .IN1(n3641), .IN2(n11720), .IN3(n3646), .QN(n11715) );
  INVX0 U11927 ( .INP(n3642), .ZN(n11720) );
  NAND2X0 U11928 ( .IN1(n3524), .IN2(n10240), .QN(n3642) );
  INVX0 U11929 ( .INP(n3003), .ZN(n10240) );
  NAND3X0 U11930 ( .IN1(g110), .IN2(n8596), .IN3(g1657), .QN(n3641) );
  NAND2X0 U11931 ( .IN1(n11721), .IN2(g1664), .QN(n11714) );
  NAND3X0 U11932 ( .IN1(n10991), .IN2(n11722), .IN3(n11723), .QN(n11721) );
  NAND2X0 U11933 ( .IN1(n3003), .IN2(n8918), .QN(n11723) );
  NAND2X0 U11934 ( .IN1(n3653), .IN2(n811), .QN(n3003) );
  INVX0 U11935 ( .INP(n11724), .ZN(n811) );
  NAND2X0 U11936 ( .IN1(n11725), .IN2(n11726), .QN(n11724) );
  XOR2X1 U11937 ( .IN1(n8052), .IN2(g73), .Q(n11726) );
  XOR2X1 U11938 ( .IN1(n8051), .IN2(g72), .Q(n11725) );
  NAND2X0 U11939 ( .IN1(n8905), .IN2(n1782), .QN(n10991) );
  INVX0 U11940 ( .INP(n2760), .ZN(n1782) );
  NAND4X0 U11941 ( .IN1(n11727), .IN2(n11728), .IN3(n11729), .IN4(n11730), 
        .QN(g32989) );
  NAND2X0 U11942 ( .IN1(n11731), .IN2(g1657), .QN(n11729) );
  NAND2X0 U11943 ( .IN1(n3646), .IN2(test_so94), .QN(n11728) );
  NAND2X0 U11944 ( .IN1(n9044), .IN2(g1664), .QN(n11727) );
  NAND3X0 U11945 ( .IN1(n11732), .IN2(n11733), .IN3(n11730), .QN(g32988) );
  NAND2X0 U11946 ( .IN1(n11731), .IN2(test_so94), .QN(n11733) );
  NAND2X0 U11947 ( .IN1(n11722), .IN2(g1624), .QN(n11732) );
  NAND4X0 U11948 ( .IN1(n11734), .IN2(n11735), .IN3(n11736), .IN4(n11730), 
        .QN(g32987) );
  INVX0 U11949 ( .INP(n3648), .ZN(n11730) );
  NAND3X0 U11950 ( .IN1(n5525), .IN2(n11737), .IN3(n3646), .QN(n11736) );
  NAND2X0 U11951 ( .IN1(n11731), .IN2(g1624), .QN(n11735) );
  NAND2X0 U11952 ( .IN1(n9044), .IN2(g1632), .QN(n11734) );
  NAND3X0 U11953 ( .IN1(n11738), .IN2(n11739), .IN3(n11740), .QN(g32986) );
  NAND3X0 U11954 ( .IN1(n11303), .IN2(n8172), .IN3(n11741), .QN(n11740) );
  INVX0 U11955 ( .INP(n11742), .ZN(n11303) );
  NAND3X0 U11956 ( .IN1(n11742), .IN2(g1373), .IN3(n8880), .QN(n11739) );
  NAND2X0 U11957 ( .IN1(n198), .IN2(n11743), .QN(n11742) );
  NAND2X0 U11958 ( .IN1(n8156), .IN2(n11305), .QN(n11743) );
  INVX0 U11959 ( .INP(n11744), .ZN(n198) );
  NAND2X0 U11960 ( .IN1(n9044), .IN2(g1367), .QN(n11738) );
  NOR2X0 U11961 ( .IN1(n5730), .IN2(n11745), .QN(g32985) );
  NOR2X0 U11962 ( .IN1(n8954), .IN2(n11746), .QN(n11745) );
  NOR2X0 U11963 ( .IN1(n9698), .IN2(n11312), .QN(n11746) );
  NAND2X0 U11964 ( .IN1(n3662), .IN2(g1270), .QN(n11312) );
  NAND3X0 U11965 ( .IN1(n11747), .IN2(n11748), .IN3(n11749), .QN(g32984) );
  NAND2X0 U11966 ( .IN1(n9044), .IN2(g1263), .QN(n11749) );
  NAND3X0 U11967 ( .IN1(n11311), .IN2(n11750), .IN3(g1270), .QN(n11748) );
  INVX0 U11968 ( .INP(n3662), .ZN(n11750) );
  NAND2X0 U11969 ( .IN1(n5716), .IN2(n3662), .QN(n11747) );
  NAND3X0 U11970 ( .IN1(n11751), .IN2(n11752), .IN3(n11753), .QN(g32983) );
  NAND3X0 U11971 ( .IN1(n11317), .IN2(n8174), .IN3(n11754), .QN(n11753) );
  INVX0 U11972 ( .INP(n11755), .ZN(n11317) );
  NAND3X0 U11973 ( .IN1(n11755), .IN2(g1030), .IN3(n8880), .QN(n11752) );
  NAND2X0 U11974 ( .IN1(n542), .IN2(n11756), .QN(n11755) );
  NAND2X0 U11975 ( .IN1(n8157), .IN2(n11319), .QN(n11756) );
  INVX0 U11976 ( .INP(n11757), .ZN(n542) );
  NAND2X0 U11977 ( .IN1(n9044), .IN2(g1024), .QN(n11751) );
  NOR2X0 U11978 ( .IN1(n5731), .IN2(n11758), .QN(g32982) );
  NOR2X0 U11979 ( .IN1(n8954), .IN2(n11759), .QN(n11758) );
  NOR2X0 U11980 ( .IN1(n9697), .IN2(n11326), .QN(n11759) );
  NAND2X0 U11981 ( .IN1(n3671), .IN2(g925), .QN(n11326) );
  NAND3X0 U11982 ( .IN1(n11760), .IN2(n11761), .IN3(n11762), .QN(g32981) );
  NAND2X0 U11983 ( .IN1(n9043), .IN2(g918), .QN(n11762) );
  NAND3X0 U11984 ( .IN1(n11325), .IN2(n11763), .IN3(g925), .QN(n11761) );
  INVX0 U11985 ( .INP(n3671), .ZN(n11763) );
  NAND2X0 U11986 ( .IN1(n5725), .IN2(n3671), .QN(n11760) );
  NOR3X0 U11987 ( .IN1(n8926), .IN2(n11764), .IN3(n11765), .QN(g32980) );
  NOR2X0 U11988 ( .IN1(n11766), .IN2(n10042), .QN(n11765) );
  INVX0 U11989 ( .INP(n2644), .ZN(n10042) );
  NOR2X0 U11990 ( .IN1(n10041), .IN2(g854), .QN(n11764) );
  INVX0 U11991 ( .INP(n11766), .ZN(n10041) );
  NAND4X0 U11992 ( .IN1(n5632), .IN2(g376), .IN3(g8719), .IN4(g370), .QN(
        n11766) );
  NAND3X0 U11993 ( .IN1(n11767), .IN2(n11768), .IN3(n11769), .QN(g32979) );
  NAND2X0 U11994 ( .IN1(test_so2), .IN2(n9055), .QN(n11769) );
  NAND3X0 U11995 ( .IN1(n2404), .IN2(n11770), .IN3(g758), .QN(n11768) );
  INVX0 U11996 ( .INP(n3272), .ZN(n11770) );
  NAND2X0 U11997 ( .IN1(n3272), .IN2(n5331), .QN(n11767) );
  NAND3X0 U11998 ( .IN1(n11771), .IN2(n11772), .IN3(n11773), .QN(g32978) );
  NAND2X0 U11999 ( .IN1(n9043), .IN2(g582), .QN(n11773) );
  NAND3X0 U12000 ( .IN1(n2421), .IN2(n11774), .IN3(g590), .QN(n11772) );
  INVX0 U12001 ( .INP(n3274), .ZN(n11774) );
  NAND2X0 U12002 ( .IN1(n3274), .IN2(n5472), .QN(n11771) );
  NAND3X0 U12003 ( .IN1(n11775), .IN2(n11776), .IN3(n11777), .QN(g32977) );
  NAND2X0 U12004 ( .IN1(test_so51), .IN2(n9055), .QN(n11777) );
  NAND3X0 U12005 ( .IN1(n8568), .IN2(n11778), .IN3(g291), .QN(n11776) );
  NAND2X0 U12006 ( .IN1(n53), .IN2(n5679), .QN(n11775) );
  INVX0 U12007 ( .INP(n11778), .ZN(n53) );
  NAND3X0 U12008 ( .IN1(test_so51), .IN2(n11779), .IN3(test_so55), .QN(n11778)
         );
  NAND3X0 U12009 ( .IN1(n11780), .IN2(n11781), .IN3(n11782), .QN(g32976) );
  NAND2X0 U12010 ( .IN1(n9043), .IN2(g164), .QN(n11782) );
  NAND3X0 U12011 ( .IN1(n10217), .IN2(n11783), .IN3(g150), .QN(n11781) );
  INVX0 U12012 ( .INP(n3281), .ZN(n11783) );
  NAND2X0 U12013 ( .IN1(n3281), .IN2(n5676), .QN(n11780) );
  NOR4X0 U12014 ( .IN1(n11784), .IN2(n11785), .IN3(n11786), .IN4(n11787), .QN(
        g32185) );
  NOR2X0 U12015 ( .IN1(n8546), .IN2(n8616), .QN(n11787) );
  NOR2X0 U12016 ( .IN1(n8460), .IN2(n8459), .QN(n11786) );
  INVX0 U12017 ( .INP(n11788), .ZN(n11785) );
  NAND2X0 U12018 ( .IN1(g2965), .IN2(test_so22), .QN(n11788) );
  NAND4X0 U12019 ( .IN1(n11789), .IN2(n11790), .IN3(n11791), .IN4(n11792), 
        .QN(n11784) );
  NAND2X0 U12020 ( .IN1(g2975), .IN2(g2970), .QN(n11792) );
  NAND2X0 U12021 ( .IN1(g2950), .IN2(g2955), .QN(n11791) );
  NAND2X0 U12022 ( .IN1(g2912), .IN2(g2917), .QN(n11790) );
  NAND2X0 U12023 ( .IN1(g2922), .IN2(g2927), .QN(n11789) );
  NAND4X0 U12024 ( .IN1(n11793), .IN2(n11794), .IN3(n11795), .IN4(n11796), 
        .QN(g31904) );
  NAND4X0 U12025 ( .IN1(n11797), .IN2(n11798), .IN3(n11475), .IN4(g5033), .QN(
        n11796) );
  NAND2X0 U12026 ( .IN1(n8518), .IN2(n11799), .QN(n11795) );
  INVX0 U12027 ( .INP(n11798), .ZN(n11799) );
  NAND2X0 U12028 ( .IN1(n9043), .IN2(g5029), .QN(n11794) );
  NAND2X0 U12029 ( .IN1(n11800), .IN2(n8918), .QN(n11793) );
  NAND4X0 U12030 ( .IN1(n11801), .IN2(n11473), .IN3(n11802), .IN4(n11803), 
        .QN(g31903) );
  NAND4X0 U12031 ( .IN1(n11804), .IN2(n11805), .IN3(n11475), .IN4(g5052), .QN(
        n11803) );
  INVX0 U12032 ( .INP(n11806), .ZN(n11805) );
  INVX0 U12033 ( .INP(n11476), .ZN(n11804) );
  NAND2X0 U12034 ( .IN1(n5607), .IN2(n11476), .QN(n11802) );
  NOR2X0 U12035 ( .IN1(n11807), .IN2(n5578), .QN(n11476) );
  NAND3X0 U12036 ( .IN1(n11806), .IN2(n8871), .IN3(n5607), .QN(n11473) );
  NAND2X0 U12037 ( .IN1(n9042), .IN2(g5046), .QN(n11801) );
  NAND3X0 U12038 ( .IN1(n11808), .IN2(n11809), .IN3(n11810), .QN(g31902) );
  NAND2X0 U12039 ( .IN1(n11811), .IN2(n8918), .QN(n11810) );
  INVX0 U12040 ( .INP(n11797), .ZN(n11811) );
  NAND4X0 U12041 ( .IN1(n11475), .IN2(g5029), .IN3(n11812), .IN4(n11813), .QN(
        n11809) );
  NAND2X0 U12042 ( .IN1(n5369), .IN2(g5022), .QN(n11813) );
  NAND2X0 U12043 ( .IN1(g5016), .IN2(g5062), .QN(n11812) );
  NAND2X0 U12044 ( .IN1(n11814), .IN2(g5016), .QN(n11808) );
  NAND2X0 U12045 ( .IN1(n11815), .IN2(n8918), .QN(n11814) );
  NAND2X0 U12046 ( .IN1(n5601), .IN2(g5062), .QN(n11815) );
  NAND4X0 U12047 ( .IN1(n11816), .IN2(n11817), .IN3(n11818), .IN4(n11819), 
        .QN(g31901) );
  NAND4X0 U12048 ( .IN1(n11820), .IN2(n11807), .IN3(n11475), .IN4(g5046), .QN(
        n11819) );
  NAND2X0 U12049 ( .IN1(n11821), .IN2(n5578), .QN(n11818) );
  INVX0 U12050 ( .INP(n11807), .ZN(n11821) );
  NAND3X0 U12051 ( .IN1(g5041), .IN2(g5037), .IN3(n11822), .QN(n11807) );
  NAND2X0 U12052 ( .IN1(n9042), .IN2(g5041), .QN(n11817) );
  NAND2X0 U12053 ( .IN1(n11806), .IN2(n8918), .QN(n11816) );
  NOR2X0 U12054 ( .IN1(n11820), .IN2(g5046), .QN(n11806) );
  NAND3X0 U12055 ( .IN1(n5605), .IN2(n11800), .IN3(n5611), .QN(n11820) );
  NAND3X0 U12056 ( .IN1(n11823), .IN2(n11824), .IN3(n11825), .QN(g31900) );
  NAND2X0 U12057 ( .IN1(n11826), .IN2(n5605), .QN(n11825) );
  INVX0 U12058 ( .INP(n11827), .ZN(n11826) );
  NAND4X0 U12059 ( .IN1(n11828), .IN2(g5041), .IN3(n11475), .IN4(n5611), .QN(
        n11824) );
  NAND2X0 U12060 ( .IN1(n11829), .IN2(g5037), .QN(n11823) );
  NAND3X0 U12061 ( .IN1(n11830), .IN2(n11831), .IN3(n8880), .QN(n11829) );
  NAND3X0 U12062 ( .IN1(n11832), .IN2(n11833), .IN3(g5041), .QN(n11831) );
  INVX0 U12063 ( .INP(n11834), .ZN(n11832) );
  NAND2X0 U12064 ( .IN1(n5605), .IN2(n11822), .QN(n11830) );
  NAND4X0 U12065 ( .IN1(n11835), .IN2(n11827), .IN3(n11836), .IN4(n11837), 
        .QN(g31899) );
  NAND4X0 U12066 ( .IN1(n11828), .IN2(n11833), .IN3(n11475), .IN4(g5037), .QN(
        n11837) );
  INVX0 U12067 ( .INP(n11822), .ZN(n11833) );
  INVX0 U12068 ( .INP(n11800), .ZN(n11828) );
  NAND2X0 U12069 ( .IN1(n5611), .IN2(n11822), .QN(n11836) );
  NOR2X0 U12070 ( .IN1(n11798), .IN2(n8518), .QN(n11822) );
  NAND3X0 U12071 ( .IN1(g5029), .IN2(g5062), .IN3(g5016), .QN(n11798) );
  NAND3X0 U12072 ( .IN1(n11800), .IN2(n8871), .IN3(n5611), .QN(n11827) );
  NOR2X0 U12073 ( .IN1(g5033), .IN2(n11797), .QN(n11800) );
  NAND3X0 U12074 ( .IN1(n5369), .IN2(g5022), .IN3(n5601), .QN(n11797) );
  NAND2X0 U12075 ( .IN1(n9042), .IN2(g5033), .QN(n11835) );
  NAND3X0 U12076 ( .IN1(n11838), .IN2(n11839), .IN3(n11840), .QN(g31898) );
  NAND3X0 U12077 ( .IN1(n11475), .IN2(n11841), .IN3(n5369), .QN(n11840) );
  NOR2X0 U12078 ( .IN1(n11834), .IN2(n8941), .QN(n11475) );
  NAND2X0 U12079 ( .IN1(n11842), .IN2(n11843), .QN(n11834) );
  NAND3X0 U12080 ( .IN1(n11844), .IN2(g5016), .IN3(n8880), .QN(n11839) );
  INVX0 U12081 ( .INP(n11841), .ZN(n11844) );
  NAND2X0 U12082 ( .IN1(n8498), .IN2(n8496), .QN(n11841) );
  NAND2X0 U12083 ( .IN1(n9042), .IN2(g5022), .QN(n11838) );
  NAND3X0 U12084 ( .IN1(n11845), .IN2(n10920), .IN3(n11846), .QN(g31897) );
  NAND2X0 U12085 ( .IN1(n11484), .IN2(g4575), .QN(n10920) );
  NAND2X0 U12086 ( .IN1(n9042), .IN2(g4423), .QN(n11845) );
  NAND3X0 U12087 ( .IN1(n11847), .IN2(n10925), .IN3(n11846), .QN(g31896) );
  INVX0 U12088 ( .INP(n11848), .ZN(n11846) );
  NAND2X0 U12089 ( .IN1(n11849), .IN2(n11850), .QN(n11848) );
  NAND2X0 U12090 ( .IN1(n11484), .IN2(n11851), .QN(n11850) );
  NAND2X0 U12091 ( .IN1(g72), .IN2(g73), .QN(n11851) );
  NAND2X0 U12092 ( .IN1(n10926), .IN2(g4372), .QN(n11849) );
  INVX0 U12093 ( .INP(n11852), .ZN(n10926) );
  NAND2X0 U12094 ( .IN1(n11484), .IN2(test_so100), .QN(n10925) );
  NOR2X0 U12095 ( .IN1(n8950), .IN2(n5670), .QN(n11484) );
  NAND2X0 U12096 ( .IN1(n9042), .IN2(g4477), .QN(n11847) );
  NAND3X0 U12097 ( .IN1(n11853), .IN2(n11854), .IN3(n11495), .QN(g31894) );
  NAND2X0 U12098 ( .IN1(n9041), .IN2(g4093), .QN(n11854) );
  NAND2X0 U12099 ( .IN1(n11855), .IN2(n8918), .QN(n11853) );
  XOR2X1 U12100 ( .IN1(n11499), .IN2(g4098), .Q(n11855) );
  NOR2X0 U12101 ( .IN1(n3729), .IN2(n5340), .QN(n11499) );
  NAND2X0 U12102 ( .IN1(n11856), .IN2(g4087), .QN(n3729) );
  NAND2X0 U12103 ( .IN1(n11857), .IN2(n11858), .QN(g31872) );
  NAND2X0 U12104 ( .IN1(n11859), .IN2(n3730), .QN(n11858) );
  XOR2X1 U12105 ( .IN1(g2748), .IN2(n11860), .Q(n11859) );
  NOR2X0 U12106 ( .IN1(n5349), .IN2(n3506), .QN(n11860) );
  NAND2X0 U12107 ( .IN1(n9041), .IN2(g2741), .QN(n11857) );
  NAND3X0 U12108 ( .IN1(n11861), .IN2(n11862), .IN3(n11863), .QN(g31871) );
  NAND2X0 U12109 ( .IN1(n3733), .IN2(n11741), .QN(n11863) );
  NAND2X0 U12110 ( .IN1(n9041), .IN2(g1361), .QN(n11862) );
  NAND3X0 U12111 ( .IN1(n11744), .IN2(g1367), .IN3(n8880), .QN(n11861) );
  NAND2X0 U12112 ( .IN1(n199), .IN2(n11864), .QN(n11744) );
  NAND2X0 U12113 ( .IN1(n8171), .IN2(n11305), .QN(n11864) );
  INVX0 U12114 ( .INP(n11865), .ZN(n199) );
  NAND3X0 U12115 ( .IN1(n11866), .IN2(n11867), .IN3(n11868), .QN(g31870) );
  NAND2X0 U12116 ( .IN1(n9041), .IN2(g1259), .QN(n11868) );
  NAND3X0 U12117 ( .IN1(n11311), .IN2(n11869), .IN3(g1263), .QN(n11867) );
  INVX0 U12118 ( .INP(n3664), .ZN(n11869) );
  NAND2X0 U12119 ( .IN1(n3664), .IN2(n5674), .QN(n11866) );
  NAND3X0 U12120 ( .IN1(n11870), .IN2(n11871), .IN3(n11872), .QN(g31869) );
  NAND2X0 U12121 ( .IN1(n3738), .IN2(n11754), .QN(n11872) );
  NAND2X0 U12122 ( .IN1(n9041), .IN2(g1018), .QN(n11871) );
  NAND3X0 U12123 ( .IN1(n11757), .IN2(g1024), .IN3(n8880), .QN(n11870) );
  NAND2X0 U12124 ( .IN1(n543), .IN2(n11873), .QN(n11757) );
  NAND2X0 U12125 ( .IN1(n8173), .IN2(n11319), .QN(n11873) );
  INVX0 U12126 ( .INP(n11874), .ZN(n543) );
  NAND3X0 U12127 ( .IN1(n11875), .IN2(n11876), .IN3(n11877), .QN(g31868) );
  NAND2X0 U12128 ( .IN1(n9040), .IN2(g914), .QN(n11877) );
  NAND3X0 U12129 ( .IN1(n11325), .IN2(n11878), .IN3(g918), .QN(n11876) );
  INVX0 U12130 ( .INP(n3673), .ZN(n11878) );
  NAND2X0 U12131 ( .IN1(n3673), .IN2(n5673), .QN(n11875) );
  NAND3X0 U12132 ( .IN1(n11879), .IN2(n11880), .IN3(n11881), .QN(g31867) );
  NAND2X0 U12133 ( .IN1(n9040), .IN2(g744), .QN(n11881) );
  NAND3X0 U12134 ( .IN1(n2404), .IN2(test_so2), .IN3(n11882), .QN(n11880) );
  INVX0 U12135 ( .INP(n3682), .ZN(n11882) );
  NAND2X0 U12136 ( .IN1(n3682), .IN2(n5471), .QN(n11879) );
  NAND3X0 U12137 ( .IN1(n11883), .IN2(n11884), .IN3(n11885), .QN(g31866) );
  NAND2X0 U12138 ( .IN1(n9040), .IN2(g577), .QN(n11885) );
  NAND3X0 U12139 ( .IN1(n2421), .IN2(n11886), .IN3(g582), .QN(n11884) );
  INVX0 U12140 ( .INP(n3684), .ZN(n11886) );
  NAND2X0 U12141 ( .IN1(n3684), .IN2(n5552), .QN(n11883) );
  NAND2X0 U12142 ( .IN1(n11887), .IN2(n11888), .QN(g31865) );
  NAND2X0 U12143 ( .IN1(test_so55), .IN2(n11889), .QN(n11888) );
  NAND2X0 U12144 ( .IN1(n11890), .IN2(n8918), .QN(n11889) );
  NAND2X0 U12145 ( .IN1(n11779), .IN2(n8631), .QN(n11890) );
  INVX0 U12146 ( .INP(n11891), .ZN(n11779) );
  NAND3X0 U12147 ( .IN1(n8568), .IN2(test_so51), .IN3(n8607), .QN(n11887) );
  NAND3X0 U12148 ( .IN1(n11892), .IN2(n11893), .IN3(n11894), .QN(g31864) );
  NAND2X0 U12149 ( .IN1(test_so73), .IN2(n8926), .QN(n11894) );
  NAND3X0 U12150 ( .IN1(n10217), .IN2(n11895), .IN3(g164), .QN(n11893) );
  NAND2X0 U12151 ( .IN1(n56), .IN2(n5561), .QN(n11892) );
  INVX0 U12152 ( .INP(n11895), .ZN(n56) );
  NAND3X0 U12153 ( .IN1(n11896), .IN2(n11897), .IN3(test_so73), .QN(n11895) );
  INVX0 U12154 ( .INP(n11898), .ZN(n11896) );
  NAND2X0 U12155 ( .IN1(n11899), .IN2(n11900), .QN(g31793) );
  NAND2X0 U12156 ( .IN1(n11901), .IN2(n9727), .QN(n11900) );
  INVX0 U12157 ( .INP(n11902), .ZN(n9727) );
  NAND2X0 U12158 ( .IN1(n11903), .IN2(n8909), .QN(n11901) );
  NAND2X0 U12159 ( .IN1(n9726), .IN2(n11904), .QN(n11903) );
  NAND2X0 U12160 ( .IN1(n11905), .IN2(n11906), .QN(n11904) );
  NAND3X0 U12161 ( .IN1(n11907), .IN2(n11908), .IN3(n8071), .QN(n11906) );
  NAND2X0 U12162 ( .IN1(g6509), .IN2(n11909), .QN(n11908) );
  NAND4X0 U12163 ( .IN1(n8180), .IN2(n8179), .IN3(n8111), .IN4(n11910), .QN(
        n11905) );
  NAND2X0 U12164 ( .IN1(n11911), .IN2(n11912), .QN(n11910) );
  NAND3X0 U12165 ( .IN1(n11913), .IN2(n11914), .IN3(n8071), .QN(n11911) );
  NAND2X0 U12166 ( .IN1(n11915), .IN2(g6163), .QN(n11914) );
  NAND2X0 U12167 ( .IN1(g5817), .IN2(g5471), .QN(n11913) );
  NAND3X0 U12168 ( .IN1(n11916), .IN2(n11917), .IN3(n9728), .QN(n11899) );
  NOR4X0 U12169 ( .IN1(g5124), .IN2(n11912), .IN3(g6509), .IN4(n11909), .QN(
        n9728) );
  NAND2X0 U12170 ( .IN1(n8180), .IN2(n8179), .QN(n11909) );
  INVX0 U12171 ( .INP(n11907), .ZN(n11912) );
  NOR2X0 U12172 ( .IN1(g6163), .IN2(n11915), .QN(n11907) );
  NAND2X0 U12173 ( .IN1(n8080), .IN2(n8073), .QN(n11915) );
  NAND2X0 U12174 ( .IN1(n11902), .IN2(n11918), .QN(n11917) );
  INVX0 U12175 ( .INP(n9726), .ZN(n11918) );
  NOR2X0 U12176 ( .IN1(g3115), .IN2(g3466), .QN(n9726) );
  NAND2X0 U12177 ( .IN1(g3466), .IN2(g3115), .QN(n11916) );
  NAND2X0 U12178 ( .IN1(g113), .IN2(g2868), .QN(g31665) );
  NAND2X0 U12179 ( .IN1(g113), .IN2(g2873), .QN(g31656) );
  NAND3X0 U12180 ( .IN1(n11919), .IN2(n11920), .IN3(n11921), .QN(g30563) );
  NAND2X0 U12181 ( .IN1(n9040), .IN2(g6653), .QN(n11921) );
  NAND2X0 U12182 ( .IN1(n11922), .IN2(g6657), .QN(n11920) );
  NAND2X0 U12183 ( .IN1(n3765), .IN2(n10839), .QN(n11919) );
  NAND3X0 U12184 ( .IN1(n11923), .IN2(n11924), .IN3(n11925), .QN(g30562) );
  NAND2X0 U12185 ( .IN1(n11926), .IN2(n3765), .QN(n11925) );
  INVX0 U12186 ( .INP(n11927), .ZN(n11926) );
  NAND3X0 U12187 ( .IN1(n11927), .IN2(g6605), .IN3(n8881), .QN(n11924) );
  NAND2X0 U12188 ( .IN1(n11366), .IN2(g6561), .QN(n11927) );
  NAND2X0 U12189 ( .IN1(n9040), .IN2(g6649), .QN(n11923) );
  NAND3X0 U12190 ( .IN1(n11928), .IN2(n11929), .IN3(n11930), .QN(g30561) );
  NAND2X0 U12191 ( .IN1(n11931), .IN2(n3765), .QN(n11930) );
  INVX0 U12192 ( .INP(n11364), .ZN(n11931) );
  NAND3X0 U12193 ( .IN1(n11364), .IN2(g6597), .IN3(n8881), .QN(n11929) );
  NAND2X0 U12194 ( .IN1(n11932), .IN2(g6561), .QN(n11364) );
  NAND2X0 U12195 ( .IN1(n9040), .IN2(g6645), .QN(n11928) );
  NAND3X0 U12196 ( .IN1(n11933), .IN2(n11934), .IN3(n11935), .QN(g30560) );
  NAND2X0 U12197 ( .IN1(n11936), .IN2(n3765), .QN(n11935) );
  INVX0 U12198 ( .INP(n11937), .ZN(n11936) );
  NAND3X0 U12199 ( .IN1(n11937), .IN2(g6589), .IN3(n8881), .QN(n11934) );
  NAND2X0 U12200 ( .IN1(n11938), .IN2(g6561), .QN(n11937) );
  NAND2X0 U12201 ( .IN1(n9039), .IN2(g6641), .QN(n11933) );
  NAND3X0 U12202 ( .IN1(n11939), .IN2(n11940), .IN3(n11941), .QN(g30559) );
  NAND2X0 U12203 ( .IN1(n3774), .IN2(n11942), .QN(n11941) );
  NAND2X0 U12204 ( .IN1(n9039), .IN2(g6637), .QN(n11940) );
  NAND3X0 U12205 ( .IN1(n11943), .IN2(g6653), .IN3(n8881), .QN(n11939) );
  NAND2X0 U12206 ( .IN1(n11942), .IN2(n11375), .QN(n11943) );
  NAND3X0 U12207 ( .IN1(n11944), .IN2(n11945), .IN3(n11946), .QN(g30558) );
  NAND2X0 U12208 ( .IN1(n3774), .IN2(n11366), .QN(n11946) );
  NAND2X0 U12209 ( .IN1(n9039), .IN2(g6633), .QN(n11945) );
  NAND3X0 U12210 ( .IN1(n11947), .IN2(g6649), .IN3(n8881), .QN(n11944) );
  NAND2X0 U12211 ( .IN1(n11366), .IN2(n11375), .QN(n11947) );
  NAND3X0 U12212 ( .IN1(n11948), .IN2(n11949), .IN3(n11950), .QN(g30557) );
  NAND2X0 U12213 ( .IN1(n3774), .IN2(n11932), .QN(n11950) );
  NAND2X0 U12214 ( .IN1(n9039), .IN2(g6629), .QN(n11949) );
  NAND3X0 U12215 ( .IN1(n11951), .IN2(g6645), .IN3(n8881), .QN(n11948) );
  NAND2X0 U12216 ( .IN1(n11932), .IN2(n11375), .QN(n11951) );
  NAND3X0 U12217 ( .IN1(n11952), .IN2(n11953), .IN3(n11954), .QN(g30556) );
  NAND2X0 U12218 ( .IN1(n3774), .IN2(n11938), .QN(n11954) );
  NAND2X0 U12219 ( .IN1(n9039), .IN2(g6625), .QN(n11953) );
  NAND3X0 U12220 ( .IN1(n11955), .IN2(g6641), .IN3(n8881), .QN(n11952) );
  NAND2X0 U12221 ( .IN1(n11938), .IN2(n11375), .QN(n11955) );
  INVX0 U12222 ( .INP(n750), .ZN(n11375) );
  NAND2X0 U12223 ( .IN1(g6549), .IN2(g6555), .QN(n750) );
  NAND3X0 U12224 ( .IN1(n11956), .IN2(n11957), .IN3(n11958), .QN(g30555) );
  NAND2X0 U12225 ( .IN1(n3780), .IN2(n11942), .QN(n11958) );
  NAND2X0 U12226 ( .IN1(n9039), .IN2(g6621), .QN(n11957) );
  NAND3X0 U12227 ( .IN1(n11959), .IN2(g6637), .IN3(n8881), .QN(n11956) );
  NAND2X0 U12228 ( .IN1(n11942), .IN2(n11380), .QN(n11959) );
  NAND3X0 U12229 ( .IN1(n11960), .IN2(n11961), .IN3(n11962), .QN(g30554) );
  NAND2X0 U12230 ( .IN1(n3780), .IN2(n11366), .QN(n11962) );
  NAND2X0 U12231 ( .IN1(n9039), .IN2(g6617), .QN(n11961) );
  NAND3X0 U12232 ( .IN1(n11963), .IN2(g6633), .IN3(n8881), .QN(n11960) );
  NAND2X0 U12233 ( .IN1(n11366), .IN2(n11380), .QN(n11963) );
  NAND3X0 U12234 ( .IN1(n11964), .IN2(n11965), .IN3(n11966), .QN(g30553) );
  NAND2X0 U12235 ( .IN1(n3780), .IN2(n11932), .QN(n11966) );
  NAND2X0 U12236 ( .IN1(n9038), .IN2(g6613), .QN(n11965) );
  NAND3X0 U12237 ( .IN1(n11967), .IN2(g6629), .IN3(n8881), .QN(n11964) );
  NAND2X0 U12238 ( .IN1(n11932), .IN2(n11380), .QN(n11967) );
  NAND3X0 U12239 ( .IN1(n11968), .IN2(n11969), .IN3(n11970), .QN(g30552) );
  NAND2X0 U12240 ( .IN1(n3780), .IN2(n11938), .QN(n11970) );
  NAND2X0 U12241 ( .IN1(n9038), .IN2(g6609), .QN(n11969) );
  NAND3X0 U12242 ( .IN1(n11971), .IN2(g6625), .IN3(n8882), .QN(n11968) );
  NAND2X0 U12243 ( .IN1(n11938), .IN2(n11380), .QN(n11971) );
  INVX0 U12244 ( .INP(n752), .ZN(n11380) );
  NAND2X0 U12245 ( .IN1(n5571), .IN2(g6555), .QN(n752) );
  NAND3X0 U12246 ( .IN1(n11972), .IN2(n11973), .IN3(n11974), .QN(g30551) );
  NAND2X0 U12247 ( .IN1(n3785), .IN2(n11942), .QN(n11974) );
  NAND2X0 U12248 ( .IN1(n9038), .IN2(g6601), .QN(n11973) );
  NAND3X0 U12249 ( .IN1(n11975), .IN2(g6621), .IN3(n8882), .QN(n11972) );
  NAND2X0 U12250 ( .IN1(n11942), .IN2(n11976), .QN(n11975) );
  INVX0 U12251 ( .INP(n1409), .ZN(n11942) );
  NAND3X0 U12252 ( .IN1(n11977), .IN2(n11978), .IN3(n11979), .QN(g30550) );
  NAND2X0 U12253 ( .IN1(n3785), .IN2(n11366), .QN(n11979) );
  NAND2X0 U12254 ( .IN1(n9038), .IN2(g6593), .QN(n11978) );
  NAND3X0 U12255 ( .IN1(n11980), .IN2(g6617), .IN3(n8882), .QN(n11977) );
  NAND2X0 U12256 ( .IN1(n11366), .IN2(n11976), .QN(n11980) );
  INVX0 U12257 ( .INP(n1401), .ZN(n11366) );
  NAND2X0 U12258 ( .IN1(n5386), .IN2(g6573), .QN(n1401) );
  NAND3X0 U12259 ( .IN1(n11981), .IN2(n11982), .IN3(n11983), .QN(g30549) );
  NAND2X0 U12260 ( .IN1(n3785), .IN2(n11932), .QN(n11983) );
  NAND2X0 U12261 ( .IN1(test_so71), .IN2(n9055), .QN(n11982) );
  NAND3X0 U12262 ( .IN1(n11984), .IN2(g6613), .IN3(n8882), .QN(n11981) );
  NAND2X0 U12263 ( .IN1(n11932), .IN2(n11976), .QN(n11984) );
  INVX0 U12264 ( .INP(n1405), .ZN(n11932) );
  NAND2X0 U12265 ( .IN1(n5563), .IN2(g6565), .QN(n1405) );
  NAND3X0 U12266 ( .IN1(n11985), .IN2(n11986), .IN3(n11987), .QN(g30548) );
  NAND2X0 U12267 ( .IN1(n3785), .IN2(n11938), .QN(n11987) );
  NAND2X0 U12268 ( .IN1(n9038), .IN2(g6581), .QN(n11986) );
  NAND3X0 U12269 ( .IN1(n11988), .IN2(g6609), .IN3(n8882), .QN(n11985) );
  NAND2X0 U12270 ( .IN1(n11938), .IN2(n11976), .QN(n11988) );
  INVX0 U12271 ( .INP(n751), .ZN(n11976) );
  NAND2X0 U12272 ( .IN1(n8495), .IN2(g6549), .QN(n751) );
  INVX0 U12273 ( .INP(n1403), .ZN(n11938) );
  NAND2X0 U12274 ( .IN1(n5386), .IN2(n5563), .QN(n1403) );
  NAND3X0 U12275 ( .IN1(n11989), .IN2(n11990), .IN3(n11991), .QN(g30547) );
  NAND2X0 U12276 ( .IN1(n9038), .IN2(g6605), .QN(n11991) );
  NAND3X0 U12277 ( .IN1(n8896), .IN2(g6601), .IN3(n11992), .QN(n11990) );
  INVX0 U12278 ( .INP(n3790), .ZN(n11992) );
  NAND2X0 U12279 ( .IN1(n3790), .IN2(n3765), .QN(n11989) );
  NAND3X0 U12280 ( .IN1(n11993), .IN2(n11994), .IN3(n11995), .QN(g30546) );
  NAND2X0 U12281 ( .IN1(n9038), .IN2(g6597), .QN(n11995) );
  NAND3X0 U12282 ( .IN1(n8896), .IN2(g6593), .IN3(n11996), .QN(n11994) );
  INVX0 U12283 ( .INP(n3793), .ZN(n11996) );
  NAND2X0 U12284 ( .IN1(n3793), .IN2(n3765), .QN(n11993) );
  NAND3X0 U12285 ( .IN1(n11997), .IN2(n11998), .IN3(n11999), .QN(g30545) );
  NAND2X0 U12286 ( .IN1(n9037), .IN2(g6589), .QN(n11999) );
  NAND3X0 U12287 ( .IN1(test_so71), .IN2(n8870), .IN3(n12000), .QN(n11998) );
  INVX0 U12288 ( .INP(n3795), .ZN(n12000) );
  NAND2X0 U12289 ( .IN1(n3795), .IN2(n3765), .QN(n11997) );
  NAND3X0 U12290 ( .IN1(n12001), .IN2(n12002), .IN3(n12003), .QN(g30544) );
  NAND2X0 U12291 ( .IN1(n9037), .IN2(g6573), .QN(n12003) );
  NAND3X0 U12292 ( .IN1(n8896), .IN2(g6581), .IN3(n12004), .QN(n12002) );
  INVX0 U12293 ( .INP(n3797), .ZN(n12004) );
  NAND2X0 U12294 ( .IN1(n3797), .IN2(n3765), .QN(n12001) );
  NOR2X0 U12295 ( .IN1(g6549), .IN2(n11372), .QN(g30543) );
  NAND3X0 U12296 ( .IN1(n11362), .IN2(n8870), .IN3(n5646), .QN(n11372) );
  NAND2X0 U12297 ( .IN1(n3799), .IN2(n10829), .QN(n11362) );
  NAND3X0 U12298 ( .IN1(n12005), .IN2(n12006), .IN3(n12007), .QN(g30542) );
  NAND2X0 U12299 ( .IN1(n9037), .IN2(g6307), .QN(n12007) );
  NAND2X0 U12300 ( .IN1(n12008), .IN2(g6311), .QN(n12006) );
  NAND2X0 U12301 ( .IN1(n12009), .IN2(n3765), .QN(n12005) );
  NAND3X0 U12302 ( .IN1(n12010), .IN2(n12011), .IN3(n12012), .QN(g30541) );
  NAND2X0 U12303 ( .IN1(n12013), .IN2(n3765), .QN(n12012) );
  INVX0 U12304 ( .INP(n12014), .ZN(n12013) );
  NAND3X0 U12305 ( .IN1(n12014), .IN2(g6259), .IN3(n8882), .QN(n12011) );
  NAND2X0 U12306 ( .IN1(n11388), .IN2(g6215), .QN(n12014) );
  NAND2X0 U12307 ( .IN1(n9037), .IN2(g6303), .QN(n12010) );
  NAND3X0 U12308 ( .IN1(n12015), .IN2(n12016), .IN3(n12017), .QN(g30540) );
  NAND2X0 U12309 ( .IN1(n12018), .IN2(n3765), .QN(n12017) );
  INVX0 U12310 ( .INP(n11386), .ZN(n12018) );
  NAND3X0 U12311 ( .IN1(n11386), .IN2(g6251), .IN3(n8882), .QN(n12016) );
  NAND2X0 U12312 ( .IN1(n12019), .IN2(g6215), .QN(n11386) );
  NAND2X0 U12313 ( .IN1(n9037), .IN2(g6299), .QN(n12015) );
  NAND3X0 U12314 ( .IN1(n12020), .IN2(n12021), .IN3(n12022), .QN(g30539) );
  NAND2X0 U12315 ( .IN1(n12023), .IN2(n3765), .QN(n12022) );
  INVX0 U12316 ( .INP(n12024), .ZN(n12023) );
  NAND3X0 U12317 ( .IN1(n12024), .IN2(g6243), .IN3(n8882), .QN(n12021) );
  NAND2X0 U12318 ( .IN1(n12025), .IN2(g6215), .QN(n12024) );
  NAND2X0 U12319 ( .IN1(n9037), .IN2(g6295), .QN(n12020) );
  NAND3X0 U12320 ( .IN1(n12026), .IN2(n12027), .IN3(n12028), .QN(g30538) );
  NAND2X0 U12321 ( .IN1(n3808), .IN2(n12029), .QN(n12028) );
  NAND2X0 U12322 ( .IN1(n9037), .IN2(g6291), .QN(n12027) );
  NAND3X0 U12323 ( .IN1(n12030), .IN2(g6307), .IN3(n8882), .QN(n12026) );
  NAND2X0 U12324 ( .IN1(n11397), .IN2(n12029), .QN(n12030) );
  NAND3X0 U12325 ( .IN1(n12031), .IN2(n12032), .IN3(n12033), .QN(g30537) );
  NAND2X0 U12326 ( .IN1(n3808), .IN2(n11388), .QN(n12033) );
  NAND2X0 U12327 ( .IN1(n9036), .IN2(g6287), .QN(n12032) );
  NAND3X0 U12328 ( .IN1(n12034), .IN2(g6303), .IN3(n8882), .QN(n12031) );
  NAND2X0 U12329 ( .IN1(n11397), .IN2(n11388), .QN(n12034) );
  NAND3X0 U12330 ( .IN1(n12035), .IN2(n12036), .IN3(n12037), .QN(g30536) );
  NAND2X0 U12331 ( .IN1(n3808), .IN2(n12019), .QN(n12037) );
  NAND2X0 U12332 ( .IN1(n9036), .IN2(g6283), .QN(n12036) );
  NAND3X0 U12333 ( .IN1(n12038), .IN2(g6299), .IN3(n8882), .QN(n12035) );
  NAND2X0 U12334 ( .IN1(n11397), .IN2(n12019), .QN(n12038) );
  NAND3X0 U12335 ( .IN1(n12039), .IN2(n12040), .IN3(n12041), .QN(g30535) );
  NAND2X0 U12336 ( .IN1(n3808), .IN2(n12025), .QN(n12041) );
  NAND2X0 U12337 ( .IN1(n9036), .IN2(g6279), .QN(n12040) );
  NAND3X0 U12338 ( .IN1(n12042), .IN2(g6295), .IN3(n8882), .QN(n12039) );
  NAND2X0 U12339 ( .IN1(n11397), .IN2(n12025), .QN(n12042) );
  INVX0 U12340 ( .INP(n1009), .ZN(n11397) );
  NAND2X0 U12341 ( .IN1(g6203), .IN2(g6209), .QN(n1009) );
  NAND3X0 U12342 ( .IN1(n12043), .IN2(n12044), .IN3(n12045), .QN(g30534) );
  NAND2X0 U12343 ( .IN1(n3814), .IN2(n12029), .QN(n12045) );
  NAND2X0 U12344 ( .IN1(n9036), .IN2(g6275), .QN(n12044) );
  NAND3X0 U12345 ( .IN1(n12046), .IN2(g6291), .IN3(n8883), .QN(n12043) );
  NAND2X0 U12346 ( .IN1(n11402), .IN2(n12029), .QN(n12046) );
  NAND3X0 U12347 ( .IN1(n12047), .IN2(n12048), .IN3(n12049), .QN(g30533) );
  NAND2X0 U12348 ( .IN1(n3814), .IN2(n11388), .QN(n12049) );
  NAND2X0 U12349 ( .IN1(n9036), .IN2(g6271), .QN(n12048) );
  NAND3X0 U12350 ( .IN1(n12050), .IN2(g6287), .IN3(n8883), .QN(n12047) );
  NAND2X0 U12351 ( .IN1(n11402), .IN2(n11388), .QN(n12050) );
  NAND3X0 U12352 ( .IN1(n12051), .IN2(n12052), .IN3(n12053), .QN(g30532) );
  NAND2X0 U12353 ( .IN1(n3814), .IN2(n12019), .QN(n12053) );
  NAND2X0 U12354 ( .IN1(n9036), .IN2(g6267), .QN(n12052) );
  NAND3X0 U12355 ( .IN1(n12054), .IN2(g6283), .IN3(n8883), .QN(n12051) );
  NAND2X0 U12356 ( .IN1(n11402), .IN2(n12019), .QN(n12054) );
  NAND3X0 U12357 ( .IN1(n12055), .IN2(n12056), .IN3(n12057), .QN(g30531) );
  NAND2X0 U12358 ( .IN1(n3814), .IN2(n12025), .QN(n12057) );
  NAND2X0 U12359 ( .IN1(n9036), .IN2(g6263), .QN(n12056) );
  NAND3X0 U12360 ( .IN1(n12058), .IN2(g6279), .IN3(n8883), .QN(n12055) );
  NAND2X0 U12361 ( .IN1(n11402), .IN2(n12025), .QN(n12058) );
  INVX0 U12362 ( .INP(n1010), .ZN(n11402) );
  NAND2X0 U12363 ( .IN1(n5574), .IN2(g6209), .QN(n1010) );
  NAND3X0 U12364 ( .IN1(n12059), .IN2(n12060), .IN3(n12061), .QN(g30530) );
  NAND2X0 U12365 ( .IN1(n3819), .IN2(n12029), .QN(n12061) );
  NAND2X0 U12366 ( .IN1(n9035), .IN2(g6255), .QN(n12060) );
  NAND3X0 U12367 ( .IN1(n12062), .IN2(g6275), .IN3(n8883), .QN(n12059) );
  NAND2X0 U12368 ( .IN1(n12063), .IN2(n12029), .QN(n12062) );
  NAND3X0 U12369 ( .IN1(n12064), .IN2(n12065), .IN3(n12066), .QN(g30529) );
  NAND2X0 U12370 ( .IN1(n3819), .IN2(n11388), .QN(n12066) );
  NAND2X0 U12371 ( .IN1(n9035), .IN2(g6247), .QN(n12065) );
  NAND3X0 U12372 ( .IN1(n12067), .IN2(g6271), .IN3(n8883), .QN(n12064) );
  NAND2X0 U12373 ( .IN1(n12063), .IN2(n11388), .QN(n12067) );
  INVX0 U12374 ( .INP(n46), .ZN(n11388) );
  NAND2X0 U12375 ( .IN1(n5385), .IN2(g6227), .QN(n46) );
  NAND3X0 U12376 ( .IN1(n12068), .IN2(n12069), .IN3(n12070), .QN(g30528) );
  NAND2X0 U12377 ( .IN1(n3819), .IN2(n12019), .QN(n12070) );
  NAND2X0 U12378 ( .IN1(n9035), .IN2(g6239), .QN(n12069) );
  NAND3X0 U12379 ( .IN1(n12071), .IN2(g6267), .IN3(n8883), .QN(n12068) );
  NAND2X0 U12380 ( .IN1(n12063), .IN2(n12019), .QN(n12071) );
  INVX0 U12381 ( .INP(n42), .ZN(n12019) );
  NAND2X0 U12382 ( .IN1(n5568), .IN2(g6219), .QN(n42) );
  NAND3X0 U12383 ( .IN1(n12072), .IN2(n12073), .IN3(n12074), .QN(g30527) );
  NAND2X0 U12384 ( .IN1(n3819), .IN2(n12025), .QN(n12074) );
  NAND2X0 U12385 ( .IN1(n9035), .IN2(g6235), .QN(n12073) );
  NAND3X0 U12386 ( .IN1(n12075), .IN2(g6263), .IN3(n8871), .QN(n12072) );
  NAND2X0 U12387 ( .IN1(n12063), .IN2(n12025), .QN(n12075) );
  INVX0 U12388 ( .INP(n44), .ZN(n12025) );
  NAND2X0 U12389 ( .IN1(n5568), .IN2(n5385), .QN(n44) );
  INVX0 U12390 ( .INP(n1011), .ZN(n12063) );
  NAND2X0 U12391 ( .IN1(n8491), .IN2(g6203), .QN(n1011) );
  NAND3X0 U12392 ( .IN1(n12076), .IN2(n12077), .IN3(n12078), .QN(g30526) );
  NAND2X0 U12393 ( .IN1(n9035), .IN2(g6259), .QN(n12078) );
  NAND3X0 U12394 ( .IN1(n8898), .IN2(g6255), .IN3(n12079), .QN(n12077) );
  INVX0 U12395 ( .INP(n3824), .ZN(n12079) );
  NAND2X0 U12396 ( .IN1(n3824), .IN2(n3765), .QN(n12076) );
  NAND3X0 U12397 ( .IN1(n12080), .IN2(n12081), .IN3(n12082), .QN(g30525) );
  NAND2X0 U12398 ( .IN1(n9035), .IN2(g6251), .QN(n12082) );
  NAND3X0 U12399 ( .IN1(n8897), .IN2(g6247), .IN3(n12083), .QN(n12081) );
  INVX0 U12400 ( .INP(n3827), .ZN(n12083) );
  NAND2X0 U12401 ( .IN1(n3827), .IN2(n3765), .QN(n12080) );
  NAND3X0 U12402 ( .IN1(n12084), .IN2(n12085), .IN3(n12086), .QN(g30524) );
  NAND2X0 U12403 ( .IN1(n9035), .IN2(g6243), .QN(n12086) );
  NAND3X0 U12404 ( .IN1(n8898), .IN2(g6239), .IN3(n12087), .QN(n12085) );
  INVX0 U12405 ( .INP(n3829), .ZN(n12087) );
  NAND2X0 U12406 ( .IN1(n3829), .IN2(n3765), .QN(n12084) );
  NAND3X0 U12407 ( .IN1(n12088), .IN2(n12089), .IN3(n12090), .QN(g30523) );
  NAND2X0 U12408 ( .IN1(n9034), .IN2(g6227), .QN(n12090) );
  NAND3X0 U12409 ( .IN1(n8897), .IN2(g6235), .IN3(n12091), .QN(n12089) );
  INVX0 U12410 ( .INP(n3831), .ZN(n12091) );
  NAND2X0 U12411 ( .IN1(n3831), .IN2(n3765), .QN(n12088) );
  NOR2X0 U12412 ( .IN1(g6203), .IN2(n11394), .QN(g30522) );
  NAND3X0 U12413 ( .IN1(n11384), .IN2(n8869), .IN3(n5651), .QN(n11394) );
  NAND3X0 U12414 ( .IN1(g4093), .IN2(g4087), .IN3(n3833), .QN(n11384) );
  NAND3X0 U12415 ( .IN1(n12092), .IN2(n12093), .IN3(n12094), .QN(g30521) );
  NAND2X0 U12416 ( .IN1(n9034), .IN2(g5961), .QN(n12094) );
  NAND2X0 U12417 ( .IN1(test_so13), .IN2(n12095), .QN(n12093) );
  NAND2X0 U12418 ( .IN1(n12096), .IN2(n3765), .QN(n12092) );
  NAND3X0 U12419 ( .IN1(n12097), .IN2(n12098), .IN3(n12099), .QN(g30520) );
  NAND2X0 U12420 ( .IN1(n12100), .IN2(n3765), .QN(n12099) );
  INVX0 U12421 ( .INP(n12101), .ZN(n12100) );
  NAND3X0 U12422 ( .IN1(n12101), .IN2(g5913), .IN3(n8877), .QN(n12098) );
  NAND2X0 U12423 ( .IN1(n11410), .IN2(g5869), .QN(n12101) );
  NAND2X0 U12424 ( .IN1(n9034), .IN2(g5957), .QN(n12097) );
  NAND3X0 U12425 ( .IN1(n12102), .IN2(n12103), .IN3(n12104), .QN(g30519) );
  NAND2X0 U12426 ( .IN1(n12105), .IN2(n3765), .QN(n12104) );
  INVX0 U12427 ( .INP(n11408), .ZN(n12105) );
  NAND3X0 U12428 ( .IN1(n11408), .IN2(g5905), .IN3(n8881), .QN(n12103) );
  NAND2X0 U12429 ( .IN1(n12106), .IN2(g5869), .QN(n11408) );
  NAND2X0 U12430 ( .IN1(n9034), .IN2(g5953), .QN(n12102) );
  NAND3X0 U12431 ( .IN1(n12107), .IN2(n12108), .IN3(n12109), .QN(g30518) );
  NAND2X0 U12432 ( .IN1(n12110), .IN2(n3765), .QN(n12109) );
  INVX0 U12433 ( .INP(n12111), .ZN(n12110) );
  NAND3X0 U12434 ( .IN1(n12111), .IN2(g5897), .IN3(n8881), .QN(n12108) );
  NAND2X0 U12435 ( .IN1(n12112), .IN2(g5869), .QN(n12111) );
  NAND2X0 U12436 ( .IN1(n9034), .IN2(g5949), .QN(n12107) );
  NAND3X0 U12437 ( .IN1(n12113), .IN2(n12114), .IN3(n12115), .QN(g30517) );
  NAND2X0 U12438 ( .IN1(n3842), .IN2(n12116), .QN(n12115) );
  NAND2X0 U12439 ( .IN1(n9034), .IN2(g5945), .QN(n12114) );
  NAND3X0 U12440 ( .IN1(n12117), .IN2(g5961), .IN3(n8880), .QN(n12113) );
  NAND2X0 U12441 ( .IN1(n11419), .IN2(n12116), .QN(n12117) );
  NAND3X0 U12442 ( .IN1(n12118), .IN2(n12119), .IN3(n12120), .QN(g30516) );
  NAND2X0 U12443 ( .IN1(n3842), .IN2(n11410), .QN(n12120) );
  NAND2X0 U12444 ( .IN1(n9034), .IN2(g5941), .QN(n12119) );
  NAND3X0 U12445 ( .IN1(n12121), .IN2(g5957), .IN3(n8880), .QN(n12118) );
  NAND2X0 U12446 ( .IN1(n11419), .IN2(n11410), .QN(n12121) );
  NAND3X0 U12447 ( .IN1(n12122), .IN2(n12123), .IN3(n12124), .QN(g30515) );
  NAND2X0 U12448 ( .IN1(n3842), .IN2(n12106), .QN(n12124) );
  NAND2X0 U12449 ( .IN1(n9033), .IN2(g5937), .QN(n12123) );
  NAND3X0 U12450 ( .IN1(n12125), .IN2(g5953), .IN3(n8880), .QN(n12122) );
  NAND2X0 U12451 ( .IN1(n11419), .IN2(n12106), .QN(n12125) );
  NAND3X0 U12452 ( .IN1(n12126), .IN2(n12127), .IN3(n12128), .QN(g30514) );
  NAND2X0 U12453 ( .IN1(n3842), .IN2(n12112), .QN(n12128) );
  NAND2X0 U12454 ( .IN1(n9033), .IN2(g5933), .QN(n12127) );
  NAND3X0 U12455 ( .IN1(n12129), .IN2(g5949), .IN3(n8880), .QN(n12126) );
  NAND2X0 U12456 ( .IN1(n11419), .IN2(n12112), .QN(n12129) );
  INVX0 U12457 ( .INP(n1073), .ZN(n11419) );
  NAND2X0 U12458 ( .IN1(g5857), .IN2(g5863), .QN(n1073) );
  NAND3X0 U12459 ( .IN1(n12130), .IN2(n12131), .IN3(n12132), .QN(g30513) );
  NAND2X0 U12460 ( .IN1(n3848), .IN2(n12116), .QN(n12132) );
  NAND2X0 U12461 ( .IN1(n9033), .IN2(g5929), .QN(n12131) );
  NAND3X0 U12462 ( .IN1(n12133), .IN2(g5945), .IN3(n8880), .QN(n12130) );
  NAND2X0 U12463 ( .IN1(n11424), .IN2(n12116), .QN(n12133) );
  NAND3X0 U12464 ( .IN1(n12134), .IN2(n12135), .IN3(n12136), .QN(g30512) );
  NAND2X0 U12465 ( .IN1(n3848), .IN2(n11410), .QN(n12136) );
  NAND2X0 U12466 ( .IN1(n9033), .IN2(g5925), .QN(n12135) );
  NAND3X0 U12467 ( .IN1(n12137), .IN2(g5941), .IN3(n8880), .QN(n12134) );
  NAND2X0 U12468 ( .IN1(n11424), .IN2(n11410), .QN(n12137) );
  NAND3X0 U12469 ( .IN1(n12138), .IN2(n12139), .IN3(n12140), .QN(g30511) );
  NAND2X0 U12470 ( .IN1(n3848), .IN2(n12106), .QN(n12140) );
  NAND2X0 U12471 ( .IN1(n9033), .IN2(g5921), .QN(n12139) );
  NAND3X0 U12472 ( .IN1(n12141), .IN2(g5937), .IN3(n8879), .QN(n12138) );
  NAND2X0 U12473 ( .IN1(n11424), .IN2(n12106), .QN(n12141) );
  NAND3X0 U12474 ( .IN1(n12142), .IN2(n12143), .IN3(n12144), .QN(g30510) );
  NAND2X0 U12475 ( .IN1(n3848), .IN2(n12112), .QN(n12144) );
  NAND2X0 U12476 ( .IN1(test_so28), .IN2(n9053), .QN(n12143) );
  NAND3X0 U12477 ( .IN1(n12145), .IN2(g5933), .IN3(n8879), .QN(n12142) );
  NAND2X0 U12478 ( .IN1(n11424), .IN2(n12112), .QN(n12145) );
  INVX0 U12479 ( .INP(n1074), .ZN(n11424) );
  NAND2X0 U12480 ( .IN1(n5573), .IN2(g5863), .QN(n1074) );
  NAND3X0 U12481 ( .IN1(n12146), .IN2(n12147), .IN3(n12148), .QN(g30509) );
  NAND2X0 U12482 ( .IN1(n3853), .IN2(n12116), .QN(n12148) );
  NAND2X0 U12483 ( .IN1(n9033), .IN2(g5909), .QN(n12147) );
  NAND3X0 U12484 ( .IN1(n12149), .IN2(g5929), .IN3(n8879), .QN(n12146) );
  NAND2X0 U12485 ( .IN1(n12150), .IN2(n12116), .QN(n12149) );
  NAND3X0 U12486 ( .IN1(n12151), .IN2(n12152), .IN3(n12153), .QN(g30508) );
  NAND2X0 U12487 ( .IN1(n3853), .IN2(n11410), .QN(n12153) );
  NAND2X0 U12488 ( .IN1(n9033), .IN2(g5901), .QN(n12152) );
  NAND3X0 U12489 ( .IN1(n12154), .IN2(g5925), .IN3(n8879), .QN(n12151) );
  NAND2X0 U12490 ( .IN1(n12150), .IN2(n11410), .QN(n12154) );
  INVX0 U12491 ( .INP(n716), .ZN(n11410) );
  NAND2X0 U12492 ( .IN1(n5388), .IN2(test_so36), .QN(n716) );
  NAND3X0 U12493 ( .IN1(n12155), .IN2(n12156), .IN3(n12157), .QN(g30507) );
  NAND2X0 U12494 ( .IN1(n3853), .IN2(n12106), .QN(n12157) );
  NAND2X0 U12495 ( .IN1(n9032), .IN2(g5893), .QN(n12156) );
  NAND3X0 U12496 ( .IN1(n12158), .IN2(g5921), .IN3(n8879), .QN(n12155) );
  NAND2X0 U12497 ( .IN1(n12150), .IN2(n12106), .QN(n12158) );
  INVX0 U12498 ( .INP(n712), .ZN(n12106) );
  NAND2X0 U12499 ( .IN1(g5873), .IN2(n8599), .QN(n712) );
  NAND3X0 U12500 ( .IN1(n12159), .IN2(n12160), .IN3(n12161), .QN(g30506) );
  NAND2X0 U12501 ( .IN1(n3853), .IN2(n12112), .QN(n12161) );
  NAND2X0 U12502 ( .IN1(n9032), .IN2(g5889), .QN(n12160) );
  NAND3X0 U12503 ( .IN1(test_so28), .IN2(n12162), .IN3(n8879), .QN(n12159) );
  NAND2X0 U12504 ( .IN1(n12150), .IN2(n12112), .QN(n12162) );
  INVX0 U12505 ( .INP(n714), .ZN(n12112) );
  NAND2X0 U12506 ( .IN1(n5388), .IN2(n8599), .QN(n714) );
  INVX0 U12507 ( .INP(n1075), .ZN(n12150) );
  NAND2X0 U12508 ( .IN1(n8493), .IN2(g5857), .QN(n1075) );
  NAND3X0 U12509 ( .IN1(n12163), .IN2(n12164), .IN3(n12165), .QN(g30505) );
  NAND2X0 U12510 ( .IN1(n9032), .IN2(g5913), .QN(n12165) );
  NAND3X0 U12511 ( .IN1(n8894), .IN2(g5909), .IN3(n12166), .QN(n12164) );
  INVX0 U12512 ( .INP(n3858), .ZN(n12166) );
  NAND2X0 U12513 ( .IN1(n3858), .IN2(n3765), .QN(n12163) );
  NAND3X0 U12514 ( .IN1(n12167), .IN2(n12168), .IN3(n12169), .QN(g30504) );
  NAND2X0 U12515 ( .IN1(n9032), .IN2(g5905), .QN(n12169) );
  NAND3X0 U12516 ( .IN1(n8894), .IN2(g5901), .IN3(n12170), .QN(n12168) );
  INVX0 U12517 ( .INP(n3861), .ZN(n12170) );
  NAND2X0 U12518 ( .IN1(n3861), .IN2(n3765), .QN(n12167) );
  NAND3X0 U12519 ( .IN1(n12171), .IN2(n12172), .IN3(n12173), .QN(g30503) );
  NAND2X0 U12520 ( .IN1(n9032), .IN2(g5897), .QN(n12173) );
  NAND3X0 U12521 ( .IN1(n8894), .IN2(g5893), .IN3(n12174), .QN(n12172) );
  INVX0 U12522 ( .INP(n3863), .ZN(n12174) );
  NAND2X0 U12523 ( .IN1(n3863), .IN2(n3765), .QN(n12171) );
  NAND3X0 U12524 ( .IN1(n12175), .IN2(n12176), .IN3(n12177), .QN(g30502) );
  NAND2X0 U12525 ( .IN1(test_so36), .IN2(n9052), .QN(n12177) );
  NAND3X0 U12526 ( .IN1(n8896), .IN2(g5889), .IN3(n12178), .QN(n12176) );
  INVX0 U12527 ( .INP(n3865), .ZN(n12178) );
  NAND2X0 U12528 ( .IN1(n3865), .IN2(n3765), .QN(n12175) );
  NOR2X0 U12529 ( .IN1(g5857), .IN2(n11416), .QN(g30501) );
  NAND3X0 U12530 ( .IN1(n11406), .IN2(n8870), .IN3(n5649), .QN(n11416) );
  NAND3X0 U12531 ( .IN1(n5480), .IN2(g4093), .IN3(n3833), .QN(n11406) );
  NAND3X0 U12532 ( .IN1(n12179), .IN2(n12180), .IN3(n12181), .QN(g30500) );
  NAND2X0 U12533 ( .IN1(n9032), .IN2(g5615), .QN(n12181) );
  NAND2X0 U12534 ( .IN1(n12182), .IN2(g5619), .QN(n12180) );
  NAND2X0 U12535 ( .IN1(n3765), .IN2(n10823), .QN(n12179) );
  NAND3X0 U12536 ( .IN1(n12183), .IN2(n12184), .IN3(n12185), .QN(g30499) );
  NAND2X0 U12537 ( .IN1(n12186), .IN2(n3765), .QN(n12185) );
  INVX0 U12538 ( .INP(n12187), .ZN(n12186) );
  NAND3X0 U12539 ( .IN1(n12187), .IN2(g5567), .IN3(n8879), .QN(n12184) );
  NAND2X0 U12540 ( .IN1(n11432), .IN2(g5523), .QN(n12187) );
  NAND2X0 U12541 ( .IN1(n9032), .IN2(g5611), .QN(n12183) );
  NAND3X0 U12542 ( .IN1(n12188), .IN2(n12189), .IN3(n12190), .QN(g30498) );
  NAND2X0 U12543 ( .IN1(n12191), .IN2(n3765), .QN(n12190) );
  INVX0 U12544 ( .INP(n11430), .ZN(n12191) );
  NAND3X0 U12545 ( .IN1(test_so6), .IN2(n11430), .IN3(n8879), .QN(n12189) );
  NAND2X0 U12546 ( .IN1(n12192), .IN2(g5523), .QN(n11430) );
  NAND2X0 U12547 ( .IN1(n9031), .IN2(g5607), .QN(n12188) );
  NAND3X0 U12548 ( .IN1(n12193), .IN2(n12194), .IN3(n12195), .QN(g30497) );
  NAND2X0 U12549 ( .IN1(n12196), .IN2(n3765), .QN(n12195) );
  INVX0 U12550 ( .INP(n12197), .ZN(n12196) );
  NAND3X0 U12551 ( .IN1(n12197), .IN2(g5551), .IN3(n8879), .QN(n12194) );
  NAND2X0 U12552 ( .IN1(n12198), .IN2(g5523), .QN(n12197) );
  NAND2X0 U12553 ( .IN1(n9031), .IN2(g5603), .QN(n12193) );
  NAND3X0 U12554 ( .IN1(n12199), .IN2(n12200), .IN3(n12201), .QN(g30496) );
  NAND2X0 U12555 ( .IN1(n3875), .IN2(n12202), .QN(n12201) );
  NAND2X0 U12556 ( .IN1(n9031), .IN2(g5599), .QN(n12200) );
  NAND3X0 U12557 ( .IN1(n12203), .IN2(g5615), .IN3(n8879), .QN(n12199) );
  NAND2X0 U12558 ( .IN1(n11441), .IN2(n12202), .QN(n12203) );
  NAND3X0 U12559 ( .IN1(n12204), .IN2(n12205), .IN3(n12206), .QN(g30495) );
  NAND2X0 U12560 ( .IN1(n3875), .IN2(n11432), .QN(n12206) );
  NAND2X0 U12561 ( .IN1(n9031), .IN2(g5595), .QN(n12205) );
  NAND3X0 U12562 ( .IN1(n12207), .IN2(g5611), .IN3(n8879), .QN(n12204) );
  NAND2X0 U12563 ( .IN1(n11441), .IN2(n11432), .QN(n12207) );
  NAND3X0 U12564 ( .IN1(n12208), .IN2(n12209), .IN3(n12210), .QN(g30494) );
  NAND2X0 U12565 ( .IN1(n3875), .IN2(n12192), .QN(n12210) );
  NAND2X0 U12566 ( .IN1(test_so5), .IN2(n9052), .QN(n12209) );
  NAND3X0 U12567 ( .IN1(n12211), .IN2(g5607), .IN3(n8878), .QN(n12208) );
  NAND2X0 U12568 ( .IN1(n11441), .IN2(n12192), .QN(n12211) );
  NAND3X0 U12569 ( .IN1(n12212), .IN2(n12213), .IN3(n12214), .QN(g30493) );
  NAND2X0 U12570 ( .IN1(n3875), .IN2(n12198), .QN(n12214) );
  NAND2X0 U12571 ( .IN1(n9031), .IN2(g5587), .QN(n12213) );
  NAND3X0 U12572 ( .IN1(n12215), .IN2(g5603), .IN3(n8878), .QN(n12212) );
  NAND2X0 U12573 ( .IN1(n11441), .IN2(n12198), .QN(n12215) );
  INVX0 U12574 ( .INP(n494), .ZN(n11441) );
  NAND2X0 U12575 ( .IN1(g5511), .IN2(g5517), .QN(n494) );
  NAND3X0 U12576 ( .IN1(n12216), .IN2(n12217), .IN3(n12218), .QN(g30492) );
  NAND2X0 U12577 ( .IN1(n3881), .IN2(n12202), .QN(n12218) );
  NAND2X0 U12578 ( .IN1(n9031), .IN2(g5583), .QN(n12217) );
  NAND3X0 U12579 ( .IN1(n12219), .IN2(g5599), .IN3(n8878), .QN(n12216) );
  NAND2X0 U12580 ( .IN1(n11446), .IN2(n12202), .QN(n12219) );
  NAND3X0 U12581 ( .IN1(n12220), .IN2(n12221), .IN3(n12222), .QN(g30491) );
  NAND2X0 U12582 ( .IN1(n3881), .IN2(n11432), .QN(n12222) );
  NAND2X0 U12583 ( .IN1(n9031), .IN2(g5579), .QN(n12221) );
  NAND3X0 U12584 ( .IN1(n12223), .IN2(g5595), .IN3(n8878), .QN(n12220) );
  NAND2X0 U12585 ( .IN1(n11446), .IN2(n11432), .QN(n12223) );
  NAND3X0 U12586 ( .IN1(n12224), .IN2(n12225), .IN3(n12226), .QN(g30490) );
  NAND2X0 U12587 ( .IN1(n3881), .IN2(n12192), .QN(n12226) );
  NAND2X0 U12588 ( .IN1(n9030), .IN2(g5575), .QN(n12225) );
  NAND3X0 U12589 ( .IN1(test_so5), .IN2(n12227), .IN3(n8878), .QN(n12224) );
  NAND2X0 U12590 ( .IN1(n11446), .IN2(n12192), .QN(n12227) );
  NAND3X0 U12591 ( .IN1(n12228), .IN2(n12229), .IN3(n12230), .QN(g30489) );
  NAND2X0 U12592 ( .IN1(n3881), .IN2(n12198), .QN(n12230) );
  NAND2X0 U12593 ( .IN1(n9030), .IN2(g5571), .QN(n12229) );
  NAND3X0 U12594 ( .IN1(n12231), .IN2(g5587), .IN3(n8878), .QN(n12228) );
  NAND2X0 U12595 ( .IN1(n11446), .IN2(n12198), .QN(n12231) );
  INVX0 U12596 ( .INP(n496), .ZN(n11446) );
  NAND2X0 U12597 ( .IN1(n5575), .IN2(g5517), .QN(n496) );
  NAND3X0 U12598 ( .IN1(n12232), .IN2(n12233), .IN3(n12234), .QN(g30488) );
  NAND2X0 U12599 ( .IN1(n3886), .IN2(n12202), .QN(n12234) );
  NAND2X0 U12600 ( .IN1(n9030), .IN2(g5563), .QN(n12233) );
  NAND3X0 U12601 ( .IN1(n12235), .IN2(g5583), .IN3(n8878), .QN(n12232) );
  NAND2X0 U12602 ( .IN1(n12236), .IN2(n12202), .QN(n12235) );
  INVX0 U12603 ( .INP(n939), .ZN(n12202) );
  NAND3X0 U12604 ( .IN1(n12237), .IN2(n12238), .IN3(n12239), .QN(g30487) );
  NAND2X0 U12605 ( .IN1(n3886), .IN2(n11432), .QN(n12239) );
  NAND2X0 U12606 ( .IN1(n9030), .IN2(g5555), .QN(n12238) );
  NAND3X0 U12607 ( .IN1(n12240), .IN2(g5579), .IN3(n8878), .QN(n12237) );
  NAND2X0 U12608 ( .IN1(n12236), .IN2(n11432), .QN(n12240) );
  INVX0 U12609 ( .INP(n935), .ZN(n11432) );
  NAND2X0 U12610 ( .IN1(n5389), .IN2(g5535), .QN(n935) );
  NAND3X0 U12611 ( .IN1(n12241), .IN2(n12242), .IN3(n12243), .QN(g30486) );
  NAND2X0 U12612 ( .IN1(n3886), .IN2(n12192), .QN(n12243) );
  NAND2X0 U12613 ( .IN1(n9030), .IN2(g5547), .QN(n12242) );
  NAND3X0 U12614 ( .IN1(n12244), .IN2(g5575), .IN3(n8878), .QN(n12241) );
  NAND2X0 U12615 ( .IN1(n12236), .IN2(n12192), .QN(n12244) );
  INVX0 U12616 ( .INP(n937), .ZN(n12192) );
  NAND2X0 U12617 ( .IN1(n5566), .IN2(g5527), .QN(n937) );
  NAND3X0 U12618 ( .IN1(n12245), .IN2(n12246), .IN3(n12247), .QN(g30485) );
  NAND2X0 U12619 ( .IN1(n3886), .IN2(n12198), .QN(n12247) );
  NAND2X0 U12620 ( .IN1(n9030), .IN2(g5543), .QN(n12246) );
  NAND3X0 U12621 ( .IN1(n12248), .IN2(g5571), .IN3(n8878), .QN(n12245) );
  NAND2X0 U12622 ( .IN1(n12236), .IN2(n12198), .QN(n12248) );
  INVX0 U12623 ( .INP(n936), .ZN(n12198) );
  NAND2X0 U12624 ( .IN1(n5389), .IN2(n5566), .QN(n936) );
  INVX0 U12625 ( .INP(n495), .ZN(n12236) );
  NAND2X0 U12626 ( .IN1(n8492), .IN2(g5511), .QN(n495) );
  NAND3X0 U12627 ( .IN1(n12249), .IN2(n12250), .IN3(n12251), .QN(g30484) );
  NAND2X0 U12628 ( .IN1(n9030), .IN2(g5567), .QN(n12251) );
  NAND3X0 U12629 ( .IN1(n8896), .IN2(g5563), .IN3(n12252), .QN(n12250) );
  INVX0 U12630 ( .INP(n3891), .ZN(n12252) );
  NAND2X0 U12631 ( .IN1(n3891), .IN2(n3765), .QN(n12249) );
  NAND3X0 U12632 ( .IN1(n12253), .IN2(n12254), .IN3(n12255), .QN(g30483) );
  NAND2X0 U12633 ( .IN1(test_so6), .IN2(n9051), .QN(n12255) );
  NAND3X0 U12634 ( .IN1(n8895), .IN2(g5555), .IN3(n12256), .QN(n12254) );
  INVX0 U12635 ( .INP(n3894), .ZN(n12256) );
  NAND2X0 U12636 ( .IN1(n3894), .IN2(n3765), .QN(n12253) );
  NAND3X0 U12637 ( .IN1(n12257), .IN2(n12258), .IN3(n12259), .QN(g30482) );
  NAND2X0 U12638 ( .IN1(n9029), .IN2(g5551), .QN(n12259) );
  NAND3X0 U12639 ( .IN1(n8895), .IN2(g5547), .IN3(n12260), .QN(n12258) );
  INVX0 U12640 ( .INP(n3896), .ZN(n12260) );
  NAND2X0 U12641 ( .IN1(n3896), .IN2(n3765), .QN(n12257) );
  NAND3X0 U12642 ( .IN1(n12261), .IN2(n12262), .IN3(n12263), .QN(g30481) );
  NAND2X0 U12643 ( .IN1(n9029), .IN2(g5535), .QN(n12263) );
  NAND3X0 U12644 ( .IN1(n8895), .IN2(g5543), .IN3(n12264), .QN(n12262) );
  INVX0 U12645 ( .INP(n3898), .ZN(n12264) );
  NAND2X0 U12646 ( .IN1(n3898), .IN2(n3765), .QN(n12261) );
  NOR2X0 U12647 ( .IN1(g5511), .IN2(n11438), .QN(g30480) );
  NAND3X0 U12648 ( .IN1(n11428), .IN2(n8870), .IN3(n5647), .QN(n11438) );
  NAND2X0 U12649 ( .IN1(n3833), .IN2(n10824), .QN(n11428) );
  NAND3X0 U12650 ( .IN1(n12265), .IN2(n12266), .IN3(n12267), .QN(g30479) );
  NAND2X0 U12651 ( .IN1(n9040), .IN2(g5268), .QN(n12267) );
  NAND2X0 U12652 ( .IN1(n12268), .IN2(g5272), .QN(n12266) );
  NAND2X0 U12653 ( .IN1(n3765), .IN2(g32975), .QN(n12265) );
  NAND3X0 U12654 ( .IN1(n12269), .IN2(n12270), .IN3(n12271), .QN(g30478) );
  NAND2X0 U12655 ( .IN1(n12272), .IN2(n3765), .QN(n12271) );
  INVX0 U12656 ( .INP(n12273), .ZN(n12272) );
  NAND3X0 U12657 ( .IN1(n12273), .IN2(g5220), .IN3(n8878), .QN(n12270) );
  NAND2X0 U12658 ( .IN1(n11454), .IN2(g5176), .QN(n12273) );
  NAND2X0 U12659 ( .IN1(n9029), .IN2(g5264), .QN(n12269) );
  NAND3X0 U12660 ( .IN1(n12274), .IN2(n12275), .IN3(n12276), .QN(g30477) );
  NAND2X0 U12661 ( .IN1(n12277), .IN2(n3765), .QN(n12276) );
  INVX0 U12662 ( .INP(n11452), .ZN(n12277) );
  NAND3X0 U12663 ( .IN1(n11452), .IN2(g5212), .IN3(n8877), .QN(n12275) );
  NAND2X0 U12664 ( .IN1(n12278), .IN2(g5176), .QN(n11452) );
  NAND2X0 U12665 ( .IN1(n9029), .IN2(g5260), .QN(n12274) );
  NAND3X0 U12666 ( .IN1(n12279), .IN2(n12280), .IN3(n12281), .QN(g30476) );
  NAND2X0 U12667 ( .IN1(n12282), .IN2(n3765), .QN(n12281) );
  INVX0 U12668 ( .INP(n12283), .ZN(n12282) );
  NAND3X0 U12669 ( .IN1(n12283), .IN2(g5204), .IN3(n8877), .QN(n12280) );
  NAND2X0 U12670 ( .IN1(n12284), .IN2(g5176), .QN(n12283) );
  NAND2X0 U12671 ( .IN1(n9029), .IN2(g5256), .QN(n12279) );
  NAND3X0 U12672 ( .IN1(n12285), .IN2(n12286), .IN3(n12287), .QN(g30475) );
  NAND2X0 U12673 ( .IN1(n3908), .IN2(n12288), .QN(n12287) );
  NAND2X0 U12674 ( .IN1(n9029), .IN2(g5252), .QN(n12286) );
  NAND3X0 U12675 ( .IN1(n12289), .IN2(g5268), .IN3(n8877), .QN(n12285) );
  NAND2X0 U12676 ( .IN1(n12288), .IN2(n11463), .QN(n12289) );
  NAND3X0 U12677 ( .IN1(n12290), .IN2(n12291), .IN3(n12292), .QN(g30474) );
  NAND2X0 U12678 ( .IN1(n3908), .IN2(n11454), .QN(n12292) );
  NAND2X0 U12679 ( .IN1(n9028), .IN2(g5248), .QN(n12291) );
  NAND3X0 U12680 ( .IN1(n12293), .IN2(g5264), .IN3(n8877), .QN(n12290) );
  NAND2X0 U12681 ( .IN1(n11454), .IN2(n11463), .QN(n12293) );
  NAND3X0 U12682 ( .IN1(n12294), .IN2(n12295), .IN3(n12296), .QN(g30473) );
  NAND2X0 U12683 ( .IN1(n3908), .IN2(n12278), .QN(n12296) );
  NAND2X0 U12684 ( .IN1(n9028), .IN2(g5244), .QN(n12295) );
  NAND3X0 U12685 ( .IN1(n12297), .IN2(g5260), .IN3(n8872), .QN(n12294) );
  NAND2X0 U12686 ( .IN1(n12278), .IN2(n11463), .QN(n12297) );
  NAND3X0 U12687 ( .IN1(n12298), .IN2(n12299), .IN3(n12300), .QN(g30472) );
  NAND2X0 U12688 ( .IN1(n3908), .IN2(n12284), .QN(n12300) );
  NAND2X0 U12689 ( .IN1(n9028), .IN2(g5240), .QN(n12299) );
  NAND3X0 U12690 ( .IN1(n12301), .IN2(g5256), .IN3(n8871), .QN(n12298) );
  NAND2X0 U12691 ( .IN1(n12284), .IN2(n11463), .QN(n12301) );
  INVX0 U12692 ( .INP(n744), .ZN(n11463) );
  NAND2X0 U12693 ( .IN1(g5164), .IN2(g5170), .QN(n744) );
  NAND3X0 U12694 ( .IN1(n12302), .IN2(n12303), .IN3(n12304), .QN(g30471) );
  NAND2X0 U12695 ( .IN1(n3914), .IN2(n12288), .QN(n12304) );
  NAND2X0 U12696 ( .IN1(n9028), .IN2(g5236), .QN(n12303) );
  NAND3X0 U12697 ( .IN1(n12305), .IN2(g5252), .IN3(n8872), .QN(n12302) );
  NAND2X0 U12698 ( .IN1(n12288), .IN2(n11468), .QN(n12305) );
  NAND3X0 U12699 ( .IN1(n12306), .IN2(n12307), .IN3(n12308), .QN(g30470) );
  NAND2X0 U12700 ( .IN1(n3914), .IN2(n11454), .QN(n12308) );
  NAND2X0 U12701 ( .IN1(n9028), .IN2(g5232), .QN(n12307) );
  NAND3X0 U12702 ( .IN1(n12309), .IN2(g5248), .IN3(n8872), .QN(n12306) );
  NAND2X0 U12703 ( .IN1(n11454), .IN2(n11468), .QN(n12309) );
  NAND3X0 U12704 ( .IN1(n12310), .IN2(n12311), .IN3(n12312), .QN(g30469) );
  NAND2X0 U12705 ( .IN1(n3914), .IN2(n12278), .QN(n12312) );
  NAND2X0 U12706 ( .IN1(test_so82), .IN2(n8951), .QN(n12311) );
  NAND3X0 U12707 ( .IN1(n12313), .IN2(g5244), .IN3(n8873), .QN(n12310) );
  NAND2X0 U12708 ( .IN1(n12278), .IN2(n11468), .QN(n12313) );
  NAND3X0 U12709 ( .IN1(n12314), .IN2(n12315), .IN3(n12316), .QN(g30468) );
  NAND2X0 U12710 ( .IN1(n3914), .IN2(n12284), .QN(n12316) );
  NAND2X0 U12711 ( .IN1(n9028), .IN2(g5224), .QN(n12315) );
  NAND3X0 U12712 ( .IN1(n12317), .IN2(g5240), .IN3(n8872), .QN(n12314) );
  NAND2X0 U12713 ( .IN1(n12284), .IN2(n11468), .QN(n12317) );
  INVX0 U12714 ( .INP(n746), .ZN(n11468) );
  NAND2X0 U12715 ( .IN1(n5570), .IN2(g5170), .QN(n746) );
  NAND3X0 U12716 ( .IN1(n12318), .IN2(n12319), .IN3(n12320), .QN(g30467) );
  NAND2X0 U12717 ( .IN1(n3919), .IN2(n12288), .QN(n12320) );
  NAND2X0 U12718 ( .IN1(n9028), .IN2(g5216), .QN(n12319) );
  NAND3X0 U12719 ( .IN1(n12321), .IN2(g5236), .IN3(n8873), .QN(n12318) );
  NAND2X0 U12720 ( .IN1(n12288), .IN2(n12322), .QN(n12321) );
  INVX0 U12721 ( .INP(n214), .ZN(n12288) );
  NAND3X0 U12722 ( .IN1(n12323), .IN2(n12324), .IN3(n12325), .QN(g30466) );
  NAND2X0 U12723 ( .IN1(n3919), .IN2(n11454), .QN(n12325) );
  NAND2X0 U12724 ( .IN1(n9027), .IN2(g5208), .QN(n12324) );
  NAND3X0 U12725 ( .IN1(n12326), .IN2(g5232), .IN3(n8872), .QN(n12323) );
  NAND2X0 U12726 ( .IN1(n11454), .IN2(n12322), .QN(n12326) );
  INVX0 U12727 ( .INP(n209), .ZN(n11454) );
  NAND2X0 U12728 ( .IN1(n5384), .IN2(g5188), .QN(n209) );
  NAND3X0 U12729 ( .IN1(n12327), .IN2(n12328), .IN3(n12329), .QN(g30465) );
  NAND2X0 U12730 ( .IN1(n3919), .IN2(n12278), .QN(n12329) );
  NAND2X0 U12731 ( .IN1(n9027), .IN2(g5200), .QN(n12328) );
  NAND3X0 U12732 ( .IN1(test_so82), .IN2(n12330), .IN3(n8872), .QN(n12327) );
  NAND2X0 U12733 ( .IN1(n12278), .IN2(n12322), .QN(n12330) );
  INVX0 U12734 ( .INP(n205), .ZN(n12278) );
  NAND2X0 U12735 ( .IN1(n5567), .IN2(g5180), .QN(n205) );
  NAND3X0 U12736 ( .IN1(n12331), .IN2(n12332), .IN3(n12333), .QN(g30464) );
  NAND2X0 U12737 ( .IN1(n3919), .IN2(n12284), .QN(n12333) );
  NAND2X0 U12738 ( .IN1(n9027), .IN2(g5196), .QN(n12332) );
  NAND3X0 U12739 ( .IN1(n12334), .IN2(g5224), .IN3(n8872), .QN(n12331) );
  NAND2X0 U12740 ( .IN1(n12284), .IN2(n12322), .QN(n12334) );
  INVX0 U12741 ( .INP(n745), .ZN(n12322) );
  NAND2X0 U12742 ( .IN1(n8489), .IN2(g5164), .QN(n745) );
  INVX0 U12743 ( .INP(n207), .ZN(n12284) );
  NAND2X0 U12744 ( .IN1(n5567), .IN2(n5384), .QN(n207) );
  NAND3X0 U12745 ( .IN1(n12335), .IN2(n12336), .IN3(n12337), .QN(g30463) );
  NAND2X0 U12746 ( .IN1(n9027), .IN2(g5220), .QN(n12337) );
  NAND3X0 U12747 ( .IN1(n8897), .IN2(g5216), .IN3(n12338), .QN(n12336) );
  INVX0 U12748 ( .INP(n3924), .ZN(n12338) );
  NAND2X0 U12749 ( .IN1(n3924), .IN2(n3765), .QN(n12335) );
  NAND3X0 U12750 ( .IN1(n12339), .IN2(n12340), .IN3(n12341), .QN(g30462) );
  NAND2X0 U12751 ( .IN1(n9027), .IN2(g5212), .QN(n12341) );
  NAND3X0 U12752 ( .IN1(n8897), .IN2(g5208), .IN3(n12342), .QN(n12340) );
  INVX0 U12753 ( .INP(n3927), .ZN(n12342) );
  NAND2X0 U12754 ( .IN1(n3927), .IN2(n3765), .QN(n12339) );
  NAND3X0 U12755 ( .IN1(n12343), .IN2(n12344), .IN3(n12345), .QN(g30461) );
  NAND2X0 U12756 ( .IN1(n9027), .IN2(g5204), .QN(n12345) );
  NAND3X0 U12757 ( .IN1(n8897), .IN2(g5200), .IN3(n12346), .QN(n12344) );
  INVX0 U12758 ( .INP(n3929), .ZN(n12346) );
  NAND2X0 U12759 ( .IN1(n3929), .IN2(n3765), .QN(n12343) );
  NAND3X0 U12760 ( .IN1(n12347), .IN2(n12348), .IN3(n12349), .QN(g30460) );
  NAND2X0 U12761 ( .IN1(n9027), .IN2(g5188), .QN(n12349) );
  NAND3X0 U12762 ( .IN1(n8897), .IN2(g5196), .IN3(n12350), .QN(n12348) );
  INVX0 U12763 ( .INP(n3931), .ZN(n12350) );
  NAND2X0 U12764 ( .IN1(n3931), .IN2(n3765), .QN(n12347) );
  NOR2X0 U12765 ( .IN1(g5164), .IN2(n11460), .QN(g30459) );
  NAND3X0 U12766 ( .IN1(n11450), .IN2(n8871), .IN3(n5650), .QN(n11460) );
  NAND2X0 U12767 ( .IN1(n3833), .IN2(n10829), .QN(n11450) );
  INVX0 U12768 ( .INP(n10053), .ZN(n10829) );
  NAND3X0 U12769 ( .IN1(n12351), .IN2(n12352), .IN3(n8873), .QN(g30458) );
  NAND2X0 U12770 ( .IN1(n12353), .IN2(g113), .QN(n12352) );
  INVX0 U12771 ( .INP(n12354), .ZN(n12353) );
  NAND2X0 U12772 ( .IN1(n12354), .IN2(g4507), .QN(n12351) );
  NAND2X0 U12773 ( .IN1(n5765), .IN2(g4473), .QN(n12354) );
  NAND2X0 U12774 ( .IN1(n12355), .IN2(n12356), .QN(g30457) );
  NAND2X0 U12775 ( .IN1(n9026), .IN2(g4122), .QN(n12356) );
  NAND2X0 U12776 ( .IN1(n12357), .IN2(n8916), .QN(n12355) );
  NAND2X0 U12777 ( .IN1(n12358), .IN2(n12359), .QN(n12357) );
  NAND2X0 U12778 ( .IN1(n12360), .IN2(n5981), .QN(n12359) );
  XNOR2X1 U12779 ( .IN1(g126), .IN2(n12361), .Q(n12360) );
  NAND2X0 U12780 ( .IN1(n12362), .IN2(n5983), .QN(n12358) );
  XNOR2X1 U12781 ( .IN1(g115), .IN2(n12363), .Q(n12362) );
  NAND3X0 U12782 ( .IN1(n12364), .IN2(n12365), .IN3(n12366), .QN(g30456) );
  NAND2X0 U12783 ( .IN1(n9026), .IN2(g4087), .QN(n12366) );
  NAND3X0 U12784 ( .IN1(n10824), .IN2(g4169), .IN3(n11856), .QN(n12365) );
  NAND2X0 U12785 ( .IN1(n3941), .IN2(n12367), .QN(n12364) );
  NAND3X0 U12786 ( .IN1(n12368), .IN2(n12369), .IN3(n12370), .QN(g30455) );
  NAND2X0 U12787 ( .IN1(n9029), .IN2(g3961), .QN(n12370) );
  NAND2X0 U12788 ( .IN1(n12371), .IN2(g3965), .QN(n12369) );
  NAND2X0 U12789 ( .IN1(n12372), .IN2(n3765), .QN(n12368) );
  NAND3X0 U12790 ( .IN1(n12373), .IN2(n12374), .IN3(n12375), .QN(g30454) );
  NAND2X0 U12791 ( .IN1(n12376), .IN2(n3765), .QN(n12375) );
  INVX0 U12792 ( .INP(n12377), .ZN(n12376) );
  NAND3X0 U12793 ( .IN1(n12377), .IN2(g3913), .IN3(n8873), .QN(n12374) );
  NAND2X0 U12794 ( .IN1(test_so33), .IN2(n11507), .QN(n12377) );
  NAND2X0 U12795 ( .IN1(n8983), .IN2(g3957), .QN(n12373) );
  NAND3X0 U12796 ( .IN1(n12378), .IN2(n12379), .IN3(n12380), .QN(g30453) );
  NAND2X0 U12797 ( .IN1(n12381), .IN2(n3765), .QN(n12380) );
  INVX0 U12798 ( .INP(n11505), .ZN(n12381) );
  NAND3X0 U12799 ( .IN1(n11505), .IN2(g3905), .IN3(n8873), .QN(n12379) );
  NAND2X0 U12800 ( .IN1(test_so33), .IN2(n12382), .QN(n11505) );
  NAND2X0 U12801 ( .IN1(n8969), .IN2(g3953), .QN(n12378) );
  NAND3X0 U12802 ( .IN1(n12383), .IN2(n12384), .IN3(n12385), .QN(g30452) );
  NAND2X0 U12803 ( .IN1(n12386), .IN2(n3765), .QN(n12385) );
  INVX0 U12804 ( .INP(n12387), .ZN(n12386) );
  NAND3X0 U12805 ( .IN1(n12387), .IN2(g3897), .IN3(n8873), .QN(n12384) );
  NAND2X0 U12806 ( .IN1(test_so33), .IN2(n12388), .QN(n12387) );
  NAND2X0 U12807 ( .IN1(test_so65), .IN2(n8952), .QN(n12383) );
  NAND3X0 U12808 ( .IN1(n12389), .IN2(n12390), .IN3(n12391), .QN(g30451) );
  NAND2X0 U12809 ( .IN1(n3951), .IN2(n12392), .QN(n12391) );
  NAND2X0 U12810 ( .IN1(n8969), .IN2(g3945), .QN(n12390) );
  NAND3X0 U12811 ( .IN1(n12393), .IN2(g3961), .IN3(n8873), .QN(n12389) );
  NAND2X0 U12812 ( .IN1(n11516), .IN2(n12392), .QN(n12393) );
  NAND3X0 U12813 ( .IN1(n12394), .IN2(n12395), .IN3(n12396), .QN(g30450) );
  NAND2X0 U12814 ( .IN1(n3951), .IN2(n11507), .QN(n12396) );
  NAND2X0 U12815 ( .IN1(n8970), .IN2(g3941), .QN(n12395) );
  NAND3X0 U12816 ( .IN1(n12397), .IN2(g3957), .IN3(n8873), .QN(n12394) );
  NAND2X0 U12817 ( .IN1(n11516), .IN2(n11507), .QN(n12397) );
  NAND3X0 U12818 ( .IN1(n12398), .IN2(n12399), .IN3(n12400), .QN(g30449) );
  NAND2X0 U12819 ( .IN1(n3951), .IN2(n12382), .QN(n12400) );
  NAND2X0 U12820 ( .IN1(n8970), .IN2(g3937), .QN(n12399) );
  NAND3X0 U12821 ( .IN1(n12401), .IN2(g3953), .IN3(n8874), .QN(n12398) );
  NAND2X0 U12822 ( .IN1(n11516), .IN2(n12382), .QN(n12401) );
  NAND3X0 U12823 ( .IN1(n12402), .IN2(n12403), .IN3(n12404), .QN(g30448) );
  NAND2X0 U12824 ( .IN1(n3951), .IN2(n12388), .QN(n12404) );
  NAND2X0 U12825 ( .IN1(n8970), .IN2(g3933), .QN(n12403) );
  NAND3X0 U12826 ( .IN1(test_so65), .IN2(n12405), .IN3(n8874), .QN(n12402) );
  NAND2X0 U12827 ( .IN1(n11516), .IN2(n12388), .QN(n12405) );
  INVX0 U12828 ( .INP(n1135), .ZN(n11516) );
  NAND2X0 U12829 ( .IN1(g3857), .IN2(g3863), .QN(n1135) );
  NAND3X0 U12830 ( .IN1(n12406), .IN2(n12407), .IN3(n12408), .QN(g30447) );
  NAND2X0 U12831 ( .IN1(n3957), .IN2(n12392), .QN(n12408) );
  NAND2X0 U12832 ( .IN1(n8970), .IN2(g3929), .QN(n12407) );
  NAND3X0 U12833 ( .IN1(n12409), .IN2(g3945), .IN3(n8874), .QN(n12406) );
  NAND2X0 U12834 ( .IN1(n11521), .IN2(n12392), .QN(n12409) );
  NAND3X0 U12835 ( .IN1(n12410), .IN2(n12411), .IN3(n12412), .QN(g30446) );
  NAND2X0 U12836 ( .IN1(n3957), .IN2(n11507), .QN(n12412) );
  NAND2X0 U12837 ( .IN1(n8971), .IN2(g3925), .QN(n12411) );
  NAND3X0 U12838 ( .IN1(n12413), .IN2(g3941), .IN3(n8874), .QN(n12410) );
  NAND2X0 U12839 ( .IN1(n11521), .IN2(n11507), .QN(n12413) );
  NAND3X0 U12840 ( .IN1(n12414), .IN2(n12415), .IN3(n12416), .QN(g30445) );
  NAND2X0 U12841 ( .IN1(n3957), .IN2(n12382), .QN(n12416) );
  NAND2X0 U12842 ( .IN1(n8971), .IN2(g3921), .QN(n12415) );
  NAND3X0 U12843 ( .IN1(n12417), .IN2(g3937), .IN3(n8874), .QN(n12414) );
  NAND2X0 U12844 ( .IN1(n11521), .IN2(n12382), .QN(n12417) );
  NAND3X0 U12845 ( .IN1(n12418), .IN2(n12419), .IN3(n12420), .QN(g30444) );
  NAND2X0 U12846 ( .IN1(n3957), .IN2(n12388), .QN(n12420) );
  NAND2X0 U12847 ( .IN1(n8971), .IN2(g3917), .QN(n12419) );
  NAND3X0 U12848 ( .IN1(n12421), .IN2(g3933), .IN3(n8874), .QN(n12418) );
  NAND2X0 U12849 ( .IN1(n11521), .IN2(n12388), .QN(n12421) );
  INVX0 U12850 ( .INP(n1136), .ZN(n11521) );
  NAND2X0 U12851 ( .IN1(n5572), .IN2(g3863), .QN(n1136) );
  NAND3X0 U12852 ( .IN1(n12422), .IN2(n12423), .IN3(n12424), .QN(g30443) );
  NAND2X0 U12853 ( .IN1(n3962), .IN2(n12392), .QN(n12424) );
  NAND2X0 U12854 ( .IN1(n8971), .IN2(g3909), .QN(n12423) );
  NAND3X0 U12855 ( .IN1(n12425), .IN2(g3929), .IN3(n8874), .QN(n12422) );
  NAND2X0 U12856 ( .IN1(n12426), .IN2(n12392), .QN(n12425) );
  NAND3X0 U12857 ( .IN1(n12427), .IN2(n12428), .IN3(n12429), .QN(g30442) );
  NAND2X0 U12858 ( .IN1(n3962), .IN2(n11507), .QN(n12429) );
  NAND2X0 U12859 ( .IN1(n8972), .IN2(g3901), .QN(n12428) );
  NAND3X0 U12860 ( .IN1(n12430), .IN2(g3925), .IN3(n8875), .QN(n12427) );
  NAND2X0 U12861 ( .IN1(n12426), .IN2(n11507), .QN(n12430) );
  INVX0 U12862 ( .INP(n830), .ZN(n11507) );
  NAND2X0 U12863 ( .IN1(n5387), .IN2(g3881), .QN(n830) );
  NAND3X0 U12864 ( .IN1(n12431), .IN2(n12432), .IN3(n12433), .QN(g30441) );
  NAND2X0 U12865 ( .IN1(n3962), .IN2(n12382), .QN(n12433) );
  NAND2X0 U12866 ( .IN1(n8972), .IN2(g3893), .QN(n12432) );
  NAND3X0 U12867 ( .IN1(n12434), .IN2(g3921), .IN3(n8875), .QN(n12431) );
  NAND2X0 U12868 ( .IN1(n12426), .IN2(n12382), .QN(n12434) );
  INVX0 U12869 ( .INP(n826), .ZN(n12382) );
  NAND2X0 U12870 ( .IN1(n5564), .IN2(g3873), .QN(n826) );
  NAND3X0 U12871 ( .IN1(n12435), .IN2(n12436), .IN3(n12437), .QN(g30440) );
  NAND2X0 U12872 ( .IN1(n3962), .IN2(n12388), .QN(n12437) );
  NAND2X0 U12873 ( .IN1(test_so24), .IN2(n9051), .QN(n12436) );
  NAND3X0 U12874 ( .IN1(n12438), .IN2(g3917), .IN3(n8875), .QN(n12435) );
  NAND2X0 U12875 ( .IN1(n12426), .IN2(n12388), .QN(n12438) );
  INVX0 U12876 ( .INP(n828), .ZN(n12388) );
  NAND2X0 U12877 ( .IN1(n5564), .IN2(n5387), .QN(n828) );
  INVX0 U12878 ( .INP(n1137), .ZN(n12426) );
  NAND2X0 U12879 ( .IN1(n8494), .IN2(g3857), .QN(n1137) );
  NAND3X0 U12880 ( .IN1(n12439), .IN2(n12440), .IN3(n12441), .QN(g30439) );
  NAND2X0 U12881 ( .IN1(n8972), .IN2(g3913), .QN(n12441) );
  NAND3X0 U12882 ( .IN1(n8895), .IN2(g3909), .IN3(n12442), .QN(n12440) );
  INVX0 U12883 ( .INP(n3967), .ZN(n12442) );
  NAND2X0 U12884 ( .IN1(n3967), .IN2(n3765), .QN(n12439) );
  NAND3X0 U12885 ( .IN1(n12443), .IN2(n12444), .IN3(n12445), .QN(g30438) );
  NAND2X0 U12886 ( .IN1(n8973), .IN2(g3905), .QN(n12445) );
  NAND3X0 U12887 ( .IN1(n8895), .IN2(g3901), .IN3(n12446), .QN(n12444) );
  INVX0 U12888 ( .INP(n3970), .ZN(n12446) );
  NAND2X0 U12889 ( .IN1(n3970), .IN2(n3765), .QN(n12443) );
  NAND3X0 U12890 ( .IN1(n12447), .IN2(n12448), .IN3(n12449), .QN(g30437) );
  NAND2X0 U12891 ( .IN1(n8973), .IN2(g3897), .QN(n12449) );
  NAND3X0 U12892 ( .IN1(n8895), .IN2(g3893), .IN3(n12450), .QN(n12448) );
  INVX0 U12893 ( .INP(n3972), .ZN(n12450) );
  NAND2X0 U12894 ( .IN1(n3972), .IN2(n3765), .QN(n12447) );
  NAND3X0 U12895 ( .IN1(n12451), .IN2(n12452), .IN3(n12453), .QN(g30436) );
  NAND2X0 U12896 ( .IN1(n8973), .IN2(g3881), .QN(n12453) );
  NAND3X0 U12897 ( .IN1(test_so24), .IN2(n8871), .IN3(n12454), .QN(n12452) );
  INVX0 U12898 ( .INP(n3974), .ZN(n12454) );
  NAND2X0 U12899 ( .IN1(n3974), .IN2(n3765), .QN(n12451) );
  NOR2X0 U12900 ( .IN1(g3857), .IN2(n11513), .QN(g30435) );
  NAND3X0 U12901 ( .IN1(n8895), .IN2(n8594), .IN3(n11503), .QN(n11513) );
  NAND3X0 U12902 ( .IN1(g4093), .IN2(g4087), .IN3(n3799), .QN(n11503) );
  NAND3X0 U12903 ( .IN1(n12455), .IN2(n12456), .IN3(n12457), .QN(g30434) );
  NAND2X0 U12904 ( .IN1(n8973), .IN2(g3610), .QN(n12457) );
  NAND2X0 U12905 ( .IN1(n12458), .IN2(g3614), .QN(n12456) );
  NAND2X0 U12906 ( .IN1(n12459), .IN2(n3765), .QN(n12455) );
  NAND3X0 U12907 ( .IN1(n12460), .IN2(n12461), .IN3(n12462), .QN(g30433) );
  NAND2X0 U12908 ( .IN1(n12463), .IN2(n3765), .QN(n12462) );
  INVX0 U12909 ( .INP(n12464), .ZN(n12463) );
  NAND3X0 U12910 ( .IN1(n12464), .IN2(g3562), .IN3(n8875), .QN(n12461) );
  NAND2X0 U12911 ( .IN1(n11529), .IN2(g3518), .QN(n12464) );
  NAND2X0 U12912 ( .IN1(n8973), .IN2(g3606), .QN(n12460) );
  NAND3X0 U12913 ( .IN1(n12465), .IN2(n12466), .IN3(n12467), .QN(g30432) );
  NAND2X0 U12914 ( .IN1(n12468), .IN2(n3765), .QN(n12467) );
  INVX0 U12915 ( .INP(n11527), .ZN(n12468) );
  NAND3X0 U12916 ( .IN1(n11527), .IN2(g3554), .IN3(n8875), .QN(n12466) );
  NAND2X0 U12917 ( .IN1(n12469), .IN2(g3518), .QN(n11527) );
  NAND2X0 U12918 ( .IN1(test_so43), .IN2(n8961), .QN(n12465) );
  NAND3X0 U12919 ( .IN1(n12470), .IN2(n12471), .IN3(n12472), .QN(g30431) );
  NAND2X0 U12920 ( .IN1(n12473), .IN2(n3765), .QN(n12472) );
  INVX0 U12921 ( .INP(n12474), .ZN(n12473) );
  NAND3X0 U12922 ( .IN1(n12474), .IN2(g3546), .IN3(n8875), .QN(n12471) );
  NAND2X0 U12923 ( .IN1(n12475), .IN2(g3518), .QN(n12474) );
  NAND2X0 U12924 ( .IN1(n8974), .IN2(g3598), .QN(n12470) );
  NAND3X0 U12925 ( .IN1(n12476), .IN2(n12477), .IN3(n12478), .QN(g30430) );
  NAND2X0 U12926 ( .IN1(n3984), .IN2(n12479), .QN(n12478) );
  NAND2X0 U12927 ( .IN1(n8974), .IN2(g3594), .QN(n12477) );
  NAND3X0 U12928 ( .IN1(n12480), .IN2(g3610), .IN3(n8875), .QN(n12476) );
  NAND2X0 U12929 ( .IN1(n12479), .IN2(n11538), .QN(n12480) );
  NAND3X0 U12930 ( .IN1(n12481), .IN2(n12482), .IN3(n12483), .QN(g30429) );
  NAND2X0 U12931 ( .IN1(n3984), .IN2(n11529), .QN(n12483) );
  NAND2X0 U12932 ( .IN1(n8974), .IN2(g3590), .QN(n12482) );
  NAND3X0 U12933 ( .IN1(n12484), .IN2(g3606), .IN3(n8876), .QN(n12481) );
  NAND2X0 U12934 ( .IN1(n11529), .IN2(n11538), .QN(n12484) );
  NAND3X0 U12935 ( .IN1(n12485), .IN2(n12486), .IN3(n12487), .QN(g30428) );
  NAND2X0 U12936 ( .IN1(n3984), .IN2(n12469), .QN(n12487) );
  NAND2X0 U12937 ( .IN1(n8975), .IN2(g3586), .QN(n12486) );
  NAND3X0 U12938 ( .IN1(test_so43), .IN2(n12488), .IN3(n8876), .QN(n12485) );
  NAND2X0 U12939 ( .IN1(n12469), .IN2(n11538), .QN(n12488) );
  NAND3X0 U12940 ( .IN1(n12489), .IN2(n12490), .IN3(n12491), .QN(g30427) );
  NAND2X0 U12941 ( .IN1(n3984), .IN2(n12475), .QN(n12491) );
  NAND2X0 U12942 ( .IN1(n8975), .IN2(g3582), .QN(n12490) );
  NAND3X0 U12943 ( .IN1(n12492), .IN2(g3598), .IN3(n8876), .QN(n12489) );
  NAND2X0 U12944 ( .IN1(n12475), .IN2(n11538), .QN(n12492) );
  INVX0 U12945 ( .INP(n99), .ZN(n11538) );
  NAND2X0 U12946 ( .IN1(g3506), .IN2(g3512), .QN(n99) );
  NAND3X0 U12947 ( .IN1(n12493), .IN2(n12494), .IN3(n12495), .QN(g30426) );
  NAND2X0 U12948 ( .IN1(n3990), .IN2(n12479), .QN(n12495) );
  NAND2X0 U12949 ( .IN1(n8975), .IN2(g3578), .QN(n12494) );
  NAND3X0 U12950 ( .IN1(n12496), .IN2(g3594), .IN3(n8876), .QN(n12493) );
  NAND2X0 U12951 ( .IN1(n11543), .IN2(n12479), .QN(n12496) );
  NAND3X0 U12952 ( .IN1(n12497), .IN2(n12498), .IN3(n12499), .QN(g30425) );
  NAND2X0 U12953 ( .IN1(n3990), .IN2(n11529), .QN(n12499) );
  NAND2X0 U12954 ( .IN1(n8976), .IN2(g3574), .QN(n12498) );
  NAND3X0 U12955 ( .IN1(n12500), .IN2(g3590), .IN3(n8876), .QN(n12497) );
  NAND2X0 U12956 ( .IN1(n11543), .IN2(n11529), .QN(n12500) );
  NAND3X0 U12957 ( .IN1(n12501), .IN2(n12502), .IN3(n12503), .QN(g30424) );
  NAND2X0 U12958 ( .IN1(n3990), .IN2(n12469), .QN(n12503) );
  NAND2X0 U12959 ( .IN1(n8976), .IN2(g3570), .QN(n12502) );
  NAND3X0 U12960 ( .IN1(n12504), .IN2(g3586), .IN3(n8876), .QN(n12501) );
  NAND2X0 U12961 ( .IN1(n11543), .IN2(n12469), .QN(n12504) );
  NAND3X0 U12962 ( .IN1(n12505), .IN2(n12506), .IN3(n12507), .QN(g30423) );
  NAND2X0 U12963 ( .IN1(n3990), .IN2(n12475), .QN(n12507) );
  NAND2X0 U12964 ( .IN1(n8976), .IN2(g3566), .QN(n12506) );
  NAND3X0 U12965 ( .IN1(n12508), .IN2(g3582), .IN3(n8876), .QN(n12505) );
  NAND2X0 U12966 ( .IN1(n11543), .IN2(n12475), .QN(n12508) );
  INVX0 U12967 ( .INP(n100), .ZN(n11543) );
  NAND2X0 U12968 ( .IN1(n5576), .IN2(g3512), .QN(n100) );
  NAND3X0 U12969 ( .IN1(n12509), .IN2(n12510), .IN3(n12511), .QN(g30422) );
  NAND2X0 U12970 ( .IN1(n3995), .IN2(n12479), .QN(n12511) );
  NAND2X0 U12971 ( .IN1(n8977), .IN2(g3558), .QN(n12510) );
  NAND3X0 U12972 ( .IN1(n12512), .IN2(g3578), .IN3(n8876), .QN(n12509) );
  NAND2X0 U12973 ( .IN1(n12513), .IN2(n12479), .QN(n12512) );
  NAND3X0 U12974 ( .IN1(n12514), .IN2(n12515), .IN3(n12516), .QN(g30421) );
  NAND2X0 U12975 ( .IN1(n3995), .IN2(n11529), .QN(n12516) );
  NAND2X0 U12976 ( .IN1(n8977), .IN2(g3550), .QN(n12515) );
  NAND3X0 U12977 ( .IN1(n12517), .IN2(g3574), .IN3(n8876), .QN(n12514) );
  NAND2X0 U12978 ( .IN1(n12513), .IN2(n11529), .QN(n12517) );
  INVX0 U12979 ( .INP(n429), .ZN(n11529) );
  NAND2X0 U12980 ( .IN1(n5383), .IN2(g3530), .QN(n429) );
  NAND3X0 U12981 ( .IN1(n12518), .IN2(n12519), .IN3(n12520), .QN(g30420) );
  NAND2X0 U12982 ( .IN1(n3995), .IN2(n12469), .QN(n12520) );
  NAND2X0 U12983 ( .IN1(n8971), .IN2(g3542), .QN(n12519) );
  NAND3X0 U12984 ( .IN1(n12521), .IN2(g3570), .IN3(n8877), .QN(n12518) );
  NAND2X0 U12985 ( .IN1(n12513), .IN2(n12469), .QN(n12521) );
  INVX0 U12986 ( .INP(n433), .ZN(n12469) );
  NAND2X0 U12987 ( .IN1(n5569), .IN2(g3522), .QN(n433) );
  NAND3X0 U12988 ( .IN1(n12522), .IN2(n12523), .IN3(n12524), .QN(g30419) );
  NAND2X0 U12989 ( .IN1(n3995), .IN2(n12475), .QN(n12524) );
  NAND2X0 U12990 ( .IN1(n8978), .IN2(g3538), .QN(n12523) );
  NAND3X0 U12991 ( .IN1(n12525), .IN2(g3566), .IN3(n8877), .QN(n12522) );
  NAND2X0 U12992 ( .IN1(n12513), .IN2(n12475), .QN(n12525) );
  INVX0 U12993 ( .INP(n431), .ZN(n12475) );
  NAND2X0 U12994 ( .IN1(n5383), .IN2(n5569), .QN(n431) );
  INVX0 U12995 ( .INP(n101), .ZN(n12513) );
  NAND2X0 U12996 ( .IN1(n8490), .IN2(g3506), .QN(n101) );
  NAND3X0 U12997 ( .IN1(n12526), .IN2(n12527), .IN3(n12528), .QN(g30418) );
  NAND2X0 U12998 ( .IN1(n8978), .IN2(g3562), .QN(n12528) );
  NAND3X0 U12999 ( .IN1(n8897), .IN2(g3558), .IN3(n12529), .QN(n12527) );
  INVX0 U13000 ( .INP(n4000), .ZN(n12529) );
  NAND2X0 U13001 ( .IN1(n4000), .IN2(n3765), .QN(n12526) );
  NAND3X0 U13002 ( .IN1(n12530), .IN2(n12531), .IN3(n12532), .QN(g30417) );
  NAND2X0 U13003 ( .IN1(n8978), .IN2(g3554), .QN(n12532) );
  NAND3X0 U13004 ( .IN1(n8897), .IN2(g3550), .IN3(n12533), .QN(n12531) );
  INVX0 U13005 ( .INP(n4003), .ZN(n12533) );
  NAND2X0 U13006 ( .IN1(n4003), .IN2(n3765), .QN(n12530) );
  NAND3X0 U13007 ( .IN1(n12534), .IN2(n12535), .IN3(n12536), .QN(g30416) );
  NAND2X0 U13008 ( .IN1(n8978), .IN2(g3546), .QN(n12536) );
  NAND3X0 U13009 ( .IN1(n8897), .IN2(g3542), .IN3(n12537), .QN(n12535) );
  INVX0 U13010 ( .INP(n4005), .ZN(n12537) );
  NAND2X0 U13011 ( .IN1(n4005), .IN2(n3765), .QN(n12534) );
  NAND3X0 U13012 ( .IN1(n12538), .IN2(n12539), .IN3(n12540), .QN(g30415) );
  NAND2X0 U13013 ( .IN1(n8978), .IN2(g3530), .QN(n12540) );
  NAND3X0 U13014 ( .IN1(n8897), .IN2(g3538), .IN3(n12541), .QN(n12539) );
  INVX0 U13015 ( .INP(n4007), .ZN(n12541) );
  NAND2X0 U13016 ( .IN1(n4007), .IN2(n3765), .QN(n12538) );
  NOR2X0 U13017 ( .IN1(g3506), .IN2(n11535), .QN(g30414) );
  NAND3X0 U13018 ( .IN1(n11525), .IN2(n8869), .IN3(n5645), .QN(n11535) );
  NAND3X0 U13019 ( .IN1(n5480), .IN2(g4093), .IN3(n3799), .QN(n11525) );
  NAND3X0 U13020 ( .IN1(n12542), .IN2(n12543), .IN3(n12544), .QN(g30413) );
  NAND2X0 U13021 ( .IN1(test_so84), .IN2(n9052), .QN(n12544) );
  NAND2X0 U13022 ( .IN1(n12545), .IN2(g3263), .QN(n12543) );
  NAND2X0 U13023 ( .IN1(n3765), .IN2(n10834), .QN(n12542) );
  NAND3X0 U13024 ( .IN1(n12546), .IN2(n12547), .IN3(n12548), .QN(g30412) );
  NAND2X0 U13025 ( .IN1(n12549), .IN2(n3765), .QN(n12548) );
  INVX0 U13026 ( .INP(n12550), .ZN(n12549) );
  NAND3X0 U13027 ( .IN1(n12550), .IN2(g3211), .IN3(n8883), .QN(n12547) );
  NAND2X0 U13028 ( .IN1(n12551), .IN2(g3167), .QN(n12550) );
  NAND2X0 U13029 ( .IN1(n8979), .IN2(g3255), .QN(n12546) );
  NAND3X0 U13030 ( .IN1(n12552), .IN2(n12553), .IN3(n12554), .QN(g30411) );
  NAND2X0 U13031 ( .IN1(n12555), .IN2(n3765), .QN(n12554) );
  INVX0 U13032 ( .INP(n11550), .ZN(n12555) );
  NAND3X0 U13033 ( .IN1(n11550), .IN2(g3203), .IN3(n8877), .QN(n12553) );
  NAND2X0 U13034 ( .IN1(n12556), .IN2(g3167), .QN(n11550) );
  NAND2X0 U13035 ( .IN1(n8979), .IN2(g3251), .QN(n12552) );
  NAND3X0 U13036 ( .IN1(n12557), .IN2(n12558), .IN3(n12559), .QN(g30410) );
  NAND2X0 U13037 ( .IN1(n12560), .IN2(n3765), .QN(n12559) );
  INVX0 U13038 ( .INP(n12561), .ZN(n12560) );
  NAND3X0 U13039 ( .IN1(test_so88), .IN2(n12561), .IN3(n8877), .QN(n12558) );
  NAND2X0 U13040 ( .IN1(n12562), .IN2(g3167), .QN(n12561) );
  NAND2X0 U13041 ( .IN1(n8979), .IN2(g3247), .QN(n12557) );
  NAND3X0 U13042 ( .IN1(n12563), .IN2(n12564), .IN3(n12565), .QN(g30409) );
  NAND2X0 U13043 ( .IN1(n4015), .IN2(n12566), .QN(n12565) );
  NAND2X0 U13044 ( .IN1(n8979), .IN2(g3243), .QN(n12564) );
  NAND3X0 U13045 ( .IN1(test_so84), .IN2(n12567), .IN3(n8877), .QN(n12563) );
  NAND2X0 U13046 ( .IN1(n11557), .IN2(n12566), .QN(n12567) );
  NAND3X0 U13047 ( .IN1(n12568), .IN2(n12569), .IN3(n12570), .QN(g30408) );
  NAND2X0 U13048 ( .IN1(n4015), .IN2(n12551), .QN(n12570) );
  NAND2X0 U13049 ( .IN1(n8979), .IN2(g3239), .QN(n12569) );
  NAND3X0 U13050 ( .IN1(n12571), .IN2(g3255), .IN3(n8877), .QN(n12568) );
  NAND2X0 U13051 ( .IN1(n11557), .IN2(n12551), .QN(n12571) );
  NAND3X0 U13052 ( .IN1(n12572), .IN2(n12573), .IN3(n12574), .QN(g30407) );
  NAND2X0 U13053 ( .IN1(n4015), .IN2(n12556), .QN(n12574) );
  NAND2X0 U13054 ( .IN1(n8980), .IN2(g3235), .QN(n12573) );
  NAND3X0 U13055 ( .IN1(n12575), .IN2(g3251), .IN3(n8893), .QN(n12572) );
  NAND2X0 U13056 ( .IN1(n11557), .IN2(n12556), .QN(n12575) );
  NAND3X0 U13057 ( .IN1(n12576), .IN2(n12577), .IN3(n12578), .QN(g30406) );
  NAND2X0 U13058 ( .IN1(n4015), .IN2(n12562), .QN(n12578) );
  NAND2X0 U13059 ( .IN1(n8980), .IN2(g3231), .QN(n12577) );
  NAND3X0 U13060 ( .IN1(n12579), .IN2(g3247), .IN3(n8890), .QN(n12576) );
  NAND2X0 U13061 ( .IN1(n11557), .IN2(n12562), .QN(n12579) );
  INVX0 U13062 ( .INP(n112), .ZN(n11557) );
  NAND2X0 U13063 ( .IN1(g3155), .IN2(g3161), .QN(n112) );
  NAND3X0 U13064 ( .IN1(n12580), .IN2(n12581), .IN3(n12582), .QN(g30405) );
  NAND2X0 U13065 ( .IN1(n4022), .IN2(n12566), .QN(n12582) );
  NAND2X0 U13066 ( .IN1(n8980), .IN2(g3227), .QN(n12581) );
  NAND3X0 U13067 ( .IN1(n12583), .IN2(g3243), .IN3(n8890), .QN(n12580) );
  NAND2X0 U13068 ( .IN1(n11563), .IN2(n12566), .QN(n12583) );
  NAND3X0 U13069 ( .IN1(n12584), .IN2(n12585), .IN3(n12586), .QN(g30404) );
  NAND2X0 U13070 ( .IN1(n4022), .IN2(n12551), .QN(n12586) );
  NAND2X0 U13071 ( .IN1(n8980), .IN2(g3223), .QN(n12585) );
  NAND3X0 U13072 ( .IN1(n12587), .IN2(g3239), .IN3(n8890), .QN(n12584) );
  NAND2X0 U13073 ( .IN1(n11563), .IN2(n12551), .QN(n12587) );
  NAND3X0 U13074 ( .IN1(n12588), .IN2(n12589), .IN3(n12590), .QN(g30403) );
  NAND2X0 U13075 ( .IN1(n4022), .IN2(n12556), .QN(n12590) );
  NAND2X0 U13076 ( .IN1(n8981), .IN2(g3219), .QN(n12589) );
  NAND3X0 U13077 ( .IN1(n12591), .IN2(g3235), .IN3(n8890), .QN(n12588) );
  NAND2X0 U13078 ( .IN1(n11563), .IN2(n12556), .QN(n12591) );
  NAND3X0 U13079 ( .IN1(n12592), .IN2(n12593), .IN3(n12594), .QN(g30402) );
  NAND2X0 U13080 ( .IN1(n4022), .IN2(n12562), .QN(n12594) );
  NAND2X0 U13081 ( .IN1(n8981), .IN2(g3215), .QN(n12593) );
  NAND3X0 U13082 ( .IN1(n12595), .IN2(g3231), .IN3(n8891), .QN(n12592) );
  NAND2X0 U13083 ( .IN1(n11563), .IN2(n12562), .QN(n12595) );
  INVX0 U13084 ( .INP(n114), .ZN(n11563) );
  NAND2X0 U13085 ( .IN1(n5366), .IN2(g3161), .QN(n114) );
  NAND3X0 U13086 ( .IN1(n12596), .IN2(n12597), .IN3(n12598), .QN(g30401) );
  NAND2X0 U13087 ( .IN1(n4027), .IN2(n12566), .QN(n12598) );
  NAND2X0 U13088 ( .IN1(n8981), .IN2(g3207), .QN(n12597) );
  NAND3X0 U13089 ( .IN1(n12599), .IN2(g3227), .IN3(n8891), .QN(n12596) );
  NAND2X0 U13090 ( .IN1(n12600), .IN2(n12566), .QN(n12599) );
  INVX0 U13091 ( .INP(n530), .ZN(n12566) );
  NAND3X0 U13092 ( .IN1(n12601), .IN2(n12602), .IN3(n12603), .QN(g30400) );
  NAND2X0 U13093 ( .IN1(n4027), .IN2(n12551), .QN(n12603) );
  NAND2X0 U13094 ( .IN1(n8981), .IN2(g3199), .QN(n12602) );
  NAND3X0 U13095 ( .IN1(n12604), .IN2(g3223), .IN3(n8891), .QN(n12601) );
  NAND2X0 U13096 ( .IN1(n12600), .IN2(n12551), .QN(n12604) );
  INVX0 U13097 ( .INP(n526), .ZN(n12551) );
  NAND2X0 U13098 ( .IN1(n5603), .IN2(g3179), .QN(n526) );
  NAND3X0 U13099 ( .IN1(n12605), .IN2(n12606), .IN3(n12607), .QN(g30399) );
  NAND2X0 U13100 ( .IN1(n4027), .IN2(n12556), .QN(n12607) );
  NAND2X0 U13101 ( .IN1(n8981), .IN2(g3191), .QN(n12606) );
  NAND3X0 U13102 ( .IN1(n12608), .IN2(g3219), .IN3(n8891), .QN(n12605) );
  NAND2X0 U13103 ( .IN1(n12600), .IN2(n12556), .QN(n12608) );
  INVX0 U13104 ( .INP(n528), .ZN(n12556) );
  NAND2X0 U13105 ( .IN1(n5390), .IN2(g3171), .QN(n528) );
  NAND3X0 U13106 ( .IN1(n12609), .IN2(n12610), .IN3(n12611), .QN(g30398) );
  NAND2X0 U13107 ( .IN1(n4027), .IN2(n12562), .QN(n12611) );
  NAND2X0 U13108 ( .IN1(n8982), .IN2(g3187), .QN(n12610) );
  NAND3X0 U13109 ( .IN1(n12612), .IN2(g3215), .IN3(n8892), .QN(n12609) );
  NAND2X0 U13110 ( .IN1(n12600), .IN2(n12562), .QN(n12612) );
  INVX0 U13111 ( .INP(n527), .ZN(n12562) );
  NAND2X0 U13112 ( .IN1(n5603), .IN2(n5390), .QN(n527) );
  INVX0 U13113 ( .INP(n113), .ZN(n12600) );
  NAND2X0 U13114 ( .IN1(n8475), .IN2(g3155), .QN(n113) );
  NAND3X0 U13115 ( .IN1(n12613), .IN2(n12614), .IN3(n12615), .QN(g30397) );
  NAND2X0 U13116 ( .IN1(n8982), .IN2(g3211), .QN(n12615) );
  NAND3X0 U13117 ( .IN1(n8894), .IN2(g3207), .IN3(n12616), .QN(n12614) );
  INVX0 U13118 ( .INP(n4032), .ZN(n12616) );
  NAND2X0 U13119 ( .IN1(n4032), .IN2(n3765), .QN(n12613) );
  NAND3X0 U13120 ( .IN1(n12617), .IN2(n12618), .IN3(n12619), .QN(g30396) );
  NAND2X0 U13121 ( .IN1(n8982), .IN2(g3203), .QN(n12619) );
  NAND3X0 U13122 ( .IN1(n8894), .IN2(g3199), .IN3(n12620), .QN(n12618) );
  INVX0 U13123 ( .INP(n4035), .ZN(n12620) );
  NAND2X0 U13124 ( .IN1(n4035), .IN2(n3765), .QN(n12617) );
  NAND3X0 U13125 ( .IN1(n12621), .IN2(n12622), .IN3(n12623), .QN(g30395) );
  NAND2X0 U13126 ( .IN1(test_so88), .IN2(n9053), .QN(n12623) );
  NAND3X0 U13127 ( .IN1(n8893), .IN2(g3191), .IN3(n12624), .QN(n12622) );
  INVX0 U13128 ( .INP(n4037), .ZN(n12624) );
  NAND2X0 U13129 ( .IN1(n4037), .IN2(n3765), .QN(n12621) );
  NAND3X0 U13130 ( .IN1(n12625), .IN2(n12626), .IN3(n12627), .QN(g30394) );
  NAND2X0 U13131 ( .IN1(n8983), .IN2(g3179), .QN(n12627) );
  NAND3X0 U13132 ( .IN1(n8896), .IN2(g3187), .IN3(n12628), .QN(n12626) );
  INVX0 U13133 ( .INP(n4039), .ZN(n12628) );
  NAND2X0 U13134 ( .IN1(n4039), .IN2(n3765), .QN(n12625) );
  NOR3X0 U13135 ( .IN1(n11558), .IN2(n8925), .IN3(g3155), .QN(g30393) );
  NAND2X0 U13136 ( .IN1(n5652), .IN2(n11549), .QN(n11558) );
  NAND2X0 U13137 ( .IN1(n3799), .IN2(n10824), .QN(n11549) );
  NAND2X0 U13138 ( .IN1(n12629), .IN2(n12630), .QN(g30392) );
  NAND2X0 U13139 ( .IN1(n8983), .IN2(g2803), .QN(n12630) );
  NAND2X0 U13140 ( .IN1(n12631), .IN2(n12632), .QN(g30391) );
  NAND2X0 U13141 ( .IN1(n8983), .IN2(g2771), .QN(n12632) );
  NAND2X0 U13142 ( .IN1(n12629), .IN2(n12633), .QN(g30390) );
  NAND2X0 U13143 ( .IN1(g2834), .IN2(n9054), .QN(n12633) );
  NAND2X0 U13144 ( .IN1(n12634), .IN2(n8914), .QN(n12629) );
  NAND2X0 U13145 ( .IN1(n12635), .IN2(n12636), .QN(n12634) );
  NAND4X0 U13146 ( .IN1(n12637), .IN2(n12638), .IN3(n12639), .IN4(n12640), 
        .QN(n12636) );
  NOR2X0 U13147 ( .IN1(n12641), .IN2(n12642), .QN(n12639) );
  NOR2X0 U13148 ( .IN1(n12643), .IN2(g2236), .QN(n12642) );
  NOR2X0 U13149 ( .IN1(n1249), .IN2(g2370), .QN(n12641) );
  NAND2X0 U13150 ( .IN1(n8512), .IN2(n12644), .QN(n12638) );
  NAND2X0 U13151 ( .IN1(n8484), .IN2(n12645), .QN(n12637) );
  NAND4X0 U13152 ( .IN1(n12646), .IN2(n12647), .IN3(n12648), .IN4(n12649), 
        .QN(n12635) );
  NOR2X0 U13153 ( .IN1(n12650), .IN2(n12651), .QN(n12648) );
  NOR2X0 U13154 ( .IN1(n5545), .IN2(n12643), .QN(n12651) );
  NOR2X0 U13155 ( .IN1(n5379), .IN2(n1249), .QN(n12650) );
  NAND2X0 U13156 ( .IN1(n12644), .IN2(g2819), .QN(n12647) );
  NAND2X0 U13157 ( .IN1(n12645), .IN2(g2815), .QN(n12646) );
  NAND2X0 U13158 ( .IN1(n12631), .IN2(n12652), .QN(g30389) );
  NAND2X0 U13159 ( .IN1(g2831), .IN2(n9054), .QN(n12652) );
  NAND2X0 U13160 ( .IN1(n12653), .IN2(n8914), .QN(n12631) );
  NAND2X0 U13161 ( .IN1(n12654), .IN2(n12655), .QN(n12653) );
  NAND4X0 U13162 ( .IN1(n12656), .IN2(n12657), .IN3(n12658), .IN4(n12640), 
        .QN(n12655) );
  NOR2X0 U13163 ( .IN1(n12659), .IN2(n12660), .QN(n12658) );
  NOR2X0 U13164 ( .IN1(n12643), .IN2(g1677), .QN(n12660) );
  NOR2X0 U13165 ( .IN1(n1249), .IN2(g1811), .QN(n12659) );
  NAND2X0 U13166 ( .IN1(n8513), .IN2(n12644), .QN(n12657) );
  NAND2X0 U13167 ( .IN1(n12645), .IN2(n8633), .QN(n12656) );
  NAND4X0 U13168 ( .IN1(n12661), .IN2(n12662), .IN3(n12663), .IN4(n12649), 
        .QN(n12654) );
  INVX0 U13169 ( .INP(n12640), .ZN(n12649) );
  NAND3X0 U13170 ( .IN1(n3653), .IN2(n12664), .IN3(n5600), .QN(n12640) );
  NOR3X0 U13171 ( .IN1(g2741), .IN2(test_so30), .IN3(g2748), .QN(n3653) );
  NOR2X0 U13172 ( .IN1(n12665), .IN2(n12666), .QN(n12663) );
  NOR2X0 U13173 ( .IN1(n5544), .IN2(n12643), .QN(n12666) );
  NOR2X0 U13174 ( .IN1(n5378), .IN2(n1249), .QN(n12665) );
  NAND2X0 U13175 ( .IN1(n12644), .IN2(g2787), .QN(n12662) );
  NAND2X0 U13176 ( .IN1(n12645), .IN2(g2783), .QN(n12661) );
  NAND2X0 U13177 ( .IN1(n12667), .IN2(n12668), .QN(g30388) );
  NAND2X0 U13178 ( .IN1(n12669), .IN2(n3730), .QN(n12668) );
  XOR2X1 U13179 ( .IN1(n3506), .IN2(n5349), .Q(n12669) );
  NAND2X0 U13180 ( .IN1(n12670), .IN2(g2735), .QN(n3506) );
  NAND2X0 U13181 ( .IN1(n8983), .IN2(g2735), .QN(n12667) );
  NAND3X0 U13182 ( .IN1(n12671), .IN2(n12672), .IN3(n12673), .QN(g30387) );
  INVX0 U13183 ( .INP(n12674), .ZN(n12673) );
  NOR2X0 U13184 ( .IN1(n12675), .IN2(n15224), .QN(n12674) );
  INVX0 U13185 ( .INP(n12676), .ZN(n12672) );
  NOR2X0 U13186 ( .IN1(n12677), .IN2(n5777), .QN(n12676) );
  NOR2X0 U13187 ( .IN1(n12678), .IN2(n8943), .QN(n12677) );
  NOR2X0 U13188 ( .IN1(n12679), .IN2(n5457), .QN(n12678) );
  NAND3X0 U13189 ( .IN1(n12680), .IN2(n5457), .IN3(n5777), .QN(n12671) );
  NAND2X0 U13190 ( .IN1(n12681), .IN2(n12682), .QN(g30386) );
  INVX0 U13191 ( .INP(n12683), .ZN(n12682) );
  NOR2X0 U13192 ( .IN1(n12675), .IN2(n5777), .QN(n12683) );
  NAND2X0 U13193 ( .IN1(n12675), .IN2(g2675), .QN(n12681) );
  NAND3X0 U13194 ( .IN1(n12684), .IN2(n12685), .IN3(n12686), .QN(g30385) );
  NAND2X0 U13195 ( .IN1(n8967), .IN2(g2657), .QN(n12686) );
  INVX0 U13196 ( .INP(n12687), .ZN(n12685) );
  NOR2X0 U13197 ( .IN1(n12675), .IN2(n5418), .QN(n12687) );
  NAND2X0 U13198 ( .IN1(n12679), .IN2(n8914), .QN(n12675) );
  NAND2X0 U13199 ( .IN1(n12680), .IN2(n5418), .QN(n12684) );
  NAND3X0 U13200 ( .IN1(n12688), .IN2(n12689), .IN3(n12690), .QN(g30384) );
  NAND2X0 U13201 ( .IN1(n8983), .IN2(g2652), .QN(n12690) );
  NAND3X0 U13202 ( .IN1(n3517), .IN2(n12691), .IN3(n8574), .QN(n12689) );
  XOR2X1 U13203 ( .IN1(n8231), .IN2(n8106), .Q(n12691) );
  NAND2X0 U13204 ( .IN1(n12692), .IN2(g2657), .QN(n12688) );
  NAND2X0 U13205 ( .IN1(n11575), .IN2(n12693), .QN(n12692) );
  NAND2X0 U13206 ( .IN1(n8902), .IN2(n11587), .QN(n12693) );
  NAND2X0 U13207 ( .IN1(n12694), .IN2(n12695), .QN(g30383) );
  NAND2X0 U13208 ( .IN1(test_so66), .IN2(n9054), .QN(n12695) );
  NAND2X0 U13209 ( .IN1(n12696), .IN2(n8914), .QN(n12694) );
  NAND2X0 U13210 ( .IN1(n12697), .IN2(n12698), .QN(n12696) );
  NAND2X0 U13211 ( .IN1(test_so34), .IN2(n12699), .QN(n12698) );
  NAND2X0 U13212 ( .IN1(n12700), .IN2(n12701), .QN(n12697) );
  NAND2X0 U13213 ( .IN1(n5351), .IN2(g2599), .QN(n12701) );
  INVX0 U13214 ( .INP(n12699), .ZN(n12700) );
  NAND3X0 U13215 ( .IN1(n12702), .IN2(g2610), .IN3(n5508), .QN(n12699) );
  NAND3X0 U13216 ( .IN1(n12703), .IN2(n12704), .IN3(n12705), .QN(g30382) );
  NAND2X0 U13217 ( .IN1(n12706), .IN2(n9295), .QN(n12705) );
  INVX0 U13218 ( .INP(n12707), .ZN(n12704) );
  NOR2X0 U13219 ( .IN1(n12708), .IN2(n5782), .QN(n12707) );
  NOR2X0 U13220 ( .IN1(n12709), .IN2(n8938), .QN(n12708) );
  NOR2X0 U13221 ( .IN1(n12710), .IN2(n5461), .QN(n12709) );
  NAND3X0 U13222 ( .IN1(n12711), .IN2(n5461), .IN3(n5782), .QN(n12703) );
  NAND2X0 U13223 ( .IN1(n12712), .IN2(n12713), .QN(g30381) );
  INVX0 U13224 ( .INP(n12714), .ZN(n12713) );
  NOR2X0 U13225 ( .IN1(n12715), .IN2(n5782), .QN(n12714) );
  NAND2X0 U13226 ( .IN1(n12715), .IN2(g2541), .QN(n12712) );
  NAND3X0 U13227 ( .IN1(n12716), .IN2(n12717), .IN3(n12718), .QN(g30380) );
  NAND2X0 U13228 ( .IN1(n8983), .IN2(g2523), .QN(n12718) );
  NAND2X0 U13229 ( .IN1(n12706), .IN2(g2527), .QN(n12717) );
  INVX0 U13230 ( .INP(n12715), .ZN(n12706) );
  NAND2X0 U13231 ( .IN1(n12710), .IN2(n8914), .QN(n12715) );
  NAND2X0 U13232 ( .IN1(n12711), .IN2(n5420), .QN(n12716) );
  NAND3X0 U13233 ( .IN1(n12719), .IN2(n12720), .IN3(n12721), .QN(g30379) );
  NAND2X0 U13234 ( .IN1(n8982), .IN2(g2518), .QN(n12721) );
  NAND3X0 U13235 ( .IN1(n3536), .IN2(n12722), .IN3(n8580), .QN(n12720) );
  XOR2X1 U13236 ( .IN1(n8230), .IN2(n8103), .Q(n12722) );
  NAND2X0 U13237 ( .IN1(n12723), .IN2(g2523), .QN(n12719) );
  NAND2X0 U13238 ( .IN1(n11596), .IN2(n12724), .QN(n12723) );
  NAND2X0 U13239 ( .IN1(n8902), .IN2(n11608), .QN(n12724) );
  NAND2X0 U13240 ( .IN1(n12725), .IN2(n12726), .QN(g30378) );
  NAND2X0 U13241 ( .IN1(n8982), .IN2(g2441), .QN(n12726) );
  NAND2X0 U13242 ( .IN1(n12727), .IN2(n8914), .QN(n12725) );
  NAND2X0 U13243 ( .IN1(n12728), .IN2(n12729), .QN(n12727) );
  NAND2X0 U13244 ( .IN1(n12730), .IN2(g2461), .QN(n12729) );
  NAND2X0 U13245 ( .IN1(n12731), .IN2(n12732), .QN(n12728) );
  NAND2X0 U13246 ( .IN1(g2465), .IN2(n8585), .QN(n12732) );
  INVX0 U13247 ( .INP(n12730), .ZN(n12731) );
  NAND3X0 U13248 ( .IN1(n12733), .IN2(g2476), .IN3(n5509), .QN(n12730) );
  NAND3X0 U13249 ( .IN1(n12734), .IN2(n12735), .IN3(n12736), .QN(g30377) );
  NAND2X0 U13250 ( .IN1(n12737), .IN2(n9324), .QN(n12736) );
  NAND2X0 U13251 ( .IN1(test_so89), .IN2(n12738), .QN(n12735) );
  INVX0 U13252 ( .INP(n12739), .ZN(n12738) );
  NOR2X0 U13253 ( .IN1(n12740), .IN2(n8933), .QN(n12739) );
  NOR2X0 U13254 ( .IN1(n12741), .IN2(n5459), .QN(n12740) );
  NAND3X0 U13255 ( .IN1(n12742), .IN2(n5459), .IN3(n8615), .QN(n12734) );
  NAND2X0 U13256 ( .IN1(n12743), .IN2(n12744), .QN(g30376) );
  NAND2X0 U13257 ( .IN1(test_so89), .IN2(n12737), .QN(n12744) );
  NAND2X0 U13258 ( .IN1(n12745), .IN2(g2407), .QN(n12743) );
  NAND3X0 U13259 ( .IN1(n12746), .IN2(n12747), .IN3(n12748), .QN(g30375) );
  NAND2X0 U13260 ( .IN1(n8982), .IN2(g2389), .QN(n12748) );
  NAND2X0 U13261 ( .IN1(n12737), .IN2(g2393), .QN(n12747) );
  INVX0 U13262 ( .INP(n12745), .ZN(n12737) );
  NAND2X0 U13263 ( .IN1(n12741), .IN2(n8914), .QN(n12745) );
  NAND2X0 U13264 ( .IN1(n12742), .IN2(n5421), .QN(n12746) );
  NAND3X0 U13265 ( .IN1(n12749), .IN2(n12750), .IN3(n12751), .QN(g30374) );
  NAND2X0 U13266 ( .IN1(n8982), .IN2(g2384), .QN(n12751) );
  NAND3X0 U13267 ( .IN1(n3555), .IN2(n12752), .IN3(n8576), .QN(n12750) );
  XOR2X1 U13268 ( .IN1(n8225), .IN2(n8102), .Q(n12752) );
  NAND2X0 U13269 ( .IN1(n12753), .IN2(g2389), .QN(n12749) );
  NAND2X0 U13270 ( .IN1(n11617), .IN2(n12754), .QN(n12753) );
  NAND2X0 U13271 ( .IN1(n8902), .IN2(n11629), .QN(n12754) );
  NAND2X0 U13272 ( .IN1(n12755), .IN2(n12756), .QN(g30373) );
  NAND2X0 U13273 ( .IN1(n8981), .IN2(g2307), .QN(n12756) );
  NAND2X0 U13274 ( .IN1(n12757), .IN2(n8914), .QN(n12755) );
  NAND2X0 U13275 ( .IN1(n12758), .IN2(n12759), .QN(n12757) );
  NAND2X0 U13276 ( .IN1(n12760), .IN2(g2327), .QN(n12759) );
  NAND2X0 U13277 ( .IN1(n12761), .IN2(n12762), .QN(n12758) );
  NAND2X0 U13278 ( .IN1(n5353), .IN2(g2331), .QN(n12762) );
  INVX0 U13279 ( .INP(n12760), .ZN(n12761) );
  NAND3X0 U13280 ( .IN1(n12763), .IN2(test_so21), .IN3(n5511), .QN(n12760) );
  NAND3X0 U13281 ( .IN1(n12764), .IN2(n12765), .IN3(n12766), .QN(g30372) );
  INVX0 U13282 ( .INP(n12767), .ZN(n12766) );
  NOR2X0 U13283 ( .IN1(n12768), .IN2(n15229), .QN(n12767) );
  INVX0 U13284 ( .INP(n12769), .ZN(n12765) );
  NOR2X0 U13285 ( .IN1(n12770), .IN2(n5778), .QN(n12769) );
  NOR2X0 U13286 ( .IN1(n12771), .IN2(n8932), .QN(n12770) );
  NOR2X0 U13287 ( .IN1(n12772), .IN2(n5458), .QN(n12771) );
  NAND3X0 U13288 ( .IN1(n12773), .IN2(n5458), .IN3(n5778), .QN(n12764) );
  NAND2X0 U13289 ( .IN1(n12774), .IN2(n12775), .QN(g30371) );
  INVX0 U13290 ( .INP(n12776), .ZN(n12775) );
  NOR2X0 U13291 ( .IN1(n12768), .IN2(n5778), .QN(n12776) );
  NAND2X0 U13292 ( .IN1(n12768), .IN2(g2273), .QN(n12774) );
  NAND3X0 U13293 ( .IN1(n12777), .IN2(n12778), .IN3(n12779), .QN(g30370) );
  NAND2X0 U13294 ( .IN1(n8981), .IN2(g2255), .QN(n12779) );
  INVX0 U13295 ( .INP(n12780), .ZN(n12778) );
  NOR2X0 U13296 ( .IN1(n12768), .IN2(n5419), .QN(n12780) );
  NAND2X0 U13297 ( .IN1(n12772), .IN2(n8914), .QN(n12768) );
  NAND2X0 U13298 ( .IN1(n12773), .IN2(n5419), .QN(n12777) );
  NAND3X0 U13299 ( .IN1(n12781), .IN2(n12782), .IN3(n12783), .QN(g30369) );
  NAND2X0 U13300 ( .IN1(n8980), .IN2(g2250), .QN(n12783) );
  NAND3X0 U13301 ( .IN1(n3574), .IN2(n12784), .IN3(n8581), .QN(n12782) );
  XOR2X1 U13302 ( .IN1(n8221), .IN2(n8105), .Q(n12784) );
  NAND2X0 U13303 ( .IN1(n12785), .IN2(g2255), .QN(n12781) );
  NAND2X0 U13304 ( .IN1(n11638), .IN2(n12786), .QN(n12785) );
  NAND2X0 U13305 ( .IN1(n8902), .IN2(n11650), .QN(n12786) );
  NAND2X0 U13306 ( .IN1(n12787), .IN2(n12788), .QN(g30368) );
  NAND2X0 U13307 ( .IN1(n8980), .IN2(g2173), .QN(n12788) );
  NAND2X0 U13308 ( .IN1(n12789), .IN2(n8914), .QN(n12787) );
  NAND2X0 U13309 ( .IN1(n12790), .IN2(n12791), .QN(n12789) );
  NAND2X0 U13310 ( .IN1(n12792), .IN2(g2193), .QN(n12791) );
  NAND2X0 U13311 ( .IN1(n12793), .IN2(n12794), .QN(n12790) );
  NAND2X0 U13312 ( .IN1(n5356), .IN2(g2197), .QN(n12794) );
  INVX0 U13313 ( .INP(n12792), .ZN(n12793) );
  NAND3X0 U13314 ( .IN1(n12795), .IN2(g2208), .IN3(n5512), .QN(n12792) );
  NAND3X0 U13315 ( .IN1(n12796), .IN2(n12797), .IN3(n12798), .QN(g30367) );
  NAND2X0 U13316 ( .IN1(n12799), .IN2(g2126), .QN(n12798) );
  INVX0 U13317 ( .INP(n12800), .ZN(n12797) );
  NOR2X0 U13318 ( .IN1(n12801), .IN2(n5784), .QN(n12800) );
  NOR2X0 U13319 ( .IN1(n12802), .IN2(n8931), .QN(n12801) );
  NOR2X0 U13320 ( .IN1(n12803), .IN2(n5463), .QN(n12802) );
  NAND3X0 U13321 ( .IN1(n12804), .IN2(n5463), .IN3(n5784), .QN(n12796) );
  NAND2X0 U13322 ( .IN1(n12805), .IN2(n12806), .QN(g30366) );
  INVX0 U13323 ( .INP(n12807), .ZN(n12806) );
  NOR2X0 U13324 ( .IN1(n12808), .IN2(n5784), .QN(n12807) );
  NAND2X0 U13325 ( .IN1(n12808), .IN2(g2116), .QN(n12805) );
  NAND3X0 U13326 ( .IN1(n12809), .IN2(n12810), .IN3(n12811), .QN(g30365) );
  NAND2X0 U13327 ( .IN1(n8980), .IN2(g2098), .QN(n12811) );
  NAND2X0 U13328 ( .IN1(n12799), .IN2(g2102), .QN(n12810) );
  INVX0 U13329 ( .INP(n12808), .ZN(n12799) );
  NAND2X0 U13330 ( .IN1(n12803), .IN2(n8914), .QN(n12808) );
  NAND2X0 U13331 ( .IN1(n12804), .IN2(n5666), .QN(n12809) );
  NAND3X0 U13332 ( .IN1(n12812), .IN2(n12813), .IN3(n12814), .QN(g30364) );
  NAND2X0 U13333 ( .IN1(test_so78), .IN2(n9055), .QN(n12814) );
  NAND3X0 U13334 ( .IN1(n8583), .IN2(n3593), .IN3(n12815), .QN(n12813) );
  XOR2X1 U13335 ( .IN1(g2089), .IN2(test_so78), .Q(n12815) );
  NAND2X0 U13336 ( .IN1(n12816), .IN2(g2098), .QN(n12812) );
  NAND2X0 U13337 ( .IN1(n11659), .IN2(n12817), .QN(n12816) );
  NAND2X0 U13338 ( .IN1(n8902), .IN2(n11671), .QN(n12817) );
  NAND2X0 U13339 ( .IN1(n12818), .IN2(n12819), .QN(g30363) );
  NAND2X0 U13340 ( .IN1(n8979), .IN2(g2016), .QN(n12819) );
  NAND2X0 U13341 ( .IN1(n12820), .IN2(n8914), .QN(n12818) );
  NAND2X0 U13342 ( .IN1(n12821), .IN2(n12822), .QN(n12820) );
  NAND2X0 U13343 ( .IN1(test_so59), .IN2(n12823), .QN(n12822) );
  NAND2X0 U13344 ( .IN1(n12824), .IN2(n12825), .QN(n12821) );
  NAND2X0 U13345 ( .IN1(n5355), .IN2(g2040), .QN(n12825) );
  INVX0 U13346 ( .INP(n12823), .ZN(n12824) );
  NAND3X0 U13347 ( .IN1(n12826), .IN2(g2051), .IN3(n5507), .QN(n12823) );
  NAND3X0 U13348 ( .IN1(n12827), .IN2(n12828), .IN3(n12829), .QN(g30362) );
  NAND2X0 U13349 ( .IN1(n12830), .IN2(g1992), .QN(n12829) );
  INVX0 U13350 ( .INP(n12831), .ZN(n12828) );
  NOR2X0 U13351 ( .IN1(n12832), .IN2(n5783), .QN(n12831) );
  NOR2X0 U13352 ( .IN1(n12833), .IN2(n8931), .QN(n12832) );
  NOR2X0 U13353 ( .IN1(n12834), .IN2(n5462), .QN(n12833) );
  NAND3X0 U13354 ( .IN1(n12835), .IN2(n5462), .IN3(n5783), .QN(n12827) );
  NAND2X0 U13355 ( .IN1(n12836), .IN2(n12837), .QN(g30361) );
  INVX0 U13356 ( .INP(n12838), .ZN(n12837) );
  NOR2X0 U13357 ( .IN1(n12839), .IN2(n5783), .QN(n12838) );
  NAND2X0 U13358 ( .IN1(n12839), .IN2(g1982), .QN(n12836) );
  NAND3X0 U13359 ( .IN1(n12840), .IN2(n12841), .IN3(n12842), .QN(g30360) );
  NAND2X0 U13360 ( .IN1(n8979), .IN2(g1964), .QN(n12842) );
  NAND2X0 U13361 ( .IN1(n12830), .IN2(g1968), .QN(n12841) );
  INVX0 U13362 ( .INP(n12839), .ZN(n12830) );
  NAND2X0 U13363 ( .IN1(n12834), .IN2(n8914), .QN(n12839) );
  NAND2X0 U13364 ( .IN1(n12835), .IN2(n5664), .QN(n12840) );
  NAND3X0 U13365 ( .IN1(n12843), .IN2(n12844), .IN3(n12845), .QN(g30359) );
  NAND2X0 U13366 ( .IN1(n8978), .IN2(g1959), .QN(n12845) );
  NAND3X0 U13367 ( .IN1(n3611), .IN2(n12846), .IN3(n8573), .QN(n12844) );
  XOR2X1 U13368 ( .IN1(n8229), .IN2(n8099), .Q(n12846) );
  NAND2X0 U13369 ( .IN1(n12847), .IN2(g1964), .QN(n12843) );
  NAND2X0 U13370 ( .IN1(n11680), .IN2(n12848), .QN(n12847) );
  NAND2X0 U13371 ( .IN1(n8902), .IN2(n11692), .QN(n12848) );
  NAND2X0 U13372 ( .IN1(n12849), .IN2(n12850), .QN(g30358) );
  NAND2X0 U13373 ( .IN1(n8978), .IN2(g1882), .QN(n12850) );
  NAND2X0 U13374 ( .IN1(n12851), .IN2(n8913), .QN(n12849) );
  NAND2X0 U13375 ( .IN1(n12852), .IN2(n12853), .QN(n12851) );
  NAND2X0 U13376 ( .IN1(n12854), .IN2(g1902), .QN(n12853) );
  NAND2X0 U13377 ( .IN1(n12855), .IN2(n12856), .QN(n12852) );
  NAND2X0 U13378 ( .IN1(g1906), .IN2(n8586), .QN(n12856) );
  INVX0 U13379 ( .INP(n12854), .ZN(n12855) );
  NAND3X0 U13380 ( .IN1(n12857), .IN2(g1917), .IN3(n5510), .QN(n12854) );
  NAND3X0 U13381 ( .IN1(n12858), .IN2(n12859), .IN3(n12860), .QN(g30357) );
  INVX0 U13382 ( .INP(n12861), .ZN(n12860) );
  NOR2X0 U13383 ( .IN1(n12862), .IN2(n5892), .QN(n12861) );
  INVX0 U13384 ( .INP(n12863), .ZN(n12859) );
  NOR2X0 U13385 ( .IN1(n12864), .IN2(n5785), .QN(n12863) );
  NOR2X0 U13386 ( .IN1(n12865), .IN2(n8939), .QN(n12864) );
  NOR2X0 U13387 ( .IN1(n12866), .IN2(n5464), .QN(n12865) );
  NAND3X0 U13388 ( .IN1(n12867), .IN2(n5464), .IN3(n5785), .QN(n12858) );
  NAND2X0 U13389 ( .IN1(n12868), .IN2(n12869), .QN(g30356) );
  INVX0 U13390 ( .INP(n12870), .ZN(n12869) );
  NOR2X0 U13391 ( .IN1(n12862), .IN2(n5785), .QN(n12870) );
  NAND2X0 U13392 ( .IN1(n12862), .IN2(g1848), .QN(n12868) );
  NAND3X0 U13393 ( .IN1(n12871), .IN2(n12872), .IN3(n12873), .QN(g30355) );
  NAND2X0 U13394 ( .IN1(n8977), .IN2(g1830), .QN(n12873) );
  INVX0 U13395 ( .INP(n12874), .ZN(n12872) );
  NOR2X0 U13396 ( .IN1(n12862), .IN2(n5665), .QN(n12874) );
  NAND2X0 U13397 ( .IN1(n12866), .IN2(n8913), .QN(n12862) );
  NAND2X0 U13398 ( .IN1(n12867), .IN2(n5665), .QN(n12871) );
  NAND3X0 U13399 ( .IN1(n12875), .IN2(n12876), .IN3(n12877), .QN(g30354) );
  NAND2X0 U13400 ( .IN1(n8977), .IN2(g1825), .QN(n12877) );
  NAND3X0 U13401 ( .IN1(n3628), .IN2(n12878), .IN3(n8579), .QN(n12876) );
  XOR2X1 U13402 ( .IN1(n8223), .IN2(n8100), .Q(n12878) );
  NAND2X0 U13403 ( .IN1(n12879), .IN2(g1830), .QN(n12875) );
  NAND2X0 U13404 ( .IN1(n11701), .IN2(n12880), .QN(n12879) );
  NAND2X0 U13405 ( .IN1(n8902), .IN2(n11713), .QN(n12880) );
  NAND2X0 U13406 ( .IN1(n12881), .IN2(n12882), .QN(g30353) );
  NAND2X0 U13407 ( .IN1(n8977), .IN2(g1748), .QN(n12882) );
  NAND2X0 U13408 ( .IN1(n12883), .IN2(n8913), .QN(n12881) );
  NAND2X0 U13409 ( .IN1(n12884), .IN2(n12885), .QN(n12883) );
  NAND2X0 U13410 ( .IN1(n12886), .IN2(g1768), .QN(n12885) );
  NAND2X0 U13411 ( .IN1(n12887), .IN2(n12888), .QN(n12884) );
  NAND2X0 U13412 ( .IN1(n5352), .IN2(g1772), .QN(n12888) );
  INVX0 U13413 ( .INP(n12886), .ZN(n12887) );
  NAND3X0 U13414 ( .IN1(n12889), .IN2(g1783), .IN3(n5359), .QN(n12886) );
  NAND3X0 U13415 ( .IN1(n12890), .IN2(n12891), .IN3(n12892), .QN(g30352) );
  NAND2X0 U13416 ( .IN1(n12893), .IN2(n9236), .QN(n12892) );
  NAND2X0 U13417 ( .IN1(n12894), .IN2(g1720), .QN(n12891) );
  NAND2X0 U13418 ( .IN1(n12895), .IN2(n8913), .QN(n12894) );
  NAND2X0 U13419 ( .IN1(n12896), .IN2(g1714), .QN(n12895) );
  NAND4X0 U13420 ( .IN1(n5460), .IN2(n8899), .IN3(n12896), .IN4(n5780), .QN(
        n12890) );
  NAND2X0 U13421 ( .IN1(n12897), .IN2(n12898), .QN(g30351) );
  NAND2X0 U13422 ( .IN1(n12893), .IN2(g1720), .QN(n12898) );
  INVX0 U13423 ( .INP(n12899), .ZN(n12897) );
  NOR2X0 U13424 ( .IN1(n12893), .IN2(n5460), .QN(n12899) );
  NAND3X0 U13425 ( .IN1(n12900), .IN2(n12901), .IN3(n12902), .QN(g30350) );
  NAND2X0 U13426 ( .IN1(n12893), .IN2(g1700), .QN(n12902) );
  NOR2X0 U13427 ( .IN1(n12896), .IN2(n8928), .QN(n12893) );
  NAND3X0 U13428 ( .IN1(n12896), .IN2(n5417), .IN3(n8893), .QN(n12901) );
  NAND2X0 U13429 ( .IN1(n8977), .IN2(g1696), .QN(n12900) );
  NAND3X0 U13430 ( .IN1(n12903), .IN2(n12904), .IN3(n12905), .QN(g30349) );
  NAND2X0 U13431 ( .IN1(n8976), .IN2(g1691), .QN(n12905) );
  NAND3X0 U13432 ( .IN1(n3646), .IN2(n12906), .IN3(n8582), .QN(n12904) );
  XOR2X1 U13433 ( .IN1(n8227), .IN2(n8104), .Q(n12906) );
  NAND2X0 U13434 ( .IN1(n12907), .IN2(g1696), .QN(n12903) );
  NAND2X0 U13435 ( .IN1(n11722), .IN2(n12908), .QN(n12907) );
  NAND2X0 U13436 ( .IN1(n8902), .IN2(n11737), .QN(n12908) );
  NAND3X0 U13437 ( .IN1(n12909), .IN2(n12910), .IN3(n12911), .QN(g30348) );
  NAND2X0 U13438 ( .IN1(n8976), .IN2(g1612), .QN(n12911) );
  NAND3X0 U13439 ( .IN1(g25167), .IN2(n11297), .IN3(n3646), .QN(n12910) );
  NAND2X0 U13440 ( .IN1(n5362), .IN2(g1636), .QN(n11297) );
  NAND2X0 U13441 ( .IN1(n12912), .IN2(g1632), .QN(n12909) );
  NAND2X0 U13442 ( .IN1(n11722), .IN2(n12913), .QN(n12912) );
  NAND2X0 U13443 ( .IN1(n10231), .IN2(n8913), .QN(n12913) );
  NAND2X0 U13444 ( .IN1(n12914), .IN2(n12915), .QN(g30347) );
  NAND3X0 U13445 ( .IN1(n12916), .IN2(n12917), .IN3(n12918), .QN(n12915) );
  NAND2X0 U13446 ( .IN1(n12919), .IN2(n12920), .QN(n12916) );
  INVX0 U13447 ( .INP(n12921), .ZN(n12920) );
  NAND2X0 U13448 ( .IN1(n8902), .IN2(g1413), .QN(n12919) );
  NAND2X0 U13449 ( .IN1(n8976), .IN2(g1542), .QN(n12914) );
  NAND2X0 U13450 ( .IN1(n12922), .IN2(n12923), .QN(g30346) );
  NAND2X0 U13451 ( .IN1(n8976), .IN2(g1536), .QN(n12923) );
  NAND3X0 U13452 ( .IN1(n12918), .IN2(n12924), .IN3(n8892), .QN(n12922) );
  XOR2X1 U13453 ( .IN1(n8487), .IN2(n12925), .Q(n12924) );
  NAND2X0 U13454 ( .IN1(n12926), .IN2(n12927), .QN(g30345) );
  NAND2X0 U13455 ( .IN1(n12928), .IN2(n8913), .QN(n12927) );
  NAND2X0 U13456 ( .IN1(n12918), .IN2(n11097), .QN(n12928) );
  INVX0 U13457 ( .INP(n12929), .ZN(n12918) );
  NAND2X0 U13458 ( .IN1(n12930), .IN2(g1514), .QN(n12926) );
  NAND2X0 U13459 ( .IN1(n12931), .IN2(n8913), .QN(n12930) );
  XOR2X1 U13460 ( .IN1(test_so49), .IN2(n5302), .Q(n12931) );
  NOR2X0 U13461 ( .IN1(n8949), .IN2(n12932), .QN(g30344) );
  NOR2X0 U13462 ( .IN1(n12929), .IN2(n12933), .QN(n12932) );
  XOR2X1 U13463 ( .IN1(n5364), .IN2(n5302), .Q(n12933) );
  NAND2X0 U13464 ( .IN1(n12934), .IN2(n12935), .QN(n12929) );
  NAND2X0 U13465 ( .IN1(n4172), .IN2(n12936), .QN(n12935) );
  INVX0 U13466 ( .INP(n12937), .ZN(n4172) );
  NAND4X0 U13467 ( .IN1(n8307), .IN2(n4895), .IN3(n12938), .IN4(g1521), .QN(
        n12937) );
  NAND3X0 U13468 ( .IN1(n12939), .IN2(n12940), .IN3(n12941), .QN(g30343) );
  NAND2X0 U13469 ( .IN1(n4175), .IN2(n11741), .QN(n12941) );
  NAND2X0 U13470 ( .IN1(n8975), .IN2(g1345), .QN(n12940) );
  NAND3X0 U13471 ( .IN1(n11865), .IN2(g1361), .IN3(n8893), .QN(n12939) );
  NAND2X0 U13472 ( .IN1(n12942), .IN2(n12943), .QN(n11865) );
  NAND2X0 U13473 ( .IN1(n8165), .IN2(n11305), .QN(n12943) );
  INVX0 U13474 ( .INP(n12944), .ZN(n11305) );
  NAND3X0 U13475 ( .IN1(n12945), .IN2(n12946), .IN3(n12947), .QN(g30342) );
  NAND2X0 U13476 ( .IN1(n8975), .IN2(g1256), .QN(n12947) );
  NAND3X0 U13477 ( .IN1(n11311), .IN2(n12948), .IN3(g1259), .QN(n12946) );
  INVX0 U13478 ( .INP(n3736), .ZN(n12948) );
  NAND2X0 U13479 ( .IN1(n3736), .IN2(n5553), .QN(n12945) );
  NAND2X0 U13480 ( .IN1(n12949), .IN2(n12950), .QN(g30341) );
  NAND3X0 U13481 ( .IN1(n12951), .IN2(n12952), .IN3(n12953), .QN(n12950) );
  NAND2X0 U13482 ( .IN1(n12954), .IN2(n12955), .QN(n12951) );
  INVX0 U13483 ( .INP(n12956), .ZN(n12955) );
  NAND2X0 U13484 ( .IN1(n8902), .IN2(g1070), .QN(n12954) );
  NAND2X0 U13485 ( .IN1(n8975), .IN2(g1199), .QN(n12949) );
  NAND2X0 U13486 ( .IN1(n12957), .IN2(n12958), .QN(g30340) );
  NAND2X0 U13487 ( .IN1(n8975), .IN2(g1193), .QN(n12958) );
  NAND3X0 U13488 ( .IN1(n12953), .IN2(n12959), .IN3(n8892), .QN(n12957) );
  XOR2X1 U13489 ( .IN1(n12960), .IN2(n8486), .Q(n12959) );
  NAND2X0 U13490 ( .IN1(n12961), .IN2(n12962), .QN(g30339) );
  NAND2X0 U13491 ( .IN1(n12963), .IN2(n8915), .QN(n12962) );
  NAND2X0 U13492 ( .IN1(n12953), .IN2(n11257), .QN(n12963) );
  INVX0 U13493 ( .INP(n12964), .ZN(n12953) );
  NAND2X0 U13494 ( .IN1(n12965), .IN2(g1171), .QN(n12961) );
  NAND2X0 U13495 ( .IN1(n12966), .IN2(n8923), .QN(n12965) );
  XOR2X1 U13496 ( .IN1(g1183), .IN2(n5304), .Q(n12966) );
  NOR2X0 U13497 ( .IN1(n8948), .IN2(n12967), .QN(g30338) );
  NOR2X0 U13498 ( .IN1(n12964), .IN2(n12968), .QN(n12967) );
  XOR2X1 U13499 ( .IN1(n5363), .IN2(n5304), .Q(n12968) );
  NAND2X0 U13500 ( .IN1(n12969), .IN2(n12970), .QN(n12964) );
  NAND2X0 U13501 ( .IN1(n4190), .IN2(n12971), .QN(n12970) );
  INVX0 U13502 ( .INP(n12972), .ZN(n4190) );
  NAND4X0 U13503 ( .IN1(n5642), .IN2(n4920), .IN3(n12973), .IN4(g1178), .QN(
        n12972) );
  NAND3X0 U13504 ( .IN1(n12974), .IN2(n12975), .IN3(n12976), .QN(g30337) );
  NAND2X0 U13505 ( .IN1(n4193), .IN2(n11754), .QN(n12976) );
  NAND2X0 U13506 ( .IN1(n8974), .IN2(g1002), .QN(n12975) );
  NAND3X0 U13507 ( .IN1(n11874), .IN2(g1018), .IN3(n8889), .QN(n12974) );
  NAND2X0 U13508 ( .IN1(n12977), .IN2(n12978), .QN(n11874) );
  NAND2X0 U13509 ( .IN1(n8166), .IN2(n11319), .QN(n12978) );
  NAND3X0 U13510 ( .IN1(n12979), .IN2(n12980), .IN3(n12981), .QN(g30336) );
  NAND2X0 U13511 ( .IN1(n8974), .IN2(g911), .QN(n12981) );
  NAND3X0 U13512 ( .IN1(n11325), .IN2(n12982), .IN3(g914), .QN(n12980) );
  INVX0 U13513 ( .INP(n3741), .ZN(n12982) );
  NAND2X0 U13514 ( .IN1(n3741), .IN2(n5560), .QN(n12979) );
  NAND3X0 U13515 ( .IN1(n12983), .IN2(n12984), .IN3(n12985), .QN(g30335) );
  NAND2X0 U13516 ( .IN1(test_so60), .IN2(n8947), .QN(n12985) );
  NAND3X0 U13517 ( .IN1(n2404), .IN2(n12986), .IN3(g744), .QN(n12984) );
  NAND2X0 U13518 ( .IN1(n55), .IN2(n5470), .QN(n12983) );
  INVX0 U13519 ( .INP(n12986), .ZN(n55) );
  NAND3X0 U13520 ( .IN1(test_so60), .IN2(n4198), .IN3(n12987), .QN(n12986) );
  NAND2X0 U13521 ( .IN1(n8514), .IN2(g11678), .QN(n4198) );
  NAND3X0 U13522 ( .IN1(n12988), .IN2(n12989), .IN3(n12990), .QN(g30334) );
  NAND2X0 U13523 ( .IN1(n8974), .IN2(g586), .QN(n12990) );
  NAND3X0 U13524 ( .IN1(n2421), .IN2(n12991), .IN3(g577), .QN(n12989) );
  INVX0 U13525 ( .INP(n3745), .ZN(n12991) );
  NAND2X0 U13526 ( .IN1(n3745), .IN2(n5294), .QN(n12988) );
  NAND2X0 U13527 ( .IN1(n12992), .IN2(n12993), .QN(g30333) );
  NAND2X0 U13528 ( .IN1(n10217), .IN2(n12994), .QN(n12993) );
  XOR2X1 U13529 ( .IN1(test_so73), .IN2(n11897), .Q(n12994) );
  NOR2X0 U13530 ( .IN1(n11898), .IN2(n8931), .QN(n10217) );
  NAND3X0 U13531 ( .IN1(n12995), .IN2(g691), .IN3(n12996), .QN(n11898) );
  NAND2X0 U13532 ( .IN1(n11897), .IN2(n12997), .QN(n12996) );
  NAND2X0 U13533 ( .IN1(n12998), .IN2(n8593), .QN(n12997) );
  INVX0 U13534 ( .INP(n12999), .ZN(n11897) );
  NAND2X0 U13535 ( .IN1(n8974), .IN2(g142), .QN(n12992) );
  NAND3X0 U13536 ( .IN1(n13000), .IN2(n13001), .IN3(n13002), .QN(g29309) );
  NAND2X0 U13537 ( .IN1(n3765), .IN2(n13003), .QN(n13002) );
  NAND2X0 U13538 ( .IN1(g6541), .IN2(n13004), .QN(n13003) );
  INVX0 U13539 ( .INP(n10839), .ZN(n13004) );
  NAND3X0 U13540 ( .IN1(n13005), .IN2(g6541), .IN3(n11922), .QN(n13000) );
  NAND3X0 U13541 ( .IN1(n13006), .IN2(n13007), .IN3(n13008), .QN(g29308) );
  NAND2X0 U13542 ( .IN1(n8973), .IN2(g6523), .QN(n13008) );
  NAND2X0 U13543 ( .IN1(n13009), .IN2(g6527), .QN(n13007) );
  NAND2X0 U13544 ( .IN1(n5659), .IN2(n13010), .QN(n13006) );
  NAND3X0 U13545 ( .IN1(n13011), .IN2(n13012), .IN3(n13013), .QN(g29307) );
  NAND2X0 U13546 ( .IN1(n13009), .IN2(g6523), .QN(n13013) );
  NAND2X0 U13547 ( .IN1(n13014), .IN2(g6519), .QN(n13012) );
  NAND2X0 U13548 ( .IN1(n13015), .IN2(n8923), .QN(n13014) );
  NAND2X0 U13549 ( .IN1(n13016), .IN2(g6513), .QN(n13015) );
  NAND3X0 U13550 ( .IN1(n5426), .IN2(n13010), .IN3(n5806), .QN(n13011) );
  NAND2X0 U13551 ( .IN1(n13017), .IN2(n13018), .QN(g29306) );
  NAND2X0 U13552 ( .IN1(n13009), .IN2(g6519), .QN(n13018) );
  NAND2X0 U13553 ( .IN1(n13019), .IN2(g6513), .QN(n13017) );
  INVX0 U13554 ( .INP(n13009), .ZN(n13019) );
  NAND3X0 U13555 ( .IN1(n13020), .IN2(n13021), .IN3(n13022), .QN(g29305) );
  NAND2X0 U13556 ( .IN1(n13009), .IN2(g6509), .QN(n13022) );
  NOR2X0 U13557 ( .IN1(n13016), .IN2(n8943), .QN(n13009) );
  NAND2X0 U13558 ( .IN1(n13023), .IN2(g6500), .QN(n13021) );
  NAND2X0 U13559 ( .IN1(n13024), .IN2(n8923), .QN(n13023) );
  NAND2X0 U13560 ( .IN1(n8138), .IN2(n13016), .QN(n13024) );
  NAND3X0 U13561 ( .IN1(n13010), .IN2(g6505), .IN3(n5748), .QN(n13020) );
  INVX0 U13562 ( .INP(n13025), .ZN(n13010) );
  NAND2X0 U13563 ( .IN1(n13016), .IN2(n8923), .QN(n13025) );
  NOR2X0 U13564 ( .IN1(n13026), .IN2(n8575), .QN(n13016) );
  NAND2X0 U13565 ( .IN1(n13027), .IN2(n13028), .QN(g29304) );
  NAND2X0 U13566 ( .IN1(n8973), .IN2(g6505), .QN(n13028) );
  NAND2X0 U13567 ( .IN1(n13029), .IN2(n8923), .QN(n13027) );
  NAND2X0 U13568 ( .IN1(n13030), .IN2(n13031), .QN(n13029) );
  NAND2X0 U13569 ( .IN1(n8575), .IN2(g6500), .QN(n13031) );
  NAND2X0 U13570 ( .IN1(n13032), .IN2(n10850), .QN(n13030) );
  XNOR2X1 U13571 ( .IN1(n13033), .IN2(n13034), .Q(n13032) );
  NAND2X0 U13572 ( .IN1(g6500), .IN2(n13026), .QN(n13033) );
  NAND3X0 U13573 ( .IN1(g6727), .IN2(g17722), .IN3(n9216), .QN(n13026) );
  NAND3X0 U13574 ( .IN1(n13035), .IN2(n13001), .IN3(n13036), .QN(g29303) );
  NAND2X0 U13575 ( .IN1(n3765), .IN2(n13037), .QN(n13036) );
  NAND2X0 U13576 ( .IN1(g6195), .IN2(n10828), .QN(n13037) );
  NAND3X0 U13577 ( .IN1(n13005), .IN2(g6195), .IN3(n12008), .QN(n13035) );
  NAND3X0 U13578 ( .IN1(n13038), .IN2(n13039), .IN3(n13040), .QN(g29302) );
  NAND2X0 U13579 ( .IN1(n8972), .IN2(g6177), .QN(n13040) );
  NAND2X0 U13580 ( .IN1(n13041), .IN2(g6181), .QN(n13039) );
  NAND2X0 U13581 ( .IN1(n5667), .IN2(n13042), .QN(n13038) );
  NAND3X0 U13582 ( .IN1(n13043), .IN2(n13044), .IN3(n13045), .QN(g29301) );
  NAND2X0 U13583 ( .IN1(n13041), .IN2(g6177), .QN(n13045) );
  NAND2X0 U13584 ( .IN1(n13046), .IN2(g6173), .QN(n13044) );
  NAND2X0 U13585 ( .IN1(n13047), .IN2(n8923), .QN(n13046) );
  NAND2X0 U13586 ( .IN1(n13048), .IN2(g6167), .QN(n13047) );
  NAND3X0 U13587 ( .IN1(n5430), .IN2(n13042), .IN3(n5810), .QN(n13043) );
  NAND2X0 U13588 ( .IN1(n13049), .IN2(n13050), .QN(g29300) );
  NAND2X0 U13589 ( .IN1(n13041), .IN2(g6173), .QN(n13050) );
  NAND2X0 U13590 ( .IN1(n13051), .IN2(g6167), .QN(n13049) );
  INVX0 U13591 ( .INP(n13041), .ZN(n13051) );
  NAND3X0 U13592 ( .IN1(n13052), .IN2(n13053), .IN3(n13054), .QN(g29299) );
  NAND2X0 U13593 ( .IN1(n13041), .IN2(g6163), .QN(n13054) );
  NOR2X0 U13594 ( .IN1(n13048), .IN2(n8929), .QN(n13041) );
  NAND2X0 U13595 ( .IN1(n13055), .IN2(g6154), .QN(n13053) );
  NAND2X0 U13596 ( .IN1(n13056), .IN2(n8923), .QN(n13055) );
  NAND2X0 U13597 ( .IN1(n8137), .IN2(n13048), .QN(n13056) );
  NAND3X0 U13598 ( .IN1(n13042), .IN2(g6159), .IN3(n5747), .QN(n13052) );
  INVX0 U13599 ( .INP(n13057), .ZN(n13042) );
  NAND2X0 U13600 ( .IN1(n13048), .IN2(n8923), .QN(n13057) );
  NOR2X0 U13601 ( .IN1(n13058), .IN2(n10868), .QN(n13048) );
  NAND2X0 U13602 ( .IN1(n13059), .IN2(n13060), .QN(g29298) );
  NAND2X0 U13603 ( .IN1(n8972), .IN2(g6159), .QN(n13060) );
  NAND2X0 U13604 ( .IN1(n13061), .IN2(n8923), .QN(n13059) );
  NAND2X0 U13605 ( .IN1(n13062), .IN2(n13063), .QN(n13061) );
  NAND2X0 U13606 ( .IN1(n10868), .IN2(g6154), .QN(n13063) );
  NAND2X0 U13607 ( .IN1(n13064), .IN2(n10862), .QN(n13062) );
  XNOR2X1 U13608 ( .IN1(n13065), .IN2(n13066), .Q(n13064) );
  NAND2X0 U13609 ( .IN1(g6154), .IN2(n13058), .QN(n13065) );
  NAND3X0 U13610 ( .IN1(n10063), .IN2(g17685), .IN3(test_so69), .QN(n13058) );
  NAND3X0 U13611 ( .IN1(n13067), .IN2(n13001), .IN3(n13068), .QN(g29297) );
  NAND2X0 U13612 ( .IN1(n3765), .IN2(n13069), .QN(n13068) );
  NAND2X0 U13613 ( .IN1(g5849), .IN2(n10827), .QN(n13069) );
  NAND3X0 U13614 ( .IN1(n13005), .IN2(g5849), .IN3(n12095), .QN(n13067) );
  NAND3X0 U13615 ( .IN1(n13070), .IN2(n13071), .IN3(n13072), .QN(g29296) );
  NAND2X0 U13616 ( .IN1(n8972), .IN2(g5831), .QN(n13072) );
  NAND2X0 U13617 ( .IN1(n13073), .IN2(g5835), .QN(n13071) );
  NAND2X0 U13618 ( .IN1(n5663), .IN2(n13074), .QN(n13070) );
  NAND3X0 U13619 ( .IN1(n13075), .IN2(n13076), .IN3(n13077), .QN(g29295) );
  NAND2X0 U13620 ( .IN1(n13073), .IN2(g5831), .QN(n13077) );
  NAND2X0 U13621 ( .IN1(n13078), .IN2(g5827), .QN(n13076) );
  NAND2X0 U13622 ( .IN1(n13079), .IN2(n8923), .QN(n13078) );
  NAND2X0 U13623 ( .IN1(n13080), .IN2(g5821), .QN(n13079) );
  NAND3X0 U13624 ( .IN1(n5429), .IN2(n13074), .IN3(n5809), .QN(n13075) );
  NAND2X0 U13625 ( .IN1(n13081), .IN2(n13082), .QN(g29294) );
  NAND2X0 U13626 ( .IN1(n13073), .IN2(g5827), .QN(n13082) );
  NAND2X0 U13627 ( .IN1(n13083), .IN2(g5821), .QN(n13081) );
  INVX0 U13628 ( .INP(n13073), .ZN(n13083) );
  NAND3X0 U13629 ( .IN1(n13084), .IN2(n13085), .IN3(n13086), .QN(g29293) );
  NAND2X0 U13630 ( .IN1(n13073), .IN2(g5817), .QN(n13086) );
  NOR2X0 U13631 ( .IN1(n13080), .IN2(n8930), .QN(n13073) );
  NAND2X0 U13632 ( .IN1(n13087), .IN2(g5808), .QN(n13085) );
  NAND2X0 U13633 ( .IN1(n13088), .IN2(n8923), .QN(n13087) );
  NAND2X0 U13634 ( .IN1(n8139), .IN2(n13080), .QN(n13088) );
  NAND3X0 U13635 ( .IN1(n13074), .IN2(g5813), .IN3(n5749), .QN(n13084) );
  INVX0 U13636 ( .INP(n13089), .ZN(n13074) );
  NAND2X0 U13637 ( .IN1(n13080), .IN2(n8923), .QN(n13089) );
  NOR2X0 U13638 ( .IN1(n13090), .IN2(n10884), .QN(n13080) );
  NAND2X0 U13639 ( .IN1(n13091), .IN2(n13092), .QN(g29292) );
  NAND2X0 U13640 ( .IN1(n8972), .IN2(g5813), .QN(n13092) );
  NAND2X0 U13641 ( .IN1(n13093), .IN2(n8923), .QN(n13091) );
  NAND2X0 U13642 ( .IN1(n13094), .IN2(n13095), .QN(n13093) );
  NAND2X0 U13643 ( .IN1(n10884), .IN2(g5808), .QN(n13095) );
  NAND2X0 U13644 ( .IN1(n13096), .IN2(n10878), .QN(n13094) );
  XNOR2X1 U13645 ( .IN1(n13097), .IN2(n13098), .Q(n13096) );
  NAND2X0 U13646 ( .IN1(g5808), .IN2(n13090), .QN(n13097) );
  NAND3X0 U13647 ( .IN1(g6035), .IN2(g17646), .IN3(n10068), .QN(n13090) );
  NAND3X0 U13648 ( .IN1(n13099), .IN2(n13001), .IN3(n13100), .QN(g29291) );
  NAND2X0 U13649 ( .IN1(n3765), .IN2(n13101), .QN(n13100) );
  NAND2X0 U13650 ( .IN1(g5503), .IN2(n13102), .QN(n13101) );
  INVX0 U13651 ( .INP(n10823), .ZN(n13102) );
  NAND3X0 U13652 ( .IN1(n13005), .IN2(g5503), .IN3(n12182), .QN(n13099) );
  NAND3X0 U13653 ( .IN1(n13103), .IN2(n13104), .IN3(n13105), .QN(g29290) );
  NAND2X0 U13654 ( .IN1(n8971), .IN2(g5485), .QN(n13105) );
  NAND2X0 U13655 ( .IN1(n13106), .IN2(g5489), .QN(n13104) );
  NAND2X0 U13656 ( .IN1(n5660), .IN2(n13107), .QN(n13103) );
  NAND3X0 U13657 ( .IN1(n13108), .IN2(n13109), .IN3(n13110), .QN(g29289) );
  NAND2X0 U13658 ( .IN1(n13106), .IN2(g5485), .QN(n13110) );
  NAND2X0 U13659 ( .IN1(n13111), .IN2(g5481), .QN(n13109) );
  NAND2X0 U13660 ( .IN1(n13112), .IN2(n8923), .QN(n13111) );
  NAND2X0 U13661 ( .IN1(n13113), .IN2(g5475), .QN(n13112) );
  NAND3X0 U13662 ( .IN1(n5425), .IN2(n13107), .IN3(n5805), .QN(n13108) );
  NAND2X0 U13663 ( .IN1(n13114), .IN2(n13115), .QN(g29288) );
  NAND2X0 U13664 ( .IN1(n13106), .IN2(g5481), .QN(n13115) );
  NAND2X0 U13665 ( .IN1(n13116), .IN2(g5475), .QN(n13114) );
  INVX0 U13666 ( .INP(n13106), .ZN(n13116) );
  NAND3X0 U13667 ( .IN1(n13117), .IN2(n13118), .IN3(n13119), .QN(g29287) );
  NAND2X0 U13668 ( .IN1(n13106), .IN2(g5471), .QN(n13119) );
  NOR2X0 U13669 ( .IN1(n13113), .IN2(n8932), .QN(n13106) );
  NAND2X0 U13670 ( .IN1(n13120), .IN2(g5462), .QN(n13118) );
  NAND2X0 U13671 ( .IN1(n13121), .IN2(n8922), .QN(n13120) );
  NAND2X0 U13672 ( .IN1(n8124), .IN2(n13113), .QN(n13121) );
  NAND3X0 U13673 ( .IN1(n13107), .IN2(g5467), .IN3(n5744), .QN(n13117) );
  INVX0 U13674 ( .INP(n13122), .ZN(n13107) );
  NAND2X0 U13675 ( .IN1(n13113), .IN2(n8922), .QN(n13122) );
  NOR2X0 U13676 ( .IN1(n13123), .IN2(n10900), .QN(n13113) );
  NAND2X0 U13677 ( .IN1(n13124), .IN2(n13125), .QN(g29286) );
  NAND2X0 U13678 ( .IN1(n8971), .IN2(g5467), .QN(n13125) );
  NAND2X0 U13679 ( .IN1(n13126), .IN2(n8922), .QN(n13124) );
  NAND2X0 U13680 ( .IN1(n13127), .IN2(n13128), .QN(n13126) );
  NAND2X0 U13681 ( .IN1(n10900), .IN2(g5462), .QN(n13128) );
  NAND2X0 U13682 ( .IN1(n13129), .IN2(n10894), .QN(n13127) );
  XNOR2X1 U13683 ( .IN1(n13130), .IN2(n13131), .Q(n13129) );
  NAND2X0 U13684 ( .IN1(g5462), .IN2(n13123), .QN(n13130) );
  NAND3X0 U13685 ( .IN1(g5689), .IN2(g17604), .IN3(n10076), .QN(n13123) );
  NAND3X0 U13686 ( .IN1(n13132), .IN2(n13001), .IN3(n13133), .QN(g29285) );
  NAND2X0 U13687 ( .IN1(n3765), .IN2(n13134), .QN(n13133) );
  NAND2X0 U13688 ( .IN1(g5156), .IN2(n13135), .QN(n13134) );
  INVX0 U13689 ( .INP(g32975), .ZN(n13135) );
  NAND3X0 U13690 ( .IN1(n13005), .IN2(g5156), .IN3(n12268), .QN(n13132) );
  NAND3X0 U13691 ( .IN1(n13136), .IN2(n13137), .IN3(n13138), .QN(g29284) );
  NAND2X0 U13692 ( .IN1(n8970), .IN2(g5138), .QN(n13138) );
  NAND2X0 U13693 ( .IN1(n13139), .IN2(g5142), .QN(n13137) );
  NAND2X0 U13694 ( .IN1(n5658), .IN2(n13140), .QN(n13136) );
  NAND3X0 U13695 ( .IN1(n13141), .IN2(n13142), .IN3(n13143), .QN(g29283) );
  NAND2X0 U13696 ( .IN1(n13139), .IN2(g5138), .QN(n13143) );
  NAND2X0 U13697 ( .IN1(n13144), .IN2(g5134), .QN(n13142) );
  NAND2X0 U13698 ( .IN1(n13145), .IN2(n8922), .QN(n13144) );
  NAND2X0 U13699 ( .IN1(test_so96), .IN2(n13146), .QN(n13145) );
  NAND3X0 U13700 ( .IN1(n13140), .IN2(n8601), .IN3(n5807), .QN(n13141) );
  NAND2X0 U13701 ( .IN1(n13147), .IN2(n13148), .QN(g29282) );
  NAND2X0 U13702 ( .IN1(n13139), .IN2(g5134), .QN(n13148) );
  NAND2X0 U13703 ( .IN1(test_so96), .IN2(n13149), .QN(n13147) );
  INVX0 U13704 ( .INP(n13139), .ZN(n13149) );
  NAND3X0 U13705 ( .IN1(n13150), .IN2(n13151), .IN3(n13152), .QN(g29281) );
  NAND2X0 U13706 ( .IN1(n13139), .IN2(g5124), .QN(n13152) );
  NOR2X0 U13707 ( .IN1(n13146), .IN2(n8942), .QN(n13139) );
  NAND2X0 U13708 ( .IN1(n13153), .IN2(g5115), .QN(n13151) );
  NAND2X0 U13709 ( .IN1(n13154), .IN2(n8922), .QN(n13153) );
  NAND2X0 U13710 ( .IN1(n8123), .IN2(n13146), .QN(n13154) );
  NAND3X0 U13711 ( .IN1(n13140), .IN2(g5120), .IN3(n5743), .QN(n13150) );
  INVX0 U13712 ( .INP(n13155), .ZN(n13140) );
  NAND2X0 U13713 ( .IN1(n13146), .IN2(n8922), .QN(n13155) );
  NOR2X0 U13714 ( .IN1(n13156), .IN2(n8570), .QN(n13146) );
  NAND2X0 U13715 ( .IN1(n13157), .IN2(n13158), .QN(g29280) );
  NAND2X0 U13716 ( .IN1(n8970), .IN2(g5120), .QN(n13158) );
  NAND2X0 U13717 ( .IN1(n13159), .IN2(n8922), .QN(n13157) );
  NAND2X0 U13718 ( .IN1(n13160), .IN2(n13161), .QN(n13159) );
  NAND2X0 U13719 ( .IN1(n8570), .IN2(g5115), .QN(n13161) );
  NAND2X0 U13720 ( .IN1(n13162), .IN2(g33959), .QN(n13160) );
  XNOR2X1 U13721 ( .IN1(n13163), .IN2(n13164), .Q(n13162) );
  NAND2X0 U13722 ( .IN1(g5115), .IN2(n13156), .QN(n13163) );
  NAND3X0 U13723 ( .IN1(g31860), .IN2(g17577), .IN3(test_so10), .QN(n13156) );
  NAND2X0 U13724 ( .IN1(n13165), .IN2(n13166), .QN(g29275) );
  NAND2X0 U13725 ( .IN1(n13167), .IN2(n12367), .QN(n13166) );
  XOR2X1 U13726 ( .IN1(n11856), .IN2(g4087), .Q(n13167) );
  NOR2X0 U13727 ( .IN1(n8598), .IN2(n13168), .QN(n11856) );
  NAND2X0 U13728 ( .IN1(test_so11), .IN2(n8946), .QN(n13165) );
  NAND3X0 U13729 ( .IN1(n13169), .IN2(n13001), .IN3(n13170), .QN(g29274) );
  NAND2X0 U13730 ( .IN1(n3765), .IN2(n13171), .QN(n13170) );
  NAND2X0 U13731 ( .IN1(g3849), .IN2(n10838), .QN(n13171) );
  NAND3X0 U13732 ( .IN1(n13005), .IN2(g3849), .IN3(n12371), .QN(n13169) );
  NAND3X0 U13733 ( .IN1(n13172), .IN2(n13173), .IN3(n13174), .QN(g29273) );
  NAND2X0 U13734 ( .IN1(n8970), .IN2(g3831), .QN(n13174) );
  NAND2X0 U13735 ( .IN1(n13175), .IN2(g3835), .QN(n13173) );
  NAND2X0 U13736 ( .IN1(n5662), .IN2(n13176), .QN(n13172) );
  NAND3X0 U13737 ( .IN1(n13177), .IN2(n13178), .IN3(n13179), .QN(g29272) );
  NAND2X0 U13738 ( .IN1(n13175), .IN2(g3831), .QN(n13179) );
  NAND2X0 U13739 ( .IN1(n13180), .IN2(g3827), .QN(n13178) );
  NAND2X0 U13740 ( .IN1(n13181), .IN2(n8922), .QN(n13180) );
  NAND2X0 U13741 ( .IN1(n13182), .IN2(g3821), .QN(n13181) );
  NAND3X0 U13742 ( .IN1(n5428), .IN2(n13176), .IN3(n5808), .QN(n13177) );
  NAND2X0 U13743 ( .IN1(n13183), .IN2(n13184), .QN(g29271) );
  NAND2X0 U13744 ( .IN1(n13175), .IN2(g3827), .QN(n13184) );
  NAND2X0 U13745 ( .IN1(n13185), .IN2(g3821), .QN(n13183) );
  INVX0 U13746 ( .INP(n13175), .ZN(n13185) );
  NOR2X0 U13747 ( .IN1(n13182), .IN2(n8930), .QN(n13175) );
  NAND3X0 U13748 ( .IN1(n13186), .IN2(n13187), .IN3(n13188), .QN(g29270) );
  NAND2X0 U13749 ( .IN1(n11902), .IN2(n13189), .QN(n13188) );
  NOR2X0 U13750 ( .IN1(n8949), .IN2(n8072), .QN(n11902) );
  NAND2X0 U13751 ( .IN1(n13190), .IN2(g3808), .QN(n13187) );
  NAND2X0 U13752 ( .IN1(n13191), .IN2(n8922), .QN(n13190) );
  NAND2X0 U13753 ( .IN1(n8125), .IN2(n13182), .QN(n13191) );
  NAND3X0 U13754 ( .IN1(n13176), .IN2(g3813), .IN3(n5745), .QN(n13186) );
  NOR2X0 U13755 ( .IN1(n13189), .IN2(n8929), .QN(n13176) );
  INVX0 U13756 ( .INP(n13182), .ZN(n13189) );
  NOR2X0 U13757 ( .IN1(n13192), .IN2(n10939), .QN(n13182) );
  NAND2X0 U13758 ( .IN1(n13193), .IN2(n13194), .QN(g29269) );
  NAND2X0 U13759 ( .IN1(n8969), .IN2(g3813), .QN(n13194) );
  NAND2X0 U13760 ( .IN1(n13195), .IN2(n8922), .QN(n13193) );
  NAND2X0 U13761 ( .IN1(n13196), .IN2(n13197), .QN(n13195) );
  NAND2X0 U13762 ( .IN1(n10939), .IN2(g3808), .QN(n13197) );
  NAND2X0 U13763 ( .IN1(n13198), .IN2(n10933), .QN(n13196) );
  XNOR2X1 U13764 ( .IN1(n13199), .IN2(n13200), .Q(n13198) );
  NAND2X0 U13765 ( .IN1(g3808), .IN2(n13192), .QN(n13199) );
  NAND3X0 U13766 ( .IN1(g4040), .IN2(g16693), .IN3(n10064), .QN(n13192) );
  NAND3X0 U13767 ( .IN1(n13201), .IN2(n13001), .IN3(n13202), .QN(g29268) );
  NAND2X0 U13768 ( .IN1(n3765), .IN2(n13203), .QN(n13202) );
  NAND2X0 U13769 ( .IN1(g3498), .IN2(n10837), .QN(n13203) );
  NAND3X0 U13770 ( .IN1(n13005), .IN2(g3498), .IN3(n12458), .QN(n13201) );
  NAND3X0 U13771 ( .IN1(n13204), .IN2(n13205), .IN3(n13206), .QN(g29267) );
  NAND2X0 U13772 ( .IN1(n8969), .IN2(g3480), .QN(n13206) );
  NAND2X0 U13773 ( .IN1(n13207), .IN2(g3484), .QN(n13205) );
  NAND2X0 U13774 ( .IN1(n5668), .IN2(n13208), .QN(n13204) );
  NAND3X0 U13775 ( .IN1(n13209), .IN2(n13210), .IN3(n13211), .QN(g29266) );
  NAND2X0 U13776 ( .IN1(n13207), .IN2(g3480), .QN(n13211) );
  NAND2X0 U13777 ( .IN1(n13212), .IN2(g3476), .QN(n13210) );
  NAND2X0 U13778 ( .IN1(n13213), .IN2(n8922), .QN(n13212) );
  NAND2X0 U13779 ( .IN1(n13214), .IN2(g3470), .QN(n13213) );
  NAND3X0 U13780 ( .IN1(n5424), .IN2(n13208), .IN3(n5786), .QN(n13209) );
  NAND2X0 U13781 ( .IN1(n13215), .IN2(n13216), .QN(g29265) );
  NAND2X0 U13782 ( .IN1(n13207), .IN2(g3476), .QN(n13216) );
  NAND2X0 U13783 ( .IN1(n13217), .IN2(g3470), .QN(n13215) );
  INVX0 U13784 ( .INP(n13207), .ZN(n13217) );
  NAND3X0 U13785 ( .IN1(n13218), .IN2(n13219), .IN3(n13220), .QN(g29264) );
  NAND2X0 U13786 ( .IN1(n13207), .IN2(g3466), .QN(n13220) );
  NOR2X0 U13787 ( .IN1(n13214), .IN2(n8933), .QN(n13207) );
  NAND2X0 U13788 ( .IN1(test_so4), .IN2(n13221), .QN(n13219) );
  NAND2X0 U13789 ( .IN1(n13222), .IN2(n8922), .QN(n13221) );
  NAND2X0 U13790 ( .IN1(n8126), .IN2(n13214), .QN(n13222) );
  NAND3X0 U13791 ( .IN1(n13208), .IN2(g3462), .IN3(n8611), .QN(n13218) );
  INVX0 U13792 ( .INP(n13223), .ZN(n13208) );
  NAND2X0 U13793 ( .IN1(n13214), .IN2(n8922), .QN(n13223) );
  NOR2X0 U13794 ( .IN1(n13224), .IN2(n10955), .QN(n13214) );
  NAND2X0 U13795 ( .IN1(n13225), .IN2(n13226), .QN(g29263) );
  NAND2X0 U13796 ( .IN1(n8969), .IN2(g3462), .QN(n13226) );
  NAND2X0 U13797 ( .IN1(n13227), .IN2(n8922), .QN(n13225) );
  NAND2X0 U13798 ( .IN1(n13228), .IN2(n13229), .QN(n13227) );
  NAND2X0 U13799 ( .IN1(test_so4), .IN2(n10955), .QN(n13229) );
  NAND2X0 U13800 ( .IN1(n13230), .IN2(n10949), .QN(n13228) );
  XNOR2X1 U13801 ( .IN1(n13231), .IN2(n13232), .Q(n13230) );
  NAND2X0 U13802 ( .IN1(test_so4), .IN2(n13224), .QN(n13231) );
  NAND3X0 U13803 ( .IN1(g3689), .IN2(g16656), .IN3(n10069), .QN(n13224) );
  NAND3X0 U13804 ( .IN1(n13233), .IN2(n13001), .IN3(n13234), .QN(g29262) );
  NAND2X0 U13805 ( .IN1(n3765), .IN2(n13235), .QN(n13234) );
  NAND2X0 U13806 ( .IN1(g3147), .IN2(n13236), .QN(n13235) );
  INVX0 U13807 ( .INP(n10834), .ZN(n13236) );
  NAND2X0 U13808 ( .IN1(n3765), .IN2(n13005), .QN(n13001) );
  NAND3X0 U13809 ( .IN1(n13005), .IN2(g3147), .IN3(n12545), .QN(n13233) );
  INVX0 U13810 ( .INP(n4210), .ZN(n13005) );
  NAND2X0 U13811 ( .IN1(n8511), .IN2(g4180), .QN(n4210) );
  NAND3X0 U13812 ( .IN1(n13237), .IN2(n13238), .IN3(n13239), .QN(g29261) );
  NAND2X0 U13813 ( .IN1(n8969), .IN2(g3129), .QN(n13239) );
  NAND2X0 U13814 ( .IN1(n13240), .IN2(g3133), .QN(n13238) );
  NAND2X0 U13815 ( .IN1(n5661), .IN2(n13241), .QN(n13237) );
  NAND3X0 U13816 ( .IN1(n13242), .IN2(n13243), .IN3(n13244), .QN(g29260) );
  NAND2X0 U13817 ( .IN1(n13240), .IN2(g3129), .QN(n13244) );
  NAND2X0 U13818 ( .IN1(n13245), .IN2(g3125), .QN(n13243) );
  NAND2X0 U13819 ( .IN1(n13246), .IN2(n8922), .QN(n13245) );
  NAND2X0 U13820 ( .IN1(n13247), .IN2(g3119), .QN(n13246) );
  NAND3X0 U13821 ( .IN1(n5423), .IN2(n13241), .IN3(n5781), .QN(n13242) );
  NAND2X0 U13822 ( .IN1(n13248), .IN2(n13249), .QN(g29259) );
  NAND2X0 U13823 ( .IN1(n13240), .IN2(g3125), .QN(n13249) );
  NAND2X0 U13824 ( .IN1(n13250), .IN2(g3119), .QN(n13248) );
  INVX0 U13825 ( .INP(n13240), .ZN(n13250) );
  NAND3X0 U13826 ( .IN1(n13251), .IN2(n13252), .IN3(n13253), .QN(g29258) );
  NAND2X0 U13827 ( .IN1(n13240), .IN2(g3115), .QN(n13253) );
  NOR2X0 U13828 ( .IN1(n13247), .IN2(n8934), .QN(n13240) );
  NAND2X0 U13829 ( .IN1(n13254), .IN2(g3106), .QN(n13252) );
  NAND2X0 U13830 ( .IN1(n13255), .IN2(n8922), .QN(n13254) );
  NAND2X0 U13831 ( .IN1(n8122), .IN2(n13247), .QN(n13255) );
  NAND3X0 U13832 ( .IN1(n13241), .IN2(g3111), .IN3(n5742), .QN(n13251) );
  INVX0 U13833 ( .INP(n13256), .ZN(n13241) );
  NAND2X0 U13834 ( .IN1(n13247), .IN2(n8922), .QN(n13256) );
  NOR2X0 U13835 ( .IN1(n13257), .IN2(n10966), .QN(n13247) );
  NAND2X0 U13836 ( .IN1(n13258), .IN2(n13259), .QN(g29257) );
  NAND2X0 U13837 ( .IN1(n8968), .IN2(g3111), .QN(n13259) );
  NAND2X0 U13838 ( .IN1(n13260), .IN2(n8922), .QN(n13258) );
  NAND2X0 U13839 ( .IN1(n13261), .IN2(n13262), .QN(n13260) );
  NAND2X0 U13840 ( .IN1(n10966), .IN2(g3106), .QN(n13262) );
  NAND2X0 U13841 ( .IN1(n13263), .IN2(n10969), .QN(n13261) );
  XNOR2X1 U13842 ( .IN1(n13264), .IN2(n13265), .Q(n13263) );
  NAND2X0 U13843 ( .IN1(g3106), .IN2(n13257), .QN(n13264) );
  NAND3X0 U13844 ( .IN1(g3338), .IN2(g16624), .IN3(n10077), .QN(n13257) );
  NAND4X0 U13845 ( .IN1(n13266), .IN2(n9200), .IN3(n13267), .IN4(n13268), .QN(
        g29256) );
  NAND3X0 U13846 ( .IN1(n13269), .IN2(g2735), .IN3(n8889), .QN(n13268) );
  INVX0 U13847 ( .INP(n12670), .ZN(n13269) );
  NAND2X0 U13848 ( .IN1(n8968), .IN2(g2729), .QN(n13267) );
  NAND2X0 U13849 ( .IN1(n5600), .IN2(n12670), .QN(n13266) );
  NOR2X0 U13850 ( .IN1(n13270), .IN2(n8186), .QN(n12670) );
  NAND2X0 U13851 ( .IN1(n13271), .IN2(n13272), .QN(g29255) );
  NAND2X0 U13852 ( .IN1(n13273), .IN2(g2652), .QN(n13272) );
  NAND2X0 U13853 ( .IN1(n11575), .IN2(n13274), .QN(n13273) );
  NAND2X0 U13854 ( .IN1(n4379), .IN2(n8922), .QN(n13274) );
  NAND2X0 U13855 ( .IN1(n13275), .IN2(g2638), .QN(n13271) );
  INVX0 U13856 ( .INP(n13276), .ZN(n13275) );
  NOR2X0 U13857 ( .IN1(n13277), .IN2(n8935), .QN(n13276) );
  NOR2X0 U13858 ( .IN1(n11572), .IN2(n9228), .QN(n13277) );
  NOR2X0 U13859 ( .IN1(n8231), .IN2(n8574), .QN(n9228) );
  NAND4X0 U13860 ( .IN1(n13278), .IN2(n13279), .IN3(n13280), .IN4(n13281), 
        .QN(g29254) );
  NAND2X0 U13861 ( .IN1(n12680), .IN2(g2567), .QN(n13281) );
  NOR2X0 U13862 ( .IN1(n12679), .IN2(n8935), .QN(n12680) );
  NAND3X0 U13863 ( .IN1(g2587), .IN2(g2619), .IN3(n12702), .QN(n12679) );
  INVX0 U13864 ( .INP(n11572), .ZN(n12702) );
  NAND2X0 U13865 ( .IN1(n3517), .IN2(n13282), .QN(n13280) );
  NAND3X0 U13866 ( .IN1(n13283), .IN2(n13284), .IN3(n13285), .QN(n13282) );
  NAND2X0 U13867 ( .IN1(n8574), .IN2(g2563), .QN(n13285) );
  INVX0 U13868 ( .INP(n11587), .ZN(n8574) );
  NAND2X0 U13869 ( .IN1(n5372), .IN2(g2610), .QN(n11587) );
  NAND2X0 U13870 ( .IN1(n5508), .IN2(n13286), .QN(n13284) );
  NAND2X0 U13871 ( .IN1(n13287), .IN2(n13288), .QN(n13286) );
  NAND2X0 U13872 ( .IN1(test_so66), .IN2(n5372), .QN(n13288) );
  NAND2X0 U13873 ( .IN1(g2583), .IN2(g2610), .QN(n13287) );
  NAND2X0 U13874 ( .IN1(n8482), .IN2(n13289), .QN(n13283) );
  NAND2X0 U13875 ( .IN1(n13290), .IN2(n13291), .QN(n13289) );
  NAND2X0 U13876 ( .IN1(test_so61), .IN2(g2587), .QN(n13291) );
  NAND2X0 U13877 ( .IN1(g2619), .IN2(g2571), .QN(n13290) );
  NOR2X0 U13878 ( .IN1(n11572), .IN2(n8935), .QN(n3517) );
  NAND2X0 U13879 ( .IN1(n11581), .IN2(g2638), .QN(n13279) );
  INVX0 U13880 ( .INP(n11575), .ZN(n11581) );
  NAND2X0 U13881 ( .IN1(n11572), .IN2(n8921), .QN(n11575) );
  NAND3X0 U13882 ( .IN1(n13292), .IN2(n13293), .IN3(n12644), .QN(n11572) );
  NAND2X0 U13883 ( .IN1(n12664), .IN2(g2819), .QN(n13292) );
  NAND2X0 U13884 ( .IN1(n8968), .IN2(g2619), .QN(n13278) );
  NAND2X0 U13885 ( .IN1(n13294), .IN2(n13295), .QN(g29253) );
  NAND2X0 U13886 ( .IN1(n13296), .IN2(g2518), .QN(n13295) );
  NAND2X0 U13887 ( .IN1(n11596), .IN2(n13297), .QN(n13296) );
  NAND2X0 U13888 ( .IN1(n4391), .IN2(n8921), .QN(n13297) );
  NAND2X0 U13889 ( .IN1(n13298), .IN2(g2504), .QN(n13294) );
  INVX0 U13890 ( .INP(n13299), .ZN(n13298) );
  NOR2X0 U13891 ( .IN1(n13300), .IN2(n8935), .QN(n13299) );
  NOR2X0 U13892 ( .IN1(n11593), .IN2(n9227), .QN(n13300) );
  NOR2X0 U13893 ( .IN1(n8230), .IN2(n8580), .QN(n9227) );
  NAND4X0 U13894 ( .IN1(n13301), .IN2(n13302), .IN3(n13303), .IN4(n13304), 
        .QN(g29252) );
  NAND2X0 U13895 ( .IN1(n12711), .IN2(g2433), .QN(n13304) );
  NOR2X0 U13896 ( .IN1(n12710), .IN2(n8935), .QN(n12711) );
  NAND3X0 U13897 ( .IN1(g2453), .IN2(g2485), .IN3(n12733), .QN(n12710) );
  INVX0 U13898 ( .INP(n11593), .ZN(n12733) );
  NAND2X0 U13899 ( .IN1(n3536), .IN2(n13305), .QN(n13303) );
  NAND3X0 U13900 ( .IN1(n13306), .IN2(n13307), .IN3(n13308), .QN(n13305) );
  NAND2X0 U13901 ( .IN1(n8580), .IN2(g2429), .QN(n13308) );
  INVX0 U13902 ( .INP(n11608), .ZN(n8580) );
  NAND2X0 U13903 ( .IN1(n5373), .IN2(g2476), .QN(n11608) );
  NAND2X0 U13904 ( .IN1(n5509), .IN2(n13309), .QN(n13307) );
  NAND2X0 U13905 ( .IN1(n13310), .IN2(n13311), .QN(n13309) );
  NAND2X0 U13906 ( .IN1(n5373), .IN2(g2441), .QN(n13311) );
  NAND2X0 U13907 ( .IN1(g2449), .IN2(g2476), .QN(n13310) );
  NAND2X0 U13908 ( .IN1(n8481), .IN2(n13312), .QN(n13306) );
  NAND2X0 U13909 ( .IN1(n13313), .IN2(n13314), .QN(n13312) );
  NAND2X0 U13910 ( .IN1(g2453), .IN2(n9274), .QN(n13314) );
  NAND2X0 U13911 ( .IN1(g2485), .IN2(g2437), .QN(n13313) );
  NOR2X0 U13912 ( .IN1(n11593), .IN2(n8936), .QN(n3536) );
  NAND2X0 U13913 ( .IN1(n11602), .IN2(g2504), .QN(n13302) );
  INVX0 U13914 ( .INP(n11596), .ZN(n11602) );
  NAND2X0 U13915 ( .IN1(n11593), .IN2(n8921), .QN(n11596) );
  NAND3X0 U13916 ( .IN1(n13315), .IN2(n13293), .IN3(n12645), .QN(n11593) );
  NAND2X0 U13917 ( .IN1(n12664), .IN2(g2815), .QN(n13315) );
  NAND2X0 U13918 ( .IN1(n8968), .IN2(g2485), .QN(n13301) );
  NAND2X0 U13919 ( .IN1(n13316), .IN2(n13317), .QN(g29251) );
  NAND2X0 U13920 ( .IN1(n13318), .IN2(g2384), .QN(n13317) );
  NAND2X0 U13921 ( .IN1(n11617), .IN2(n13319), .QN(n13318) );
  NAND2X0 U13922 ( .IN1(n4402), .IN2(n8921), .QN(n13319) );
  NAND2X0 U13923 ( .IN1(n13320), .IN2(g2370), .QN(n13316) );
  INVX0 U13924 ( .INP(n13321), .ZN(n13320) );
  NOR2X0 U13925 ( .IN1(n13322), .IN2(n8936), .QN(n13321) );
  NOR2X0 U13926 ( .IN1(n11614), .IN2(n9226), .QN(n13322) );
  NOR2X0 U13927 ( .IN1(n8225), .IN2(n8576), .QN(n9226) );
  NAND4X0 U13928 ( .IN1(n13323), .IN2(n13324), .IN3(n13325), .IN4(n13326), 
        .QN(g29250) );
  NAND2X0 U13929 ( .IN1(n12742), .IN2(g2299), .QN(n13326) );
  NOR2X0 U13930 ( .IN1(n12741), .IN2(n8936), .QN(n12742) );
  NAND3X0 U13931 ( .IN1(g2319), .IN2(g2351), .IN3(n12763), .QN(n12741) );
  INVX0 U13932 ( .INP(n11614), .ZN(n12763) );
  NAND2X0 U13933 ( .IN1(n3555), .IN2(n13327), .QN(n13325) );
  NAND3X0 U13934 ( .IN1(n13328), .IN2(n13329), .IN3(n13330), .QN(n13327) );
  NAND2X0 U13935 ( .IN1(n8576), .IN2(g2295), .QN(n13330) );
  INVX0 U13936 ( .INP(n11629), .ZN(n8576) );
  NAND2X0 U13937 ( .IN1(test_so21), .IN2(n5375), .QN(n11629) );
  NAND2X0 U13938 ( .IN1(n5511), .IN2(n13331), .QN(n13329) );
  NAND2X0 U13939 ( .IN1(n13332), .IN2(n13333), .QN(n13331) );
  NAND2X0 U13940 ( .IN1(n5375), .IN2(g2307), .QN(n13333) );
  NAND2X0 U13941 ( .IN1(test_so21), .IN2(g2315), .QN(n13332) );
  NAND2X0 U13942 ( .IN1(n13334), .IN2(n8591), .QN(n13328) );
  NAND2X0 U13943 ( .IN1(n13335), .IN2(n13336), .QN(n13334) );
  NAND2X0 U13944 ( .IN1(g2319), .IN2(n9314), .QN(n13336) );
  NAND2X0 U13945 ( .IN1(g2351), .IN2(g2303), .QN(n13335) );
  NOR2X0 U13946 ( .IN1(n11614), .IN2(n8936), .QN(n3555) );
  NAND2X0 U13947 ( .IN1(n11623), .IN2(g2370), .QN(n13324) );
  INVX0 U13948 ( .INP(n11617), .ZN(n11623) );
  NAND2X0 U13949 ( .IN1(n11614), .IN2(n8921), .QN(n11617) );
  NAND3X0 U13950 ( .IN1(n13293), .IN2(n13337), .IN3(n13338), .QN(n11614) );
  NAND2X0 U13951 ( .IN1(n12664), .IN2(g2807), .QN(n13338) );
  NAND2X0 U13952 ( .IN1(n8968), .IN2(g2351), .QN(n13323) );
  NAND2X0 U13953 ( .IN1(n13339), .IN2(n13340), .QN(g29249) );
  NAND2X0 U13954 ( .IN1(n13341), .IN2(g2250), .QN(n13340) );
  NAND2X0 U13955 ( .IN1(n11638), .IN2(n13342), .QN(n13341) );
  NAND2X0 U13956 ( .IN1(n4414), .IN2(n8921), .QN(n13342) );
  NAND2X0 U13957 ( .IN1(n13343), .IN2(g2236), .QN(n13339) );
  INVX0 U13958 ( .INP(n13344), .ZN(n13343) );
  NOR2X0 U13959 ( .IN1(n13345), .IN2(n8937), .QN(n13344) );
  NOR2X0 U13960 ( .IN1(n11635), .IN2(n9225), .QN(n13345) );
  NOR2X0 U13961 ( .IN1(n8221), .IN2(n8581), .QN(n9225) );
  NAND4X0 U13962 ( .IN1(n13346), .IN2(n13347), .IN3(n13348), .IN4(n13349), 
        .QN(g29248) );
  NAND2X0 U13963 ( .IN1(n12773), .IN2(g2165), .QN(n13349) );
  NOR2X0 U13964 ( .IN1(n12772), .IN2(n8937), .QN(n12773) );
  NAND3X0 U13965 ( .IN1(g2185), .IN2(g2217), .IN3(n12795), .QN(n12772) );
  INVX0 U13966 ( .INP(n11635), .ZN(n12795) );
  NAND2X0 U13967 ( .IN1(n3574), .IN2(n13350), .QN(n13348) );
  NAND3X0 U13968 ( .IN1(n13351), .IN2(n13352), .IN3(n13353), .QN(n13350) );
  NAND2X0 U13969 ( .IN1(n8581), .IN2(g2161), .QN(n13353) );
  INVX0 U13970 ( .INP(n11650), .ZN(n8581) );
  NAND2X0 U13971 ( .IN1(n5376), .IN2(g2208), .QN(n11650) );
  NAND2X0 U13972 ( .IN1(n5512), .IN2(n13354), .QN(n13352) );
  NAND2X0 U13973 ( .IN1(n13355), .IN2(n13356), .QN(n13354) );
  NAND2X0 U13974 ( .IN1(n5376), .IN2(g2173), .QN(n13356) );
  NAND2X0 U13975 ( .IN1(g2181), .IN2(g2208), .QN(n13355) );
  NAND2X0 U13976 ( .IN1(n8479), .IN2(n13357), .QN(n13351) );
  NAND2X0 U13977 ( .IN1(n13358), .IN2(n13359), .QN(n13357) );
  NAND2X0 U13978 ( .IN1(g2185), .IN2(n9352), .QN(n13359) );
  NAND2X0 U13979 ( .IN1(g2217), .IN2(g2169), .QN(n13358) );
  NOR2X0 U13980 ( .IN1(n11635), .IN2(n8938), .QN(n3574) );
  NAND2X0 U13981 ( .IN1(n11644), .IN2(g2236), .QN(n13347) );
  INVX0 U13982 ( .INP(n11638), .ZN(n11644) );
  NAND2X0 U13983 ( .IN1(n11635), .IN2(n8921), .QN(n11638) );
  NAND3X0 U13984 ( .IN1(n13360), .IN2(n13293), .IN3(n13361), .QN(n11635) );
  NAND2X0 U13985 ( .IN1(n12664), .IN2(g2803), .QN(n13360) );
  NAND2X0 U13986 ( .IN1(n8968), .IN2(g2217), .QN(n13346) );
  NAND2X0 U13987 ( .IN1(n13362), .IN2(n13363), .QN(g29247) );
  NAND2X0 U13988 ( .IN1(n13364), .IN2(g2079), .QN(n13363) );
  NAND2X0 U13989 ( .IN1(n13365), .IN2(n8921), .QN(n13364) );
  NAND2X0 U13990 ( .IN1(n12826), .IN2(n9346), .QN(n13365) );
  NAND2X0 U13991 ( .IN1(test_so78), .IN2(n11671), .QN(n9346) );
  NAND2X0 U13992 ( .IN1(test_so78), .IN2(n13366), .QN(n13362) );
  NAND2X0 U13993 ( .IN1(n11659), .IN2(n13367), .QN(n13366) );
  NAND2X0 U13994 ( .IN1(n4425), .IN2(n8921), .QN(n13367) );
  NAND4X0 U13995 ( .IN1(n13368), .IN2(n13369), .IN3(n13370), .IN4(n13371), 
        .QN(g29246) );
  NAND2X0 U13996 ( .IN1(n12804), .IN2(g2008), .QN(n13371) );
  NOR2X0 U13997 ( .IN1(n12803), .IN2(n8938), .QN(n12804) );
  NAND3X0 U13998 ( .IN1(g2028), .IN2(g2060), .IN3(n12826), .QN(n12803) );
  INVX0 U13999 ( .INP(n11656), .ZN(n12826) );
  NAND2X0 U14000 ( .IN1(n3593), .IN2(n13372), .QN(n13370) );
  NAND3X0 U14001 ( .IN1(n13373), .IN2(n13374), .IN3(n13375), .QN(n13372) );
  NAND2X0 U14002 ( .IN1(n8583), .IN2(g2004), .QN(n13375) );
  INVX0 U14003 ( .INP(n11671), .ZN(n8583) );
  NAND2X0 U14004 ( .IN1(n5371), .IN2(g2051), .QN(n11671) );
  NAND2X0 U14005 ( .IN1(n5507), .IN2(n13376), .QN(n13374) );
  NAND2X0 U14006 ( .IN1(n13377), .IN2(n13378), .QN(n13376) );
  NAND2X0 U14007 ( .IN1(n5371), .IN2(g2016), .QN(n13378) );
  NAND2X0 U14008 ( .IN1(g2024), .IN2(g2051), .QN(n13377) );
  NAND2X0 U14009 ( .IN1(n8483), .IN2(n13379), .QN(n13373) );
  NAND2X0 U14010 ( .IN1(n13380), .IN2(n13381), .QN(n13379) );
  NAND2X0 U14011 ( .IN1(g2028), .IN2(n9312), .QN(n13381) );
  NAND2X0 U14012 ( .IN1(g2060), .IN2(g2012), .QN(n13380) );
  NOR2X0 U14013 ( .IN1(n11656), .IN2(n8938), .QN(n3593) );
  NAND2X0 U14014 ( .IN1(n11665), .IN2(g2079), .QN(n13369) );
  INVX0 U14015 ( .INP(n11659), .ZN(n11665) );
  NAND2X0 U14016 ( .IN1(n11656), .IN2(n8921), .QN(n11659) );
  NAND3X0 U14017 ( .IN1(n13382), .IN2(n13293), .IN3(n12644), .QN(n11656) );
  NAND2X0 U14018 ( .IN1(n12664), .IN2(g2787), .QN(n13382) );
  NAND2X0 U14019 ( .IN1(n8967), .IN2(g2060), .QN(n13368) );
  NAND2X0 U14020 ( .IN1(n13383), .IN2(n13384), .QN(g29245) );
  NAND2X0 U14021 ( .IN1(n13385), .IN2(g1959), .QN(n13384) );
  NAND2X0 U14022 ( .IN1(n11680), .IN2(n13386), .QN(n13385) );
  NAND2X0 U14023 ( .IN1(n4436), .IN2(n8921), .QN(n13386) );
  NAND2X0 U14024 ( .IN1(test_so53), .IN2(n13387), .QN(n13383) );
  INVX0 U14025 ( .INP(n13388), .ZN(n13387) );
  NOR2X0 U14026 ( .IN1(n13389), .IN2(n8939), .QN(n13388) );
  NOR2X0 U14027 ( .IN1(n11677), .IN2(n9224), .QN(n13389) );
  NOR2X0 U14028 ( .IN1(n8229), .IN2(n8573), .QN(n9224) );
  NAND4X0 U14029 ( .IN1(n13390), .IN2(n13391), .IN3(n13392), .IN4(n13393), 
        .QN(g29244) );
  NAND2X0 U14030 ( .IN1(n12835), .IN2(g1874), .QN(n13393) );
  NOR2X0 U14031 ( .IN1(n12834), .IN2(n8939), .QN(n12835) );
  NAND3X0 U14032 ( .IN1(g1894), .IN2(g1926), .IN3(n12857), .QN(n12834) );
  INVX0 U14033 ( .INP(n11677), .ZN(n12857) );
  NAND2X0 U14034 ( .IN1(n3611), .IN2(n13394), .QN(n13392) );
  NAND3X0 U14035 ( .IN1(n13395), .IN2(n13396), .IN3(n13397), .QN(n13394) );
  NAND2X0 U14036 ( .IN1(n8573), .IN2(g1870), .QN(n13397) );
  INVX0 U14037 ( .INP(n11692), .ZN(n8573) );
  NAND2X0 U14038 ( .IN1(n5374), .IN2(g1917), .QN(n11692) );
  NAND2X0 U14039 ( .IN1(n5510), .IN2(n13398), .QN(n13396) );
  NAND2X0 U14040 ( .IN1(n13399), .IN2(n13400), .QN(n13398) );
  NAND2X0 U14041 ( .IN1(n5374), .IN2(g1882), .QN(n13400) );
  NAND2X0 U14042 ( .IN1(g1890), .IN2(g1917), .QN(n13399) );
  NAND2X0 U14043 ( .IN1(n8480), .IN2(n13401), .QN(n13395) );
  NAND2X0 U14044 ( .IN1(n13402), .IN2(n13403), .QN(n13401) );
  NAND2X0 U14045 ( .IN1(g1894), .IN2(n9280), .QN(n13403) );
  NAND2X0 U14046 ( .IN1(g1926), .IN2(g1878), .QN(n13402) );
  NOR2X0 U14047 ( .IN1(n11677), .IN2(n8939), .QN(n3611) );
  NAND2X0 U14048 ( .IN1(n11686), .IN2(test_so53), .QN(n13391) );
  INVX0 U14049 ( .INP(n11680), .ZN(n11686) );
  NAND2X0 U14050 ( .IN1(n11677), .IN2(n8921), .QN(n11680) );
  NAND3X0 U14051 ( .IN1(n13404), .IN2(n13293), .IN3(n12645), .QN(n11677) );
  NAND2X0 U14052 ( .IN1(n12664), .IN2(g2783), .QN(n13404) );
  NAND2X0 U14053 ( .IN1(n8967), .IN2(g1926), .QN(n13390) );
  NAND2X0 U14054 ( .IN1(n13405), .IN2(n13406), .QN(g29243) );
  NAND2X0 U14055 ( .IN1(n13407), .IN2(g1825), .QN(n13406) );
  NAND2X0 U14056 ( .IN1(n11701), .IN2(n13408), .QN(n13407) );
  NAND2X0 U14057 ( .IN1(n4447), .IN2(n8921), .QN(n13408) );
  NAND2X0 U14058 ( .IN1(n13409), .IN2(g1811), .QN(n13405) );
  INVX0 U14059 ( .INP(n13410), .ZN(n13409) );
  NOR2X0 U14060 ( .IN1(n13411), .IN2(n8940), .QN(n13410) );
  NOR2X0 U14061 ( .IN1(n11698), .IN2(n9223), .QN(n13411) );
  NOR2X0 U14062 ( .IN1(n8223), .IN2(n8579), .QN(n9223) );
  NAND4X0 U14063 ( .IN1(n13412), .IN2(n13413), .IN3(n13414), .IN4(n13415), 
        .QN(g29242) );
  NAND2X0 U14064 ( .IN1(n12867), .IN2(g1740), .QN(n13415) );
  NOR2X0 U14065 ( .IN1(n12866), .IN2(n8940), .QN(n12867) );
  NAND3X0 U14066 ( .IN1(g1792), .IN2(g1760), .IN3(n12889), .QN(n12866) );
  INVX0 U14067 ( .INP(n11698), .ZN(n12889) );
  NAND2X0 U14068 ( .IN1(n3628), .IN2(n13416), .QN(n13414) );
  NAND3X0 U14069 ( .IN1(n13417), .IN2(n13418), .IN3(n13419), .QN(n13416) );
  NAND2X0 U14070 ( .IN1(n8579), .IN2(g1736), .QN(n13419) );
  INVX0 U14071 ( .INP(n11713), .ZN(n8579) );
  NAND2X0 U14072 ( .IN1(n5602), .IN2(g1783), .QN(n11713) );
  NAND2X0 U14073 ( .IN1(n5359), .IN2(n13420), .QN(n13418) );
  NAND2X0 U14074 ( .IN1(n13421), .IN2(n13422), .QN(n13420) );
  NAND2X0 U14075 ( .IN1(g1783), .IN2(g1756), .QN(n13422) );
  NAND2X0 U14076 ( .IN1(n5602), .IN2(g1748), .QN(n13421) );
  NAND2X0 U14077 ( .IN1(n5596), .IN2(n13423), .QN(n13417) );
  NAND2X0 U14078 ( .IN1(n13424), .IN2(n13425), .QN(n13423) );
  NAND2X0 U14079 ( .IN1(g1792), .IN2(g1744), .QN(n13425) );
  NAND2X0 U14080 ( .IN1(g1760), .IN2(g1752), .QN(n13424) );
  NOR2X0 U14081 ( .IN1(n11698), .IN2(n8941), .QN(n3628) );
  NAND2X0 U14082 ( .IN1(n11707), .IN2(g1811), .QN(n13413) );
  INVX0 U14083 ( .INP(n11701), .ZN(n11707) );
  NAND2X0 U14084 ( .IN1(n11698), .IN2(n8921), .QN(n11701) );
  NAND3X0 U14085 ( .IN1(n13293), .IN2(n13337), .IN3(n13426), .QN(n11698) );
  NAND2X0 U14086 ( .IN1(n12664), .IN2(g2775), .QN(n13426) );
  INVX0 U14087 ( .INP(n1249), .ZN(n13337) );
  NAND2X0 U14088 ( .IN1(n5465), .IN2(g2715), .QN(n1249) );
  NAND2X0 U14089 ( .IN1(n8968), .IN2(g1792), .QN(n13412) );
  NAND2X0 U14090 ( .IN1(n13427), .IN2(n13428), .QN(g29241) );
  NAND2X0 U14091 ( .IN1(n13429), .IN2(g1691), .QN(n13428) );
  NAND2X0 U14092 ( .IN1(n11722), .IN2(n13430), .QN(n13429) );
  NAND2X0 U14093 ( .IN1(n4458), .IN2(n8921), .QN(n13430) );
  NAND2X0 U14094 ( .IN1(n13431), .IN2(g1677), .QN(n13427) );
  INVX0 U14095 ( .INP(n13432), .ZN(n13431) );
  NOR2X0 U14096 ( .IN1(n13433), .IN2(n8941), .QN(n13432) );
  NOR2X0 U14097 ( .IN1(n11719), .IN2(n9222), .QN(n13433) );
  NOR2X0 U14098 ( .IN1(n8227), .IN2(n8582), .QN(n9222) );
  NAND4X0 U14099 ( .IN1(n13434), .IN2(n13435), .IN3(n13436), .IN4(n13437), 
        .QN(g29240) );
  NAND2X0 U14100 ( .IN1(n3646), .IN2(n13438), .QN(n13437) );
  NAND4X0 U14101 ( .IN1(n13439), .IN2(n13440), .IN3(n13441), .IN4(n13442), 
        .QN(n13438) );
  NAND3X0 U14102 ( .IN1(n5370), .IN2(g1612), .IN3(n5525), .QN(n13442) );
  NAND2X0 U14103 ( .IN1(n13443), .IN2(n8596), .QN(n13441) );
  NAND2X0 U14104 ( .IN1(n13444), .IN2(n13445), .QN(n13443) );
  NAND2X0 U14105 ( .IN1(g1624), .IN2(n9303), .QN(n13445) );
  NAND2X0 U14106 ( .IN1(g1657), .IN2(g1608), .QN(n13444) );
  NAND2X0 U14107 ( .IN1(g25167), .IN2(g1620), .QN(n13440) );
  NAND2X0 U14108 ( .IN1(n8582), .IN2(g1600), .QN(n13439) );
  INVX0 U14109 ( .INP(n11737), .ZN(n8582) );
  NAND2X0 U14110 ( .IN1(test_so94), .IN2(n5370), .QN(n11737) );
  NOR2X0 U14111 ( .IN1(n11719), .IN2(n8942), .QN(n3646) );
  NAND2X0 U14112 ( .IN1(n12896), .IN2(g1604), .QN(n13436) );
  NOR3X0 U14113 ( .IN1(n5370), .IN2(n5525), .IN3(n11719), .QN(n12896) );
  NAND2X0 U14114 ( .IN1(n11731), .IN2(g1677), .QN(n13435) );
  INVX0 U14115 ( .INP(n11722), .ZN(n11731) );
  NAND2X0 U14116 ( .IN1(n11719), .IN2(n8921), .QN(n11722) );
  NAND3X0 U14117 ( .IN1(n13446), .IN2(n13293), .IN3(n13361), .QN(n11719) );
  INVX0 U14118 ( .INP(n12643), .ZN(n13361) );
  NAND2X0 U14119 ( .IN1(n5465), .IN2(n5299), .QN(n12643) );
  NAND2X0 U14120 ( .IN1(n12664), .IN2(n13447), .QN(n13293) );
  INVX0 U14121 ( .INP(n4388), .ZN(n13447) );
  NAND2X0 U14122 ( .IN1(n12664), .IN2(g2771), .QN(n13446) );
  INVX0 U14123 ( .INP(n10030), .ZN(n12664) );
  NAND2X0 U14124 ( .IN1(n8186), .IN2(n5301), .QN(n10030) );
  NAND2X0 U14125 ( .IN1(n8967), .IN2(g1657), .QN(n13434) );
  NAND3X0 U14126 ( .IN1(n13448), .IN2(n13449), .IN3(n13450), .QN(g29239) );
  NAND3X0 U14127 ( .IN1(n13451), .IN2(n12936), .IN3(n13452), .QN(n13450) );
  NAND2X0 U14128 ( .IN1(n8966), .IN2(g1478), .QN(n13449) );
  NAND3X0 U14129 ( .IN1(n13453), .IN2(g1454), .IN3(n8889), .QN(n13448) );
  NAND2X0 U14130 ( .IN1(n13454), .IN2(n13455), .QN(n13453) );
  INVX0 U14131 ( .INP(n13451), .ZN(n13455) );
  XNOR2X1 U14132 ( .IN1(g1448), .IN2(n13456), .Q(n13451) );
  NAND3X0 U14133 ( .IN1(n13457), .IN2(n13458), .IN3(n13459), .QN(g29238) );
  NAND2X0 U14134 ( .IN1(n13460), .IN2(g1484), .QN(n13459) );
  NAND2X0 U14135 ( .IN1(n8967), .IN2(g1472), .QN(n13458) );
  NAND3X0 U14136 ( .IN1(n13461), .IN2(n13462), .IN3(n8889), .QN(n13457) );
  NAND2X0 U14137 ( .IN1(n5865), .IN2(n13463), .QN(n13462) );
  NAND3X0 U14138 ( .IN1(n8440), .IN2(n5850), .IN3(n13464), .QN(n13463) );
  XOR2X1 U14139 ( .IN1(g1300), .IN2(n13465), .Q(n13461) );
  INVX0 U14140 ( .INP(n13456), .ZN(n13465) );
  NAND3X0 U14141 ( .IN1(n13466), .IN2(n13467), .IN3(n13468), .QN(g29237) );
  NAND3X0 U14142 ( .IN1(n13452), .IN2(n13469), .IN3(n13470), .QN(n13468) );
  NAND2X0 U14143 ( .IN1(n8966), .IN2(g1448), .QN(n13467) );
  NAND3X0 U14144 ( .IN1(n13471), .IN2(g1467), .IN3(n8888), .QN(n13466) );
  NAND3X0 U14145 ( .IN1(n13472), .IN2(g13272), .IN3(n13469), .QN(n13471) );
  INVX0 U14146 ( .INP(n13470), .ZN(n13472) );
  XNOR2X1 U14147 ( .IN1(g1472), .IN2(n13456), .Q(n13470) );
  NAND3X0 U14148 ( .IN1(n13473), .IN2(n13474), .IN3(n13475), .QN(g29236) );
  NAND4X0 U14149 ( .IN1(n13476), .IN2(n13452), .IN3(g1514), .IN4(n8608), .QN(
        n13475) );
  NOR4X0 U14150 ( .IN1(g1442), .IN2(g1489), .IN3(n8927), .IN4(n8521), .QN(
        n13452) );
  NAND2X0 U14151 ( .IN1(n8967), .IN2(g1442), .QN(n13474) );
  NAND3X0 U14152 ( .IN1(n13477), .IN2(g1437), .IN3(n8888), .QN(n13473) );
  NAND2X0 U14153 ( .IN1(n13478), .IN2(n13479), .QN(n13477) );
  INVX0 U14154 ( .INP(n13476), .ZN(n13479) );
  XNOR2X1 U14155 ( .IN1(g1478), .IN2(n13456), .Q(n13476) );
  NAND2X0 U14156 ( .IN1(n9698), .IN2(DFF_1092_n1), .QN(n13456) );
  INVX0 U14157 ( .INP(n9768), .ZN(n9698) );
  NAND3X0 U14158 ( .IN1(n13480), .IN2(n13481), .IN3(n13482), .QN(g29235) );
  NAND2X0 U14159 ( .IN1(n8966), .IN2(g1252), .QN(n13482) );
  NAND3X0 U14160 ( .IN1(n11311), .IN2(n13483), .IN3(g1256), .QN(n13481) );
  INVX0 U14161 ( .INP(n4178), .ZN(n13483) );
  NAND2X0 U14162 ( .IN1(n4178), .IN2(n5558), .QN(n13480) );
  NAND3X0 U14163 ( .IN1(n13484), .IN2(n13485), .IN3(n13486), .QN(g29234) );
  NAND3X0 U14164 ( .IN1(n13487), .IN2(n12971), .IN3(n13488), .QN(n13486) );
  NAND2X0 U14165 ( .IN1(n8966), .IN2(g1135), .QN(n13485) );
  NAND3X0 U14166 ( .IN1(test_so90), .IN2(n13489), .IN3(n8888), .QN(n13484) );
  NAND2X0 U14167 ( .IN1(n13490), .IN2(n13491), .QN(n13489) );
  INVX0 U14168 ( .INP(n13487), .ZN(n13491) );
  XOR2X1 U14169 ( .IN1(n13492), .IN2(n5478), .Q(n13487) );
  NAND3X0 U14170 ( .IN1(n13493), .IN2(n13494), .IN3(n13495), .QN(g29233) );
  NAND2X0 U14171 ( .IN1(n13496), .IN2(g1141), .QN(n13495) );
  NAND2X0 U14172 ( .IN1(n8967), .IN2(g1129), .QN(n13494) );
  NAND3X0 U14173 ( .IN1(n13497), .IN2(n13498), .IN3(n8888), .QN(n13493) );
  NAND2X0 U14174 ( .IN1(n5691), .IN2(n13499), .QN(n13498) );
  NAND3X0 U14175 ( .IN1(n5851), .IN2(n8588), .IN3(n13500), .QN(n13499) );
  XOR2X1 U14176 ( .IN1(n13492), .IN2(n5341), .Q(n13497) );
  NAND3X0 U14177 ( .IN1(n13501), .IN2(n13502), .IN3(n13503), .QN(g29232) );
  NAND3X0 U14178 ( .IN1(n13488), .IN2(n11219), .IN3(n13504), .QN(n13503) );
  NAND2X0 U14179 ( .IN1(n8966), .IN2(g1105), .QN(n13502) );
  NAND3X0 U14180 ( .IN1(n13505), .IN2(g1124), .IN3(n8888), .QN(n13501) );
  NAND3X0 U14181 ( .IN1(n13506), .IN2(g13259), .IN3(n11219), .QN(n13505) );
  INVX0 U14182 ( .INP(n13504), .ZN(n13506) );
  XOR2X1 U14183 ( .IN1(n13492), .IN2(n5329), .Q(n13504) );
  NAND3X0 U14184 ( .IN1(n13507), .IN2(n13508), .IN3(n13509), .QN(g29231) );
  NAND3X0 U14185 ( .IN1(n13488), .IN2(n11350), .IN3(n13510), .QN(n13509) );
  NOR4X0 U14186 ( .IN1(g1146), .IN2(n8926), .IN3(n8527), .IN4(test_so7), .QN(
        n13488) );
  NAND2X0 U14187 ( .IN1(test_so7), .IN2(n8964), .QN(n13508) );
  NAND3X0 U14188 ( .IN1(n13511), .IN2(g1094), .IN3(n8888), .QN(n13507) );
  NAND3X0 U14189 ( .IN1(n13512), .IN2(g13259), .IN3(n11350), .QN(n13511) );
  INVX0 U14190 ( .INP(n13510), .ZN(n13512) );
  XOR2X1 U14191 ( .IN1(n13492), .IN2(n5328), .Q(n13510) );
  NAND2X0 U14192 ( .IN1(n9697), .IN2(DFF_24_n1), .QN(n13492) );
  INVX0 U14193 ( .INP(n13513), .ZN(n9697) );
  NAND3X0 U14194 ( .IN1(n13514), .IN2(n13515), .IN3(n13516), .QN(g29230) );
  NAND2X0 U14195 ( .IN1(n8977), .IN2(g907), .QN(n13516) );
  NAND3X0 U14196 ( .IN1(n11325), .IN2(n13517), .IN3(g911), .QN(n13515) );
  INVX0 U14197 ( .INP(n4196), .ZN(n13517) );
  NAND2X0 U14198 ( .IN1(n4196), .IN2(n5559), .QN(n13514) );
  NAND3X0 U14199 ( .IN1(n13518), .IN2(n13519), .IN3(n13520), .QN(g29229) );
  NAND2X0 U14200 ( .IN1(n9044), .IN2(g827), .QN(n13520) );
  NAND2X0 U14201 ( .IN1(n4517), .IN2(g723), .QN(n13519) );
  NAND3X0 U14202 ( .IN1(n4516), .IN2(n13521), .IN3(n5826), .QN(n13518) );
  NAND2X0 U14203 ( .IN1(n13522), .IN2(n13523), .QN(g29228) );
  NAND2X0 U14204 ( .IN1(n2404), .IN2(n13524), .QN(n13523) );
  XOR2X1 U14205 ( .IN1(test_so60), .IN2(n12987), .Q(n13524) );
  NOR2X0 U14206 ( .IN1(n12995), .IN2(n13525), .QN(n12987) );
  NOR2X0 U14207 ( .IN1(g11678), .IN2(n8627), .QN(n13525) );
  INVX0 U14208 ( .INP(n13526), .ZN(n13522) );
  NOR2X0 U14209 ( .IN1(n8900), .IN2(n8514), .QN(n13526) );
  NAND3X0 U14210 ( .IN1(n13527), .IN2(n13528), .IN3(n13529), .QN(g29227) );
  NAND2X0 U14211 ( .IN1(n9043), .IN2(g676), .QN(n13529) );
  NAND3X0 U14212 ( .IN1(n4523), .IN2(n13530), .IN3(n8603), .QN(n13528) );
  NAND2X0 U14213 ( .IN1(n4524), .IN2(test_so70), .QN(n13527) );
  NAND3X0 U14214 ( .IN1(n13531), .IN2(n13532), .IN3(n13533), .QN(g29226) );
  NAND2X0 U14215 ( .IN1(n9038), .IN2(g671), .QN(n13533) );
  NAND3X0 U14216 ( .IN1(n4525), .IN2(n13534), .IN3(g676), .QN(n13532) );
  INVX0 U14217 ( .INP(n4526), .ZN(n13534) );
  NAND3X0 U14218 ( .IN1(n4526), .IN2(n13530), .IN3(n5751), .QN(n13531) );
  NAND2X0 U14219 ( .IN1(n13535), .IN2(n13536), .QN(g29225) );
  NAND2X0 U14220 ( .IN1(n13537), .IN2(n4525), .QN(n13536) );
  INVX0 U14221 ( .INP(n13538), .ZN(n4525) );
  NAND2X0 U14222 ( .IN1(n13530), .IN2(n8920), .QN(n13538) );
  NOR2X0 U14223 ( .IN1(n5821), .IN2(n13539), .QN(n13530) );
  NOR4X0 U14224 ( .IN1(n4535), .IN2(n13540), .IN3(n8569), .IN4(n8158), .QN(
        n13539) );
  XNOR2X1 U14225 ( .IN1(g655), .IN2(n8552), .Q(n4535) );
  XOR2X1 U14226 ( .IN1(n8569), .IN2(n8079), .Q(n13537) );
  INVX0 U14227 ( .INP(n13541), .ZN(n8569) );
  NAND2X0 U14228 ( .IN1(n9037), .IN2(g667), .QN(n13535) );
  NAND3X0 U14229 ( .IN1(n13542), .IN2(n13543), .IN3(n13544), .QN(g29224) );
  NAND2X0 U14230 ( .IN1(n9046), .IN2(g572), .QN(n13544) );
  NAND3X0 U14231 ( .IN1(n2421), .IN2(n13545), .IN3(g586), .QN(n13543) );
  INVX0 U14232 ( .INP(n4201), .ZN(n13545) );
  NAND2X0 U14233 ( .IN1(n4201), .IN2(n5336), .QN(n13542) );
  NAND3X0 U14234 ( .IN1(n13546), .IN2(n13547), .IN3(n13548), .QN(g29223) );
  NAND2X0 U14235 ( .IN1(n13549), .IN2(n5708), .QN(n13548) );
  NAND2X0 U14236 ( .IN1(n8998), .IN2(g482), .QN(n13547) );
  NAND2X0 U14237 ( .IN1(n13550), .IN2(n8920), .QN(n13546) );
  NAND2X0 U14238 ( .IN1(n13551), .IN2(n13552), .QN(n13550) );
  NAND2X0 U14239 ( .IN1(n13553), .IN2(g490), .QN(n13552) );
  INVX0 U14240 ( .INP(n13549), .ZN(n13553) );
  NOR2X0 U14241 ( .IN1(n13554), .IN2(n5820), .QN(n13549) );
  NAND3X0 U14242 ( .IN1(n13555), .IN2(n13556), .IN3(n13557), .QN(g29222) );
  NAND2X0 U14243 ( .IN1(n13558), .IN2(g411), .QN(n13557) );
  NAND2X0 U14244 ( .IN1(n13559), .IN2(g417), .QN(n13556) );
  NAND2X0 U14245 ( .IN1(n13560), .IN2(n8920), .QN(n13559) );
  INVX0 U14246 ( .INP(n13561), .ZN(n13560) );
  NOR2X0 U14247 ( .IN1(n13562), .IN2(n3676), .QN(n13561) );
  NAND3X0 U14248 ( .IN1(n13563), .IN2(n3676), .IN3(n5358), .QN(n13555) );
  XOR2X1 U14249 ( .IN1(g417), .IN2(n13564), .Q(n3676) );
  NOR2X0 U14250 ( .IN1(n13565), .IN2(n13566), .QN(n13564) );
  NOR2X0 U14251 ( .IN1(g392), .IN2(n13567), .QN(n13566) );
  NOR2X0 U14252 ( .IN1(n13568), .IN2(n13569), .QN(n13567) );
  NOR2X0 U14253 ( .IN1(n8509), .IN2(n8164), .QN(n13569) );
  NOR2X0 U14254 ( .IN1(n8507), .IN2(g405), .QN(n13568) );
  NOR2X0 U14255 ( .IN1(n8510), .IN2(n13570), .QN(n13565) );
  NOR2X0 U14256 ( .IN1(n13571), .IN2(n13572), .QN(n13570) );
  NOR2X0 U14257 ( .IN1(n8164), .IN2(g405), .QN(n13572) );
  NOR2X0 U14258 ( .IN1(n8509), .IN2(n8508), .QN(n13571) );
  NAND3X0 U14259 ( .IN1(n13573), .IN2(n13574), .IN3(n13575), .QN(g28105) );
  NAND2X0 U14260 ( .IN1(n10857), .IN2(g5011), .QN(n13575) );
  NAND2X0 U14261 ( .IN1(n8998), .IN2(g6657), .QN(n13574) );
  NAND3X0 U14262 ( .IN1(n13034), .IN2(n10850), .IN3(n8888), .QN(n13573) );
  NAND2X0 U14263 ( .IN1(n13576), .IN2(n13577), .QN(n13034) );
  NAND2X0 U14264 ( .IN1(n5531), .IN2(n13578), .QN(n13577) );
  NAND4X0 U14265 ( .IN1(n13579), .IN2(n13580), .IN3(n13581), .IN4(n13582), 
        .QN(n13578) );
  NOR3X0 U14266 ( .IN1(n13583), .IN2(n13584), .IN3(n13585), .QN(n13582) );
  NOR2X0 U14267 ( .IN1(n13586), .IN2(n8592), .QN(n13585) );
  NOR2X0 U14268 ( .IN1(n13587), .IN2(n13588), .QN(n13586) );
  NOR2X0 U14269 ( .IN1(n8333), .IN2(n13589), .QN(n13587) );
  NOR2X0 U14270 ( .IN1(test_so80), .IN2(n13590), .QN(n13584) );
  NOR2X0 U14271 ( .IN1(n13591), .IN2(n13592), .QN(n13583) );
  NOR2X0 U14272 ( .IN1(n13593), .IN2(n13594), .QN(n13591) );
  NOR2X0 U14273 ( .IN1(n8392), .IN2(n8391), .QN(n13594) );
  NOR2X0 U14274 ( .IN1(n8390), .IN2(n8389), .QN(n13593) );
  NAND2X0 U14275 ( .IN1(n9214), .IN2(n13595), .QN(n13581) );
  NAND2X0 U14276 ( .IN1(n13596), .IN2(n13597), .QN(n13595) );
  NAND2X0 U14277 ( .IN1(g6723), .IN2(g6605), .QN(n13597) );
  NAND2X0 U14278 ( .IN1(g13099), .IN2(g6593), .QN(n13596) );
  NAND3X0 U14279 ( .IN1(g14749), .IN2(g6633), .IN3(n9215), .QN(n13580) );
  NAND3X0 U14280 ( .IN1(g17871), .IN2(g6617), .IN3(n9216), .QN(n13579) );
  NAND2X0 U14281 ( .IN1(n13598), .IN2(g6727), .QN(n13576) );
  NAND4X0 U14282 ( .IN1(n13599), .IN2(n13600), .IN3(n13601), .IN4(n13602), 
        .QN(n13598) );
  INVX0 U14283 ( .INP(n13603), .ZN(n13602) );
  NAND3X0 U14284 ( .IN1(n13604), .IN2(n13605), .IN3(n13606), .QN(n13603) );
  NAND2X0 U14285 ( .IN1(n13607), .IN2(test_so80), .QN(n13606) );
  NAND2X0 U14286 ( .IN1(n13608), .IN2(n13590), .QN(n13607) );
  INVX0 U14287 ( .INP(n13609), .ZN(n13590) );
  NAND3X0 U14288 ( .IN1(n13610), .IN2(n13611), .IN3(n13612), .QN(n13609) );
  NAND3X0 U14289 ( .IN1(g14828), .IN2(g6613), .IN3(n9214), .QN(n13612) );
  NAND3X0 U14290 ( .IN1(g17688), .IN2(g6645), .IN3(n9215), .QN(n13611) );
  NAND3X0 U14291 ( .IN1(g17778), .IN2(g6629), .IN3(n9216), .QN(n13610) );
  NAND2X0 U14292 ( .IN1(n9217), .IN2(test_so71), .QN(n13608) );
  NAND2X0 U14293 ( .IN1(n8592), .IN2(n13588), .QN(n13605) );
  NAND3X0 U14294 ( .IN1(n13613), .IN2(n13614), .IN3(n13615), .QN(n13588) );
  NAND3X0 U14295 ( .IN1(g6637), .IN2(g17778), .IN3(n9217), .QN(n13615) );
  NAND3X0 U14296 ( .IN1(g14828), .IN2(g6621), .IN3(n9215), .QN(n13614) );
  NAND3X0 U14297 ( .IN1(g6653), .IN2(g17688), .IN3(n9214), .QN(n13613) );
  NAND2X0 U14298 ( .IN1(n13616), .IN2(n9216), .QN(n13604) );
  INVX0 U14299 ( .INP(n13589), .ZN(n9216) );
  NAND2X0 U14300 ( .IN1(g6741), .IN2(g6682), .QN(n13589) );
  INVX0 U14301 ( .INP(n13617), .ZN(n13616) );
  NOR2X0 U14302 ( .IN1(n13618), .IN2(n13619), .QN(n13617) );
  NOR2X0 U14303 ( .IN1(n8389), .IN2(n8202), .QN(n13619) );
  NOR2X0 U14304 ( .IN1(n8391), .IN2(n8201), .QN(n13618) );
  NAND2X0 U14305 ( .IN1(n9215), .IN2(n13620), .QN(n13601) );
  NAND2X0 U14306 ( .IN1(n13621), .IN2(n13622), .QN(n13620) );
  NAND2X0 U14307 ( .IN1(g6589), .IN2(g6723), .QN(n13622) );
  NAND2X0 U14308 ( .IN1(g6581), .IN2(g13099), .QN(n13621) );
  NOR2X0 U14309 ( .IN1(g6682), .IN2(g6741), .QN(n9215) );
  NAND3X0 U14310 ( .IN1(g14749), .IN2(g6625), .IN3(n9214), .QN(n13600) );
  NOR2X0 U14311 ( .IN1(g6741), .IN2(n5590), .QN(n9214) );
  NAND3X0 U14312 ( .IN1(g6609), .IN2(g17871), .IN3(n9217), .QN(n13599) );
  INVX0 U14313 ( .INP(n13592), .ZN(n9217) );
  NAND2X0 U14314 ( .IN1(n5590), .IN2(g6741), .QN(n13592) );
  NAND3X0 U14315 ( .IN1(n13623), .IN2(n13624), .IN3(n13625), .QN(g28102) );
  NAND2X0 U14316 ( .IN1(n10873), .IN2(g4826), .QN(n13625) );
  NAND2X0 U14317 ( .IN1(n8998), .IN2(g6311), .QN(n13624) );
  NAND3X0 U14318 ( .IN1(n10862), .IN2(n13066), .IN3(n8888), .QN(n13623) );
  NAND2X0 U14319 ( .IN1(n13626), .IN2(n13627), .QN(n13066) );
  NAND2X0 U14320 ( .IN1(test_so69), .IN2(n13628), .QN(n13627) );
  NAND4X0 U14321 ( .IN1(n13629), .IN2(n13630), .IN3(n13631), .IN4(n13632), 
        .QN(n13628) );
  NOR3X0 U14322 ( .IN1(n13633), .IN2(n13634), .IN3(n13635), .QN(n13632) );
  NOR2X0 U14323 ( .IN1(n5437), .IN2(n13636), .QN(n13635) );
  NOR2X0 U14324 ( .IN1(n13637), .IN2(n13638), .QN(n13636) );
  INVX0 U14325 ( .INP(n13639), .ZN(n13637) );
  NAND2X0 U14326 ( .IN1(g6239), .IN2(n10864), .QN(n13639) );
  INVX0 U14327 ( .INP(n13640), .ZN(n13634) );
  NAND2X0 U14328 ( .IN1(n13641), .IN2(n5437), .QN(n13640) );
  NOR2X0 U14329 ( .IN1(n13642), .IN2(n13643), .QN(n13633) );
  NOR2X0 U14330 ( .IN1(n13644), .IN2(n13645), .QN(n13642) );
  NOR2X0 U14331 ( .IN1(n8399), .IN2(n8209), .QN(n13645) );
  NOR2X0 U14332 ( .IN1(n8401), .IN2(n8208), .QN(n13644) );
  NAND2X0 U14333 ( .IN1(n13646), .IN2(n13647), .QN(n13631) );
  NAND2X0 U14334 ( .IN1(n13648), .IN2(n13649), .QN(n13647) );
  NAND2X0 U14335 ( .IN1(g6243), .IN2(g6377), .QN(n13649) );
  NAND2X0 U14336 ( .IN1(g6235), .IN2(g13085), .QN(n13648) );
  NAND3X0 U14337 ( .IN1(g6263), .IN2(g17845), .IN3(n10864), .QN(n13630) );
  NAND3X0 U14338 ( .IN1(g14705), .IN2(g6279), .IN3(n10869), .QN(n13629) );
  NAND2X0 U14339 ( .IN1(n13650), .IN2(n8614), .QN(n13626) );
  NAND4X0 U14340 ( .IN1(n13651), .IN2(n13652), .IN3(n13653), .IN4(n13654), 
        .QN(n13650) );
  NOR3X0 U14341 ( .IN1(n13655), .IN2(n13656), .IN3(n13657), .QN(n13654) );
  NOR2X0 U14342 ( .IN1(n5437), .IN2(n13658), .QN(n13657) );
  NOR2X0 U14343 ( .IN1(n13659), .IN2(n13641), .QN(n13658) );
  NAND3X0 U14344 ( .IN1(n13660), .IN2(n13661), .IN3(n13662), .QN(n13641) );
  NAND3X0 U14345 ( .IN1(g6307), .IN2(g17649), .IN3(n10869), .QN(n13662) );
  NAND3X0 U14346 ( .IN1(g6291), .IN2(g17760), .IN3(n10864), .QN(n13661) );
  NAND3X0 U14347 ( .IN1(g14779), .IN2(g6275), .IN3(n13646), .QN(n13660) );
  NOR2X0 U14348 ( .IN1(n8339), .IN2(n13643), .QN(n13659) );
  INVX0 U14349 ( .INP(n13663), .ZN(n13656) );
  NAND2X0 U14350 ( .IN1(n13638), .IN2(n5437), .QN(n13663) );
  NAND3X0 U14351 ( .IN1(n13664), .IN2(n13665), .IN3(n13666), .QN(n13638) );
  NAND3X0 U14352 ( .IN1(g17760), .IN2(g6283), .IN3(n10063), .QN(n13666) );
  NAND3X0 U14353 ( .IN1(g17649), .IN2(g6299), .IN3(n13646), .QN(n13665) );
  NAND3X0 U14354 ( .IN1(g14779), .IN2(g6267), .IN3(n10869), .QN(n13664) );
  NOR2X0 U14355 ( .IN1(n13667), .IN2(n13668), .QN(n13655) );
  NOR2X0 U14356 ( .IN1(n13669), .IN2(n13670), .QN(n13667) );
  NOR2X0 U14357 ( .IN1(n8429), .IN2(n8428), .QN(n13670) );
  NOR2X0 U14358 ( .IN1(n8427), .IN2(n8426), .QN(n13669) );
  NAND2X0 U14359 ( .IN1(n10864), .IN2(n13671), .QN(n13653) );
  NAND2X0 U14360 ( .IN1(n13672), .IN2(n13673), .QN(n13671) );
  NAND2X0 U14361 ( .IN1(g17743), .IN2(g6303), .QN(n13673) );
  NAND2X0 U14362 ( .IN1(g17685), .IN2(g6251), .QN(n13672) );
  NAND3X0 U14363 ( .IN1(g14705), .IN2(g6287), .IN3(n13646), .QN(n13652) );
  NAND3X0 U14364 ( .IN1(g17845), .IN2(g6271), .IN3(n10063), .QN(n13651) );
  NAND3X0 U14365 ( .IN1(n13674), .IN2(n13675), .IN3(n13676), .QN(g28099) );
  NAND2X0 U14366 ( .IN1(n10889), .IN2(g4831), .QN(n13676) );
  NAND2X0 U14367 ( .IN1(test_so13), .IN2(n8959), .QN(n13675) );
  NAND3X0 U14368 ( .IN1(n10878), .IN2(n13098), .IN3(n8888), .QN(n13674) );
  NAND2X0 U14369 ( .IN1(n13677), .IN2(n13678), .QN(n13098) );
  NAND2X0 U14370 ( .IN1(n5528), .IN2(n13679), .QN(n13678) );
  NAND4X0 U14371 ( .IN1(n13680), .IN2(n13681), .IN3(n13682), .IN4(n13683), 
        .QN(n13679) );
  NOR3X0 U14372 ( .IN1(n13684), .IN2(n13685), .IN3(n13686), .QN(n13683) );
  NOR2X0 U14373 ( .IN1(n5432), .IN2(n13687), .QN(n13686) );
  NOR2X0 U14374 ( .IN1(n13688), .IN2(n13689), .QN(n13687) );
  NOR2X0 U14375 ( .IN1(n8324), .IN2(n13690), .QN(n13688) );
  INVX0 U14376 ( .INP(n13691), .ZN(n13685) );
  NAND2X0 U14377 ( .IN1(n13692), .IN2(n5432), .QN(n13691) );
  NOR2X0 U14378 ( .IN1(n13693), .IN2(n13694), .QN(n13684) );
  NOR2X0 U14379 ( .IN1(n13695), .IN2(n13696), .QN(n13693) );
  NOR2X0 U14380 ( .IN1(n8409), .IN2(n8408), .QN(n13696) );
  NOR2X0 U14381 ( .IN1(n8407), .IN2(n8406), .QN(n13695) );
  NAND2X0 U14382 ( .IN1(n10880), .IN2(n13697), .QN(n13682) );
  NAND2X0 U14383 ( .IN1(n13698), .IN2(n13699), .QN(n13697) );
  NAND2X0 U14384 ( .IN1(g17715), .IN2(g5957), .QN(n13699) );
  NAND2X0 U14385 ( .IN1(g17646), .IN2(g5905), .QN(n13698) );
  NAND3X0 U14386 ( .IN1(g14673), .IN2(g5941), .IN3(n13700), .QN(n13681) );
  NAND3X0 U14387 ( .IN1(g17819), .IN2(g5925), .IN3(n10068), .QN(n13680) );
  NAND2X0 U14388 ( .IN1(n13701), .IN2(g6035), .QN(n13677) );
  NAND4X0 U14389 ( .IN1(n13702), .IN2(n13703), .IN3(n13704), .IN4(n13705), 
        .QN(n13701) );
  NOR3X0 U14390 ( .IN1(n13706), .IN2(n13707), .IN3(n13708), .QN(n13705) );
  NOR2X0 U14391 ( .IN1(n5432), .IN2(n13709), .QN(n13708) );
  NOR2X0 U14392 ( .IN1(n13710), .IN2(n13692), .QN(n13709) );
  NAND3X0 U14393 ( .IN1(n13711), .IN2(n13712), .IN3(n13713), .QN(n13692) );
  NAND3X0 U14394 ( .IN1(g17739), .IN2(g5937), .IN3(n10068), .QN(n13713) );
  NAND3X0 U14395 ( .IN1(g17607), .IN2(g5953), .IN3(n13700), .QN(n13712) );
  NAND3X0 U14396 ( .IN1(g14738), .IN2(g5921), .IN3(n10885), .QN(n13711) );
  INVX0 U14397 ( .INP(n13714), .ZN(n13710) );
  NAND2X0 U14398 ( .IN1(g5893), .IN2(n10880), .QN(n13714) );
  INVX0 U14399 ( .INP(n13715), .ZN(n13707) );
  NAND2X0 U14400 ( .IN1(n13689), .IN2(n5432), .QN(n13715) );
  NAND3X0 U14401 ( .IN1(n13716), .IN2(n13717), .IN3(n13718), .QN(n13689) );
  NAND3X0 U14402 ( .IN1(g5961), .IN2(g17607), .IN3(n10885), .QN(n13718) );
  NAND3X0 U14403 ( .IN1(g5945), .IN2(g17739), .IN3(n10880), .QN(n13717) );
  NAND3X0 U14404 ( .IN1(g14738), .IN2(g5929), .IN3(n13700), .QN(n13716) );
  NOR2X0 U14405 ( .IN1(n13719), .IN2(n13690), .QN(n13706) );
  NOR2X0 U14406 ( .IN1(n13720), .IN2(n13721), .QN(n13719) );
  NOR2X0 U14407 ( .IN1(n8377), .IN2(n8626), .QN(n13721) );
  NOR2X0 U14408 ( .IN1(n8375), .IN2(n8216), .QN(n13720) );
  NAND2X0 U14409 ( .IN1(n13700), .IN2(n13722), .QN(n13704) );
  NAND2X0 U14410 ( .IN1(n13723), .IN2(n13724), .QN(n13722) );
  NAND2X0 U14411 ( .IN1(g5897), .IN2(g6031), .QN(n13724) );
  NAND2X0 U14412 ( .IN1(g5889), .IN2(g13068), .QN(n13723) );
  NAND3X0 U14413 ( .IN1(n10880), .IN2(g17819), .IN3(test_so28), .QN(n13703) );
  NAND3X0 U14414 ( .IN1(g14673), .IN2(g5933), .IN3(n10885), .QN(n13702) );
  NAND3X0 U14415 ( .IN1(n13725), .IN2(n13726), .IN3(n13727), .QN(g28096) );
  NAND2X0 U14416 ( .IN1(n10905), .IN2(g4821), .QN(n13727) );
  NAND2X0 U14417 ( .IN1(n8998), .IN2(g5619), .QN(n13726) );
  NAND3X0 U14418 ( .IN1(n10894), .IN2(n13131), .IN3(n8888), .QN(n13725) );
  NAND2X0 U14419 ( .IN1(n13728), .IN2(n13729), .QN(n13131) );
  NAND2X0 U14420 ( .IN1(n5529), .IN2(n13730), .QN(n13729) );
  NAND4X0 U14421 ( .IN1(n13731), .IN2(n13732), .IN3(n13733), .IN4(n13734), 
        .QN(n13730) );
  NOR3X0 U14422 ( .IN1(n13735), .IN2(n13736), .IN3(n13737), .QN(n13734) );
  NOR2X0 U14423 ( .IN1(n5439), .IN2(n13738), .QN(n13737) );
  NOR2X0 U14424 ( .IN1(n13739), .IN2(n13740), .QN(n13738) );
  NOR2X0 U14425 ( .IN1(n8327), .IN2(n13741), .QN(n13739) );
  INVX0 U14426 ( .INP(n13742), .ZN(n13736) );
  NAND2X0 U14427 ( .IN1(n13743), .IN2(n5439), .QN(n13742) );
  NOR2X0 U14428 ( .IN1(n13744), .IN2(n13745), .QN(n13735) );
  NOR2X0 U14429 ( .IN1(n13746), .IN2(n13747), .QN(n13744) );
  NOR2X0 U14430 ( .IN1(n8413), .IN2(n8412), .QN(n13747) );
  NOR2X0 U14431 ( .IN1(n8411), .IN2(n8410), .QN(n13746) );
  NAND2X0 U14432 ( .IN1(n10896), .IN2(n13748), .QN(n13733) );
  NAND2X0 U14433 ( .IN1(n13749), .IN2(n13750), .QN(n13748) );
  NAND2X0 U14434 ( .IN1(g17678), .IN2(g5611), .QN(n13750) );
  NAND2X0 U14435 ( .IN1(test_so6), .IN2(g17604), .QN(n13749) );
  NAND3X0 U14436 ( .IN1(g14635), .IN2(g5595), .IN3(n13751), .QN(n13732) );
  NAND3X0 U14437 ( .IN1(g17813), .IN2(g5579), .IN3(n10076), .QN(n13731) );
  NAND2X0 U14438 ( .IN1(n13752), .IN2(g5689), .QN(n13728) );
  NAND4X0 U14439 ( .IN1(n13753), .IN2(n13754), .IN3(n13755), .IN4(n13756), 
        .QN(n13752) );
  NOR3X0 U14440 ( .IN1(n13757), .IN2(n13758), .IN3(n13759), .QN(n13756) );
  NOR2X0 U14441 ( .IN1(n5439), .IN2(n13760), .QN(n13759) );
  NOR2X0 U14442 ( .IN1(n13761), .IN2(n13743), .QN(n13760) );
  NAND3X0 U14443 ( .IN1(n13762), .IN2(n13763), .IN3(n13764), .QN(n13743) );
  NAND3X0 U14444 ( .IN1(n10076), .IN2(g17711), .IN3(test_so5), .QN(n13764) );
  NAND3X0 U14445 ( .IN1(g17580), .IN2(g5607), .IN3(n13751), .QN(n13763) );
  NAND3X0 U14446 ( .IN1(g14694), .IN2(g5575), .IN3(n10901), .QN(n13762) );
  INVX0 U14447 ( .INP(n13765), .ZN(n13761) );
  NAND2X0 U14448 ( .IN1(g5547), .IN2(n10896), .QN(n13765) );
  INVX0 U14449 ( .INP(n13766), .ZN(n13758) );
  NAND2X0 U14450 ( .IN1(n13740), .IN2(n5439), .QN(n13766) );
  NAND3X0 U14451 ( .IN1(n13767), .IN2(n13768), .IN3(n13769), .QN(n13740) );
  NAND3X0 U14452 ( .IN1(g5615), .IN2(g17580), .IN3(n10901), .QN(n13769) );
  NAND3X0 U14453 ( .IN1(g5599), .IN2(g17711), .IN3(n10896), .QN(n13768) );
  NAND3X0 U14454 ( .IN1(g14694), .IN2(g5583), .IN3(n13751), .QN(n13767) );
  NOR2X0 U14455 ( .IN1(n13770), .IN2(n13741), .QN(n13757) );
  NOR2X0 U14456 ( .IN1(n13771), .IN2(n13772), .QN(n13770) );
  NOR2X0 U14457 ( .IN1(n8380), .IN2(n8198), .QN(n13772) );
  NOR2X0 U14458 ( .IN1(n8382), .IN2(n8197), .QN(n13771) );
  NAND2X0 U14459 ( .IN1(n13751), .IN2(n13773), .QN(n13755) );
  NAND2X0 U14460 ( .IN1(n13774), .IN2(n13775), .QN(n13773) );
  NAND2X0 U14461 ( .IN1(g5551), .IN2(g5685), .QN(n13775) );
  NAND2X0 U14462 ( .IN1(g5543), .IN2(g13049), .QN(n13774) );
  NAND3X0 U14463 ( .IN1(g5571), .IN2(g17813), .IN3(n10896), .QN(n13754) );
  NAND3X0 U14464 ( .IN1(g14635), .IN2(g5587), .IN3(n10901), .QN(n13753) );
  NAND3X0 U14465 ( .IN1(n13776), .IN2(n13777), .IN3(n13778), .QN(g28093) );
  NAND2X0 U14466 ( .IN1(n10917), .IN2(g29220), .QN(n13778) );
  NAND2X0 U14467 ( .IN1(n8998), .IN2(g5272), .QN(n13777) );
  NAND3X0 U14468 ( .IN1(n13164), .IN2(g33959), .IN3(n8888), .QN(n13776) );
  NAND2X0 U14469 ( .IN1(n13779), .IN2(n13780), .QN(n13164) );
  NAND2X0 U14470 ( .IN1(test_so10), .IN2(n13781), .QN(n13780) );
  NAND4X0 U14471 ( .IN1(n13782), .IN2(n13783), .IN3(n13784), .IN4(n13785), 
        .QN(n13781) );
  NOR3X0 U14472 ( .IN1(n13786), .IN2(n13787), .IN3(n13788), .QN(n13785) );
  NOR2X0 U14473 ( .IN1(n5438), .IN2(n13789), .QN(n13788) );
  NOR2X0 U14474 ( .IN1(n13790), .IN2(n13791), .QN(n13789) );
  NOR2X0 U14475 ( .IN1(n8215), .IN2(n13792), .QN(n13790) );
  INVX0 U14476 ( .INP(n13793), .ZN(n13787) );
  NAND2X0 U14477 ( .IN1(n13794), .IN2(n5438), .QN(n13793) );
  NOR2X0 U14478 ( .IN1(n13795), .IN2(n13796), .QN(n13786) );
  NOR2X0 U14479 ( .IN1(n13797), .IN2(n13798), .QN(n13795) );
  NOR2X0 U14480 ( .IN1(n8370), .IN2(n8213), .QN(n13798) );
  NOR2X0 U14481 ( .IN1(n8372), .IN2(n8212), .QN(n13797) );
  NAND2X0 U14482 ( .IN1(n9208), .IN2(n13799), .QN(n13784) );
  NAND2X0 U14483 ( .IN1(n13800), .IN2(n13801), .QN(n13799) );
  NAND2X0 U14484 ( .IN1(g5339), .IN2(g5204), .QN(n13801) );
  NAND2X0 U14485 ( .IN1(g13039), .IN2(g5196), .QN(n13800) );
  NAND3X0 U14486 ( .IN1(g14597), .IN2(g5240), .IN3(n9207), .QN(n13783) );
  NAND3X0 U14487 ( .IN1(g5224), .IN2(g17787), .IN3(n9209), .QN(n13782) );
  NAND2X0 U14488 ( .IN1(n13802), .IN2(n8613), .QN(n13779) );
  NAND4X0 U14489 ( .IN1(n13803), .IN2(n13804), .IN3(n13805), .IN4(n13806), 
        .QN(n13802) );
  NOR3X0 U14490 ( .IN1(n13807), .IN2(n13808), .IN3(n13809), .QN(n13806) );
  NOR2X0 U14491 ( .IN1(n5438), .IN2(n13810), .QN(n13809) );
  NOR2X0 U14492 ( .IN1(n13811), .IN2(n13794), .QN(n13810) );
  NAND3X0 U14493 ( .IN1(n13812), .IN2(n13813), .IN3(n13814), .QN(n13794) );
  NAND3X0 U14494 ( .IN1(g5252), .IN2(g17674), .IN3(n9209), .QN(n13814) );
  INVX0 U14495 ( .INP(n13792), .ZN(n9209) );
  NAND3X0 U14496 ( .IN1(g5268), .IN2(g17519), .IN3(n9207), .QN(n13813) );
  NAND3X0 U14497 ( .IN1(g14662), .IN2(g5236), .IN3(n9208), .QN(n13812) );
  NOR2X0 U14498 ( .IN1(n8321), .IN2(n13796), .QN(n13811) );
  INVX0 U14499 ( .INP(n13815), .ZN(n13808) );
  NAND2X0 U14500 ( .IN1(n13791), .IN2(n5438), .QN(n13815) );
  NAND3X0 U14501 ( .IN1(n13816), .IN2(n13817), .IN3(n13818), .QN(n13791) );
  NAND3X0 U14502 ( .IN1(g17674), .IN2(g5244), .IN3(g31860), .QN(n13818) );
  NAND3X0 U14503 ( .IN1(n9207), .IN2(g14662), .IN3(test_so82), .QN(n13817) );
  NAND3X0 U14504 ( .IN1(g17519), .IN2(g5260), .IN3(n9208), .QN(n13816) );
  NOR2X0 U14505 ( .IN1(n13819), .IN2(n13792), .QN(n13807) );
  NAND2X0 U14506 ( .IN1(n5588), .IN2(g5357), .QN(n13792) );
  NOR2X0 U14507 ( .IN1(n13820), .IN2(n13821), .QN(n13819) );
  NOR2X0 U14508 ( .IN1(n8373), .IN2(n8372), .QN(n13821) );
  NOR2X0 U14509 ( .IN1(n8371), .IN2(n8370), .QN(n13820) );
  NAND2X0 U14510 ( .IN1(n9207), .IN2(n13822), .QN(n13805) );
  NAND2X0 U14511 ( .IN1(n13823), .IN2(n13824), .QN(n13822) );
  NAND2X0 U14512 ( .IN1(g5220), .IN2(g5339), .QN(n13824) );
  NAND2X0 U14513 ( .IN1(g5208), .IN2(g13039), .QN(n13823) );
  NOR2X0 U14514 ( .IN1(g5357), .IN2(n5588), .QN(n9207) );
  NAND3X0 U14515 ( .IN1(g14597), .IN2(g5248), .IN3(n9208), .QN(n13804) );
  NOR2X0 U14516 ( .IN1(g5297), .IN2(g5357), .QN(n9208) );
  NAND3X0 U14517 ( .IN1(g17787), .IN2(g5232), .IN3(g31860), .QN(n13803) );
  INVX0 U14518 ( .INP(n13796), .ZN(g31860) );
  NAND2X0 U14519 ( .IN1(g5357), .IN2(g5297), .QN(n13796) );
  NAND2X0 U14520 ( .IN1(n13825), .IN2(n13826), .QN(g28092) );
  NAND2X0 U14521 ( .IN1(n8998), .IN2(g5057), .QN(n13826) );
  NAND2X0 U14522 ( .IN1(n11843), .IN2(n8920), .QN(n13825) );
  NAND2X0 U14523 ( .IN1(n13827), .IN2(n13828), .QN(n11843) );
  INVX0 U14524 ( .INP(n13829), .ZN(n13828) );
  NOR3X0 U14525 ( .IN1(n5615), .IN2(n8496), .IN3(g5046), .QN(n13827) );
  NAND2X0 U14526 ( .IN1(n13830), .IN2(n13831), .QN(g28091) );
  NAND2X0 U14527 ( .IN1(n8998), .IN2(g5069), .QN(n13831) );
  NAND2X0 U14528 ( .IN1(n11842), .IN2(n8920), .QN(n13830) );
  NAND2X0 U14529 ( .IN1(n13832), .IN2(n13829), .QN(n11842) );
  NAND2X0 U14530 ( .IN1(n13833), .IN2(n13834), .QN(n13829) );
  NAND2X0 U14531 ( .IN1(g84), .IN2(g5041), .QN(n13834) );
  NAND2X0 U14532 ( .IN1(n13835), .IN2(g5052), .QN(n13833) );
  INVX0 U14533 ( .INP(g84), .ZN(n13835) );
  NOR3X0 U14534 ( .IN1(n5578), .IN2(n8498), .IN3(g5057), .QN(n13832) );
  NAND2X0 U14535 ( .IN1(n13836), .IN2(n13837), .QN(g28090) );
  NAND3X0 U14536 ( .IN1(n13838), .IN2(n8869), .IN3(n10120), .QN(n13837) );
  INVX0 U14537 ( .INP(n10118), .ZN(n10120) );
  NAND2X0 U14538 ( .IN1(n13839), .IN2(n9296), .QN(n10118) );
  NAND2X0 U14539 ( .IN1(n5770), .IN2(n13840), .QN(n13838) );
  NAND2X0 U14540 ( .IN1(n10933), .IN2(n13841), .QN(n13840) );
  NAND4X0 U14541 ( .IN1(n13842), .IN2(n13843), .IN3(n13844), .IN4(n13845), 
        .QN(n13841) );
  NAND2X0 U14542 ( .IN1(n10940), .IN2(g4045), .QN(n13845) );
  NAND2X0 U14543 ( .IN1(n8306), .IN2(n13846), .QN(n13844) );
  NAND2X0 U14544 ( .IN1(n10064), .IN2(g4049), .QN(n13843) );
  NAND2X0 U14545 ( .IN1(n8305), .IN2(n10935), .QN(n13842) );
  NAND2X0 U14546 ( .IN1(n10944), .IN2(g4961), .QN(n13836) );
  NAND2X0 U14547 ( .IN1(n13847), .IN2(n13848), .QN(g28089) );
  NAND3X0 U14548 ( .IN1(n13849), .IN2(n8869), .IN3(n10126), .QN(n13848) );
  INVX0 U14549 ( .INP(n10125), .ZN(n10126) );
  NAND2X0 U14550 ( .IN1(n13839), .IN2(n9297), .QN(n10125) );
  NAND2X0 U14551 ( .IN1(n5772), .IN2(n13850), .QN(n13849) );
  NAND2X0 U14552 ( .IN1(n10949), .IN2(n13851), .QN(n13850) );
  NAND4X0 U14553 ( .IN1(n13852), .IN2(n13853), .IN3(n13854), .IN4(n13855), 
        .QN(n13851) );
  NAND2X0 U14554 ( .IN1(n10956), .IN2(g3694), .QN(n13855) );
  NAND2X0 U14555 ( .IN1(n8302), .IN2(n13856), .QN(n13854) );
  NAND2X0 U14556 ( .IN1(n10069), .IN2(g3698), .QN(n13853) );
  NAND2X0 U14557 ( .IN1(n8301), .IN2(n10951), .QN(n13852) );
  NAND2X0 U14558 ( .IN1(n10960), .IN2(g4950), .QN(n13847) );
  NAND2X0 U14559 ( .IN1(n13857), .IN2(n13858), .QN(g28088) );
  NAND3X0 U14560 ( .IN1(n13859), .IN2(n8869), .IN3(n10134), .QN(n13858) );
  INVX0 U14561 ( .INP(n10131), .ZN(n10134) );
  NAND2X0 U14562 ( .IN1(n13839), .IN2(n9292), .QN(n10131) );
  NAND2X0 U14563 ( .IN1(n5776), .IN2(n13860), .QN(n13859) );
  NAND2X0 U14564 ( .IN1(n10969), .IN2(n13861), .QN(n13860) );
  NAND4X0 U14565 ( .IN1(n13862), .IN2(n13863), .IN3(n13864), .IN4(n13865), 
        .QN(n13861) );
  INVX0 U14566 ( .INP(n13866), .ZN(n13865) );
  NOR2X0 U14567 ( .IN1(n10970), .IN2(n8297), .QN(n13866) );
  INVX0 U14568 ( .INP(n13867), .ZN(n10970) );
  NAND2X0 U14569 ( .IN1(n8297), .IN2(n13868), .QN(n13864) );
  NAND2X0 U14570 ( .IN1(n10077), .IN2(g3347), .QN(n13863) );
  NAND2X0 U14571 ( .IN1(n8296), .IN2(n13869), .QN(n13862) );
  NAND2X0 U14572 ( .IN1(n10975), .IN2(g4939), .QN(n13857) );
  NAND2X0 U14573 ( .IN1(n13870), .IN2(n13871), .QN(g28087) );
  NAND2X0 U14574 ( .IN1(n13872), .IN2(n9749), .QN(n13871) );
  INVX0 U14575 ( .INP(n10142), .ZN(n9749) );
  NAND2X0 U14576 ( .IN1(n13839), .IN2(n9293), .QN(n10142) );
  INVX0 U14577 ( .INP(n9279), .ZN(n13839) );
  NAND3X0 U14578 ( .IN1(g4966), .IN2(n8587), .IN3(g4983), .QN(n9279) );
  NOR2X0 U14579 ( .IN1(n8957), .IN2(n13873), .QN(n13872) );
  NOR2X0 U14580 ( .IN1(n4689), .IN2(g4894), .QN(n13873) );
  NAND2X0 U14581 ( .IN1(n10857), .IN2(g4894), .QN(n13870) );
  NOR2X0 U14582 ( .IN1(n10850), .IN2(n8943), .QN(n10857) );
  INVX0 U14583 ( .INP(n8575), .ZN(n10850) );
  NAND2X0 U14584 ( .IN1(g4836), .IN2(n13874), .QN(n8575) );
  NAND3X0 U14585 ( .IN1(n13875), .IN2(g4888), .IN3(n9292), .QN(n13874) );
  NOR2X0 U14586 ( .IN1(g4899), .IN2(g4975), .QN(n9292) );
  NAND2X0 U14587 ( .IN1(n13876), .IN2(n13877), .QN(g28086) );
  NAND3X0 U14588 ( .IN1(n13878), .IN2(n8869), .IN3(n10152), .QN(n13877) );
  INVX0 U14589 ( .INP(n10150), .ZN(n10152) );
  NAND2X0 U14590 ( .IN1(n13879), .IN2(n9253), .QN(n10150) );
  NAND2X0 U14591 ( .IN1(n5769), .IN2(n13880), .QN(n13878) );
  NAND2X0 U14592 ( .IN1(n10862), .IN2(n13881), .QN(n13880) );
  NAND4X0 U14593 ( .IN1(n13882), .IN2(n13883), .IN3(n13884), .IN4(n13885), 
        .QN(n13881) );
  NAND2X0 U14594 ( .IN1(n10063), .IN2(g6390), .QN(n13885) );
  INVX0 U14595 ( .INP(n13643), .ZN(n10063) );
  NAND2X0 U14596 ( .IN1(g6395), .IN2(g6336), .QN(n13643) );
  NAND2X0 U14597 ( .IN1(n8298), .IN2(n10864), .QN(n13884) );
  NOR2X0 U14598 ( .IN1(g6336), .IN2(n5396), .QN(n10864) );
  NAND2X0 U14599 ( .IN1(n10869), .IN2(g6386), .QN(n13883) );
  INVX0 U14600 ( .INP(n13668), .ZN(n10869) );
  NAND2X0 U14601 ( .IN1(n5396), .IN2(g6336), .QN(n13668) );
  NAND2X0 U14602 ( .IN1(n8299), .IN2(n13646), .QN(n13882) );
  NOR2X0 U14603 ( .IN1(g6395), .IN2(g6336), .QN(n13646) );
  NAND2X0 U14604 ( .IN1(n10873), .IN2(g4771), .QN(n13876) );
  NOR2X0 U14605 ( .IN1(n10862), .IN2(n8943), .QN(n10873) );
  INVX0 U14606 ( .INP(n10868), .ZN(n10862) );
  NAND2X0 U14607 ( .IN1(g4688), .IN2(n13886), .QN(n10868) );
  NAND3X0 U14608 ( .IN1(n13887), .IN2(g4765), .IN3(n9256), .QN(n13886) );
  NAND2X0 U14609 ( .IN1(n13888), .IN2(n13889), .QN(g28085) );
  NAND3X0 U14610 ( .IN1(n13890), .IN2(n8869), .IN3(n10158), .QN(n13889) );
  INVX0 U14611 ( .INP(n10157), .ZN(n10158) );
  NAND2X0 U14612 ( .IN1(n13879), .IN2(n9254), .QN(n10157) );
  NAND2X0 U14613 ( .IN1(n5775), .IN2(n13891), .QN(n13890) );
  NAND2X0 U14614 ( .IN1(n10878), .IN2(n13892), .QN(n13891) );
  NAND4X0 U14615 ( .IN1(n13893), .IN2(n13894), .IN3(n13895), .IN4(n13896), 
        .QN(n13892) );
  NAND2X0 U14616 ( .IN1(n10880), .IN2(n8610), .QN(n13896) );
  NOR2X0 U14617 ( .IN1(g5990), .IN2(n8597), .QN(n10880) );
  NAND2X0 U14618 ( .IN1(test_so50), .IN2(n10068), .QN(n13895) );
  INVX0 U14619 ( .INP(n13690), .ZN(n10068) );
  NAND2X0 U14620 ( .IN1(test_so57), .IN2(g5990), .QN(n13690) );
  NAND2X0 U14621 ( .IN1(n10885), .IN2(g6040), .QN(n13894) );
  INVX0 U14622 ( .INP(n13694), .ZN(n10885) );
  NAND2X0 U14623 ( .IN1(g5990), .IN2(n8597), .QN(n13694) );
  NAND2X0 U14624 ( .IN1(n8300), .IN2(n13700), .QN(n13893) );
  NOR2X0 U14625 ( .IN1(g5990), .IN2(test_so57), .QN(n13700) );
  NAND2X0 U14626 ( .IN1(n10889), .IN2(g4760), .QN(n13888) );
  NOR2X0 U14627 ( .IN1(n10878), .IN2(n8943), .QN(n10889) );
  INVX0 U14628 ( .INP(n10884), .ZN(n10878) );
  NAND2X0 U14629 ( .IN1(g4681), .IN2(n13897), .QN(n10884) );
  NAND3X0 U14630 ( .IN1(n13887), .IN2(g4754), .IN3(n9253), .QN(n13897) );
  INVX0 U14631 ( .INP(n9263), .ZN(n9253) );
  NAND2X0 U14632 ( .IN1(n5361), .IN2(g4709), .QN(n9263) );
  NAND2X0 U14633 ( .IN1(n13898), .IN2(n13899), .QN(g28084) );
  NAND3X0 U14634 ( .IN1(n13900), .IN2(n8870), .IN3(n10166), .QN(n13899) );
  INVX0 U14635 ( .INP(n10163), .ZN(n10166) );
  NAND2X0 U14636 ( .IN1(n13879), .IN2(n9257), .QN(n10163) );
  NAND2X0 U14637 ( .IN1(n8635), .IN2(n13901), .QN(n13900) );
  NAND2X0 U14638 ( .IN1(n10894), .IN2(n13902), .QN(n13901) );
  NAND4X0 U14639 ( .IN1(n13903), .IN2(n13904), .IN3(n13905), .IN4(n13906), 
        .QN(n13902) );
  NAND2X0 U14640 ( .IN1(n10076), .IN2(g5698), .QN(n13906) );
  INVX0 U14641 ( .INP(n13741), .ZN(n10076) );
  NAND2X0 U14642 ( .IN1(g5703), .IN2(g5644), .QN(n13741) );
  NAND2X0 U14643 ( .IN1(n8303), .IN2(n10896), .QN(n13905) );
  NOR2X0 U14644 ( .IN1(g5644), .IN2(n5397), .QN(n10896) );
  NAND2X0 U14645 ( .IN1(n10901), .IN2(g5694), .QN(n13904) );
  INVX0 U14646 ( .INP(n13745), .ZN(n10901) );
  NAND2X0 U14647 ( .IN1(n5397), .IN2(g5644), .QN(n13745) );
  NAND2X0 U14648 ( .IN1(n8304), .IN2(n13751), .QN(n13903) );
  NOR2X0 U14649 ( .IN1(g5703), .IN2(g5644), .QN(n13751) );
  NAND2X0 U14650 ( .IN1(n10905), .IN2(test_so18), .QN(n13898) );
  NOR2X0 U14651 ( .IN1(n10894), .IN2(n8942), .QN(n10905) );
  INVX0 U14652 ( .INP(n10900), .ZN(n10894) );
  NAND2X0 U14653 ( .IN1(g4674), .IN2(n13907), .QN(n10900) );
  NAND3X0 U14654 ( .IN1(n13887), .IN2(g4743), .IN3(n9254), .QN(n13907) );
  INVX0 U14655 ( .INP(n9264), .ZN(n9254) );
  NAND2X0 U14656 ( .IN1(n5518), .IN2(g4785), .QN(n9264) );
  NAND2X0 U14657 ( .IN1(n13908), .IN2(n13909), .QN(g28083) );
  NAND2X0 U14658 ( .IN1(n13910), .IN2(n9752), .QN(n13909) );
  INVX0 U14659 ( .INP(n10174), .ZN(n9752) );
  NAND2X0 U14660 ( .IN1(n13879), .IN2(n9256), .QN(n10174) );
  NOR2X0 U14661 ( .IN1(n5361), .IN2(n5518), .QN(n9256) );
  INVX0 U14662 ( .INP(n9239), .ZN(n13879) );
  NAND3X0 U14663 ( .IN1(g4776), .IN2(n8595), .IN3(g4793), .QN(n9239) );
  NOR2X0 U14664 ( .IN1(n8956), .IN2(n13911), .QN(n13910) );
  NOR2X0 U14665 ( .IN1(n4708), .IN2(g4704), .QN(n13911) );
  NAND2X0 U14666 ( .IN1(n10917), .IN2(g4704), .QN(n13908) );
  NOR2X0 U14667 ( .IN1(g33959), .IN2(n8942), .QN(n10917) );
  INVX0 U14668 ( .INP(n8570), .ZN(g33959) );
  NAND2X0 U14669 ( .IN1(g4646), .IN2(n13912), .QN(n8570) );
  NAND3X0 U14670 ( .IN1(n9257), .IN2(g4698), .IN3(n13887), .QN(n13912) );
  NOR4X0 U14671 ( .IN1(g4793), .IN2(n10296), .IN3(n5707), .IN4(test_so29), 
        .QN(n13887) );
  NAND3X0 U14672 ( .IN1(g4669), .IN2(g4659), .IN3(test_so19), .QN(n10296) );
  NOR2X0 U14673 ( .IN1(g4709), .IN2(g4785), .QN(n9257) );
  NAND2X0 U14674 ( .IN1(n13913), .IN2(n13914), .QN(g28082) );
  NAND2X0 U14675 ( .IN1(n13915), .IN2(g4521), .QN(n13914) );
  NAND2X0 U14676 ( .IN1(n13916), .IN2(n8920), .QN(n13915) );
  XOR2X1 U14677 ( .IN1(g4527), .IN2(n13917), .Q(n13916) );
  NAND3X0 U14678 ( .IN1(n9637), .IN2(n8870), .IN3(n5752), .QN(n13913) );
  INVX0 U14679 ( .INP(n13918), .ZN(n9637) );
  NAND3X0 U14680 ( .IN1(n13919), .IN2(n13920), .IN3(n13921), .QN(g28074) );
  NAND2X0 U14681 ( .IN1(n8997), .IN2(g4119), .QN(n13921) );
  NAND3X0 U14682 ( .IN1(n8895), .IN2(g4122), .IN3(n13922), .QN(n13920) );
  INVX0 U14683 ( .INP(n4714), .ZN(n13922) );
  NAND2X0 U14684 ( .IN1(n4714), .IN2(n4721), .QN(n13919) );
  NAND3X0 U14685 ( .IN1(n13923), .IN2(n13924), .IN3(n13925), .QN(g28073) );
  NAND2X0 U14686 ( .IN1(n13926), .IN2(n4721), .QN(n13925) );
  INVX0 U14687 ( .INP(n13927), .ZN(n13926) );
  NAND3X0 U14688 ( .IN1(n13927), .IN2(g4119), .IN3(n8888), .QN(n13924) );
  NAND3X0 U14689 ( .IN1(n5416), .IN2(g4057), .IN3(n4722), .QN(n13927) );
  NAND2X0 U14690 ( .IN1(n8997), .IN2(g4116), .QN(n13923) );
  NAND3X0 U14691 ( .IN1(n13928), .IN2(n13929), .IN3(n13930), .QN(g28072) );
  NAND2X0 U14692 ( .IN1(n13931), .IN2(n4721), .QN(n13930) );
  INVX0 U14693 ( .INP(n13932), .ZN(n13931) );
  NAND3X0 U14694 ( .IN1(n13932), .IN2(g4116), .IN3(n8887), .QN(n13929) );
  NAND3X0 U14695 ( .IN1(n5711), .IN2(g4064), .IN3(n4722), .QN(n13932) );
  INVX0 U14696 ( .INP(n13933), .ZN(n4722) );
  NAND2X0 U14697 ( .IN1(n8997), .IN2(g4112), .QN(n13928) );
  NAND2X0 U14698 ( .IN1(n13934), .IN2(n13935), .QN(g28071) );
  NAND2X0 U14699 ( .IN1(n13936), .IN2(g4112), .QN(n13935) );
  INVX0 U14700 ( .INP(n13937), .ZN(n13934) );
  NOR2X0 U14701 ( .IN1(n13936), .IN2(n8449), .QN(n13937) );
  NOR2X0 U14702 ( .IN1(n13938), .IN2(n8941), .QN(n13936) );
  NOR3X0 U14703 ( .IN1(g4057), .IN2(g4064), .IN3(n13933), .QN(n13938) );
  NAND4X0 U14704 ( .IN1(n8163), .IN2(n5612), .IN3(n13939), .IN4(n5350), .QN(
        n13933) );
  NOR2X0 U14705 ( .IN1(test_so11), .IN2(n10053), .QN(n13939) );
  NAND2X0 U14706 ( .IN1(n5340), .IN2(n5480), .QN(n10053) );
  NAND4X0 U14707 ( .IN1(n13940), .IN2(n11495), .IN3(n13941), .IN4(n13942), 
        .QN(g28070) );
  NAND3X0 U14708 ( .IN1(test_so11), .IN2(n13168), .IN3(n8887), .QN(n13942) );
  NAND2X0 U14709 ( .IN1(n8997), .IN2(g4082), .QN(n13941) );
  INVX0 U14710 ( .INP(n13943), .ZN(n13940) );
  NOR2X0 U14711 ( .IN1(n13168), .IN2(test_so11), .QN(n13943) );
  NAND2X0 U14712 ( .IN1(n13944), .IN2(g4082), .QN(n13168) );
  NAND3X0 U14713 ( .IN1(n13945), .IN2(n13946), .IN3(n13947), .QN(g28069) );
  NAND2X0 U14714 ( .IN1(n10944), .IN2(g4035), .QN(n13947) );
  NOR2X0 U14715 ( .IN1(n10933), .IN2(n8941), .QN(n10944) );
  NAND2X0 U14716 ( .IN1(n8997), .IN2(g3965), .QN(n13946) );
  NAND3X0 U14717 ( .IN1(n10933), .IN2(n13200), .IN3(n8887), .QN(n13945) );
  NAND2X0 U14718 ( .IN1(n13948), .IN2(n13949), .QN(n13200) );
  NAND2X0 U14719 ( .IN1(n5530), .IN2(n13950), .QN(n13949) );
  NAND4X0 U14720 ( .IN1(n13951), .IN2(n13952), .IN3(n13953), .IN4(n13954), 
        .QN(n13950) );
  NOR3X0 U14721 ( .IN1(n13955), .IN2(n13956), .IN3(n13957), .QN(n13954) );
  NOR2X0 U14722 ( .IN1(n5435), .IN2(n13958), .QN(n13957) );
  NOR2X0 U14723 ( .IN1(n13959), .IN2(n13960), .QN(n13958) );
  NOR2X0 U14724 ( .IN1(n8330), .IN2(n13961), .QN(n13959) );
  INVX0 U14725 ( .INP(n13962), .ZN(n13956) );
  NAND2X0 U14726 ( .IN1(n13963), .IN2(n5435), .QN(n13962) );
  NOR2X0 U14727 ( .IN1(n13964), .IN2(n13965), .QN(n13955) );
  NOR2X0 U14728 ( .IN1(n13966), .IN2(n13967), .QN(n13964) );
  NOR2X0 U14729 ( .IN1(n8387), .IN2(n8386), .QN(n13967) );
  NOR2X0 U14730 ( .IN1(n8385), .IN2(n8384), .QN(n13966) );
  NAND2X0 U14731 ( .IN1(n10940), .IN2(n13968), .QN(n13953) );
  NAND2X0 U14732 ( .IN1(n13969), .IN2(n13970), .QN(n13968) );
  NAND2X0 U14733 ( .IN1(g4031), .IN2(g3913), .QN(n13970) );
  NAND2X0 U14734 ( .IN1(g14518), .IN2(g3901), .QN(n13969) );
  NAND3X0 U14735 ( .IN1(g13906), .IN2(g3941), .IN3(n13846), .QN(n13952) );
  NAND3X0 U14736 ( .IN1(g16955), .IN2(g3925), .IN3(n10064), .QN(n13951) );
  NAND2X0 U14737 ( .IN1(n13971), .IN2(g4040), .QN(n13948) );
  NAND4X0 U14738 ( .IN1(n13972), .IN2(n13973), .IN3(n13974), .IN4(n13975), 
        .QN(n13971) );
  NOR3X0 U14739 ( .IN1(n13976), .IN2(n13977), .IN3(n13978), .QN(n13975) );
  NOR2X0 U14740 ( .IN1(n5435), .IN2(n13979), .QN(n13978) );
  NOR2X0 U14741 ( .IN1(n13980), .IN2(n13963), .QN(n13979) );
  NAND3X0 U14742 ( .IN1(n13981), .IN2(n13982), .IN3(n13983), .QN(n13963) );
  NAND3X0 U14743 ( .IN1(g13966), .IN2(g3921), .IN3(n10940), .QN(n13983) );
  NAND3X0 U14744 ( .IN1(g16659), .IN2(g3953), .IN3(n13846), .QN(n13982) );
  NAND3X0 U14745 ( .IN1(g16775), .IN2(g3937), .IN3(n10064), .QN(n13981) );
  INVX0 U14746 ( .INP(n13961), .ZN(n10064) );
  NOR2X0 U14747 ( .IN1(n8220), .IN2(n13965), .QN(n13980) );
  INVX0 U14748 ( .INP(n10935), .ZN(n13965) );
  INVX0 U14749 ( .INP(n13984), .ZN(n13977) );
  NAND2X0 U14750 ( .IN1(n13960), .IN2(n5435), .QN(n13984) );
  NAND3X0 U14751 ( .IN1(n13985), .IN2(n13986), .IN3(n13987), .QN(n13960) );
  NAND3X0 U14752 ( .IN1(g3945), .IN2(g16775), .IN3(n10935), .QN(n13987) );
  NAND3X0 U14753 ( .IN1(g13966), .IN2(g3929), .IN3(n13846), .QN(n13986) );
  NAND3X0 U14754 ( .IN1(g3961), .IN2(g16659), .IN3(n10940), .QN(n13985) );
  NOR2X0 U14755 ( .IN1(n13988), .IN2(n13961), .QN(n13976) );
  NAND2X0 U14756 ( .IN1(g4054), .IN2(g3990), .QN(n13961) );
  NOR2X0 U14757 ( .IN1(n13989), .IN2(n13990), .QN(n13988) );
  NOR2X0 U14758 ( .IN1(n8384), .IN2(n8618), .QN(n13990) );
  NOR2X0 U14759 ( .IN1(n8386), .IN2(n8218), .QN(n13989) );
  NAND2X0 U14760 ( .IN1(n13846), .IN2(n13991), .QN(n13974) );
  NAND2X0 U14761 ( .IN1(n13992), .IN2(n13993), .QN(n13991) );
  NAND2X0 U14762 ( .IN1(g3897), .IN2(g4031), .QN(n13993) );
  NAND2X0 U14763 ( .IN1(test_so24), .IN2(g14518), .QN(n13992) );
  NOR2X0 U14764 ( .IN1(g4054), .IN2(g3990), .QN(n13846) );
  NAND3X0 U14765 ( .IN1(g13906), .IN2(g3933), .IN3(n10940), .QN(n13973) );
  NOR2X0 U14766 ( .IN1(g4054), .IN2(n5594), .QN(n10940) );
  NAND3X0 U14767 ( .IN1(g3917), .IN2(g16955), .IN3(n10935), .QN(n13972) );
  NOR2X0 U14768 ( .IN1(g3990), .IN2(n5395), .QN(n10935) );
  INVX0 U14769 ( .INP(n10939), .ZN(n10933) );
  NAND2X0 U14770 ( .IN1(g4878), .IN2(n13994), .QN(n10939) );
  NAND3X0 U14771 ( .IN1(n13875), .IN2(g4955), .IN3(n9293), .QN(n13994) );
  NOR2X0 U14772 ( .IN1(n5360), .IN2(n5517), .QN(n9293) );
  NAND3X0 U14773 ( .IN1(n13995), .IN2(n13996), .IN3(n13997), .QN(g28066) );
  NAND2X0 U14774 ( .IN1(n10960), .IN2(g3684), .QN(n13997) );
  NOR2X0 U14775 ( .IN1(n10949), .IN2(n8940), .QN(n10960) );
  NAND2X0 U14776 ( .IN1(n8997), .IN2(g3614), .QN(n13996) );
  NAND3X0 U14777 ( .IN1(n10949), .IN2(n13232), .IN3(n8887), .QN(n13995) );
  NAND2X0 U14778 ( .IN1(n13998), .IN2(n13999), .QN(n13232) );
  NAND2X0 U14779 ( .IN1(n5532), .IN2(n14000), .QN(n13999) );
  NAND4X0 U14780 ( .IN1(n14001), .IN2(n14002), .IN3(n14003), .IN4(n14004), 
        .QN(n14000) );
  NOR3X0 U14781 ( .IN1(n14005), .IN2(n14006), .IN3(n14007), .QN(n14004) );
  NOR2X0 U14782 ( .IN1(n5433), .IN2(n14008), .QN(n14007) );
  NOR2X0 U14783 ( .IN1(n14009), .IN2(n14010), .QN(n14008) );
  NOR2X0 U14784 ( .IN1(n8336), .IN2(n14011), .QN(n14009) );
  INVX0 U14785 ( .INP(n14012), .ZN(n14006) );
  NAND2X0 U14786 ( .IN1(n14013), .IN2(n5433), .QN(n14012) );
  NOR2X0 U14787 ( .IN1(n14014), .IN2(n14015), .QN(n14005) );
  NOR2X0 U14788 ( .IN1(n14016), .IN2(n14017), .QN(n14014) );
  NOR2X0 U14789 ( .IN1(n8397), .IN2(n8396), .QN(n14017) );
  NOR2X0 U14790 ( .IN1(n8395), .IN2(n8394), .QN(n14016) );
  NAND2X0 U14791 ( .IN1(n10956), .IN2(n14018), .QN(n14003) );
  NAND2X0 U14792 ( .IN1(n14019), .IN2(n14020), .QN(n14018) );
  NAND2X0 U14793 ( .IN1(g3680), .IN2(g3562), .QN(n14020) );
  NAND2X0 U14794 ( .IN1(g14451), .IN2(g3550), .QN(n14019) );
  NAND3X0 U14795 ( .IN1(test_so26), .IN2(g3590), .IN3(n13856), .QN(n14002) );
  NAND3X0 U14796 ( .IN1(g16924), .IN2(g3574), .IN3(n10069), .QN(n14001) );
  NAND2X0 U14797 ( .IN1(n14021), .IN2(g3689), .QN(n13998) );
  NAND4X0 U14798 ( .IN1(n14022), .IN2(n14023), .IN3(n14024), .IN4(n14025), 
        .QN(n14021) );
  NOR3X0 U14799 ( .IN1(n14026), .IN2(n14027), .IN3(n14028), .QN(n14025) );
  NOR2X0 U14800 ( .IN1(n5433), .IN2(n14029), .QN(n14028) );
  NOR2X0 U14801 ( .IN1(n14030), .IN2(n14013), .QN(n14029) );
  NAND3X0 U14802 ( .IN1(n14031), .IN2(n14032), .IN3(n14033), .QN(n14013) );
  NAND3X0 U14803 ( .IN1(g13926), .IN2(g3570), .IN3(n10956), .QN(n14033) );
  NAND3X0 U14804 ( .IN1(test_so43), .IN2(g16627), .IN3(n13856), .QN(n14032) );
  NAND3X0 U14805 ( .IN1(g16744), .IN2(g3586), .IN3(n10069), .QN(n14031) );
  INVX0 U14806 ( .INP(n14011), .ZN(n10069) );
  NOR2X0 U14807 ( .IN1(n8207), .IN2(n14015), .QN(n14030) );
  INVX0 U14808 ( .INP(n10951), .ZN(n14015) );
  INVX0 U14809 ( .INP(n14034), .ZN(n14027) );
  NAND2X0 U14810 ( .IN1(n14010), .IN2(n5433), .QN(n14034) );
  NAND3X0 U14811 ( .IN1(n14035), .IN2(n14036), .IN3(n14037), .QN(n14010) );
  NAND3X0 U14812 ( .IN1(g3594), .IN2(g16744), .IN3(n10951), .QN(n14037) );
  NAND3X0 U14813 ( .IN1(g13926), .IN2(g3578), .IN3(n13856), .QN(n14036) );
  NAND3X0 U14814 ( .IN1(g3610), .IN2(g16627), .IN3(n10956), .QN(n14035) );
  NOR2X0 U14815 ( .IN1(n14038), .IN2(n14011), .QN(n14026) );
  NAND2X0 U14816 ( .IN1(g3703), .IN2(g3639), .QN(n14011) );
  NOR2X0 U14817 ( .IN1(n14039), .IN2(n14040), .QN(n14038) );
  NOR2X0 U14818 ( .IN1(n8394), .IN2(n8205), .QN(n14040) );
  NOR2X0 U14819 ( .IN1(n8396), .IN2(n8204), .QN(n14039) );
  NAND2X0 U14820 ( .IN1(n13856), .IN2(n14041), .QN(n14024) );
  NAND2X0 U14821 ( .IN1(n14042), .IN2(n14043), .QN(n14041) );
  NAND2X0 U14822 ( .IN1(g3546), .IN2(g3680), .QN(n14043) );
  NAND2X0 U14823 ( .IN1(g3538), .IN2(g14451), .QN(n14042) );
  NOR2X0 U14824 ( .IN1(g3703), .IN2(g3639), .QN(n13856) );
  NAND3X0 U14825 ( .IN1(n10956), .IN2(g3582), .IN3(test_so26), .QN(n14023) );
  NOR2X0 U14826 ( .IN1(g3703), .IN2(n5591), .QN(n10956) );
  NAND3X0 U14827 ( .IN1(g3566), .IN2(g16924), .IN3(n10951), .QN(n14022) );
  NOR2X0 U14828 ( .IN1(g3639), .IN2(n5399), .QN(n10951) );
  INVX0 U14829 ( .INP(n10955), .ZN(n10949) );
  NAND2X0 U14830 ( .IN1(g4871), .IN2(n14044), .QN(n10955) );
  NAND3X0 U14831 ( .IN1(n13875), .IN2(g4944), .IN3(n9296), .QN(n14044) );
  INVX0 U14832 ( .INP(n9304), .ZN(n9296) );
  NAND2X0 U14833 ( .IN1(n5360), .IN2(g4899), .QN(n9304) );
  NAND3X0 U14834 ( .IN1(n14045), .IN2(n14046), .IN3(n14047), .QN(g28063) );
  NAND2X0 U14835 ( .IN1(n10975), .IN2(g3333), .QN(n14047) );
  NOR2X0 U14836 ( .IN1(n10969), .IN2(n8940), .QN(n10975) );
  NAND2X0 U14837 ( .IN1(n8997), .IN2(g3263), .QN(n14046) );
  NAND3X0 U14838 ( .IN1(n10969), .IN2(n13265), .IN3(n8887), .QN(n14045) );
  NAND2X0 U14839 ( .IN1(n14048), .IN2(n14049), .QN(n13265) );
  NAND2X0 U14840 ( .IN1(n5527), .IN2(n14050), .QN(n14049) );
  NAND4X0 U14841 ( .IN1(n14051), .IN2(n14052), .IN3(n14053), .IN4(n14054), 
        .QN(n14050) );
  NOR3X0 U14842 ( .IN1(n14055), .IN2(n14056), .IN3(n14057), .QN(n14054) );
  NOR2X0 U14843 ( .IN1(n5436), .IN2(n14058), .QN(n14057) );
  NOR2X0 U14844 ( .IN1(n14059), .IN2(n14060), .QN(n14058) );
  NOR2X0 U14845 ( .IN1(n8318), .IN2(n14061), .QN(n14059) );
  INVX0 U14846 ( .INP(n14062), .ZN(n14056) );
  NAND2X0 U14847 ( .IN1(n14063), .IN2(n5436), .QN(n14062) );
  NOR2X0 U14848 ( .IN1(n14064), .IN2(n10971), .QN(n14055) );
  NOR2X0 U14849 ( .IN1(n14065), .IN2(n14066), .QN(n14064) );
  NOR2X0 U14850 ( .IN1(n8368), .IN2(n8367), .QN(n14066) );
  NOR2X0 U14851 ( .IN1(n8366), .IN2(n8365), .QN(n14065) );
  NAND2X0 U14852 ( .IN1(n13867), .IN2(n14067), .QN(n14053) );
  NAND2X0 U14853 ( .IN1(n14068), .IN2(n14069), .QN(n14067) );
  NAND2X0 U14854 ( .IN1(test_so91), .IN2(g3211), .QN(n14069) );
  NAND2X0 U14855 ( .IN1(g14421), .IN2(g3199), .QN(n14068) );
  NAND3X0 U14856 ( .IN1(g13865), .IN2(g3239), .IN3(n13868), .QN(n14052) );
  NAND3X0 U14857 ( .IN1(g16874), .IN2(g3223), .IN3(n10077), .QN(n14051) );
  NAND2X0 U14858 ( .IN1(n14070), .IN2(g3338), .QN(n14048) );
  NAND4X0 U14859 ( .IN1(n14071), .IN2(n14072), .IN3(n14073), .IN4(n14074), 
        .QN(n14070) );
  NOR3X0 U14860 ( .IN1(n14075), .IN2(n14076), .IN3(n14077), .QN(n14074) );
  NOR2X0 U14861 ( .IN1(n5436), .IN2(n14078), .QN(n14077) );
  NOR2X0 U14862 ( .IN1(n14079), .IN2(n14063), .QN(n14078) );
  NAND3X0 U14863 ( .IN1(n14080), .IN2(n14081), .IN3(n14082), .QN(n14063) );
  NAND3X0 U14864 ( .IN1(g13895), .IN2(g3219), .IN3(n13867), .QN(n14082) );
  NAND3X0 U14865 ( .IN1(g16603), .IN2(g3251), .IN3(n13868), .QN(n14081) );
  NAND3X0 U14866 ( .IN1(g16718), .IN2(g3235), .IN3(n10077), .QN(n14080) );
  INVX0 U14867 ( .INP(n14061), .ZN(n10077) );
  NOR2X0 U14868 ( .IN1(n8196), .IN2(n10971), .QN(n14079) );
  INVX0 U14869 ( .INP(n14083), .ZN(n14076) );
  NAND2X0 U14870 ( .IN1(n14060), .IN2(n5436), .QN(n14083) );
  NAND3X0 U14871 ( .IN1(n14084), .IN2(n14085), .IN3(n14086), .QN(n14060) );
  NAND3X0 U14872 ( .IN1(g3243), .IN2(g16718), .IN3(n13869), .QN(n14086) );
  NAND3X0 U14873 ( .IN1(g13895), .IN2(g3227), .IN3(n13868), .QN(n14085) );
  NAND3X0 U14874 ( .IN1(test_so84), .IN2(g16603), .IN3(n13867), .QN(n14084) );
  NOR2X0 U14875 ( .IN1(n14087), .IN2(n14061), .QN(n14075) );
  NAND2X0 U14876 ( .IN1(g3288), .IN2(g3352), .QN(n14061) );
  NOR2X0 U14877 ( .IN1(n14088), .IN2(n14089), .QN(n14087) );
  NOR2X0 U14878 ( .IN1(n8365), .IN2(n8194), .QN(n14089) );
  NOR2X0 U14879 ( .IN1(n8367), .IN2(n8193), .QN(n14088) );
  NAND2X0 U14880 ( .IN1(n13868), .IN2(n14090), .QN(n14073) );
  NAND2X0 U14881 ( .IN1(n14091), .IN2(n14092), .QN(n14090) );
  NAND2X0 U14882 ( .IN1(g3187), .IN2(g14421), .QN(n14092) );
  NAND2X0 U14883 ( .IN1(test_so91), .IN2(test_so88), .QN(n14091) );
  NOR2X0 U14884 ( .IN1(g3352), .IN2(g3288), .QN(n13868) );
  NAND3X0 U14885 ( .IN1(g13865), .IN2(g3231), .IN3(n13867), .QN(n14072) );
  NOR2X0 U14886 ( .IN1(g3352), .IN2(n5400), .QN(n13867) );
  NAND3X0 U14887 ( .IN1(g3215), .IN2(g16874), .IN3(n13869), .QN(n14071) );
  INVX0 U14888 ( .INP(n10971), .ZN(n13869) );
  NAND2X0 U14889 ( .IN1(n5400), .IN2(g3352), .QN(n10971) );
  INVX0 U14890 ( .INP(n10966), .ZN(n10969) );
  NAND2X0 U14891 ( .IN1(g4864), .IN2(n14093), .QN(n10966) );
  NAND3X0 U14892 ( .IN1(n13875), .IN2(g4933), .IN3(n9297), .QN(n14093) );
  INVX0 U14893 ( .INP(n9305), .ZN(n9297) );
  NAND2X0 U14894 ( .IN1(n5517), .IN2(g4975), .QN(n9305) );
  INVX0 U14895 ( .INP(n14094), .ZN(n13875) );
  NAND4X0 U14896 ( .IN1(n5367), .IN2(n10268), .IN3(g4966), .IN4(n8587), .QN(
        n14094) );
  NOR3X0 U14897 ( .IN1(n8556), .IN2(n8557), .IN3(n8555), .QN(n10268) );
  NAND4X0 U14898 ( .IN1(n14095), .IN2(n9200), .IN3(n14096), .IN4(n14097), .QN(
        g28060) );
  NAND3X0 U14899 ( .IN1(n13270), .IN2(g2729), .IN3(n8887), .QN(n14097) );
  NAND2X0 U14900 ( .IN1(n8996), .IN2(g2724), .QN(n14096) );
  NAND2X0 U14901 ( .IN1(n14098), .IN2(n8186), .QN(n14095) );
  INVX0 U14902 ( .INP(n13270), .ZN(n14098) );
  NAND2X0 U14903 ( .IN1(n12644), .IN2(g2724), .QN(n13270) );
  NAND3X0 U14904 ( .IN1(n14099), .IN2(n14100), .IN3(n14101), .QN(g28059) );
  NAND2X0 U14905 ( .IN1(n8996), .IN2(g1351), .QN(n14101) );
  NAND3X0 U14906 ( .IN1(n11741), .IN2(n8165), .IN3(n12942), .QN(n14100) );
  NOR2X0 U14907 ( .IN1(n12944), .IN2(n8939), .QN(n11741) );
  NAND4X0 U14908 ( .IN1(n5466), .IN2(n14102), .IN3(n14103), .IN4(n14104), .QN(
        n12944) );
  NAND2X0 U14909 ( .IN1(n14105), .IN2(n5322), .QN(n14104) );
  NAND3X0 U14910 ( .IN1(n14106), .IN2(g1351), .IN3(n14107), .QN(n14103) );
  NAND2X0 U14911 ( .IN1(n4798), .IN2(n14108), .QN(n14099) );
  INVX0 U14912 ( .INP(n12942), .ZN(n14108) );
  NAND3X0 U14913 ( .IN1(n14109), .IN2(n14110), .IN3(n14111), .QN(g28058) );
  NAND2X0 U14914 ( .IN1(test_so77), .IN2(n8953), .QN(n14111) );
  NAND3X0 U14915 ( .IN1(n11311), .IN2(n14112), .IN3(g1252), .QN(n14110) );
  INVX0 U14916 ( .INP(n4490), .ZN(n14112) );
  NAND2X0 U14917 ( .IN1(n4490), .IN2(n5554), .QN(n14109) );
  NAND3X0 U14918 ( .IN1(n14113), .IN2(n14114), .IN3(n14115), .QN(g28057) );
  NAND2X0 U14919 ( .IN1(n8996), .IN2(g1008), .QN(n14115) );
  NAND3X0 U14920 ( .IN1(n11754), .IN2(n8166), .IN3(n12977), .QN(n14114) );
  INVX0 U14921 ( .INP(n14116), .ZN(n11754) );
  NAND2X0 U14922 ( .IN1(n11319), .IN2(n8919), .QN(n14116) );
  NOR4X0 U14923 ( .IN1(n14117), .IN2(test_so20), .IN3(n14118), .IN4(n14119), 
        .QN(n11319) );
  NOR2X0 U14924 ( .IN1(n14120), .IN2(n14121), .QN(n14119) );
  NOR2X0 U14925 ( .IN1(g1008), .IN2(n14122), .QN(n14118) );
  NAND2X0 U14926 ( .IN1(n4805), .IN2(n14123), .QN(n14113) );
  NAND3X0 U14927 ( .IN1(n14124), .IN2(n14125), .IN3(n14126), .QN(g28056) );
  NAND2X0 U14928 ( .IN1(n8996), .IN2(g936), .QN(n14126) );
  NAND3X0 U14929 ( .IN1(n11325), .IN2(n14127), .IN3(g907), .QN(n14125) );
  INVX0 U14930 ( .INP(n4514), .ZN(n14127) );
  NAND2X0 U14931 ( .IN1(n4514), .IN2(n5555), .QN(n14124) );
  NAND3X0 U14932 ( .IN1(n14128), .IN2(n14129), .IN3(n14130), .QN(g28055) );
  NAND2X0 U14933 ( .IN1(n8996), .IN2(g822), .QN(n14130) );
  NAND3X0 U14934 ( .IN1(n4518), .IN2(n14131), .IN3(g827), .QN(n14129) );
  INVX0 U14935 ( .INP(n4519), .ZN(n14131) );
  NAND3X0 U14936 ( .IN1(n4519), .IN2(n13521), .IN3(n5728), .QN(n14128) );
  NAND2X0 U14937 ( .IN1(n14132), .IN2(n14133), .QN(g28054) );
  NAND2X0 U14938 ( .IN1(n14134), .IN2(g728), .QN(n14133) );
  NAND2X0 U14939 ( .IN1(n14135), .IN2(g661), .QN(n14132) );
  NAND3X0 U14940 ( .IN1(n14136), .IN2(n14137), .IN3(n14138), .QN(g28053) );
  NAND2X0 U14941 ( .IN1(n8996), .IN2(g681), .QN(n14138) );
  INVX0 U14942 ( .INP(n14139), .ZN(n14137) );
  NAND2X0 U14943 ( .IN1(n13558), .IN2(test_so87), .QN(n14136) );
  NAND2X0 U14944 ( .IN1(n14140), .IN2(n14141), .QN(g28052) );
  NAND2X0 U14945 ( .IN1(n14134), .IN2(g661), .QN(n14141) );
  NAND2X0 U14946 ( .IN1(n14135), .IN2(g718), .QN(n14140) );
  NAND2X0 U14947 ( .IN1(n14142), .IN2(n14143), .QN(g28051) );
  NAND2X0 U14948 ( .IN1(n14134), .IN2(g718), .QN(n14143) );
  NAND2X0 U14949 ( .IN1(n14135), .IN2(g655), .QN(n14142) );
  NAND2X0 U14950 ( .IN1(n14144), .IN2(n14145), .QN(g28050) );
  NAND2X0 U14951 ( .IN1(n14134), .IN2(g655), .QN(n14145) );
  NAND2X0 U14952 ( .IN1(n14135), .IN2(g650), .QN(n14144) );
  NAND3X0 U14953 ( .IN1(n14146), .IN2(n14147), .IN3(n14148), .QN(g28049) );
  NAND2X0 U14954 ( .IN1(test_so87), .IN2(n8956), .QN(n14148) );
  NAND2X0 U14955 ( .IN1(n14139), .IN2(g681), .QN(n14147) );
  NAND2X0 U14956 ( .IN1(n14134), .IN2(g650), .QN(n14146) );
  NAND3X0 U14957 ( .IN1(n14149), .IN2(n14150), .IN3(n14151), .QN(g28048) );
  NAND2X0 U14958 ( .IN1(n8996), .IN2(g29212), .QN(n14151) );
  NAND2X0 U14959 ( .IN1(n14152), .IN2(g691), .QN(n14150) );
  NAND2X0 U14960 ( .IN1(n14153), .IN2(n14154), .QN(n14152) );
  NAND3X0 U14961 ( .IN1(g703), .IN2(n8603), .IN3(n8887), .QN(n14154) );
  NAND2X0 U14962 ( .IN1(n14155), .IN2(n14156), .QN(n14149) );
  INVX0 U14963 ( .INP(n4819), .ZN(n14156) );
  NAND4X0 U14964 ( .IN1(n5520), .IN2(n5112), .IN3(n14157), .IN4(g703), .QN(
        n4819) );
  INVX0 U14965 ( .INP(n13540), .ZN(n14157) );
  NAND4X0 U14966 ( .IN1(n14158), .IN2(test_so87), .IN3(n8183), .IN4(n8182), 
        .QN(n13540) );
  XOR2X1 U14967 ( .IN1(g661), .IN2(n8192), .Q(n14158) );
  NAND2X0 U14968 ( .IN1(n14159), .IN2(n14160), .QN(g28047) );
  NAND2X0 U14969 ( .IN1(n14134), .IN2(g681), .QN(n14160) );
  NAND2X0 U14970 ( .IN1(n14135), .IN2(g645), .QN(n14159) );
  NAND2X0 U14971 ( .IN1(n14161), .IN2(n14162), .QN(g28046) );
  NAND2X0 U14972 ( .IN1(n14139), .IN2(g446), .QN(n14162) );
  NOR2X0 U14973 ( .IN1(n14163), .IN2(n8938), .QN(n14139) );
  NAND2X0 U14974 ( .IN1(n14134), .IN2(g645), .QN(n14161) );
  INVX0 U14975 ( .INP(n14135), .ZN(n14134) );
  NAND2X0 U14976 ( .IN1(n14163), .IN2(n8919), .QN(n14135) );
  NAND4X0 U14977 ( .IN1(n8539), .IN2(n14164), .IN3(n14165), .IN4(n14166), .QN(
        n14163) );
  NAND2X0 U14978 ( .IN1(n14167), .IN2(g691), .QN(n14166) );
  INVX0 U14979 ( .INP(n14168), .ZN(n14167) );
  NAND2X0 U14980 ( .IN1(n5520), .IN2(n14169), .QN(n14165) );
  NAND3X0 U14981 ( .IN1(n5629), .IN2(g417), .IN3(n8507), .QN(n14169) );
  NAND3X0 U14982 ( .IN1(n14170), .IN2(n14171), .IN3(n14172), .QN(g28045) );
  NAND2X0 U14983 ( .IN1(n8995), .IN2(g568), .QN(n14172) );
  NAND3X0 U14984 ( .IN1(n2421), .IN2(n14173), .IN3(g572), .QN(n14171) );
  INVX0 U14985 ( .INP(n4537), .ZN(n14173) );
  NAND2X0 U14986 ( .IN1(n4537), .IN2(n5337), .QN(n14170) );
  NAND2X0 U14987 ( .IN1(n14174), .IN2(n14175), .QN(g28044) );
  NAND2X0 U14988 ( .IN1(n8995), .IN2(g528), .QN(n14175) );
  NAND2X0 U14989 ( .IN1(n14176), .IN2(n8919), .QN(n14174) );
  NAND2X0 U14990 ( .IN1(n14177), .IN2(n13551), .QN(n14176) );
  XOR2X1 U14991 ( .IN1(g482), .IN2(n13554), .Q(n14177) );
  NAND2X0 U14992 ( .IN1(n14178), .IN2(n14179), .QN(n13554) );
  NAND2X0 U14993 ( .IN1(n5327), .IN2(n14180), .QN(n14179) );
  NAND2X0 U14994 ( .IN1(n14181), .IN2(n14182), .QN(g28043) );
  NAND2X0 U14995 ( .IN1(n8568), .IN2(n8607), .QN(n14182) );
  NOR2X0 U14996 ( .IN1(n11891), .IN2(n8937), .QN(n8568) );
  NAND4X0 U14997 ( .IN1(n14183), .IN2(n12995), .IN3(n9328), .IN4(g691), .QN(
        n11891) );
  NAND2X0 U14998 ( .IN1(n5627), .IN2(n14184), .QN(n9328) );
  NAND4X0 U14999 ( .IN1(n8308), .IN2(n6008), .IN3(n8309), .IN4(n14185), .QN(
        n14184) );
  NOR4X0 U15000 ( .IN1(n8189), .IN2(n8188), .IN3(n8187), .IN4(g225), .QN(
        n14185) );
  NAND4X0 U15001 ( .IN1(n14186), .IN2(n14187), .IN3(n14188), .IN4(n14189), 
        .QN(n12995) );
  NAND3X0 U15002 ( .IN1(g655), .IN2(g753), .IN3(g718), .QN(n14189) );
  NAND3X0 U15003 ( .IN1(n8551), .IN2(n8550), .IN3(n8552), .QN(n14188) );
  NAND2X0 U15004 ( .IN1(g807), .IN2(g554), .QN(n14187) );
  NAND2X0 U15005 ( .IN1(n9329), .IN2(g278), .QN(n14183) );
  NAND4X0 U15006 ( .IN1(n8188), .IN2(n8187), .IN3(n8189), .IN4(n14190), .QN(
        n9329) );
  NOR4X0 U15007 ( .IN1(n8309), .IN2(n8308), .IN3(n6008), .IN4(n5597), .QN(
        n14190) );
  NAND2X0 U15008 ( .IN1(n8995), .IN2(g278), .QN(n14181) );
  NAND3X0 U15009 ( .IN1(n5796), .IN2(n8870), .IN3(n5630), .QN(g28042) );
  NAND3X0 U15010 ( .IN1(n13513), .IN2(n8871), .IN3(n9768), .QN(g28041) );
  NAND2X0 U15011 ( .IN1(n1376), .IN2(g1536), .QN(n9768) );
  NAND2X0 U15012 ( .IN1(n4837), .IN2(g1193), .QN(n13513) );
  INVX0 U15013 ( .INP(n14191), .ZN(n4837) );
  NAND2X0 U15014 ( .IN1(n14192), .IN2(n14193), .QN(g28030) );
  NAND3X0 U15015 ( .IN1(n5861), .IN2(n14194), .IN3(n5882), .QN(n14193) );
  NAND2X0 U15016 ( .IN1(n14195), .IN2(n14196), .QN(n14194) );
  NAND2X0 U15017 ( .IN1(n14197), .IN2(n9721), .QN(n14196) );
  NAND2X0 U15018 ( .IN1(n14198), .IN2(n14199), .QN(n14197) );
  NAND3X0 U15019 ( .IN1(n5872), .IN2(n14200), .IN3(n5886), .QN(n14199) );
  NAND2X0 U15020 ( .IN1(n14201), .IN2(n14202), .QN(n14200) );
  NAND2X0 U15021 ( .IN1(n14203), .IN2(n14204), .QN(n14202) );
  NAND2X0 U15022 ( .IN1(n14205), .IN2(n14206), .QN(n14203) );
  NAND4X0 U15023 ( .IN1(n5885), .IN2(n5869), .IN3(n14207), .IN4(n14208), .QN(
        n14206) );
  NAND3X0 U15024 ( .IN1(n5874), .IN2(n14209), .IN3(n5888), .QN(n14205) );
  NAND2X0 U15025 ( .IN1(n14210), .IN2(n14211), .QN(n14209) );
  NAND3X0 U15026 ( .IN1(n5869), .IN2(n14212), .IN3(n5885), .QN(n14211) );
  NAND2X0 U15027 ( .IN1(n14213), .IN2(n14214), .QN(n14212) );
  INVX0 U15028 ( .INP(n14207), .ZN(n14214) );
  NAND2X0 U15029 ( .IN1(n14207), .IN2(n14208), .QN(n14210) );
  NAND2X0 U15030 ( .IN1(n14215), .IN2(n14204), .QN(n14198) );
  NAND2X0 U15031 ( .IN1(n9720), .IN2(n9721), .QN(n14192) );
  NAND2X0 U15032 ( .IN1(n14216), .IN2(n8919), .QN(n9721) );
  NAND2X0 U15033 ( .IN1(n5889), .IN2(n5868), .QN(n14216) );
  INVX0 U15034 ( .INP(n14195), .ZN(n9720) );
  NAND3X0 U15035 ( .IN1(n14217), .IN2(n14204), .IN3(n14215), .QN(n14195) );
  INVX0 U15036 ( .INP(n14201), .ZN(n14215) );
  NAND3X0 U15037 ( .IN1(n14207), .IN2(n14208), .IN3(n14218), .QN(n14201) );
  NAND2X0 U15038 ( .IN1(n14219), .IN2(n8919), .QN(n14218) );
  NAND4X0 U15039 ( .IN1(n5888), .IN2(n5885), .IN3(n5874), .IN4(n5869), .QN(
        n14219) );
  INVX0 U15040 ( .INP(n14213), .ZN(n14208) );
  NOR2X0 U15041 ( .IN1(n14220), .IN2(n8936), .QN(n14213) );
  NOR2X0 U15042 ( .IN1(g5831), .IN2(test_so83), .QN(n14220) );
  NAND2X0 U15043 ( .IN1(n14221), .IN2(n8919), .QN(n14207) );
  NAND2X0 U15044 ( .IN1(n5884), .IN2(n5870), .QN(n14221) );
  NAND2X0 U15045 ( .IN1(n14222), .IN2(n8919), .QN(n14204) );
  NAND2X0 U15046 ( .IN1(n5883), .IN2(n5871), .QN(n14222) );
  NAND2X0 U15047 ( .IN1(n14223), .IN2(n8919), .QN(n14217) );
  NAND2X0 U15048 ( .IN1(n5886), .IN2(n5872), .QN(n14223) );
  NAND3X0 U15049 ( .IN1(n14224), .IN2(n14225), .IN3(n11852), .QN(g26971) );
  NAND2X0 U15050 ( .IN1(n5670), .IN2(n8918), .QN(n11852) );
  NAND2X0 U15051 ( .IN1(n15223), .IN2(n8918), .QN(n14225) );
  NAND2X0 U15052 ( .IN1(n8995), .IN2(g4512), .QN(n14224) );
  NAND2X0 U15053 ( .IN1(n14226), .IN2(n14227), .QN(g26970) );
  NAND2X0 U15054 ( .IN1(n8904), .IN2(g4473), .QN(n14227) );
  NAND2X0 U15055 ( .IN1(n8995), .IN2(g4459), .QN(n14226) );
  NAND2X0 U15056 ( .IN1(n14228), .IN2(n14229), .QN(g26969) );
  NAND2X0 U15057 ( .IN1(n8995), .IN2(g4462), .QN(n14229) );
  NAND3X0 U15058 ( .IN1(n8140), .IN2(n8584), .IN3(n8887), .QN(n14228) );
  NAND2X0 U15059 ( .IN1(n14230), .IN2(n14231), .QN(g26968) );
  NAND2X0 U15060 ( .IN1(n8995), .IN2(g4558), .QN(n14230) );
  NAND2X0 U15061 ( .IN1(n14232), .IN2(n14233), .QN(g26967) );
  NAND2X0 U15062 ( .IN1(n8994), .IN2(g4561), .QN(n14232) );
  NAND2X0 U15063 ( .IN1(n14234), .IN2(n14235), .QN(g26966) );
  NAND2X0 U15064 ( .IN1(n8994), .IN2(g4555), .QN(n14234) );
  XOR2X1 U15065 ( .IN1(DFF_228_n1), .IN2(n14236), .Q(g26965) );
  NAND2X0 U15066 ( .IN1(n8904), .IN2(g10306), .QN(n14236) );
  NAND2X0 U15067 ( .IN1(n14237), .IN2(n14238), .QN(g26964) );
  NAND3X0 U15068 ( .IN1(n14239), .IN2(n14240), .IN3(n8887), .QN(n14238) );
  NAND2X0 U15069 ( .IN1(n8437), .IN2(g4521), .QN(n14240) );
  NAND2X0 U15070 ( .IN1(n5752), .IN2(n14241), .QN(n14239) );
  NAND2X0 U15071 ( .IN1(n8448), .IN2(n10305), .QN(n14241) );
  INVX0 U15072 ( .INP(n13917), .ZN(n10305) );
  NAND2X0 U15073 ( .IN1(n14242), .IN2(g4527), .QN(n14237) );
  NAND2X0 U15074 ( .IN1(n14243), .IN2(n8918), .QN(n14242) );
  NAND2X0 U15075 ( .IN1(n5752), .IN2(n13917), .QN(n14243) );
  NAND4X0 U15076 ( .IN1(test_so27), .IN2(g4483), .IN3(g4489), .IN4(g4492), 
        .QN(n13917) );
  NAND2X0 U15077 ( .IN1(n14244), .IN2(n14233), .QN(g26963) );
  NAND2X0 U15078 ( .IN1(g6750), .IN2(n8918), .QN(n14233) );
  NAND2X0 U15079 ( .IN1(n8994), .IN2(g4489), .QN(n14244) );
  NAND2X0 U15080 ( .IN1(n14231), .IN2(n14245), .QN(g26962) );
  NAND2X0 U15081 ( .IN1(test_so27), .IN2(n9051), .QN(n14245) );
  NAND2X0 U15082 ( .IN1(g6749), .IN2(n8918), .QN(n14231) );
  NAND2X0 U15083 ( .IN1(n14246), .IN2(n14235), .QN(g26961) );
  NAND2X0 U15084 ( .IN1(g6748), .IN2(n8918), .QN(n14235) );
  NAND2X0 U15085 ( .IN1(n8994), .IN2(g4483), .QN(n14246) );
  NAND2X0 U15086 ( .IN1(n14247), .IN2(n14248), .QN(g26958) );
  NAND2X0 U15087 ( .IN1(n8994), .IN2(g4455), .QN(n14248) );
  NAND2X0 U15088 ( .IN1(n14249), .IN2(n14250), .QN(g26957) );
  NAND2X0 U15089 ( .IN1(n14251), .IN2(g4434), .QN(n14250) );
  NAND2X0 U15090 ( .IN1(n14252), .IN2(n8918), .QN(n14251) );
  NAND2X0 U15091 ( .IN1(n14253), .IN2(g4392), .QN(n14252) );
  NAND2X0 U15092 ( .IN1(test_so47), .IN2(n8921), .QN(n14249) );
  NAND2X0 U15093 ( .IN1(n15225), .IN2(n14254), .QN(g26956) );
  NAND3X0 U15094 ( .IN1(n14253), .IN2(g4430), .IN3(n14255), .QN(n14254) );
  NAND2X0 U15095 ( .IN1(n14256), .IN2(n14257), .QN(g26955) );
  NAND3X0 U15096 ( .IN1(n8894), .IN2(g4392), .IN3(n14253), .QN(n14257) );
  NAND2X0 U15097 ( .IN1(n14258), .IN2(g4438), .QN(n14256) );
  NAND3X0 U15098 ( .IN1(n14259), .IN2(n14260), .IN3(n14261), .QN(g26954) );
  NAND2X0 U15099 ( .IN1(test_so47), .IN2(n9052), .QN(n14261) );
  NAND2X0 U15100 ( .IN1(n14255), .IN2(n14253), .QN(n14260) );
  INVX0 U15101 ( .INP(n14262), .ZN(n14253) );
  NAND4X0 U15102 ( .IN1(n15225), .IN2(n8442), .IN3(n14263), .IN4(DFF_1225_n1), 
        .QN(n14262) );
  NOR2X0 U15103 ( .IN1(test_so47), .IN2(g7260), .QN(n14263) );
  NAND2X0 U15104 ( .IN1(n14264), .IN2(g4438), .QN(n14259) );
  NAND2X0 U15105 ( .IN1(n14265), .IN2(n14266), .QN(g26952) );
  NAND2X0 U15106 ( .IN1(n14267), .IN2(g4430), .QN(n14266) );
  NAND2X0 U15107 ( .IN1(n8905), .IN2(g4388), .QN(n14267) );
  NAND2X0 U15108 ( .IN1(n14268), .IN2(n8907), .QN(n14265) );
  NAND2X0 U15109 ( .IN1(n14269), .IN2(n14270), .QN(n14268) );
  NAND2X0 U15110 ( .IN1(n8121), .IN2(g4388), .QN(n14270) );
  XOR2X1 U15111 ( .IN1(g4401), .IN2(n8119), .Q(n14269) );
  NAND2X0 U15112 ( .IN1(n14247), .IN2(n14271), .QN(g26950) );
  NAND2X0 U15113 ( .IN1(n8994), .IN2(g4417), .QN(n14271) );
  NAND2X0 U15114 ( .IN1(n14272), .IN2(n8906), .QN(n14247) );
  NAND2X0 U15115 ( .IN1(n14273), .IN2(n14274), .QN(n14272) );
  NAND2X0 U15116 ( .IN1(n14275), .IN2(g4392), .QN(n14274) );
  NAND2X0 U15117 ( .IN1(n14276), .IN2(n14277), .QN(g26949) );
  NAND2X0 U15118 ( .IN1(n14278), .IN2(g4401), .QN(n14277) );
  NAND2X0 U15119 ( .IN1(n14279), .IN2(n8907), .QN(n14278) );
  NAND2X0 U15120 ( .IN1(n14280), .IN2(g4392), .QN(n14279) );
  NAND2X0 U15121 ( .IN1(n8905), .IN2(g4411), .QN(n14276) );
  NAND2X0 U15122 ( .IN1(n8561), .IN2(n14281), .QN(g26948) );
  NAND3X0 U15123 ( .IN1(n14280), .IN2(g4388), .IN3(n14255), .QN(n14281) );
  NAND2X0 U15124 ( .IN1(n14282), .IN2(n14283), .QN(g26947) );
  NAND2X0 U15125 ( .IN1(n8994), .IN2(g4388), .QN(n14283) );
  NAND2X0 U15126 ( .IN1(n14284), .IN2(n8906), .QN(n14282) );
  NAND2X0 U15127 ( .IN1(n14273), .IN2(n14285), .QN(n14284) );
  NAND2X0 U15128 ( .IN1(n14286), .IN2(n14275), .QN(n14285) );
  XOR2X1 U15129 ( .IN1(n8560), .IN2(n5714), .Q(n14286) );
  NAND3X0 U15130 ( .IN1(n5710), .IN2(n14280), .IN3(n8048), .QN(n14273) );
  NAND2X0 U15131 ( .IN1(n14287), .IN2(n14288), .QN(g26946) );
  NAND3X0 U15132 ( .IN1(n8894), .IN2(g4392), .IN3(n14280), .QN(n14288) );
  NAND2X0 U15133 ( .IN1(n14258), .IN2(g4375), .QN(n14287) );
  NAND3X0 U15134 ( .IN1(n14289), .IN2(n14290), .IN3(n14291), .QN(g26945) );
  NAND2X0 U15135 ( .IN1(n8993), .IN2(g4411), .QN(n14291) );
  NAND2X0 U15136 ( .IN1(n14255), .IN2(n14280), .QN(n14290) );
  INVX0 U15137 ( .INP(n14275), .ZN(n14280) );
  NAND4X0 U15138 ( .IN1(n8561), .IN2(n8560), .IN3(n8562), .IN4(n14292), .QN(
        n14275) );
  NOR2X0 U15139 ( .IN1(g4411), .IN2(g7257), .QN(n14292) );
  NOR2X0 U15140 ( .IN1(g4392), .IN2(n8934), .QN(n14255) );
  NAND2X0 U15141 ( .IN1(n14264), .IN2(g4375), .QN(n14289) );
  INVX0 U15142 ( .INP(n14258), .ZN(n14264) );
  NAND2X0 U15143 ( .IN1(n5714), .IN2(n8907), .QN(n14258) );
  NOR2X0 U15144 ( .IN1(n8955), .IN2(n14293), .QN(g26944) );
  NOR4X0 U15145 ( .IN1(n14294), .IN2(n13918), .IN3(n8590), .IN4(n10178), .QN(
        n14293) );
  NAND2X0 U15146 ( .IN1(n14295), .IN2(n14296), .QN(n13918) );
  INVX0 U15147 ( .INP(g135), .ZN(n14296) );
  NAND3X0 U15148 ( .IN1(n14297), .IN2(n14298), .IN3(n14299), .QN(n14295) );
  NAND3X0 U15149 ( .IN1(n14300), .IN2(n5608), .IN3(n14301), .QN(n14299) );
  XOR2X1 U15150 ( .IN1(g4608), .IN2(n5539), .Q(n14301) );
  XOR2X1 U15151 ( .IN1(g4593), .IN2(n5365), .Q(n14300) );
  NAND4X0 U15152 ( .IN1(n5365), .IN2(g4593), .IN3(n5274), .IN4(g4584), .QN(
        n14298) );
  NAND3X0 U15153 ( .IN1(n5303), .IN2(g4608), .IN3(n5539), .QN(n14297) );
  NAND3X0 U15154 ( .IN1(g4340), .IN2(g4633), .IN3(g4358), .QN(n14294) );
  NAND2X0 U15155 ( .IN1(n14302), .IN2(n14303), .QN(g26940) );
  NAND2X0 U15156 ( .IN1(n8993), .IN2(g4153), .QN(n14303) );
  NAND2X0 U15157 ( .IN1(n12363), .IN2(n8908), .QN(n14302) );
  NAND2X0 U15158 ( .IN1(n14304), .IN2(n14305), .QN(n12363) );
  NAND2X0 U15159 ( .IN1(g116), .IN2(g4157), .QN(n14305) );
  NAND2X0 U15160 ( .IN1(g114), .IN2(n5983), .QN(n14304) );
  NAND2X0 U15161 ( .IN1(n14306), .IN2(n14307), .QN(g26939) );
  NAND2X0 U15162 ( .IN1(n8993), .IN2(g4104), .QN(n14307) );
  NAND2X0 U15163 ( .IN1(n12361), .IN2(n8907), .QN(n14306) );
  NAND2X0 U15164 ( .IN1(n14308), .IN2(n14309), .QN(n12361) );
  NAND2X0 U15165 ( .IN1(g124), .IN2(g4146), .QN(n14309) );
  NAND2X0 U15166 ( .IN1(g120), .IN2(n5981), .QN(n14308) );
  NAND3X0 U15167 ( .IN1(n14310), .IN2(n14311), .IN3(n11495), .QN(g26938) );
  NAND2X0 U15168 ( .IN1(n8993), .IN2(g4141), .QN(n14311) );
  NAND2X0 U15169 ( .IN1(n14312), .IN2(n8906), .QN(n14310) );
  XOR2X1 U15170 ( .IN1(n13944), .IN2(g4082), .Q(n14312) );
  NOR2X0 U15171 ( .IN1(n1242), .IN2(n5612), .QN(n13944) );
  NAND3X0 U15172 ( .IN1(n14313), .IN2(n14314), .IN3(n14315), .QN(g26934) );
  NAND2X0 U15173 ( .IN1(n4888), .IN2(g2827), .QN(n14315) );
  NAND2X0 U15174 ( .IN1(n14316), .IN2(n8636), .QN(n14314) );
  NAND2X0 U15175 ( .IN1(test_so37), .IN2(n9053), .QN(n14313) );
  NAND3X0 U15176 ( .IN1(n14317), .IN2(n14318), .IN3(n14319), .QN(g26933) );
  NAND2X0 U15177 ( .IN1(n4888), .IN2(test_so37), .QN(n14319) );
  NAND2X0 U15178 ( .IN1(n5840), .IN2(n14316), .QN(n14318) );
  NAND2X0 U15179 ( .IN1(n8993), .IN2(g2811), .QN(n14317) );
  NAND3X0 U15180 ( .IN1(n14320), .IN2(n14321), .IN3(n14322), .QN(g26932) );
  NAND2X0 U15181 ( .IN1(n4888), .IN2(g2811), .QN(n14322) );
  NAND2X0 U15182 ( .IN1(n5841), .IN2(n14316), .QN(n14321) );
  NAND2X0 U15183 ( .IN1(n8993), .IN2(g2799), .QN(n14320) );
  NAND3X0 U15184 ( .IN1(n14323), .IN2(n14324), .IN3(n14325), .QN(g26931) );
  NAND2X0 U15185 ( .IN1(n4888), .IN2(g2799), .QN(n14325) );
  NAND2X0 U15186 ( .IN1(n5839), .IN2(n14316), .QN(n14324) );
  NAND2X0 U15187 ( .IN1(n8993), .IN2(g29219), .QN(n14323) );
  NAND3X0 U15188 ( .IN1(n14326), .IN2(n14327), .IN3(n14328), .QN(g26930) );
  NAND2X0 U15189 ( .IN1(n4888), .IN2(g2795), .QN(n14328) );
  NAND2X0 U15190 ( .IN1(n14316), .IN2(n8637), .QN(n14327) );
  NAND2X0 U15191 ( .IN1(n8992), .IN2(g2791), .QN(n14326) );
  NAND3X0 U15192 ( .IN1(n14329), .IN2(n14330), .IN3(n14331), .QN(g26929) );
  NAND2X0 U15193 ( .IN1(n4888), .IN2(g2791), .QN(n14331) );
  NAND2X0 U15194 ( .IN1(n5837), .IN2(n14316), .QN(n14330) );
  NAND2X0 U15195 ( .IN1(n8992), .IN2(g2779), .QN(n14329) );
  NAND3X0 U15196 ( .IN1(n14332), .IN2(n14333), .IN3(n14334), .QN(g26928) );
  NAND2X0 U15197 ( .IN1(n4888), .IN2(g2779), .QN(n14334) );
  NAND2X0 U15198 ( .IN1(n5834), .IN2(n14316), .QN(n14333) );
  NAND2X0 U15199 ( .IN1(n8992), .IN2(g2767), .QN(n14332) );
  NAND3X0 U15200 ( .IN1(n14335), .IN2(n14336), .IN3(n14337), .QN(g26927) );
  NAND2X0 U15201 ( .IN1(n4888), .IN2(g2767), .QN(n14337) );
  NAND2X0 U15202 ( .IN1(n5836), .IN2(n14316), .QN(n14336) );
  INVX0 U15203 ( .INP(n14338), .ZN(n14316) );
  NAND3X0 U15204 ( .IN1(n14339), .IN2(n10015), .IN3(n4888), .QN(n14338) );
  NAND3X0 U15205 ( .IN1(n3505), .IN2(g2735), .IN3(test_so30), .QN(n10015) );
  NOR2X0 U15206 ( .IN1(n5349), .IN2(n5516), .QN(n3505) );
  NAND2X0 U15207 ( .IN1(n5516), .IN2(n5300), .QN(n14339) );
  NAND2X0 U15208 ( .IN1(n8992), .IN2(g2763), .QN(n14335) );
  NAND2X0 U15209 ( .IN1(n14340), .IN2(n14341), .QN(g26926) );
  NAND2X0 U15210 ( .IN1(n14342), .IN2(n3730), .QN(n14341) );
  XOR2X1 U15211 ( .IN1(g2724), .IN2(n12644), .Q(n14342) );
  NOR2X0 U15212 ( .IN1(n5299), .IN2(n5465), .QN(n12644) );
  INVX0 U15213 ( .INP(n14343), .ZN(n14340) );
  NOR2X0 U15214 ( .IN1(n8900), .IN2(n5465), .QN(n14343) );
  NAND2X0 U15215 ( .IN1(n14344), .IN2(n14345), .QN(g26925) );
  NAND2X0 U15216 ( .IN1(n8992), .IN2(g1532), .QN(n14345) );
  NAND2X0 U15217 ( .IN1(n14346), .IN2(n8907), .QN(n14344) );
  NAND2X0 U15218 ( .IN1(n12934), .IN2(n14347), .QN(n14346) );
  NAND2X0 U15219 ( .IN1(n12917), .IN2(g1536), .QN(n14347) );
  NAND2X0 U15220 ( .IN1(n12921), .IN2(g1413), .QN(n12917) );
  NOR2X0 U15221 ( .IN1(n12925), .IN2(n8487), .QN(n12921) );
  NAND3X0 U15222 ( .IN1(n14348), .IN2(g7946), .IN3(n12936), .QN(n12925) );
  INVX0 U15223 ( .INP(n11097), .ZN(n12936) );
  NAND3X0 U15224 ( .IN1(g1339), .IN2(g1521), .IN3(n8307), .QN(n14348) );
  INVX0 U15225 ( .INP(n4173), .ZN(n12934) );
  NAND2X0 U15226 ( .IN1(n14349), .IN2(n14350), .QN(g26924) );
  NAND2X0 U15227 ( .IN1(n14351), .IN2(g1437), .QN(n14350) );
  NAND2X0 U15228 ( .IN1(n14352), .IN2(n8906), .QN(n14351) );
  NAND3X0 U15229 ( .IN1(n13478), .IN2(n5289), .IN3(n14353), .QN(n14352) );
  NAND3X0 U15230 ( .IN1(n8894), .IN2(g1478), .IN3(n14354), .QN(n14349) );
  NAND3X0 U15231 ( .IN1(n13478), .IN2(g1437), .IN3(n14353), .QN(n14354) );
  NOR3X0 U15232 ( .IN1(n8521), .IN2(test_so49), .IN3(n5364), .QN(n13478) );
  NAND3X0 U15233 ( .IN1(n14355), .IN2(n14356), .IN3(n14357), .QN(g26923) );
  NAND2X0 U15234 ( .IN1(n14358), .IN2(n5290), .QN(n14357) );
  INVX0 U15235 ( .INP(n14359), .ZN(n14358) );
  NAND3X0 U15236 ( .IN1(n14359), .IN2(g1472), .IN3(n8887), .QN(n14356) );
  NAND4X0 U15237 ( .IN1(n14353), .IN2(n13469), .IN3(g1467), .IN4(g13272), .QN(
        n14359) );
  NAND2X0 U15238 ( .IN1(n8992), .IN2(g1467), .QN(n14355) );
  NAND3X0 U15239 ( .IN1(n14360), .IN2(n14361), .IN3(n14362), .QN(g26922) );
  NAND2X0 U15240 ( .IN1(n14363), .IN2(n5343), .QN(n14362) );
  INVX0 U15241 ( .INP(n14364), .ZN(n14363) );
  NAND3X0 U15242 ( .IN1(n14364), .IN2(g1448), .IN3(n8887), .QN(n14361) );
  NAND3X0 U15243 ( .IN1(n13454), .IN2(g1454), .IN3(n14353), .QN(n14364) );
  NOR2X0 U15244 ( .IN1(n11097), .IN2(n8521), .QN(n13454) );
  NAND2X0 U15245 ( .IN1(test_so49), .IN2(n5364), .QN(n11097) );
  NAND2X0 U15246 ( .IN1(n8992), .IN2(g1454), .QN(n14360) );
  NAND2X0 U15247 ( .IN1(n14365), .IN2(n14366), .QN(g26921) );
  NAND2X0 U15248 ( .IN1(n8991), .IN2(g1395), .QN(n14366) );
  NAND3X0 U15249 ( .IN1(n14367), .IN2(n8602), .IN3(n8887), .QN(n14365) );
  XNOR2X1 U15250 ( .IN1(n14368), .IN2(n8167), .Q(n14367) );
  NAND2X0 U15251 ( .IN1(n14369), .IN2(n14370), .QN(g26920) );
  NAND2X0 U15252 ( .IN1(n8991), .IN2(g1384), .QN(n14370) );
  NAND2X0 U15253 ( .IN1(n14371), .IN2(n8907), .QN(n14369) );
  NAND2X0 U15254 ( .IN1(n14372), .IN2(n14373), .QN(n14371) );
  NAND2X0 U15255 ( .IN1(n9339), .IN2(g1389), .QN(n14373) );
  NAND2X0 U15256 ( .IN1(n14374), .IN2(n14375), .QN(n9339) );
  NAND2X0 U15257 ( .IN1(n8055), .IN2(g1351), .QN(n14375) );
  NAND2X0 U15258 ( .IN1(n4913), .IN2(g1351), .QN(n14372) );
  NAND3X0 U15259 ( .IN1(n14376), .IN2(n14377), .IN3(n14378), .QN(g26919) );
  NAND2X0 U15260 ( .IN1(n8991), .IN2(g1266), .QN(n14378) );
  NAND3X0 U15261 ( .IN1(test_so77), .IN2(n11311), .IN3(n14379), .QN(n14377) );
  NAND2X0 U15262 ( .IN1(n1220), .IN2(n5556), .QN(n14376) );
  INVX0 U15263 ( .INP(n14379), .ZN(n1220) );
  NAND3X0 U15264 ( .IN1(g1249), .IN2(g1266), .IN3(g12923), .QN(n14379) );
  NAND2X0 U15265 ( .IN1(n14380), .IN2(n14381), .QN(g26918) );
  NAND2X0 U15266 ( .IN1(n8991), .IN2(g1189), .QN(n14381) );
  NAND2X0 U15267 ( .IN1(n14382), .IN2(n8907), .QN(n14380) );
  NAND2X0 U15268 ( .IN1(n12969), .IN2(n14383), .QN(n14382) );
  NAND2X0 U15269 ( .IN1(n12952), .IN2(g1193), .QN(n14383) );
  NAND2X0 U15270 ( .IN1(n12956), .IN2(g1070), .QN(n12952) );
  NOR2X0 U15271 ( .IN1(n12960), .IN2(n8486), .QN(n12956) );
  NAND3X0 U15272 ( .IN1(n14384), .IN2(g7916), .IN3(n12971), .QN(n12960) );
  INVX0 U15273 ( .INP(n11257), .ZN(n12971) );
  NAND3X0 U15274 ( .IN1(g1178), .IN2(g996), .IN3(n5642), .QN(n14384) );
  INVX0 U15275 ( .INP(n4191), .ZN(n12969) );
  NAND3X0 U15276 ( .IN1(n14385), .IN2(n14386), .IN3(n14387), .QN(g26917) );
  NAND2X0 U15277 ( .IN1(n14388), .IN2(n5328), .QN(n14387) );
  INVX0 U15278 ( .INP(n14389), .ZN(n14388) );
  NAND3X0 U15279 ( .IN1(n14389), .IN2(g1135), .IN3(n8886), .QN(n14386) );
  NAND4X0 U15280 ( .IN1(n14390), .IN2(n11350), .IN3(g1094), .IN4(g13259), .QN(
        n14389) );
  NOR2X0 U15281 ( .IN1(g1183), .IN2(n5363), .QN(n11350) );
  NAND2X0 U15282 ( .IN1(n8991), .IN2(g1094), .QN(n14385) );
  NAND3X0 U15283 ( .IN1(n14391), .IN2(n14392), .IN3(n14393), .QN(g26916) );
  NAND2X0 U15284 ( .IN1(n14394), .IN2(n5329), .QN(n14393) );
  INVX0 U15285 ( .INP(n14395), .ZN(n14394) );
  NAND3X0 U15286 ( .IN1(n14395), .IN2(g1129), .IN3(n8886), .QN(n14392) );
  NAND4X0 U15287 ( .IN1(n14390), .IN2(n11219), .IN3(g1124), .IN4(g13259), .QN(
        n14395) );
  NAND2X0 U15288 ( .IN1(n8991), .IN2(g1124), .QN(n14391) );
  NAND3X0 U15289 ( .IN1(n14396), .IN2(n14397), .IN3(n14398), .QN(g26915) );
  NAND2X0 U15290 ( .IN1(n14399), .IN2(n5478), .QN(n14398) );
  INVX0 U15291 ( .INP(n14400), .ZN(n14399) );
  NAND3X0 U15292 ( .IN1(n14400), .IN2(g1105), .IN3(n8886), .QN(n14397) );
  NAND3X0 U15293 ( .IN1(test_so90), .IN2(n13490), .IN3(n14390), .QN(n14400) );
  NOR2X0 U15294 ( .IN1(n11257), .IN2(n8527), .QN(n13490) );
  NAND2X0 U15295 ( .IN1(n5363), .IN2(g1183), .QN(n11257) );
  NAND2X0 U15296 ( .IN1(test_so90), .IN2(n9054), .QN(n14396) );
  NAND2X0 U15297 ( .IN1(n14401), .IN2(n14402), .QN(g26914) );
  NAND2X0 U15298 ( .IN1(n8991), .IN2(g1052), .QN(n14402) );
  NAND3X0 U15299 ( .IN1(n5320), .IN2(n14403), .IN3(n8886), .QN(n14401) );
  XNOR2X1 U15300 ( .IN1(n14404), .IN2(n8168), .Q(n14403) );
  NAND3X0 U15301 ( .IN1(n14405), .IN2(n14406), .IN3(n14407), .QN(g26913) );
  NAND2X0 U15302 ( .IN1(n4938), .IN2(n14408), .QN(n14407) );
  NAND2X0 U15303 ( .IN1(n8990), .IN2(g1041), .QN(n14406) );
  NAND3X0 U15304 ( .IN1(n9199), .IN2(g1046), .IN3(n8886), .QN(n14405) );
  NAND2X0 U15305 ( .IN1(n14409), .IN2(n14410), .QN(n9199) );
  NAND2X0 U15306 ( .IN1(n8054), .IN2(g1008), .QN(n14410) );
  NAND3X0 U15307 ( .IN1(n14411), .IN2(n14412), .IN3(n14413), .QN(g26912) );
  NAND2X0 U15308 ( .IN1(n8990), .IN2(g921), .QN(n14413) );
  NAND3X0 U15309 ( .IN1(n11325), .IN2(n14414), .IN3(g936), .QN(n14412) );
  NAND2X0 U15310 ( .IN1(n279), .IN2(n5557), .QN(n14411) );
  INVX0 U15311 ( .INP(n14414), .ZN(n279) );
  NAND3X0 U15312 ( .IN1(g921), .IN2(g904), .IN3(g12919), .QN(n14414) );
  XOR2X1 U15313 ( .IN1(n14415), .IN2(n5682), .Q(g26910) );
  NAND2X0 U15314 ( .IN1(n5305), .IN2(n8907), .QN(n14415) );
  NAND2X0 U15315 ( .IN1(n14416), .IN2(n14417), .QN(g26909) );
  NAND2X0 U15316 ( .IN1(n8990), .IN2(g890), .QN(n14417) );
  NAND2X0 U15317 ( .IN1(n14418), .IN2(n8907), .QN(n14416) );
  NAND2X0 U15318 ( .IN1(n14419), .IN2(n14420), .QN(n14418) );
  NAND2X0 U15319 ( .IN1(n5431), .IN2(g862), .QN(n14420) );
  NAND2X0 U15320 ( .IN1(n5305), .IN2(g896), .QN(n14419) );
  NAND3X0 U15321 ( .IN1(n14421), .IN2(n14422), .IN3(n14423), .QN(g26908) );
  NAND2X0 U15322 ( .IN1(n4945), .IN2(g446), .QN(n14423) );
  NAND2X0 U15323 ( .IN1(n14424), .IN2(g872), .QN(n14422) );
  NAND2X0 U15324 ( .IN1(n8990), .IN2(g246), .QN(n14421) );
  NAND3X0 U15325 ( .IN1(n14425), .IN2(n14426), .IN3(n14427), .QN(g26907) );
  NAND2X0 U15326 ( .IN1(n4945), .IN2(g246), .QN(n14427) );
  NAND2X0 U15327 ( .IN1(n14424), .IN2(g14167), .QN(n14426) );
  NAND2X0 U15328 ( .IN1(n8990), .IN2(g269), .QN(n14425) );
  NAND3X0 U15329 ( .IN1(n14428), .IN2(n14429), .IN3(n14430), .QN(g26906) );
  NAND2X0 U15330 ( .IN1(n4945), .IN2(g269), .QN(n14430) );
  NAND2X0 U15331 ( .IN1(n14424), .IN2(g14147), .QN(n14429) );
  NAND2X0 U15332 ( .IN1(n8990), .IN2(g239), .QN(n14428) );
  NAND3X0 U15333 ( .IN1(n14431), .IN2(n14432), .IN3(n14433), .QN(g26905) );
  NAND2X0 U15334 ( .IN1(n4945), .IN2(g239), .QN(n14433) );
  NAND2X0 U15335 ( .IN1(n14424), .IN2(g14125), .QN(n14432) );
  NAND2X0 U15336 ( .IN1(n8990), .IN2(g262), .QN(n14431) );
  NAND3X0 U15337 ( .IN1(n14434), .IN2(n14435), .IN3(n14436), .QN(g26904) );
  NAND2X0 U15338 ( .IN1(n4945), .IN2(g262), .QN(n14436) );
  NAND2X0 U15339 ( .IN1(n14424), .IN2(g14096), .QN(n14435) );
  NAND2X0 U15340 ( .IN1(n8989), .IN2(g232), .QN(n14434) );
  NAND3X0 U15341 ( .IN1(n14437), .IN2(n14438), .IN3(n14439), .QN(g26903) );
  NAND2X0 U15342 ( .IN1(n4945), .IN2(g232), .QN(n14439) );
  NAND2X0 U15343 ( .IN1(n14424), .IN2(g14217), .QN(n14438) );
  NAND2X0 U15344 ( .IN1(n8989), .IN2(g255), .QN(n14437) );
  NAND3X0 U15345 ( .IN1(n14440), .IN2(n14441), .IN3(n14442), .QN(g26902) );
  NAND2X0 U15346 ( .IN1(n4945), .IN2(g255), .QN(n14442) );
  NAND2X0 U15347 ( .IN1(n14424), .IN2(g14201), .QN(n14441) );
  NAND2X0 U15348 ( .IN1(n8989), .IN2(g225), .QN(n14440) );
  NAND3X0 U15349 ( .IN1(n14443), .IN2(n14444), .IN3(n14445), .QN(g26901) );
  NAND2X0 U15350 ( .IN1(n4945), .IN2(g225), .QN(n14445) );
  NAND2X0 U15351 ( .IN1(n14424), .IN2(g14189), .QN(n14444) );
  NOR2X0 U15352 ( .IN1(n8948), .IN2(n4946), .QN(n14424) );
  NAND3X0 U15353 ( .IN1(n5431), .IN2(g890), .IN3(n5682), .QN(n4946) );
  NAND2X0 U15354 ( .IN1(n8989), .IN2(g872), .QN(n14443) );
  NAND2X0 U15355 ( .IN1(n14446), .IN2(n14447), .QN(g26899) );
  NAND2X0 U15356 ( .IN1(n14448), .IN2(n4518), .QN(n14447) );
  XOR2X1 U15357 ( .IN1(n4814), .IN2(g822), .Q(n14448) );
  NOR3X0 U15358 ( .IN1(n5822), .IN2(n8519), .IN3(n13562), .QN(n4814) );
  NAND2X0 U15359 ( .IN1(n8989), .IN2(g832), .QN(n14446) );
  NAND2X0 U15360 ( .IN1(n14449), .IN2(n14450), .QN(g26898) );
  NAND2X0 U15361 ( .IN1(n14451), .IN2(n14452), .QN(n14450) );
  NAND2X0 U15362 ( .IN1(n14453), .IN2(n14454), .QN(n14452) );
  NAND2X0 U15363 ( .IN1(n8148), .IN2(n8908), .QN(n14454) );
  NAND2X0 U15364 ( .IN1(n14455), .IN2(g843), .QN(n14449) );
  NAND2X0 U15365 ( .IN1(n14456), .IN2(n8908), .QN(n14455) );
  NAND3X0 U15366 ( .IN1(n5733), .IN2(g837), .IN3(n14457), .QN(n14456) );
  NAND2X0 U15367 ( .IN1(n14458), .IN2(n14459), .QN(g26897) );
  NAND2X0 U15368 ( .IN1(n14460), .IN2(g753), .QN(n14459) );
  INVX0 U15369 ( .INP(n14461), .ZN(n14458) );
  NOR2X0 U15370 ( .IN1(n14460), .IN2(n5732), .QN(n14461) );
  NOR2X0 U15371 ( .IN1(n14186), .IN2(n8928), .QN(n14460) );
  NAND3X0 U15372 ( .IN1(n14462), .IN2(n14463), .IN3(n14464), .QN(g26896) );
  NAND2X0 U15373 ( .IN1(n4956), .IN2(n13541), .QN(n14464) );
  NAND2X0 U15374 ( .IN1(n14465), .IN2(g29212), .QN(n14463) );
  NAND2X0 U15375 ( .IN1(n14466), .IN2(g728), .QN(n14462) );
  INVX0 U15376 ( .INP(n14465), .ZN(n14466) );
  NOR2X0 U15377 ( .IN1(n13541), .IN2(n8929), .QN(n14465) );
  NOR4X0 U15378 ( .IN1(n13562), .IN2(n14180), .IN3(g528), .IN4(n14467), .QN(
        n13541) );
  NAND2X0 U15379 ( .IN1(n5519), .IN2(test_so54), .QN(n14467) );
  NAND3X0 U15380 ( .IN1(n14468), .IN2(n14469), .IN3(n14470), .QN(g26895) );
  NAND2X0 U15381 ( .IN1(n8989), .IN2(g562), .QN(n14470) );
  NAND3X0 U15382 ( .IN1(n2421), .IN2(n14471), .IN3(g568), .QN(n14469) );
  NAND2X0 U15383 ( .IN1(n5), .IN2(n5335), .QN(n14468) );
  INVX0 U15384 ( .INP(n14471), .ZN(n5) );
  NAND3X0 U15385 ( .IN1(n14472), .IN2(g562), .IN3(n4959), .QN(n14471) );
  NAND2X0 U15386 ( .IN1(n14473), .IN2(n14474), .QN(g26894) );
  NAND2X0 U15387 ( .IN1(n8989), .IN2(g518), .QN(n14474) );
  NAND4X0 U15388 ( .IN1(n14475), .IN2(n14476), .IN3(n13551), .IN4(n8901), .QN(
        n14473) );
  NAND2X0 U15389 ( .IN1(n14178), .IN2(g528), .QN(n14476) );
  NAND2X0 U15390 ( .IN1(n5327), .IN2(n14477), .QN(n14475) );
  NAND2X0 U15391 ( .IN1(n14178), .IN2(n14180), .QN(n14477) );
  NAND2X0 U15392 ( .IN1(g482), .IN2(g490), .QN(n14180) );
  NOR3X0 U15393 ( .IN1(g513), .IN2(n5287), .IN3(n14478), .QN(n14178) );
  NAND2X0 U15394 ( .IN1(n14479), .IN2(n14480), .QN(g26893) );
  NAND2X0 U15395 ( .IN1(n9027), .IN2(g355), .QN(n14480) );
  NAND2X0 U15396 ( .IN1(n14481), .IN2(n8907), .QN(n14479) );
  NAND2X0 U15397 ( .IN1(n14482), .IN2(n14483), .QN(n14481) );
  NAND2X0 U15398 ( .IN1(g29211), .IN2(n8609), .QN(n14483) );
  NAND2X0 U15399 ( .IN1(test_so17), .IN2(n14484), .QN(n14482) );
  NAND2X0 U15400 ( .IN1(n14485), .IN2(n14486), .QN(g26892) );
  NAND3X0 U15401 ( .IN1(n8895), .IN2(n14484), .IN3(n8609), .QN(n14486) );
  NAND2X0 U15402 ( .IN1(n8439), .IN2(n8438), .QN(n14484) );
  NAND2X0 U15403 ( .IN1(test_so17), .IN2(n9055), .QN(n14485) );
  NAND2X0 U15404 ( .IN1(n14487), .IN2(n14488), .QN(g26891) );
  NAND2X0 U15405 ( .IN1(n9018), .IN2(g347), .QN(n14488) );
  NAND3X0 U15406 ( .IN1(n8894), .IN2(g7540), .IN3(n5860), .QN(n14487) );
  NAND2X0 U15407 ( .IN1(n14489), .IN2(n14490), .QN(g26890) );
  NAND2X0 U15408 ( .IN1(n5860), .IN2(n8907), .QN(n14490) );
  NAND2X0 U15409 ( .IN1(n9017), .IN2(g333), .QN(n14489) );
  NAND2X0 U15410 ( .IN1(n14491), .IN2(n14492), .QN(g26889) );
  NAND2X0 U15411 ( .IN1(n9021), .IN2(g29211), .QN(n14492) );
  NAND4X0 U15412 ( .IN1(g329), .IN2(DFF_709_n1), .IN3(n14493), .IN4(n8901), 
        .QN(n14491) );
  NAND2X0 U15413 ( .IN1(n14494), .IN2(n14495), .QN(g26888) );
  NAND2X0 U15414 ( .IN1(n8904), .IN2(g316), .QN(n14495) );
  NAND2X0 U15415 ( .IN1(n9022), .IN2(g29216), .QN(n14494) );
  NAND3X0 U15416 ( .IN1(n14496), .IN2(n14497), .IN3(n14498), .QN(g26887) );
  NAND2X0 U15417 ( .IN1(n9026), .IN2(g336), .QN(n14497) );
  NAND3X0 U15418 ( .IN1(n5317), .IN2(g324), .IN3(n8886), .QN(n14496) );
  NAND3X0 U15419 ( .IN1(n14499), .IN2(n14500), .IN3(n14501), .QN(g26886) );
  INVX0 U15420 ( .INP(n14502), .ZN(n14501) );
  NOR2X0 U15421 ( .IN1(n14498), .IN2(n14493), .QN(n14502) );
  NAND3X0 U15422 ( .IN1(n14493), .IN2(g336), .IN3(n8886), .QN(n14500) );
  NAND2X0 U15423 ( .IN1(n9025), .IN2(g311), .QN(n14499) );
  NAND2X0 U15424 ( .IN1(n14503), .IN2(n14504), .QN(g26884) );
  NAND2X0 U15425 ( .IN1(n9035), .IN2(g329), .QN(n14504) );
  NAND2X0 U15426 ( .IN1(n14505), .IN2(n8907), .QN(n14503) );
  NAND2X0 U15427 ( .IN1(n14506), .IN2(n14507), .QN(n14505) );
  NAND4X0 U15428 ( .IN1(n5766), .IN2(n5456), .IN3(n5282), .IN4(n5317), .QN(
        n14507) );
  NAND2X0 U15429 ( .IN1(n14508), .IN2(n14509), .QN(n14506) );
  NAND3X0 U15430 ( .IN1(n14510), .IN2(n14511), .IN3(n5456), .QN(n14509) );
  NAND2X0 U15431 ( .IN1(n5824), .IN2(g311), .QN(n14511) );
  NAND2X0 U15432 ( .IN1(g305), .IN2(g336), .QN(n14510) );
  NAND2X0 U15433 ( .IN1(n14512), .IN2(n14513), .QN(g26883) );
  NAND2X0 U15434 ( .IN1(n9036), .IN2(g324), .QN(n14513) );
  NAND2X0 U15435 ( .IN1(n14508), .IN2(n8908), .QN(n14512) );
  INVX0 U15436 ( .INP(n14493), .ZN(n14508) );
  NAND2X0 U15437 ( .IN1(n14514), .IN2(n14515), .QN(n14493) );
  NAND2X0 U15438 ( .IN1(n5282), .IN2(g324), .QN(n14515) );
  NAND2X0 U15439 ( .IN1(n5827), .IN2(n5317), .QN(n14514) );
  NAND3X0 U15440 ( .IN1(n14516), .IN2(n14517), .IN3(n14498), .QN(g26882) );
  NAND2X0 U15441 ( .IN1(n8904), .IN2(g305), .QN(n14498) );
  NAND2X0 U15442 ( .IN1(n8903), .IN2(g311), .QN(n14517) );
  NAND2X0 U15443 ( .IN1(n9029), .IN2(g316), .QN(n14516) );
  NAND2X0 U15444 ( .IN1(n14518), .IN2(n14519), .QN(g26881) );
  NAND2X0 U15445 ( .IN1(g6744), .IN2(n8908), .QN(n14519) );
  NAND2X0 U15446 ( .IN1(n9030), .IN2(g305), .QN(n14518) );
  NAND3X0 U15447 ( .IN1(n9714), .IN2(n8871), .IN3(n9715), .QN(g26877) );
  NAND4X0 U15448 ( .IN1(n5620), .IN2(n5619), .IN3(n14520), .IN4(n14521), .QN(
        n9715) );
  NOR4X0 U15449 ( .IN1(test_so40), .IN2(g2357), .IN3(g2338), .IN4(g2606), .QN(
        n14521) );
  NOR2X0 U15450 ( .IN1(g2491), .IN2(g2223), .QN(n14520) );
  NAND4X0 U15451 ( .IN1(n5833), .IN2(n5832), .IN3(n14522), .IN4(n14523), .QN(
        n9714) );
  NOR4X0 U15452 ( .IN1(test_so75), .IN2(g1664), .IN3(g1913), .IN4(g1932), .QN(
        n14523) );
  NOR2X0 U15453 ( .IN1(g1779), .IN2(g2047), .QN(n14522) );
  NAND2X0 U15454 ( .IN1(n14524), .IN2(n9679), .QN(g26876) );
  NAND4X0 U15455 ( .IN1(n15228), .IN2(n5892), .IN3(n14525), .IN4(n14526), .QN(
        n9679) );
  NOR4X0 U15456 ( .IN1(g1710), .IN2(g1978), .IN3(g1844), .IN4(g2112), .QN(
        n14526) );
  NOR2X0 U15457 ( .IN1(g1992), .IN2(g2126), .QN(n14525) );
  INVX0 U15458 ( .INP(n9675), .ZN(n14524) );
  NAND2X0 U15459 ( .IN1(n14527), .IN2(n8908), .QN(n9675) );
  NAND4X0 U15460 ( .IN1(n15224), .IN2(n15229), .IN3(n14528), .IN4(n14529), 
        .QN(n14527) );
  NOR4X0 U15461 ( .IN1(test_so31), .IN2(g2671), .IN3(g2269), .IN4(g2537), .QN(
        n14529) );
  NOR2X0 U15462 ( .IN1(n9324), .IN2(n9295), .QN(n14528) );
  NAND2X0 U15463 ( .IN1(n14530), .IN2(n9680), .QN(g26875) );
  NAND4X0 U15464 ( .IN1(n5628), .IN2(n5413), .IN3(n5315), .IN4(n5280), .QN(
        n9680) );
  INVX0 U15465 ( .INP(n9676), .ZN(n14530) );
  NAND2X0 U15466 ( .IN1(n14531), .IN2(n8908), .QN(n9676) );
  NAND4X0 U15467 ( .IN1(n5631), .IN2(n5414), .IN3(n5316), .IN4(n5281), .QN(
        n14531) );
  NAND2X0 U15468 ( .IN1(n14532), .IN2(n14533), .QN(g25764) );
  NAND2X0 U15469 ( .IN1(n11922), .IN2(g6505), .QN(n14533) );
  NAND2X0 U15470 ( .IN1(n14534), .IN2(g6541), .QN(n14532) );
  NAND3X0 U15471 ( .IN1(n14535), .IN2(n14536), .IN3(n14537), .QN(g25763) );
  NAND2X0 U15472 ( .IN1(n11922), .IN2(g6537), .QN(n14537) );
  NAND2X0 U15473 ( .IN1(n14538), .IN2(g6533), .QN(n14536) );
  NAND2X0 U15474 ( .IN1(n14539), .IN2(n8908), .QN(n14538) );
  NAND2X0 U15475 ( .IN1(n10839), .IN2(g6527), .QN(n14539) );
  NAND4X0 U15476 ( .IN1(n10839), .IN2(n8899), .IN3(n5659), .IN4(n5445), .QN(
        n14535) );
  NAND2X0 U15477 ( .IN1(n14540), .IN2(n14541), .QN(g25762) );
  NAND2X0 U15478 ( .IN1(n11922), .IN2(g6533), .QN(n14541) );
  NAND2X0 U15479 ( .IN1(n14534), .IN2(g6527), .QN(n14540) );
  INVX0 U15480 ( .INP(n11922), .ZN(n14534) );
  NAND3X0 U15481 ( .IN1(n14542), .IN2(n14543), .IN3(n14544), .QN(g25761) );
  NAND2X0 U15482 ( .IN1(n11922), .IN2(g6513), .QN(n14544) );
  NOR2X0 U15483 ( .IN1(n10839), .IN2(n8928), .QN(n11922) );
  NAND3X0 U15484 ( .IN1(n5426), .IN2(n10839), .IN3(n8886), .QN(n14543) );
  NOR2X0 U15485 ( .IN1(n1409), .IN2(n5646), .QN(n10839) );
  NAND2X0 U15486 ( .IN1(g6565), .IN2(g6573), .QN(n1409) );
  NAND2X0 U15487 ( .IN1(n9032), .IN2(g6509), .QN(n14542) );
  NAND2X0 U15488 ( .IN1(n14545), .IN2(n14546), .QN(g25758) );
  NAND2X0 U15489 ( .IN1(n9028), .IN2(g6494), .QN(n14546) );
  NAND3X0 U15490 ( .IN1(n8088), .IN2(n14547), .IN3(n8886), .QN(n14545) );
  NAND2X0 U15491 ( .IN1(n5990), .IN2(n14548), .QN(n14547) );
  NAND2X0 U15492 ( .IN1(n8528), .IN2(g9743), .QN(n14548) );
  NAND2X0 U15493 ( .IN1(n14549), .IN2(n14550), .QN(g25757) );
  NAND2X0 U15494 ( .IN1(n8904), .IN2(g6727), .QN(n14550) );
  NAND2X0 U15495 ( .IN1(n8988), .IN2(g6444), .QN(n14549) );
  NOR2X0 U15496 ( .IN1(n8950), .IN2(n5563), .QN(g25756) );
  NAND2X0 U15497 ( .IN1(n14551), .IN2(n14552), .QN(g25750) );
  NAND2X0 U15498 ( .IN1(n12008), .IN2(g6159), .QN(n14552) );
  NAND2X0 U15499 ( .IN1(n14553), .IN2(g6195), .QN(n14551) );
  NAND3X0 U15500 ( .IN1(n14554), .IN2(n14555), .IN3(n14556), .QN(g25749) );
  NAND2X0 U15501 ( .IN1(n12008), .IN2(g6191), .QN(n14556) );
  NAND2X0 U15502 ( .IN1(n14557), .IN2(g6187), .QN(n14555) );
  NAND2X0 U15503 ( .IN1(n14558), .IN2(n8909), .QN(n14557) );
  NAND2X0 U15504 ( .IN1(n12009), .IN2(g6181), .QN(n14558) );
  NAND4X0 U15505 ( .IN1(n12009), .IN2(n8899), .IN3(n5667), .IN4(n5453), .QN(
        n14554) );
  NAND2X0 U15506 ( .IN1(n14559), .IN2(n14560), .QN(g25748) );
  NAND2X0 U15507 ( .IN1(n12008), .IN2(g6187), .QN(n14560) );
  NAND2X0 U15508 ( .IN1(n14553), .IN2(g6181), .QN(n14559) );
  NAND3X0 U15509 ( .IN1(n14561), .IN2(n14562), .IN3(n14563), .QN(g25747) );
  NAND2X0 U15510 ( .IN1(n12008), .IN2(g6167), .QN(n14563) );
  INVX0 U15511 ( .INP(n14553), .ZN(n12008) );
  NAND2X0 U15512 ( .IN1(n10828), .IN2(n8908), .QN(n14553) );
  NAND3X0 U15513 ( .IN1(n5430), .IN2(n12009), .IN3(n8889), .QN(n14562) );
  INVX0 U15514 ( .INP(n10828), .ZN(n12009) );
  NAND2X0 U15515 ( .IN1(n12029), .IN2(g6215), .QN(n10828) );
  INVX0 U15516 ( .INP(n51), .ZN(n12029) );
  NAND2X0 U15517 ( .IN1(g6219), .IN2(g6227), .QN(n51) );
  NAND2X0 U15518 ( .IN1(n8988), .IN2(g6163), .QN(n14561) );
  NAND2X0 U15519 ( .IN1(n14564), .IN2(n14565), .QN(g25744) );
  NAND2X0 U15520 ( .IN1(n8988), .IN2(g6148), .QN(n14565) );
  NAND3X0 U15521 ( .IN1(n8084), .IN2(n14566), .IN3(n8886), .QN(n14564) );
  NAND2X0 U15522 ( .IN1(n5988), .IN2(n14567), .QN(n14566) );
  NAND2X0 U15523 ( .IN1(test_so92), .IN2(n8529), .QN(n14567) );
  NAND2X0 U15524 ( .IN1(n14568), .IN2(n14569), .QN(g25743) );
  NAND2X0 U15525 ( .IN1(test_so69), .IN2(n8908), .QN(n14569) );
  NAND2X0 U15526 ( .IN1(n8988), .IN2(g6098), .QN(n14568) );
  NOR2X0 U15527 ( .IN1(n8951), .IN2(n5568), .QN(g25742) );
  NAND2X0 U15528 ( .IN1(n14570), .IN2(n14571), .QN(g25736) );
  NAND2X0 U15529 ( .IN1(n12095), .IN2(g5813), .QN(n14571) );
  NAND2X0 U15530 ( .IN1(n14572), .IN2(g5849), .QN(n14570) );
  NAND3X0 U15531 ( .IN1(n14573), .IN2(n14574), .IN3(n14575), .QN(g25735) );
  NAND2X0 U15532 ( .IN1(test_so83), .IN2(n12095), .QN(n14575) );
  NAND2X0 U15533 ( .IN1(n14576), .IN2(g5841), .QN(n14574) );
  NAND2X0 U15534 ( .IN1(n14577), .IN2(n8909), .QN(n14576) );
  NAND2X0 U15535 ( .IN1(n12096), .IN2(g5835), .QN(n14577) );
  NAND4X0 U15536 ( .IN1(n12096), .IN2(n8899), .IN3(n5663), .IN4(n5449), .QN(
        n14573) );
  NAND2X0 U15537 ( .IN1(n14578), .IN2(n14579), .QN(g25734) );
  NAND2X0 U15538 ( .IN1(n12095), .IN2(g5841), .QN(n14579) );
  NAND2X0 U15539 ( .IN1(n14572), .IN2(g5835), .QN(n14578) );
  NAND3X0 U15540 ( .IN1(n14580), .IN2(n14581), .IN3(n14582), .QN(g25733) );
  NAND2X0 U15541 ( .IN1(n12095), .IN2(g5821), .QN(n14582) );
  INVX0 U15542 ( .INP(n14572), .ZN(n12095) );
  NAND2X0 U15543 ( .IN1(n10827), .IN2(n8908), .QN(n14572) );
  NAND3X0 U15544 ( .IN1(n5429), .IN2(n12096), .IN3(n8886), .QN(n14581) );
  INVX0 U15545 ( .INP(n10827), .ZN(n12096) );
  NAND2X0 U15546 ( .IN1(n12116), .IN2(g5869), .QN(n10827) );
  INVX0 U15547 ( .INP(n720), .ZN(n12116) );
  NAND2X0 U15548 ( .IN1(test_so36), .IN2(g5873), .QN(n720) );
  NAND2X0 U15549 ( .IN1(n8988), .IN2(g5817), .QN(n14580) );
  NAND2X0 U15550 ( .IN1(n14583), .IN2(n14584), .QN(g25730) );
  NAND2X0 U15551 ( .IN1(n8988), .IN2(g5802), .QN(n14584) );
  NAND3X0 U15552 ( .IN1(n8095), .IN2(n14585), .IN3(n8886), .QN(n14583) );
  NAND2X0 U15553 ( .IN1(n5996), .IN2(n14586), .QN(n14585) );
  NAND2X0 U15554 ( .IN1(n8523), .IN2(g9617), .QN(n14586) );
  NAND2X0 U15555 ( .IN1(n14587), .IN2(n14588), .QN(g25729) );
  NAND2X0 U15556 ( .IN1(n8903), .IN2(g6035), .QN(n14588) );
  NAND2X0 U15557 ( .IN1(n8988), .IN2(g5752), .QN(n14587) );
  NOR2X0 U15558 ( .IN1(n8599), .IN2(n9047), .QN(g25728) );
  NAND2X0 U15559 ( .IN1(n14589), .IN2(n14590), .QN(g25722) );
  NAND2X0 U15560 ( .IN1(n12182), .IN2(g5467), .QN(n14590) );
  NAND2X0 U15561 ( .IN1(n14591), .IN2(g5503), .QN(n14589) );
  NAND3X0 U15562 ( .IN1(n14592), .IN2(n14593), .IN3(n14594), .QN(g25721) );
  NAND2X0 U15563 ( .IN1(n12182), .IN2(g5499), .QN(n14594) );
  NAND2X0 U15564 ( .IN1(n14595), .IN2(g5495), .QN(n14593) );
  NAND2X0 U15565 ( .IN1(n14596), .IN2(n8909), .QN(n14595) );
  NAND2X0 U15566 ( .IN1(n10823), .IN2(g5489), .QN(n14596) );
  NAND4X0 U15567 ( .IN1(n10823), .IN2(n8899), .IN3(n5660), .IN4(n5446), .QN(
        n14592) );
  NAND2X0 U15568 ( .IN1(n14597), .IN2(n14598), .QN(g25720) );
  NAND2X0 U15569 ( .IN1(n12182), .IN2(g5495), .QN(n14598) );
  NAND2X0 U15570 ( .IN1(n14591), .IN2(g5489), .QN(n14597) );
  INVX0 U15571 ( .INP(n12182), .ZN(n14591) );
  NAND3X0 U15572 ( .IN1(n14599), .IN2(n14600), .IN3(n14601), .QN(g25719) );
  NAND2X0 U15573 ( .IN1(n12182), .IN2(g5475), .QN(n14601) );
  NOR2X0 U15574 ( .IN1(n10823), .IN2(n9048), .QN(n12182) );
  NAND3X0 U15575 ( .IN1(n5425), .IN2(n10823), .IN3(n8885), .QN(n14600) );
  NOR2X0 U15576 ( .IN1(n939), .IN2(n5647), .QN(n10823) );
  NAND2X0 U15577 ( .IN1(g5527), .IN2(g5535), .QN(n939) );
  NAND2X0 U15578 ( .IN1(n8987), .IN2(g5471), .QN(n14599) );
  NAND2X0 U15579 ( .IN1(n14602), .IN2(n14603), .QN(g25716) );
  NAND2X0 U15580 ( .IN1(n8987), .IN2(g5456), .QN(n14603) );
  NAND3X0 U15581 ( .IN1(n14604), .IN2(n8090), .IN3(n8885), .QN(n14602) );
  NAND2X0 U15582 ( .IN1(n5992), .IN2(n14605), .QN(n14604) );
  NAND2X0 U15583 ( .IN1(n8525), .IN2(g9555), .QN(n14605) );
  NAND2X0 U15584 ( .IN1(n14606), .IN2(n14607), .QN(g25715) );
  NAND2X0 U15585 ( .IN1(n8903), .IN2(g5689), .QN(n14607) );
  NAND2X0 U15586 ( .IN1(n8987), .IN2(g5406), .QN(n14606) );
  NOR2X0 U15587 ( .IN1(n8949), .IN2(n5566), .QN(g25714) );
  NAND2X0 U15588 ( .IN1(n14608), .IN2(n14609), .QN(g25708) );
  NAND2X0 U15589 ( .IN1(n12268), .IN2(g5120), .QN(n14609) );
  NAND2X0 U15590 ( .IN1(n14610), .IN2(g5156), .QN(n14608) );
  NAND3X0 U15591 ( .IN1(n14611), .IN2(n14612), .IN3(n14613), .QN(g25707) );
  NAND2X0 U15592 ( .IN1(n12268), .IN2(g5152), .QN(n14613) );
  NAND2X0 U15593 ( .IN1(test_so98), .IN2(n14614), .QN(n14612) );
  NAND2X0 U15594 ( .IN1(n14615), .IN2(n8909), .QN(n14614) );
  NAND2X0 U15595 ( .IN1(g32975), .IN2(g5142), .QN(n14615) );
  NAND4X0 U15596 ( .IN1(g32975), .IN2(n8899), .IN3(n5658), .IN4(n8622), .QN(
        n14611) );
  NAND2X0 U15597 ( .IN1(n14616), .IN2(n14617), .QN(g25706) );
  NAND2X0 U15598 ( .IN1(test_so98), .IN2(n12268), .QN(n14617) );
  NAND2X0 U15599 ( .IN1(n14610), .IN2(g5142), .QN(n14616) );
  INVX0 U15600 ( .INP(n12268), .ZN(n14610) );
  NAND3X0 U15601 ( .IN1(n14618), .IN2(n14619), .IN3(n14620), .QN(g25705) );
  NAND2X0 U15602 ( .IN1(test_so96), .IN2(n12268), .QN(n14620) );
  NOR2X0 U15603 ( .IN1(g32975), .IN2(n8931), .QN(n12268) );
  NAND3X0 U15604 ( .IN1(g32975), .IN2(n8601), .IN3(n8885), .QN(n14619) );
  NOR2X0 U15605 ( .IN1(n214), .IN2(n5650), .QN(g32975) );
  NAND2X0 U15606 ( .IN1(g5180), .IN2(g5188), .QN(n214) );
  NAND2X0 U15607 ( .IN1(n8987), .IN2(g5124), .QN(n14618) );
  NOR2X0 U15608 ( .IN1(n8128), .IN2(n14621), .QN(g25704) );
  NOR2X0 U15609 ( .IN1(n8952), .IN2(g5069), .QN(n14621) );
  NAND2X0 U15610 ( .IN1(n14622), .IN2(n14623), .QN(g25703) );
  NAND2X0 U15611 ( .IN1(n8987), .IN2(g5112), .QN(n14623) );
  NAND3X0 U15612 ( .IN1(n5689), .IN2(n14624), .IN3(n8885), .QN(n14622) );
  NAND2X0 U15613 ( .IN1(n8496), .IN2(n14625), .QN(n14624) );
  NAND2X0 U15614 ( .IN1(n8096), .IN2(g9553), .QN(n14625) );
  NAND2X0 U15615 ( .IN1(n14626), .IN2(n14627), .QN(g25702) );
  NAND2X0 U15616 ( .IN1(test_so32), .IN2(n8925), .QN(n14627) );
  NAND3X0 U15617 ( .IN1(n5690), .IN2(n14628), .IN3(n8885), .QN(n14626) );
  NAND2X0 U15618 ( .IN1(n8498), .IN2(n14629), .QN(n14628) );
  INVX0 U15619 ( .INP(n14630), .ZN(n14629) );
  NOR2X0 U15620 ( .IN1(n5689), .IN2(test_so32), .QN(n14630) );
  NAND2X0 U15621 ( .IN1(n14631), .IN2(n14632), .QN(g25701) );
  NAND2X0 U15622 ( .IN1(test_so10), .IN2(n8909), .QN(n14632) );
  NAND2X0 U15623 ( .IN1(n8987), .IN2(g5062), .QN(n14631) );
  NOR2X0 U15624 ( .IN1(n8952), .IN2(n5567), .QN(g25700) );
  NAND3X0 U15625 ( .IN1(n14633), .IN2(n14634), .IN3(n14635), .QN(g25699) );
  NAND2X0 U15626 ( .IN1(n8987), .IN2(g5097), .QN(n14635) );
  INVX0 U15627 ( .INP(n14636), .ZN(n14634) );
  NOR3X0 U15628 ( .IN1(n8926), .IN2(n5014), .IN3(n5669), .QN(n14636) );
  NAND2X0 U15629 ( .IN1(n5014), .IN2(n5669), .QN(n14633) );
  NAND3X0 U15630 ( .IN1(n14637), .IN2(n14638), .IN3(n14639), .QN(g25698) );
  NAND2X0 U15631 ( .IN1(n8986), .IN2(g5092), .QN(n14639) );
  NAND3X0 U15632 ( .IN1(n8895), .IN2(n14640), .IN3(g5097), .QN(n14638) );
  INVX0 U15633 ( .INP(n5016), .ZN(n14640) );
  NAND2X0 U15634 ( .IN1(n5016), .IN2(n5753), .QN(n14637) );
  XOR2X1 U15635 ( .IN1(n14641), .IN2(n5681), .Q(g25697) );
  NAND2X0 U15636 ( .IN1(n8903), .IN2(g5092), .QN(n14641) );
  NAND3X0 U15637 ( .IN1(n14642), .IN2(n14643), .IN3(n14644), .QN(g25696) );
  NAND3X0 U15638 ( .IN1(n8896), .IN2(g5077), .IN3(n8128), .QN(n14644) );
  INVX0 U15639 ( .INP(n14645), .ZN(n14643) );
  NOR2X0 U15640 ( .IN1(n14646), .IN2(n5893), .QN(n14645) );
  NAND3X0 U15641 ( .IN1(n14646), .IN2(n14647), .IN3(n5893), .QN(n14642) );
  NAND2X0 U15642 ( .IN1(n8127), .IN2(g5077), .QN(n14647) );
  NOR2X0 U15643 ( .IN1(g5084), .IN2(n8932), .QN(n14646) );
  NOR2X0 U15644 ( .IN1(n5455), .IN2(n14648), .QN(g25695) );
  NOR3X0 U15645 ( .IN1(n8926), .IN2(n14649), .IN3(n14650), .QN(n14648) );
  NOR2X0 U15646 ( .IN1(g5084), .IN2(g5073), .QN(n14650) );
  NOR2X0 U15647 ( .IN1(n5681), .IN2(g5069), .QN(n14649) );
  NAND2X0 U15648 ( .IN1(n14651), .IN2(n14652), .QN(g25691) );
  NAND2X0 U15649 ( .IN1(n8577), .IN2(n14653), .QN(n14652) );
  NAND4X0 U15650 ( .IN1(n5416), .IN2(test_so11), .IN3(n5711), .IN4(n14654), 
        .QN(n14653) );
  INVX0 U15651 ( .INP(n14655), .ZN(n14654) );
  NAND4X0 U15652 ( .IN1(g4098), .IN2(n10824), .IN3(n5612), .IN4(n8163), .QN(
        n14655) );
  NOR2X0 U15653 ( .IN1(g4093), .IN2(n5480), .QN(n10824) );
  INVX0 U15654 ( .INP(n11495), .ZN(n8577) );
  NAND2X0 U15655 ( .IN1(n8986), .IN2(g4125), .QN(n14651) );
  NAND2X0 U15656 ( .IN1(n14656), .IN2(n14657), .QN(g25690) );
  NAND2X0 U15657 ( .IN1(n8986), .IN2(g4169), .QN(n14657) );
  NAND3X0 U15658 ( .IN1(n8430), .IN2(g25689), .IN3(n8885), .QN(n14656) );
  NAND3X0 U15659 ( .IN1(n14658), .IN2(n14659), .IN3(n14660), .QN(g25687) );
  NAND2X0 U15660 ( .IN1(n8986), .IN2(g4057), .QN(n14660) );
  NAND3X0 U15661 ( .IN1(n14661), .IN2(g4169), .IN3(n5612), .QN(n14659) );
  INVX0 U15662 ( .INP(n1242), .ZN(n14661) );
  NAND2X0 U15663 ( .IN1(g4057), .IN2(g4064), .QN(n1242) );
  NAND2X0 U15664 ( .IN1(n5026), .IN2(n12367), .QN(n14658) );
  NAND2X0 U15665 ( .IN1(n14662), .IN2(n14663), .QN(g25686) );
  NAND2X0 U15666 ( .IN1(n14664), .IN2(g4064), .QN(n14663) );
  NAND2X0 U15667 ( .IN1(n14665), .IN2(n8909), .QN(n14664) );
  NAND2X0 U15668 ( .IN1(n5711), .IN2(g4169), .QN(n14665) );
  NAND3X0 U15669 ( .IN1(n12367), .IN2(g4057), .IN3(n5416), .QN(n14662) );
  NOR2X0 U15670 ( .IN1(n8953), .IN2(n5729), .QN(n12367) );
  NAND3X0 U15671 ( .IN1(n14666), .IN2(n14667), .IN3(n11495), .QN(g25685) );
  NAND2X0 U15672 ( .IN1(n5729), .IN2(n8909), .QN(n11495) );
  NAND2X0 U15673 ( .IN1(n5416), .IN2(n8909), .QN(n14667) );
  NAND2X0 U15674 ( .IN1(n8986), .IN2(g4072), .QN(n14666) );
  NAND2X0 U15675 ( .IN1(n14668), .IN2(n14669), .QN(g25684) );
  NAND2X0 U15676 ( .IN1(n12371), .IN2(g3813), .QN(n14669) );
  NAND2X0 U15677 ( .IN1(n14670), .IN2(g3849), .QN(n14668) );
  NAND3X0 U15678 ( .IN1(n14671), .IN2(n14672), .IN3(n14673), .QN(g25683) );
  NAND2X0 U15679 ( .IN1(n12371), .IN2(g3845), .QN(n14673) );
  NAND2X0 U15680 ( .IN1(test_so97), .IN2(n14674), .QN(n14672) );
  NAND2X0 U15681 ( .IN1(n14675), .IN2(n8910), .QN(n14674) );
  NAND2X0 U15682 ( .IN1(n12372), .IN2(g3835), .QN(n14675) );
  NAND4X0 U15683 ( .IN1(n12372), .IN2(n8900), .IN3(n5662), .IN4(n8623), .QN(
        n14671) );
  NAND2X0 U15684 ( .IN1(n14676), .IN2(n14677), .QN(g25682) );
  NAND2X0 U15685 ( .IN1(test_so97), .IN2(n12371), .QN(n14677) );
  NAND2X0 U15686 ( .IN1(n14670), .IN2(g3835), .QN(n14676) );
  NAND3X0 U15687 ( .IN1(n14678), .IN2(n14679), .IN3(n14680), .QN(g25681) );
  NAND2X0 U15688 ( .IN1(n12371), .IN2(g3821), .QN(n14680) );
  INVX0 U15689 ( .INP(n14670), .ZN(n12371) );
  NAND2X0 U15690 ( .IN1(n10838), .IN2(n8910), .QN(n14670) );
  NAND3X0 U15691 ( .IN1(n5428), .IN2(n12372), .IN3(n8885), .QN(n14679) );
  INVX0 U15692 ( .INP(n10838), .ZN(n12372) );
  NAND2X0 U15693 ( .IN1(test_so33), .IN2(n12392), .QN(n10838) );
  INVX0 U15694 ( .INP(n835), .ZN(n12392) );
  NAND2X0 U15695 ( .IN1(g3873), .IN2(g3881), .QN(n835) );
  NAND2X0 U15696 ( .IN1(n8986), .IN2(g3817), .QN(n14678) );
  NAND2X0 U15697 ( .IN1(n14681), .IN2(n14682), .QN(g25678) );
  NAND2X0 U15698 ( .IN1(n8986), .IN2(g3802), .QN(n14682) );
  NAND3X0 U15699 ( .IN1(n8091), .IN2(n14683), .IN3(n8885), .QN(n14681) );
  NAND2X0 U15700 ( .IN1(n5994), .IN2(n14684), .QN(n14683) );
  NAND2X0 U15701 ( .IN1(n8524), .IN2(g8344), .QN(n14684) );
  NAND2X0 U15702 ( .IN1(n14685), .IN2(n14686), .QN(g25677) );
  NAND2X0 U15703 ( .IN1(n8903), .IN2(g4040), .QN(n14686) );
  NAND2X0 U15704 ( .IN1(n8985), .IN2(g3752), .QN(n14685) );
  NOR2X0 U15705 ( .IN1(n8953), .IN2(n5564), .QN(g25676) );
  NAND2X0 U15706 ( .IN1(n14687), .IN2(n14688), .QN(g25670) );
  NAND2X0 U15707 ( .IN1(n12458), .IN2(g3462), .QN(n14688) );
  NAND2X0 U15708 ( .IN1(n14689), .IN2(g3498), .QN(n14687) );
  NAND3X0 U15709 ( .IN1(n14690), .IN2(n14691), .IN3(n14692), .QN(g25669) );
  NAND2X0 U15710 ( .IN1(n12458), .IN2(g3494), .QN(n14692) );
  NAND2X0 U15711 ( .IN1(n14693), .IN2(g3490), .QN(n14691) );
  NAND2X0 U15712 ( .IN1(n14694), .IN2(n8910), .QN(n14693) );
  NAND2X0 U15713 ( .IN1(n12459), .IN2(g3484), .QN(n14694) );
  NAND4X0 U15714 ( .IN1(n12459), .IN2(n8899), .IN3(n5668), .IN4(n5454), .QN(
        n14690) );
  NAND2X0 U15715 ( .IN1(n14695), .IN2(n14696), .QN(g25668) );
  NAND2X0 U15716 ( .IN1(n12458), .IN2(g3490), .QN(n14696) );
  NAND2X0 U15717 ( .IN1(n14689), .IN2(g3484), .QN(n14695) );
  NAND3X0 U15718 ( .IN1(n14697), .IN2(n14698), .IN3(n14699), .QN(g25667) );
  NAND2X0 U15719 ( .IN1(n12458), .IN2(g3470), .QN(n14699) );
  INVX0 U15720 ( .INP(n14689), .ZN(n12458) );
  NAND2X0 U15721 ( .IN1(n10837), .IN2(n8910), .QN(n14689) );
  NAND3X0 U15722 ( .IN1(n5424), .IN2(n12459), .IN3(n8885), .QN(n14698) );
  INVX0 U15723 ( .INP(n10837), .ZN(n12459) );
  NAND2X0 U15724 ( .IN1(n12479), .IN2(g3518), .QN(n10837) );
  INVX0 U15725 ( .INP(n438), .ZN(n12479) );
  NAND2X0 U15726 ( .IN1(g3522), .IN2(g3530), .QN(n438) );
  NAND2X0 U15727 ( .IN1(n8985), .IN2(g3466), .QN(n14697) );
  NAND2X0 U15728 ( .IN1(n14700), .IN2(n14701), .QN(g25664) );
  NAND2X0 U15729 ( .IN1(n8985), .IN2(g3451), .QN(n14701) );
  NAND3X0 U15730 ( .IN1(n8074), .IN2(n14702), .IN3(n8885), .QN(n14700) );
  NAND2X0 U15731 ( .IN1(n5986), .IN2(n14703), .QN(n14702) );
  NAND2X0 U15732 ( .IN1(n8530), .IN2(g8279), .QN(n14703) );
  NAND2X0 U15733 ( .IN1(n14704), .IN2(n14705), .QN(g25663) );
  NAND2X0 U15734 ( .IN1(n8903), .IN2(g3689), .QN(n14705) );
  NAND2X0 U15735 ( .IN1(n8985), .IN2(g3401), .QN(n14704) );
  NOR2X0 U15736 ( .IN1(n8955), .IN2(n5569), .QN(g25662) );
  NAND2X0 U15737 ( .IN1(n14706), .IN2(n14707), .QN(g25656) );
  NAND2X0 U15738 ( .IN1(n12545), .IN2(g3111), .QN(n14707) );
  NAND2X0 U15739 ( .IN1(n14708), .IN2(g3147), .QN(n14706) );
  NAND3X0 U15740 ( .IN1(n14709), .IN2(n14710), .IN3(n14711), .QN(g25655) );
  NAND2X0 U15741 ( .IN1(n12545), .IN2(g3143), .QN(n14711) );
  NAND2X0 U15742 ( .IN1(n14712), .IN2(g3139), .QN(n14710) );
  NAND2X0 U15743 ( .IN1(n14713), .IN2(n8910), .QN(n14712) );
  NAND2X0 U15744 ( .IN1(n10834), .IN2(g3133), .QN(n14713) );
  NAND4X0 U15745 ( .IN1(n10834), .IN2(n8899), .IN3(n5661), .IN4(n5447), .QN(
        n14709) );
  NAND2X0 U15746 ( .IN1(n14714), .IN2(n14715), .QN(g25654) );
  NAND2X0 U15747 ( .IN1(n12545), .IN2(g3139), .QN(n14715) );
  NAND2X0 U15748 ( .IN1(n14708), .IN2(g3133), .QN(n14714) );
  INVX0 U15749 ( .INP(n12545), .ZN(n14708) );
  NAND3X0 U15750 ( .IN1(n14716), .IN2(n14717), .IN3(n14718), .QN(g25653) );
  NAND2X0 U15751 ( .IN1(n12545), .IN2(g3119), .QN(n14718) );
  NOR2X0 U15752 ( .IN1(n10834), .IN2(n8940), .QN(n12545) );
  NAND3X0 U15753 ( .IN1(n5423), .IN2(n10834), .IN3(n8885), .QN(n14717) );
  NOR2X0 U15754 ( .IN1(n530), .IN2(n5652), .QN(n10834) );
  NAND2X0 U15755 ( .IN1(g3179), .IN2(g3171), .QN(n530) );
  NAND2X0 U15756 ( .IN1(n8985), .IN2(g3115), .QN(n14716) );
  NAND2X0 U15757 ( .IN1(n14719), .IN2(n14720), .QN(g25650) );
  NAND2X0 U15758 ( .IN1(n8985), .IN2(g3100), .QN(n14720) );
  NAND3X0 U15759 ( .IN1(n8097), .IN2(n14721), .IN3(n8885), .QN(n14719) );
  NAND2X0 U15760 ( .IN1(n5998), .IN2(n14722), .QN(n14721) );
  NAND2X0 U15761 ( .IN1(n8522), .IN2(g8215), .QN(n14722) );
  NAND2X0 U15762 ( .IN1(n14723), .IN2(n14724), .QN(g25649) );
  NAND2X0 U15763 ( .IN1(n8902), .IN2(g3338), .QN(n14724) );
  NAND2X0 U15764 ( .IN1(n8985), .IN2(g3050), .QN(n14723) );
  NOR2X0 U15765 ( .IN1(n8953), .IN2(n5390), .QN(g25648) );
  NAND3X0 U15766 ( .IN1(n14725), .IN2(n14726), .IN3(n14727), .QN(g25639) );
  INVX0 U15767 ( .INP(n5045), .ZN(n14727) );
  NAND2X0 U15768 ( .IN1(n8984), .IN2(g2715), .QN(n14726) );
  NAND2X0 U15769 ( .IN1(n12645), .IN2(n8910), .QN(n14725) );
  NOR2X0 U15770 ( .IN1(g2715), .IN2(n5465), .QN(n12645) );
  NAND2X0 U15771 ( .IN1(n14728), .IN2(n14729), .QN(g25638) );
  NAND2X0 U15772 ( .IN1(n8984), .IN2(g1564), .QN(n14729) );
  NAND2X0 U15773 ( .IN1(n14730), .IN2(n8910), .QN(n14728) );
  NAND2X0 U15774 ( .IN1(n14731), .IN2(n14732), .QN(n14730) );
  NAND2X0 U15775 ( .IN1(n14733), .IN2(g1559), .QN(n14732) );
  NAND3X0 U15776 ( .IN1(n14734), .IN2(n5768), .IN3(n5441), .QN(n14731) );
  NAND2X0 U15777 ( .IN1(n14735), .IN2(n14736), .QN(g25637) );
  NAND3X0 U15778 ( .IN1(n8896), .IN2(g1554), .IN3(n14733), .QN(n14736) );
  NAND2X0 U15779 ( .IN1(n14737), .IN2(g1559), .QN(n14735) );
  NAND2X0 U15780 ( .IN1(n14738), .IN2(n8910), .QN(n14737) );
  NAND2X0 U15781 ( .IN1(n14734), .IN2(n5768), .QN(n14738) );
  NAND2X0 U15782 ( .IN1(n14739), .IN2(n14740), .QN(g25636) );
  NAND2X0 U15783 ( .IN1(n8984), .IN2(g1521), .QN(n14740) );
  NAND2X0 U15784 ( .IN1(n14741), .IN2(n8911), .QN(n14739) );
  NAND2X0 U15785 ( .IN1(n14742), .IN2(n14743), .QN(n14741) );
  NAND2X0 U15786 ( .IN1(n13469), .IN2(n12938), .QN(n14743) );
  INVX0 U15787 ( .INP(n14744), .ZN(n12938) );
  NAND2X0 U15788 ( .IN1(n14745), .IN2(g1306), .QN(n14742) );
  NAND2X0 U15789 ( .IN1(n13469), .IN2(g7946), .QN(n14745) );
  INVX0 U15790 ( .INP(n11059), .ZN(n13469) );
  NAND2X0 U15791 ( .IN1(test_so49), .IN2(g1514), .QN(n11059) );
  NAND2X0 U15792 ( .IN1(n14746), .IN2(n14747), .QN(g25635) );
  NAND2X0 U15793 ( .IN1(n14748), .IN2(g1484), .QN(n14747) );
  NAND2X0 U15794 ( .IN1(n14749), .IN2(n8911), .QN(n14748) );
  NAND3X0 U15795 ( .IN1(n5483), .IN2(n13464), .IN3(n14353), .QN(n14749) );
  NAND2X0 U15796 ( .IN1(n14750), .IN2(g1300), .QN(n14746) );
  NAND2X0 U15797 ( .IN1(n14751), .IN2(n14752), .QN(n14750) );
  NAND2X0 U15798 ( .IN1(n14753), .IN2(n8911), .QN(n14752) );
  NAND2X0 U15799 ( .IN1(n14353), .IN2(g1484), .QN(n14753) );
  NOR2X0 U15800 ( .IN1(n8440), .IN2(test_so12), .QN(n14353) );
  NOR3X0 U15801 ( .IN1(n14754), .IN2(test_so68), .IN3(n14368), .QN(g25634) );
  NOR3X0 U15802 ( .IN1(n5655), .IN2(n8501), .IN3(n14755), .QN(n14368) );
  NOR2X0 U15803 ( .IN1(n14756), .IN2(n14757), .QN(n14754) );
  NOR2X0 U15804 ( .IN1(n8501), .IN2(n8939), .QN(n14757) );
  NOR2X0 U15805 ( .IN1(n14755), .IN2(n14758), .QN(n14756) );
  NAND2X0 U15806 ( .IN1(n14759), .IN2(n14760), .QN(g25633) );
  NAND2X0 U15807 ( .IN1(n8984), .IN2(g1379), .QN(n14760) );
  NAND2X0 U15808 ( .IN1(n14761), .IN2(n8911), .QN(n14759) );
  NAND2X0 U15809 ( .IN1(n14762), .IN2(n14763), .QN(n14761) );
  NAND2X0 U15810 ( .IN1(n14764), .IN2(g1384), .QN(n14763) );
  NAND3X0 U15811 ( .IN1(n14374), .IN2(g1351), .IN3(n8055), .QN(n14762) );
  NAND2X0 U15812 ( .IN1(n14765), .IN2(n14766), .QN(g25632) );
  NAND2X0 U15813 ( .IN1(n14767), .IN2(g1312), .QN(n14766) );
  NAND2X0 U15814 ( .IN1(n14764), .IN2(n8911), .QN(n14767) );
  NAND4X0 U15815 ( .IN1(n14768), .IN2(n14769), .IN3(n8898), .IN4(g1351), .QN(
        n14765) );
  NAND2X0 U15816 ( .IN1(n14106), .IN2(n12942), .QN(n14769) );
  NAND2X0 U15817 ( .IN1(n14374), .IN2(g1389), .QN(n14768) );
  NOR2X0 U15818 ( .IN1(n8955), .IN2(n14770), .QN(g25631) );
  NOR2X0 U15819 ( .IN1(n14771), .IN2(n14772), .QN(n14770) );
  NOR2X0 U15820 ( .IN1(n5466), .IN2(n14374), .QN(n14772) );
  INVX0 U15821 ( .INP(n14773), .ZN(n14771) );
  NAND3X0 U15822 ( .IN1(n12942), .IN2(n14774), .IN3(n14775), .QN(n14773) );
  NAND2X0 U15823 ( .IN1(g1351), .IN2(n14776), .QN(n14775) );
  NAND2X0 U15824 ( .IN1(n14102), .IN2(n14106), .QN(n14776) );
  NOR2X0 U15825 ( .IN1(n8171), .IN2(n8172), .QN(n14106) );
  NAND2X0 U15826 ( .IN1(n14105), .IN2(g1389), .QN(n14102) );
  NAND2X0 U15827 ( .IN1(n4896), .IN2(n5322), .QN(n14774) );
  NAND4X0 U15828 ( .IN1(n14107), .IN2(g1367), .IN3(g1345), .IN4(g1379), .QN(
        n4896) );
  NAND2X0 U15829 ( .IN1(n14777), .IN2(n14778), .QN(g25630) );
  NAND2X0 U15830 ( .IN1(n14779), .IN2(g1249), .QN(n14778) );
  NAND2X0 U15831 ( .IN1(n14780), .IN2(n8911), .QN(n14779) );
  NAND2X0 U15832 ( .IN1(n8504), .IN2(g12923), .QN(n14780) );
  NAND2X0 U15833 ( .IN1(g24247), .IN2(g1266), .QN(n14777) );
  NAND2X0 U15834 ( .IN1(n14781), .IN2(n14782), .QN(g25629) );
  NAND2X0 U15835 ( .IN1(n8984), .IN2(g1221), .QN(n14782) );
  NAND2X0 U15836 ( .IN1(n14783), .IN2(n8911), .QN(n14781) );
  NAND2X0 U15837 ( .IN1(n14784), .IN2(n14785), .QN(n14783) );
  NAND2X0 U15838 ( .IN1(n14786), .IN2(g1216), .QN(n14785) );
  NAND3X0 U15839 ( .IN1(n14787), .IN2(n8604), .IN3(n5442), .QN(n14784) );
  NAND2X0 U15840 ( .IN1(n14788), .IN2(n14789), .QN(g25628) );
  NAND3X0 U15841 ( .IN1(n14786), .IN2(n8871), .IN3(test_so76), .QN(n14789) );
  NAND2X0 U15842 ( .IN1(n14790), .IN2(g1216), .QN(n14788) );
  NAND2X0 U15843 ( .IN1(n14791), .IN2(n8911), .QN(n14790) );
  NAND2X0 U15844 ( .IN1(n14787), .IN2(n8604), .QN(n14791) );
  NAND2X0 U15845 ( .IN1(n14792), .IN2(n14793), .QN(g25627) );
  NAND2X0 U15846 ( .IN1(n8984), .IN2(g1178), .QN(n14793) );
  NAND2X0 U15847 ( .IN1(n14794), .IN2(n8911), .QN(n14792) );
  NAND2X0 U15848 ( .IN1(n14795), .IN2(n14796), .QN(n14794) );
  NAND2X0 U15849 ( .IN1(n11219), .IN2(n12973), .QN(n14796) );
  INVX0 U15850 ( .INP(n14797), .ZN(n12973) );
  NAND2X0 U15851 ( .IN1(n14798), .IN2(g962), .QN(n14795) );
  NAND2X0 U15852 ( .IN1(n11219), .IN2(g7916), .QN(n14798) );
  NOR2X0 U15853 ( .IN1(n5599), .IN2(n5363), .QN(n11219) );
  NAND2X0 U15854 ( .IN1(n14799), .IN2(n14800), .QN(g25626) );
  NAND2X0 U15855 ( .IN1(n14801), .IN2(g1141), .QN(n14800) );
  NAND2X0 U15856 ( .IN1(n14802), .IN2(n8911), .QN(n14801) );
  NAND3X0 U15857 ( .IN1(n5341), .IN2(n13500), .IN3(n14390), .QN(n14802) );
  NAND2X0 U15858 ( .IN1(n14803), .IN2(g956), .QN(n14799) );
  NAND2X0 U15859 ( .IN1(n14804), .IN2(n14805), .QN(n14803) );
  NAND2X0 U15860 ( .IN1(n14806), .IN2(n8911), .QN(n14805) );
  NAND2X0 U15861 ( .IN1(n14390), .IN2(g1141), .QN(n14806) );
  NOR2X0 U15862 ( .IN1(g1152), .IN2(n8588), .QN(n14390) );
  NOR3X0 U15863 ( .IN1(g979), .IN2(n14404), .IN3(n14807), .QN(g25625) );
  NOR2X0 U15864 ( .IN1(n14808), .IN2(n14809), .QN(n14807) );
  NOR2X0 U15865 ( .IN1(n8502), .IN2(n8937), .QN(n14809) );
  NOR2X0 U15866 ( .IN1(n14810), .IN2(n9201), .QN(n14808) );
  NOR3X0 U15867 ( .IN1(n5654), .IN2(n8502), .IN3(n14810), .QN(n14404) );
  NAND3X0 U15868 ( .IN1(n14811), .IN2(n14812), .IN3(n14813), .QN(g25624) );
  NAND3X0 U15869 ( .IN1(n14409), .IN2(n8054), .IN3(n14408), .QN(n14813) );
  NAND3X0 U15870 ( .IN1(n14814), .IN2(g1041), .IN3(n8884), .QN(n14812) );
  NAND2X0 U15871 ( .IN1(n8984), .IN2(g1036), .QN(n14811) );
  NAND2X0 U15872 ( .IN1(n14815), .IN2(n14816), .QN(g25623) );
  NAND2X0 U15873 ( .IN1(test_so20), .IN2(n14817), .QN(n14816) );
  NAND2X0 U15874 ( .IN1(n14814), .IN2(n8911), .QN(n14817) );
  NAND2X0 U15875 ( .IN1(n14408), .IN2(n14818), .QN(n14815) );
  NAND2X0 U15876 ( .IN1(n12977), .IN2(n14819), .QN(n14818) );
  NAND2X0 U15877 ( .IN1(n14820), .IN2(n14821), .QN(n14819) );
  NAND2X0 U15878 ( .IN1(g1030), .IN2(g1018), .QN(n14820) );
  NOR2X0 U15879 ( .IN1(n8954), .IN2(n5321), .QN(n14408) );
  NOR2X0 U15880 ( .IN1(n8954), .IN2(n14822), .QN(g25622) );
  NOR2X0 U15881 ( .IN1(n14823), .IN2(n14824), .QN(n14822) );
  NOR2X0 U15882 ( .IN1(n14409), .IN2(n8612), .QN(n14824) );
  NOR2X0 U15883 ( .IN1(n14123), .IN2(n14825), .QN(n14823) );
  NOR2X0 U15884 ( .IN1(n14826), .IN2(n14827), .QN(n14825) );
  NOR2X0 U15885 ( .IN1(n4921), .IN2(g1008), .QN(n14827) );
  NAND4X0 U15886 ( .IN1(n14122), .IN2(g1024), .IN3(g1002), .IN4(g1036), .QN(
        n4921) );
  INVX0 U15887 ( .INP(n14120), .ZN(n14122) );
  NOR2X0 U15888 ( .IN1(n14117), .IN2(n14121), .QN(n14826) );
  NAND3X0 U15889 ( .IN1(g1018), .IN2(g1030), .IN3(g1008), .QN(n14121) );
  INVX0 U15890 ( .INP(n14821), .ZN(n14117) );
  NAND2X0 U15891 ( .IN1(n14120), .IN2(g1046), .QN(n14821) );
  INVX0 U15892 ( .INP(n12977), .ZN(n14123) );
  NAND2X0 U15893 ( .IN1(n14828), .IN2(n14829), .QN(g25621) );
  NAND2X0 U15894 ( .IN1(n14830), .IN2(g904), .QN(n14829) );
  NAND2X0 U15895 ( .IN1(n14831), .IN2(n8912), .QN(n14830) );
  NAND2X0 U15896 ( .IN1(n8505), .IN2(g12919), .QN(n14831) );
  NAND2X0 U15897 ( .IN1(g24231), .IN2(g921), .QN(n14828) );
  NOR2X0 U15898 ( .IN1(n5562), .IN2(n14832), .QN(g25619) );
  NOR2X0 U15899 ( .IN1(n8954), .IN2(n14833), .QN(n14832) );
  XOR2X1 U15900 ( .IN1(n14457), .IN2(g843), .Q(n14833) );
  NAND2X0 U15901 ( .IN1(n14834), .IN2(n14835), .QN(g25618) );
  NAND2X0 U15902 ( .IN1(n14836), .IN2(g817), .QN(n14835) );
  NAND2X0 U15903 ( .IN1(n14837), .IN2(n8912), .QN(n14836) );
  NAND3X0 U15904 ( .IN1(n4948), .IN2(n13521), .IN3(n8519), .QN(n14837) );
  NAND2X0 U15905 ( .IN1(n14838), .IN2(g832), .QN(n14834) );
  NAND2X0 U15906 ( .IN1(n14839), .IN2(n14840), .QN(n14838) );
  NAND2X0 U15907 ( .IN1(n13558), .IN2(n13521), .QN(n14840) );
  NAND2X0 U15908 ( .IN1(n5822), .IN2(n4518), .QN(n14839) );
  INVX0 U15909 ( .INP(n14841), .ZN(n4518) );
  NAND2X0 U15910 ( .IN1(n13521), .IN2(n8912), .QN(n14841) );
  NAND2X0 U15911 ( .IN1(n14842), .IN2(n14843), .QN(g25617) );
  NAND3X0 U15912 ( .IN1(n14844), .IN2(n14845), .IN3(n13521), .QN(n14843) );
  NAND2X0 U15913 ( .IN1(g847), .IN2(n14846), .QN(n13521) );
  NAND2X0 U15914 ( .IN1(n5733), .IN2(g837), .QN(n14846) );
  NAND2X0 U15915 ( .IN1(n14847), .IN2(g817), .QN(n14845) );
  NAND2X0 U15916 ( .IN1(n5822), .IN2(n14848), .QN(n14844) );
  NAND2X0 U15917 ( .IN1(n8998), .IN2(g812), .QN(n14842) );
  NOR2X0 U15918 ( .IN1(n8953), .IN2(n14849), .QN(g25616) );
  XOR3X1 U15919 ( .IN1(n14850), .IN2(n14851), .IN3(n14852), .Q(n14849) );
  XOR2X1 U15920 ( .IN1(n14853), .IN2(g225), .Q(n14852) );
  NOR2X0 U15921 ( .IN1(n5732), .IN2(n14186), .QN(n14853) );
  INVX0 U15922 ( .INP(n14854), .ZN(n14186) );
  NAND4X0 U15923 ( .IN1(n5327), .IN2(n14164), .IN3(n14168), .IN4(n14855), .QN(
        n14854) );
  NOR3X0 U15924 ( .IN1(g370), .IN2(g490), .IN3(g482), .QN(n14855) );
  NOR2X0 U15925 ( .IN1(g518), .IN2(test_so54), .QN(n14168) );
  XOR2X1 U15926 ( .IN1(g255), .IN2(n6008), .Q(n14851) );
  XOR3X1 U15927 ( .IN1(n8189), .IN2(n8188), .IN3(n14856), .Q(n14850) );
  XOR2X1 U15928 ( .IN1(n8309), .IN2(n8308), .Q(n14856) );
  NAND2X0 U15929 ( .IN1(n14857), .IN2(n14858), .QN(g25615) );
  NAND2X0 U15930 ( .IN1(n14859), .IN2(g667), .QN(n14858) );
  NAND2X0 U15931 ( .IN1(n14153), .IN2(g686), .QN(n14857) );
  NAND3X0 U15932 ( .IN1(n14860), .IN2(n14861), .IN3(n14862), .QN(g25614) );
  NAND2X0 U15933 ( .IN1(n8982), .IN2(g691), .QN(n14862) );
  NAND2X0 U15934 ( .IN1(n14859), .IN2(g686), .QN(n14861) );
  NAND2X0 U15935 ( .IN1(n5111), .IN2(n14863), .QN(n14860) );
  NAND2X0 U15936 ( .IN1(n14864), .IN2(n14865), .QN(g25613) );
  NAND2X0 U15937 ( .IN1(n8983), .IN2(g559), .QN(n14865) );
  NAND3X0 U15938 ( .IN1(n2421), .IN2(n14866), .IN3(n14867), .QN(n14864) );
  XOR2X1 U15939 ( .IN1(g562), .IN2(n14472), .Q(n14867) );
  INVX0 U15940 ( .INP(n14868), .ZN(n14472) );
  NAND2X0 U15941 ( .IN1(g29211), .IN2(n14869), .QN(n14868) );
  NAND2X0 U15942 ( .IN1(n8045), .IN2(g12368), .QN(n14869) );
  NAND2X0 U15943 ( .IN1(g626), .IN2(n9340), .QN(n14866) );
  NAND2X0 U15944 ( .IN1(n14870), .IN2(n14871), .QN(g25612) );
  NAND2X0 U15945 ( .IN1(n14872), .IN2(g513), .QN(n14871) );
  NAND2X0 U15946 ( .IN1(n14859), .IN2(g518), .QN(n14870) );
  NAND2X0 U15947 ( .IN1(n14873), .IN2(n14874), .QN(g25611) );
  NAND2X0 U15948 ( .IN1(n14872), .IN2(g504), .QN(n14874) );
  NAND2X0 U15949 ( .IN1(n14875), .IN2(n8912), .QN(n14872) );
  NAND2X0 U15950 ( .IN1(n14863), .IN2(n13551), .QN(n14875) );
  INVX0 U15951 ( .INP(n4962), .ZN(n13551) );
  INVX0 U15952 ( .INP(n14478), .ZN(n14863) );
  NAND2X0 U15953 ( .IN1(n14859), .IN2(g513), .QN(n14873) );
  NAND3X0 U15954 ( .IN1(n14876), .IN2(n14877), .IN3(n14878), .QN(g25610) );
  NAND2X0 U15955 ( .IN1(n14859), .IN2(g504), .QN(n14877) );
  INVX0 U15956 ( .INP(n14153), .ZN(n14859) );
  NAND2X0 U15957 ( .IN1(test_so54), .IN2(n14153), .QN(n14876) );
  NAND3X0 U15958 ( .IN1(n14879), .IN2(n14878), .IN3(n14880), .QN(g25609) );
  NAND2X0 U15959 ( .IN1(n14155), .IN2(n5287), .QN(n14880) );
  NAND2X0 U15960 ( .IN1(n4962), .IN2(n14155), .QN(n14878) );
  NOR2X0 U15961 ( .IN1(n14478), .IN2(n8933), .QN(n14155) );
  NAND2X0 U15962 ( .IN1(test_so54), .IN2(n14881), .QN(n14879) );
  NAND2X0 U15963 ( .IN1(n14153), .IN2(n14882), .QN(n14881) );
  NAND2X0 U15964 ( .IN1(n5548), .IN2(n8912), .QN(n14882) );
  NAND2X0 U15965 ( .IN1(n14478), .IN2(n8912), .QN(n14153) );
  NAND3X0 U15966 ( .IN1(g385), .IN2(g358), .IN3(n5633), .QN(n14478) );
  NAND3X0 U15967 ( .IN1(n14883), .IN2(n14884), .IN3(n14885), .QN(g25605) );
  NAND2X0 U15968 ( .IN1(n8979), .IN2(g168), .QN(n14885) );
  NAND3X0 U15969 ( .IN1(n14164), .IN2(g246), .IN3(n14886), .QN(n14884) );
  NAND2X0 U15970 ( .IN1(n14887), .IN2(g460), .QN(n14883) );
  NAND2X0 U15971 ( .IN1(n14888), .IN2(n14889), .QN(g25604) );
  NAND2X0 U15972 ( .IN1(n14887), .IN2(g452), .QN(n14889) );
  NAND2X0 U15973 ( .IN1(n14890), .IN2(g460), .QN(n14888) );
  NAND3X0 U15974 ( .IN1(n14891), .IN2(n14892), .IN3(n14893), .QN(g25602) );
  NAND2X0 U15975 ( .IN1(n8978), .IN2(g405), .QN(n14893) );
  NAND3X0 U15976 ( .IN1(n14164), .IN2(g446), .IN3(n14886), .QN(n14892) );
  NAND2X0 U15977 ( .IN1(n14887), .IN2(test_so72), .QN(n14891) );
  NAND2X0 U15978 ( .IN1(n14894), .IN2(n14895), .QN(g25601) );
  NAND2X0 U15979 ( .IN1(n14887), .IN2(g174), .QN(n14895) );
  NAND2X0 U15980 ( .IN1(test_so72), .IN2(n14890), .QN(n14894) );
  NAND2X0 U15981 ( .IN1(n14896), .IN2(n14897), .QN(g25600) );
  NAND2X0 U15982 ( .IN1(n14887), .IN2(g168), .QN(n14897) );
  INVX0 U15983 ( .INP(n14890), .ZN(n14887) );
  NAND2X0 U15984 ( .IN1(n14890), .IN2(g174), .QN(n14896) );
  NAND2X0 U15985 ( .IN1(n14898), .IN2(n8912), .QN(n14890) );
  NAND2X0 U15986 ( .IN1(n8539), .IN2(n14164), .QN(n14898) );
  INVX0 U15987 ( .INP(n1161), .ZN(n14164) );
  NAND2X0 U15988 ( .IN1(n10040), .IN2(n14899), .QN(g25599) );
  NAND2X0 U15989 ( .IN1(n8981), .IN2(g385), .QN(n14899) );
  NAND2X0 U15990 ( .IN1(n14900), .IN2(n14901), .QN(g25598) );
  NAND3X0 U15991 ( .IN1(n8896), .IN2(g385), .IN3(n1161), .QN(n14901) );
  NAND2X0 U15992 ( .IN1(n14902), .IN2(g376), .QN(n14900) );
  NAND2X0 U15993 ( .IN1(n14903), .IN2(n8912), .QN(n14902) );
  NAND2X0 U15994 ( .IN1(n1161), .IN2(g358), .QN(n14903) );
  NAND3X0 U15995 ( .IN1(g376), .IN2(g358), .IN3(g385), .QN(n1161) );
  NAND3X0 U15996 ( .IN1(n14904), .IN2(n14905), .IN3(n14906), .QN(g25597) );
  NAND2X0 U15997 ( .IN1(n14907), .IN2(n14886), .QN(n14906) );
  NOR2X0 U15998 ( .IN1(g370), .IN2(n8932), .QN(n14886) );
  INVX0 U15999 ( .INP(n10040), .ZN(n14907) );
  NAND3X0 U16000 ( .IN1(n10040), .IN2(g370), .IN3(n8884), .QN(n14905) );
  NAND3X0 U16001 ( .IN1(g376), .IN2(g8719), .IN3(g385), .QN(n10040) );
  NAND2X0 U16002 ( .IN1(n8980), .IN2(g358), .QN(n14904) );
  NAND2X0 U16003 ( .IN1(n14908), .IN2(n14909), .QN(g25596) );
  NAND2X0 U16004 ( .IN1(n8992), .IN2(g370), .QN(n14909) );
  NAND2X0 U16005 ( .IN1(n14910), .IN2(n8912), .QN(n14908) );
  XOR2X1 U16006 ( .IN1(n8190), .IN2(n5633), .Q(n14910) );
  NOR3X0 U16007 ( .IN1(g8719), .IN2(n8925), .IN3(g358), .QN(g25595) );
  NAND2X0 U16008 ( .IN1(n14911), .IN2(n14912), .QN(g25593) );
  NAND2X0 U16009 ( .IN1(n8991), .IN2(g191), .QN(n14912) );
  NAND2X0 U16010 ( .IN1(n14913), .IN2(n8912), .QN(n14911) );
  NAND2X0 U16011 ( .IN1(n14914), .IN2(n14915), .QN(n14913) );
  NAND2X0 U16012 ( .IN1(n14916), .IN2(g209), .QN(n14915) );
  NAND2X0 U16013 ( .IN1(n14917), .IN2(n14918), .QN(n14914) );
  INVX0 U16014 ( .INP(n14916), .ZN(n14918) );
  NAND2X0 U16015 ( .IN1(n14919), .IN2(n14920), .QN(g25592) );
  NAND2X0 U16016 ( .IN1(n8993), .IN2(g222), .QN(n14920) );
  NAND2X0 U16017 ( .IN1(n14921), .IN2(n8912), .QN(n14919) );
  XNOR2X1 U16018 ( .IN1(n8169), .IN2(n14922), .Q(n14921) );
  NOR2X0 U16019 ( .IN1(n14916), .IN2(n14917), .QN(n14922) );
  XOR2X1 U16020 ( .IN1(n8169), .IN2(n8170), .Q(n14917) );
  NAND2X0 U16021 ( .IN1(test_so42), .IN2(g218), .QN(n14916) );
  NAND2X0 U16022 ( .IN1(n14923), .IN2(n14924), .QN(g25591) );
  NAND2X0 U16023 ( .IN1(n8441), .IN2(n8912), .QN(n14924) );
  NAND2X0 U16024 ( .IN1(n8994), .IN2(g209), .QN(n14923) );
  NOR2X0 U16025 ( .IN1(g1636), .IN2(n5598), .QN(g25259) );
  INVX0 U16026 ( .INP(n10231), .ZN(g25167) );
  NAND2X0 U16027 ( .IN1(n5525), .IN2(test_so94), .QN(n10231) );
  NOR2X0 U16028 ( .IN1(n8433), .IN2(n14925), .QN(g24355) );
  NOR2X0 U16029 ( .IN1(n8952), .IN2(n14926), .QN(n14925) );
  NAND2X0 U16030 ( .IN1(n14927), .IN2(n14928), .QN(g24354) );
  NAND2X0 U16031 ( .IN1(n8996), .IN2(g6727), .QN(n14928) );
  NAND3X0 U16032 ( .IN1(n8432), .IN2(n14926), .IN3(n8884), .QN(n14927) );
  NAND2X0 U16033 ( .IN1(n14929), .IN2(g6727), .QN(n14926) );
  NAND2X0 U16034 ( .IN1(n14930), .IN2(n14931), .QN(g24353) );
  NAND2X0 U16035 ( .IN1(n8995), .IN2(g6723), .QN(n14931) );
  NAND2X0 U16036 ( .IN1(n14932), .IN2(n8912), .QN(n14930) );
  XOR2X1 U16037 ( .IN1(n14929), .IN2(g6727), .Q(n14932) );
  NOR4X0 U16038 ( .IN1(n8592), .IN2(n5700), .IN3(n8276), .IN4(n8290), .QN(
        n14929) );
  NOR4X0 U16039 ( .IN1(n14933), .IN2(g13099), .IN3(n14934), .IN4(n14935), .QN(
        g24352) );
  NOR2X0 U16040 ( .IN1(test_so80), .IN2(n5700), .QN(n14935) );
  NOR2X0 U16041 ( .IN1(n8290), .IN2(g14828), .QN(n14934) );
  NAND3X0 U16042 ( .IN1(n8276), .IN2(n8871), .IN3(n8391), .QN(n14933) );
  NOR2X0 U16043 ( .IN1(n8299), .IN2(n14936), .QN(g24351) );
  NOR2X0 U16044 ( .IN1(n8950), .IN2(n14937), .QN(n14936) );
  NAND2X0 U16045 ( .IN1(n14938), .IN2(n14939), .QN(g24350) );
  NAND2X0 U16046 ( .IN1(test_so69), .IN2(n9052), .QN(n14939) );
  NAND3X0 U16047 ( .IN1(n8298), .IN2(n14937), .IN3(n8884), .QN(n14938) );
  NAND2X0 U16048 ( .IN1(n14940), .IN2(test_so69), .QN(n14937) );
  NAND2X0 U16049 ( .IN1(n14941), .IN2(n14942), .QN(g24349) );
  NAND2X0 U16050 ( .IN1(n8997), .IN2(g6377), .QN(n14942) );
  NAND2X0 U16051 ( .IN1(n14943), .IN2(n8913), .QN(n14941) );
  XOR2X1 U16052 ( .IN1(test_so69), .IN2(n14940), .Q(n14943) );
  NOR4X0 U16053 ( .IN1(n5437), .IN2(n5703), .IN3(n8279), .IN4(n8294), .QN(
        n14940) );
  NOR4X0 U16054 ( .IN1(n14944), .IN2(g13085), .IN3(n14945), .IN4(n14946), .QN(
        g24348) );
  NOR2X0 U16055 ( .IN1(n5703), .IN2(g12422), .QN(n14946) );
  NOR2X0 U16056 ( .IN1(n8294), .IN2(g14779), .QN(n14945) );
  NAND3X0 U16057 ( .IN1(n8279), .IN2(n8870), .IN3(n8401), .QN(n14944) );
  NOR2X0 U16058 ( .IN1(n8300), .IN2(n14947), .QN(g24347) );
  NOR2X0 U16059 ( .IN1(n8951), .IN2(n14948), .QN(n14947) );
  NAND2X0 U16060 ( .IN1(n14949), .IN2(n14950), .QN(g24346) );
  NAND2X0 U16061 ( .IN1(n8974), .IN2(g6035), .QN(n14950) );
  NAND3X0 U16062 ( .IN1(n14948), .IN2(n8610), .IN3(n8884), .QN(n14949) );
  NAND2X0 U16063 ( .IN1(n14951), .IN2(g6035), .QN(n14948) );
  NAND2X0 U16064 ( .IN1(n14952), .IN2(n14953), .QN(g24345) );
  NAND2X0 U16065 ( .IN1(n8975), .IN2(g6031), .QN(n14953) );
  NAND2X0 U16066 ( .IN1(n14954), .IN2(n8913), .QN(n14952) );
  XOR2X1 U16067 ( .IN1(g6035), .IN2(n14951), .Q(n14954) );
  NOR4X0 U16068 ( .IN1(n5432), .IN2(n5698), .IN3(n8270), .IN4(n8285), .QN(
        n14951) );
  NOR4X0 U16069 ( .IN1(n14955), .IN2(g13068), .IN3(n14956), .IN4(n14957), .QN(
        g24344) );
  NOR2X0 U16070 ( .IN1(n5698), .IN2(g12350), .QN(n14957) );
  NOR2X0 U16071 ( .IN1(n8285), .IN2(g14738), .QN(n14956) );
  NAND3X0 U16072 ( .IN1(n8270), .IN2(n8870), .IN3(n8377), .QN(n14955) );
  NOR2X0 U16073 ( .IN1(n8304), .IN2(n14958), .QN(g24343) );
  NOR2X0 U16074 ( .IN1(n8951), .IN2(n14959), .QN(n14958) );
  NAND2X0 U16075 ( .IN1(n14960), .IN2(n14961), .QN(g24342) );
  NAND2X0 U16076 ( .IN1(n8969), .IN2(g5689), .QN(n14961) );
  NAND3X0 U16077 ( .IN1(n8303), .IN2(n14959), .IN3(n8884), .QN(n14960) );
  NAND2X0 U16078 ( .IN1(n14962), .IN2(g5689), .QN(n14959) );
  NAND2X0 U16079 ( .IN1(n14963), .IN2(n14964), .QN(g24341) );
  NAND2X0 U16080 ( .IN1(n8968), .IN2(g5685), .QN(n14964) );
  NAND2X0 U16081 ( .IN1(n14965), .IN2(n8906), .QN(n14963) );
  XOR2X1 U16082 ( .IN1(g5689), .IN2(n14962), .Q(n14965) );
  NOR4X0 U16083 ( .IN1(n5439), .IN2(n5705), .IN3(n8272), .IN4(n8287), .QN(
        n14962) );
  NOR4X0 U16084 ( .IN1(n14966), .IN2(g13049), .IN3(n14967), .IN4(n14968), .QN(
        g24340) );
  NOR2X0 U16085 ( .IN1(n5705), .IN2(g12300), .QN(n14968) );
  NOR2X0 U16086 ( .IN1(n8287), .IN2(g14694), .QN(n14967) );
  NAND3X0 U16087 ( .IN1(n8272), .IN2(n8870), .IN3(n8382), .QN(n14966) );
  NOR2X0 U16088 ( .IN1(n8435), .IN2(n14969), .QN(g24339) );
  NOR2X0 U16089 ( .IN1(n8949), .IN2(n14970), .QN(n14969) );
  NAND2X0 U16090 ( .IN1(n14971), .IN2(n14972), .QN(g24338) );
  NAND2X0 U16091 ( .IN1(test_so10), .IN2(n9052), .QN(n14972) );
  NAND3X0 U16092 ( .IN1(n8434), .IN2(n14970), .IN3(n8884), .QN(n14971) );
  NAND2X0 U16093 ( .IN1(n14973), .IN2(test_so10), .QN(n14970) );
  NAND2X0 U16094 ( .IN1(n14974), .IN2(n14975), .QN(g24337) );
  NAND2X0 U16095 ( .IN1(n8967), .IN2(g5339), .QN(n14975) );
  NAND2X0 U16096 ( .IN1(n14976), .IN2(n8912), .QN(n14974) );
  XOR2X1 U16097 ( .IN1(test_so10), .IN2(n14973), .Q(n14976) );
  NOR4X0 U16098 ( .IN1(n5438), .IN2(n5704), .IN3(n8268), .IN4(n8283), .QN(
        n14973) );
  NOR4X0 U16099 ( .IN1(n14977), .IN2(g17577), .IN3(n14978), .IN4(n14979), .QN(
        g24336) );
  NOR2X0 U16100 ( .IN1(n5704), .IN2(g12238), .QN(n14979) );
  NOR2X0 U16101 ( .IN1(n8283), .IN2(g14662), .QN(n14978) );
  NAND3X0 U16102 ( .IN1(n8268), .IN2(n8870), .IN3(n8351), .QN(n14977) );
  NAND2X0 U16103 ( .IN1(n14980), .IN2(n14981), .QN(g24335) );
  NAND3X0 U16104 ( .IN1(n5653), .IN2(g4643), .IN3(n14982), .QN(n14981) );
  INVX0 U16105 ( .INP(n14983), .ZN(n14982) );
  NAND2X0 U16106 ( .IN1(n8990), .IN2(g18881), .QN(n14980) );
  NAND2X0 U16107 ( .IN1(n14984), .IN2(n14985), .QN(g24334) );
  NAND4X0 U16108 ( .IN1(n5303), .IN2(n5365), .IN3(n14986), .IN4(n14987), .QN(
        n14985) );
  NOR4X0 U16109 ( .IN1(g4584), .IN2(g4608), .IN3(g4616), .IN4(n14983), .QN(
        n14987) );
  NAND4X0 U16110 ( .IN1(n8902), .IN2(n8590), .IN3(n5506), .IN4(n14988), .QN(
        n14983) );
  NOR3X0 U16111 ( .IN1(g4358), .IN2(g4332), .IN3(g4311), .QN(n14988) );
  NOR3X0 U16112 ( .IN1(n10178), .IN2(n5844), .IN3(n5653), .QN(n14986) );
  NAND2X0 U16113 ( .IN1(test_so3), .IN2(n5727), .QN(n10178) );
  NAND2X0 U16114 ( .IN1(n8989), .IN2(g4358), .QN(n14984) );
  NOR2X0 U16115 ( .IN1(n5710), .IN2(n8898), .QN(g24298) );
  NAND2X0 U16116 ( .IN1(n14989), .IN2(n14990), .QN(g24282) );
  NAND2X0 U16117 ( .IN1(n14991), .IN2(g4308), .QN(n14990) );
  NAND2X0 U16118 ( .IN1(n8905), .IN2(g9251), .QN(n14991) );
  NAND2X0 U16119 ( .IN1(g24281), .IN2(g9251), .QN(n14989) );
  NOR2X0 U16120 ( .IN1(g4308), .IN2(n8930), .QN(g24281) );
  NAND2X0 U16121 ( .IN1(n14992), .IN2(n14993), .QN(g24280) );
  NAND2X0 U16122 ( .IN1(n14994), .IN2(g4269), .QN(n14993) );
  NAND2X0 U16123 ( .IN1(n14995), .IN2(n8912), .QN(n14994) );
  NAND3X0 U16124 ( .IN1(g4264), .IN2(g4258), .IN3(n5764), .QN(n14995) );
  NAND2X0 U16125 ( .IN1(n14996), .IN2(g4273), .QN(n14992) );
  NAND2X0 U16126 ( .IN1(n14997), .IN2(n14998), .QN(n14996) );
  NAND2X0 U16127 ( .IN1(n5763), .IN2(n8912), .QN(n14998) );
  NAND3X0 U16128 ( .IN1(n14999), .IN2(n15000), .IN3(n15001), .QN(g24279) );
  NAND2X0 U16129 ( .IN1(n15002), .IN2(n15003), .QN(n15001) );
  NAND2X0 U16130 ( .IN1(n9003), .IN2(g4235), .QN(n15000) );
  NAND2X0 U16131 ( .IN1(n15004), .IN2(n8911), .QN(n14999) );
  NAND2X0 U16132 ( .IN1(n15005), .IN2(n15006), .QN(n15004) );
  INVX0 U16133 ( .INP(n15007), .ZN(n15006) );
  NOR3X0 U16134 ( .IN1(n15003), .IN2(n15002), .IN3(n15008), .QN(n15007) );
  NOR2X0 U16135 ( .IN1(n8232), .IN2(n5726), .QN(n15002) );
  NAND2X0 U16136 ( .IN1(n15008), .IN2(n15003), .QN(n15005) );
  INVX0 U16137 ( .INP(n15009), .ZN(n15008) );
  NAND3X0 U16138 ( .IN1(n5726), .IN2(n15010), .IN3(n8232), .QN(n15009) );
  NAND4X0 U16139 ( .IN1(n15231), .IN2(n15232), .IN3(n15230), .IN4(n15011), 
        .QN(n15010) );
  NOR4X0 U16140 ( .IN1(g8915), .IN2(g8916), .IN3(g11770), .IN4(g8920), .QN(
        n15011) );
  NOR2X0 U16141 ( .IN1(n8306), .IN2(n15012), .QN(g24278) );
  NOR2X0 U16142 ( .IN1(n8951), .IN2(n15013), .QN(n15012) );
  NAND2X0 U16143 ( .IN1(n15014), .IN2(n15015), .QN(g24277) );
  NAND2X0 U16144 ( .IN1(n8970), .IN2(g4040), .QN(n15015) );
  NAND3X0 U16145 ( .IN1(n8305), .IN2(n15013), .IN3(n8884), .QN(n15014) );
  NAND2X0 U16146 ( .IN1(n15016), .IN2(g4040), .QN(n15013) );
  NAND2X0 U16147 ( .IN1(n15017), .IN2(n15018), .QN(g24276) );
  NAND2X0 U16148 ( .IN1(n8971), .IN2(g4031), .QN(n15018) );
  NAND2X0 U16149 ( .IN1(n15019), .IN2(n8911), .QN(n15017) );
  XOR2X1 U16150 ( .IN1(g4040), .IN2(n15016), .Q(n15019) );
  NOR4X0 U16151 ( .IN1(n5435), .IN2(n5701), .IN3(n8274), .IN4(n8288), .QN(
        n15016) );
  NOR4X0 U16152 ( .IN1(n15020), .IN2(g14518), .IN3(n15021), .IN4(n15022), .QN(
        g24275) );
  NOR2X0 U16153 ( .IN1(n5701), .IN2(g11418), .QN(n15022) );
  NOR2X0 U16154 ( .IN1(n8288), .IN2(g13966), .QN(n15021) );
  NAND3X0 U16155 ( .IN1(n8274), .IN2(n8870), .IN3(n8386), .QN(n15020) );
  NOR2X0 U16156 ( .IN1(n8302), .IN2(n15023), .QN(g24274) );
  NOR2X0 U16157 ( .IN1(n8948), .IN2(n15024), .QN(n15023) );
  NAND2X0 U16158 ( .IN1(n15025), .IN2(n15026), .QN(g24273) );
  NAND2X0 U16159 ( .IN1(n8977), .IN2(g3689), .QN(n15026) );
  NAND3X0 U16160 ( .IN1(n8301), .IN2(n15024), .IN3(n8884), .QN(n15025) );
  NAND2X0 U16161 ( .IN1(n15027), .IN2(g3689), .QN(n15024) );
  NAND2X0 U16162 ( .IN1(n15028), .IN2(n15029), .QN(g24272) );
  NAND2X0 U16163 ( .IN1(n8976), .IN2(g3680), .QN(n15029) );
  NAND2X0 U16164 ( .IN1(n15030), .IN2(n8911), .QN(n15028) );
  XOR2X1 U16165 ( .IN1(g3689), .IN2(n15027), .Q(n15030) );
  NOR4X0 U16166 ( .IN1(n5433), .IN2(n5699), .IN3(n8278), .IN4(n8292), .QN(
        n15027) );
  NOR4X0 U16167 ( .IN1(n15031), .IN2(g14451), .IN3(n15032), .IN4(n15033), .QN(
        g24271) );
  NOR2X0 U16168 ( .IN1(n5699), .IN2(g11388), .QN(n15033) );
  NOR2X0 U16169 ( .IN1(n8292), .IN2(g13926), .QN(n15032) );
  NAND3X0 U16170 ( .IN1(n8278), .IN2(n8869), .IN3(n8396), .QN(n15031) );
  NOR2X0 U16171 ( .IN1(n8297), .IN2(n15034), .QN(g24270) );
  NOR2X0 U16172 ( .IN1(n8948), .IN2(n15035), .QN(n15034) );
  NAND2X0 U16173 ( .IN1(n15036), .IN2(n15037), .QN(g24269) );
  NAND2X0 U16174 ( .IN1(n8973), .IN2(g3338), .QN(n15037) );
  NAND3X0 U16175 ( .IN1(n8296), .IN2(n15035), .IN3(n8884), .QN(n15036) );
  NAND2X0 U16176 ( .IN1(n15038), .IN2(g3338), .QN(n15035) );
  NAND2X0 U16177 ( .IN1(n15039), .IN2(n15040), .QN(g24268) );
  NAND2X0 U16178 ( .IN1(test_so91), .IN2(n8962), .QN(n15040) );
  NAND2X0 U16179 ( .IN1(n15041), .IN2(n8910), .QN(n15039) );
  XOR2X1 U16180 ( .IN1(g3338), .IN2(n15038), .Q(n15041) );
  NOR4X0 U16181 ( .IN1(n5436), .IN2(n5702), .IN3(n8266), .IN4(n8281), .QN(
        n15038) );
  NOR4X0 U16182 ( .IN1(n15042), .IN2(g14421), .IN3(n15043), .IN4(n15044), .QN(
        g24267) );
  NOR2X0 U16183 ( .IN1(n5702), .IN2(g11349), .QN(n15044) );
  NOR2X0 U16184 ( .IN1(n8281), .IN2(g13895), .QN(n15043) );
  NAND3X0 U16185 ( .IN1(n8266), .IN2(n8869), .IN3(n8367), .QN(n15042) );
  NAND2X0 U16186 ( .IN1(n15045), .IN2(n15046), .QN(g24266) );
  INVX0 U16187 ( .INP(n15047), .ZN(n15046) );
  NOR2X0 U16188 ( .IN1(n8900), .IN2(n5963), .QN(n15047) );
  NAND3X0 U16189 ( .IN1(test_so9), .IN2(n8083), .IN3(n8884), .QN(n15045) );
  NAND3X0 U16190 ( .IN1(n15048), .IN2(n15049), .IN3(n9200), .QN(g24263) );
  NAND2X0 U16191 ( .IN1(n5963), .IN2(n8910), .QN(n9200) );
  NAND2X0 U16192 ( .IN1(n5299), .IN2(n8910), .QN(n15049) );
  NAND2X0 U16193 ( .IN1(n8972), .IN2(g2712), .QN(n15048) );
  NAND3X0 U16194 ( .IN1(n15050), .IN2(n15051), .IN3(n15052), .QN(g24262) );
  NAND2X0 U16195 ( .IN1(n15053), .IN2(n8443), .QN(n15052) );
  NAND3X0 U16196 ( .IN1(n15054), .IN2(g1564), .IN3(n8884), .QN(n15051) );
  INVX0 U16197 ( .INP(n15053), .ZN(n15054) );
  NAND2X0 U16198 ( .IN1(n9002), .IN2(g1548), .QN(n15050) );
  NAND2X0 U16199 ( .IN1(n14758), .IN2(n15055), .QN(g24261) );
  NAND2X0 U16200 ( .IN1(n9001), .IN2(g1585), .QN(n15055) );
  XOR2X1 U16201 ( .IN1(n15056), .IN2(n8444), .Q(g24260) );
  NAND2X0 U16202 ( .IN1(n8906), .IN2(g1548), .QN(n15056) );
  NAND2X0 U16203 ( .IN1(n14758), .IN2(n15057), .QN(g24259) );
  NAND2X0 U16204 ( .IN1(n9006), .IN2(g1579), .QN(n15057) );
  NAND2X0 U16205 ( .IN1(n15058), .IN2(n15059), .QN(g24258) );
  NAND2X0 U16206 ( .IN1(n8905), .IN2(g496), .QN(n15059) );
  NAND2X0 U16207 ( .IN1(n9005), .IN2(g1554), .QN(n15058) );
  XNOR2X1 U16208 ( .IN1(n15060), .IN2(n5616), .Q(g24257) );
  NOR2X0 U16209 ( .IN1(n15061), .IN2(n8929), .QN(n15060) );
  NAND2X0 U16210 ( .IN1(n15062), .IN2(n15063), .QN(g24256) );
  NAND2X0 U16211 ( .IN1(n8999), .IN2(g1339), .QN(n15063) );
  NAND2X0 U16212 ( .IN1(n15064), .IN2(n8909), .QN(n15062) );
  XOR2X1 U16213 ( .IN1(n15061), .IN2(n15065), .Q(n15064) );
  NAND3X0 U16214 ( .IN1(n8520), .IN2(n14755), .IN3(n8521), .QN(n15065) );
  INVX0 U16215 ( .INP(n15066), .ZN(n14755) );
  NAND3X0 U16216 ( .IN1(n5302), .IN2(n5616), .IN3(n5401), .QN(n15066) );
  NAND3X0 U16217 ( .IN1(n14374), .IN2(n15067), .IN3(n15068), .QN(n15061) );
  XOR2X1 U16218 ( .IN1(g1579), .IN2(test_so68), .Q(n15068) );
  NAND3X0 U16219 ( .IN1(n15069), .IN2(n15070), .IN3(n15071), .QN(g24255) );
  NAND2X0 U16220 ( .IN1(n11311), .IN2(g17423), .QN(n15071) );
  NAND3X0 U16221 ( .IN1(n8159), .IN2(g10527), .IN3(n8883), .QN(n15070) );
  NAND2X0 U16222 ( .IN1(n9000), .IN2(g1589), .QN(n15069) );
  INVX0 U16223 ( .INP(n15072), .ZN(g24254) );
  NAND4X0 U16224 ( .IN1(n8159), .IN2(n15073), .IN3(n8160), .IN4(n8161), .QN(
        n15072) );
  INVX0 U16225 ( .INP(n15074), .ZN(n15073) );
  NAND2X0 U16226 ( .IN1(n15075), .IN2(n8909), .QN(n15074) );
  NAND3X0 U16227 ( .IN1(n15076), .IN2(g1554), .IN3(n14734), .QN(n15075) );
  INVX0 U16228 ( .INP(n14733), .ZN(n14734) );
  NAND2X0 U16229 ( .IN1(n15053), .IN2(g1564), .QN(n14733) );
  NOR2X0 U16230 ( .IN1(n8444), .IN2(n5546), .QN(n15053) );
  NAND2X0 U16231 ( .IN1(n14374), .IN2(n15067), .QN(n15076) );
  INVX0 U16232 ( .INP(n1376), .ZN(n15067) );
  NAND2X0 U16233 ( .IN1(n5466), .IN2(n5322), .QN(n1376) );
  INVX0 U16234 ( .INP(n14764), .ZN(n14374) );
  NAND2X0 U16235 ( .IN1(n14105), .IN2(n12942), .QN(n14764) );
  NAND2X0 U16236 ( .IN1(n5616), .IN2(n8602), .QN(n12942) );
  INVX0 U16237 ( .INP(n14107), .ZN(n14105) );
  XNOR2X1 U16238 ( .IN1(g1339), .IN2(test_so68), .Q(n14107) );
  NAND2X0 U16239 ( .IN1(n15077), .IN2(n15078), .QN(g24253) );
  NAND2X0 U16240 ( .IN1(n9004), .IN2(g1306), .QN(n15078) );
  NAND2X0 U16241 ( .IN1(n15079), .IN2(n8909), .QN(n15077) );
  NAND2X0 U16242 ( .IN1(n15080), .IN2(n15081), .QN(n15079) );
  NAND2X0 U16243 ( .IN1(n5302), .IN2(g1532), .QN(n15081) );
  NAND2X0 U16244 ( .IN1(g7946), .IN2(g1521), .QN(n15080) );
  NAND2X0 U16245 ( .IN1(n15082), .IN2(n15083), .QN(g24252) );
  NAND2X0 U16246 ( .IN1(test_so49), .IN2(n8955), .QN(n15083) );
  NAND2X0 U16247 ( .IN1(n15084), .IN2(n8909), .QN(n15082) );
  NAND2X0 U16248 ( .IN1(n14744), .IN2(n15085), .QN(n15084) );
  NAND2X0 U16249 ( .IN1(n5302), .IN2(g1521), .QN(n15085) );
  NAND2X0 U16250 ( .IN1(g7946), .IN2(g1339), .QN(n14744) );
  NAND2X0 U16251 ( .IN1(n15086), .IN2(n15087), .QN(g24251) );
  NAND2X0 U16252 ( .IN1(n13460), .IN2(g1442), .QN(n15087) );
  NAND2X0 U16253 ( .IN1(test_so12), .IN2(n14751), .QN(n15086) );
  NAND2X0 U16254 ( .IN1(n15088), .IN2(n15089), .QN(g24250) );
  NAND2X0 U16255 ( .IN1(test_so12), .IN2(n13460), .QN(n15089) );
  NAND2X0 U16256 ( .IN1(n14751), .IN2(g1489), .QN(n15088) );
  NAND2X0 U16257 ( .IN1(n15090), .IN2(n15091), .QN(g24249) );
  NAND3X0 U16258 ( .IN1(n8440), .IN2(n8869), .IN3(n13464), .QN(n15091) );
  NAND2X0 U16259 ( .IN1(n15092), .IN2(g1489), .QN(n15090) );
  NAND2X0 U16260 ( .IN1(n14751), .IN2(n15093), .QN(n15092) );
  NAND2X0 U16261 ( .IN1(n8906), .IN2(n8632), .QN(n15093) );
  INVX0 U16262 ( .INP(n13460), .ZN(n14751) );
  NOR2X0 U16263 ( .IN1(n13464), .IN2(n8933), .QN(n13460) );
  NOR3X0 U16264 ( .IN1(n8521), .IN2(test_so49), .IN3(g1514), .QN(n13464) );
  NAND3X0 U16265 ( .IN1(n15094), .IN2(n15095), .IN3(n15096), .QN(g24248) );
  XNOR2X1 U16266 ( .IN1(n8167), .IN2(n15097), .Q(n15096) );
  NAND2X0 U16267 ( .IN1(n5655), .IN2(n8909), .QN(n15097) );
  NAND2X0 U16268 ( .IN1(n11311), .IN2(g1395), .QN(n15095) );
  INVX0 U16269 ( .INP(n14758), .ZN(n11311) );
  NAND2X0 U16270 ( .IN1(n5401), .IN2(n8909), .QN(n15094) );
  NOR2X0 U16271 ( .IN1(g1249), .IN2(n14758), .QN(g24247) );
  NAND2X0 U16272 ( .IN1(n8906), .IN2(g12923), .QN(n14758) );
  NAND3X0 U16273 ( .IN1(n15098), .IN2(n15099), .IN3(n15100), .QN(g24246) );
  NAND2X0 U16274 ( .IN1(n15101), .IN2(n8445), .QN(n15100) );
  NAND3X0 U16275 ( .IN1(n15102), .IN2(g1221), .IN3(n8883), .QN(n15099) );
  INVX0 U16276 ( .INP(n15101), .ZN(n15102) );
  NAND2X0 U16277 ( .IN1(n9009), .IN2(g1205), .QN(n15098) );
  NAND2X0 U16278 ( .IN1(n9201), .IN2(n15103), .QN(g24245) );
  NAND2X0 U16279 ( .IN1(n9016), .IN2(g30332), .QN(n15103) );
  XOR2X1 U16280 ( .IN1(n15104), .IN2(n8446), .Q(g24244) );
  NAND2X0 U16281 ( .IN1(n8906), .IN2(g1205), .QN(n15104) );
  NAND2X0 U16282 ( .IN1(n15105), .IN2(n15106), .QN(g24242) );
  NAND2X0 U16283 ( .IN1(n8906), .IN2(g29215), .QN(n15106) );
  NAND2X0 U16284 ( .IN1(test_so76), .IN2(n8954), .QN(n15105) );
  XNOR2X1 U16285 ( .IN1(n15107), .IN2(n5622), .Q(g24241) );
  NOR2X0 U16286 ( .IN1(n15108), .IN2(n8929), .QN(n15107) );
  NAND2X0 U16287 ( .IN1(n15109), .IN2(n15110), .QN(g24240) );
  NAND2X0 U16288 ( .IN1(n9015), .IN2(g996), .QN(n15110) );
  NAND2X0 U16289 ( .IN1(n15111), .IN2(n8909), .QN(n15109) );
  XOR2X1 U16290 ( .IN1(n15108), .IN2(n15112), .Q(n15111) );
  NAND3X0 U16291 ( .IN1(n8526), .IN2(n14810), .IN3(n8527), .QN(n15112) );
  INVX0 U16292 ( .INP(n15113), .ZN(n14810) );
  NAND3X0 U16293 ( .IN1(n5304), .IN2(n5622), .IN3(n5392), .QN(n15113) );
  NAND3X0 U16294 ( .IN1(n15114), .IN2(n14191), .IN3(n14409), .QN(n15108) );
  XOR2X1 U16295 ( .IN1(n8152), .IN2(n5320), .Q(n15114) );
  NAND3X0 U16296 ( .IN1(n15115), .IN2(n15116), .IN3(n15117), .QN(g24239) );
  INVX0 U16297 ( .INP(n15118), .ZN(n15117) );
  NOR2X0 U16298 ( .IN1(n9201), .IN2(n8155), .QN(n15118) );
  NAND3X0 U16299 ( .IN1(n8155), .IN2(g10500), .IN3(n8883), .QN(n15116) );
  NAND2X0 U16300 ( .IN1(n9014), .IN2(g1246), .QN(n15115) );
  INVX0 U16301 ( .INP(n15119), .ZN(g24238) );
  NAND4X0 U16302 ( .IN1(n15120), .IN2(n15121), .IN3(n8155), .IN4(n8150), .QN(
        n15119) );
  NOR2X0 U16303 ( .IN1(n8951), .IN2(test_so44), .QN(n15121) );
  NAND3X0 U16304 ( .IN1(test_so76), .IN2(n15122), .IN3(n14787), .QN(n15120) );
  INVX0 U16305 ( .INP(n14786), .ZN(n14787) );
  NAND2X0 U16306 ( .IN1(n15101), .IN2(g1221), .QN(n14786) );
  NOR2X0 U16307 ( .IN1(n8446), .IN2(n5547), .QN(n15101) );
  NAND2X0 U16308 ( .IN1(n14191), .IN2(n14409), .QN(n15122) );
  INVX0 U16309 ( .INP(n14814), .ZN(n14409) );
  NAND2X0 U16310 ( .IN1(n14120), .IN2(n12977), .QN(n14814) );
  NAND2X0 U16311 ( .IN1(n5622), .IN2(n5320), .QN(n12977) );
  XNOR2X1 U16312 ( .IN1(g996), .IN2(n5320), .Q(n14120) );
  NOR2X0 U16313 ( .IN1(g1008), .IN2(test_so20), .QN(n14191) );
  NAND2X0 U16314 ( .IN1(n15123), .IN2(n15124), .QN(g24237) );
  NAND2X0 U16315 ( .IN1(n9013), .IN2(g962), .QN(n15124) );
  NAND2X0 U16316 ( .IN1(n15125), .IN2(n8908), .QN(n15123) );
  NAND2X0 U16317 ( .IN1(n15126), .IN2(n15127), .QN(n15125) );
  NAND2X0 U16318 ( .IN1(n5304), .IN2(g1189), .QN(n15127) );
  NAND2X0 U16319 ( .IN1(g7916), .IN2(g1178), .QN(n15126) );
  NAND2X0 U16320 ( .IN1(n15128), .IN2(n15129), .QN(g24236) );
  NAND2X0 U16321 ( .IN1(n9012), .IN2(g1183), .QN(n15129) );
  NAND2X0 U16322 ( .IN1(n15130), .IN2(n8908), .QN(n15128) );
  NAND2X0 U16323 ( .IN1(n14797), .IN2(n15131), .QN(n15130) );
  NAND2X0 U16324 ( .IN1(n5304), .IN2(g1178), .QN(n15131) );
  NAND2X0 U16325 ( .IN1(g7916), .IN2(g996), .QN(n14797) );
  NAND2X0 U16326 ( .IN1(n15132), .IN2(n15133), .QN(g24235) );
  NAND2X0 U16327 ( .IN1(test_so7), .IN2(n13496), .QN(n15133) );
  NAND2X0 U16328 ( .IN1(n14804), .IN2(g1152), .QN(n15132) );
  NAND2X0 U16329 ( .IN1(n15134), .IN2(n15135), .QN(g24234) );
  NAND2X0 U16330 ( .IN1(n13496), .IN2(g1152), .QN(n15135) );
  NAND2X0 U16331 ( .IN1(n14804), .IN2(g1146), .QN(n15134) );
  NAND2X0 U16332 ( .IN1(n15136), .IN2(n15137), .QN(g24233) );
  NAND3X0 U16333 ( .IN1(n8897), .IN2(n8588), .IN3(n13500), .QN(n15137) );
  NAND2X0 U16334 ( .IN1(n15138), .IN2(g1146), .QN(n15136) );
  NAND2X0 U16335 ( .IN1(n14804), .IN2(n15139), .QN(n15138) );
  NAND2X0 U16336 ( .IN1(n5618), .IN2(n8908), .QN(n15139) );
  INVX0 U16337 ( .INP(n13496), .ZN(n14804) );
  NOR2X0 U16338 ( .IN1(n13500), .IN2(n8932), .QN(n13496) );
  NOR3X0 U16339 ( .IN1(g1171), .IN2(n8527), .IN3(g1183), .QN(n13500) );
  NAND3X0 U16340 ( .IN1(n15140), .IN2(n15141), .IN3(n15142), .QN(g24232) );
  XNOR2X1 U16341 ( .IN1(n8168), .IN2(n15143), .Q(n15142) );
  NAND2X0 U16342 ( .IN1(n5654), .IN2(n8907), .QN(n15143) );
  NAND2X0 U16343 ( .IN1(n11325), .IN2(g1052), .QN(n15141) );
  INVX0 U16344 ( .INP(n9201), .ZN(n11325) );
  NAND2X0 U16345 ( .IN1(n5392), .IN2(n8908), .QN(n15140) );
  NOR2X0 U16346 ( .IN1(g904), .IN2(n9201), .QN(g24231) );
  NAND2X0 U16347 ( .IN1(n8906), .IN2(g12919), .QN(n9201) );
  NAND2X0 U16348 ( .IN1(n15144), .IN2(n15145), .QN(g24216) );
  NAND2X0 U16349 ( .IN1(n13558), .IN2(g847), .QN(n15145) );
  NAND2X0 U16350 ( .IN1(n14847), .IN2(g854), .QN(n15144) );
  NAND2X0 U16351 ( .IN1(n15146), .IN2(n15147), .QN(g24215) );
  NAND2X0 U16352 ( .IN1(n15148), .IN2(g837), .QN(n15147) );
  NAND2X0 U16353 ( .IN1(n14847), .IN2(n15149), .QN(n15148) );
  NAND3X0 U16354 ( .IN1(n15150), .IN2(n8869), .IN3(n15151), .QN(n15149) );
  NAND2X0 U16355 ( .IN1(g827), .IN2(g832), .QN(n15151) );
  NAND2X0 U16356 ( .IN1(g847), .IN2(g812), .QN(n15150) );
  NAND2X0 U16357 ( .IN1(n15152), .IN2(g703), .QN(n15146) );
  NAND2X0 U16358 ( .IN1(n15153), .IN2(n8907), .QN(n15152) );
  NAND2X0 U16359 ( .IN1(n5562), .IN2(n14457), .QN(n15153) );
  NOR2X0 U16360 ( .IN1(n13562), .IN2(n5709), .QN(n14457) );
  NAND3X0 U16361 ( .IN1(n15154), .IN2(n15155), .IN3(n15156), .QN(g24214) );
  NAND2X0 U16362 ( .IN1(n15157), .IN2(g703), .QN(n15156) );
  NAND2X0 U16363 ( .IN1(n14453), .IN2(n15158), .QN(n15157) );
  NAND2X0 U16364 ( .IN1(n15159), .IN2(n8907), .QN(n15158) );
  INVX0 U16365 ( .INP(n14451), .ZN(n15159) );
  NOR2X0 U16366 ( .IN1(n5733), .IN2(n5562), .QN(n14451) );
  NOR2X0 U16367 ( .IN1(n13558), .IN2(n15160), .QN(n14453) );
  NOR2X0 U16368 ( .IN1(g847), .IN2(n8930), .QN(n15160) );
  NAND2X0 U16369 ( .IN1(n9011), .IN2(g847), .QN(n15155) );
  NAND4X0 U16370 ( .IN1(g817), .IN2(g723), .IN3(n15161), .IN4(n5709), .QN(
        n15154) );
  NOR2X0 U16371 ( .IN1(n5422), .IN2(n14848), .QN(n15161) );
  NAND2X0 U16372 ( .IN1(n15162), .IN2(n15163), .QN(g24211) );
  NAND2X0 U16373 ( .IN1(n2404), .IN2(n15164), .QN(n15163) );
  NAND2X0 U16374 ( .IN1(n8634), .IN2(g691), .QN(n15164) );
  NAND2X0 U16375 ( .IN1(n9020), .IN2(g546), .QN(n15162) );
  NOR3X0 U16376 ( .IN1(n12999), .IN2(n8925), .IN3(n15165), .QN(g24210) );
  NOR2X0 U16377 ( .IN1(n15166), .IN2(n15167), .QN(n15165) );
  NOR2X0 U16378 ( .IN1(n5606), .IN2(n5402), .QN(n15167) );
  NOR2X0 U16379 ( .IN1(n12998), .IN2(n8593), .QN(n15166) );
  NOR2X0 U16380 ( .IN1(g168), .IN2(g174), .QN(n12998) );
  NAND3X0 U16381 ( .IN1(g518), .IN2(g203), .IN3(n5548), .QN(n12999) );
  NAND2X0 U16382 ( .IN1(n15168), .IN2(n15169), .QN(g24209) );
  NAND2X0 U16383 ( .IN1(n13563), .IN2(g446), .QN(n15169) );
  NAND2X0 U16384 ( .IN1(n13558), .IN2(g417), .QN(n15168) );
  NAND3X0 U16385 ( .IN1(n15170), .IN2(n15171), .IN3(n15172), .QN(g24208) );
  NAND2X0 U16386 ( .IN1(n9019), .IN2(g424), .QN(n15172) );
  NAND2X0 U16387 ( .IN1(n13563), .IN2(g246), .QN(n15171) );
  NAND2X0 U16388 ( .IN1(n13558), .IN2(g475), .QN(n15170) );
  NAND2X0 U16389 ( .IN1(n15173), .IN2(n15174), .QN(g24207) );
  NAND2X0 U16390 ( .IN1(n13558), .IN2(g441), .QN(n15174) );
  NAND2X0 U16391 ( .IN1(n14847), .IN2(g475), .QN(n15173) );
  NAND2X0 U16392 ( .IN1(n15175), .IN2(n15176), .QN(g24206) );
  NAND2X0 U16393 ( .IN1(n13558), .IN2(g437), .QN(n15176) );
  NAND2X0 U16394 ( .IN1(n14847), .IN2(g441), .QN(n15175) );
  NAND3X0 U16395 ( .IN1(n15177), .IN2(n15178), .IN3(n15179), .QN(g24205) );
  NAND2X0 U16396 ( .IN1(n9024), .IN2(g437), .QN(n15179) );
  NAND2X0 U16397 ( .IN1(n13563), .IN2(g269), .QN(n15178) );
  NAND2X0 U16398 ( .IN1(test_so23), .IN2(n13558), .QN(n15177) );
  NAND2X0 U16399 ( .IN1(n15180), .IN2(n15181), .QN(g24204) );
  NAND2X0 U16400 ( .IN1(n13558), .IN2(g429), .QN(n15181) );
  NAND2X0 U16401 ( .IN1(test_so23), .IN2(n14847), .QN(n15180) );
  NAND2X0 U16402 ( .IN1(n15182), .IN2(n15183), .QN(g24203) );
  NAND2X0 U16403 ( .IN1(n13558), .IN2(g401), .QN(n15183) );
  NAND2X0 U16404 ( .IN1(n14847), .IN2(g429), .QN(n15182) );
  NAND2X0 U16405 ( .IN1(n15184), .IN2(n15185), .QN(g24202) );
  NAND2X0 U16406 ( .IN1(n13558), .IN2(g424), .QN(n15185) );
  NAND2X0 U16407 ( .IN1(n14847), .IN2(g411), .QN(n15184) );
  NAND2X0 U16408 ( .IN1(n15186), .IN2(n15187), .QN(g24201) );
  NAND2X0 U16409 ( .IN1(n13558), .IN2(g405), .QN(n15187) );
  NAND2X0 U16410 ( .IN1(n14847), .IN2(g392), .QN(n15186) );
  NAND3X0 U16411 ( .IN1(n15188), .IN2(n15189), .IN3(n15190), .QN(g24200) );
  NAND2X0 U16412 ( .IN1(n9023), .IN2(g401), .QN(n15190) );
  NAND3X0 U16413 ( .IN1(n5821), .IN2(g854), .IN3(n13563), .QN(n15189) );
  INVX0 U16414 ( .INP(n14848), .ZN(n13563) );
  NAND2X0 U16415 ( .IN1(n4948), .IN2(n8907), .QN(n14848) );
  NAND2X0 U16416 ( .IN1(n13558), .IN2(g392), .QN(n15188) );
  INVX0 U16417 ( .INP(n14847), .ZN(n13558) );
  NAND2X0 U16418 ( .IN1(n8905), .IN2(n13562), .QN(n14847) );
  INVX0 U16419 ( .INP(n4948), .ZN(n13562) );
  NOR2X0 U16420 ( .IN1(g22), .IN2(g25), .QN(g23190) );
  NAND2X0 U16421 ( .IN1(n15191), .IN2(n15192), .QN(g21901) );
  NAND2X0 U16422 ( .IN1(n9008), .IN2(g2946), .QN(n15192) );
  NAND2X0 U16423 ( .IN1(n15193), .IN2(n8907), .QN(n15191) );
  NAND2X0 U16424 ( .IN1(n15194), .IN2(n15195), .QN(n15193) );
  NAND2X0 U16425 ( .IN1(n5694), .IN2(g4180), .QN(n15195) );
  NAND2X0 U16426 ( .IN1(n5380), .IN2(n15196), .QN(n15194) );
  NAND2X0 U16427 ( .IN1(n5694), .IN2(n15197), .QN(n15196) );
  NAND4X0 U16428 ( .IN1(n15234), .IN2(n8177), .IN3(n15233), .IN4(n15198), .QN(
        n15197) );
  NOR4X0 U16429 ( .IN1(test_so86), .IN2(test_so39), .IN3(g8787), .IN4(g8788), 
        .QN(n15198) );
  NAND2X0 U16430 ( .IN1(n15199), .IN2(n15200), .QN(g21900) );
  NAND2X0 U16431 ( .IN1(n9007), .IN2(g4239), .QN(n15200) );
  NAND3X0 U16432 ( .IN1(n8087), .IN2(n8086), .IN3(n8883), .QN(n15199) );
  XOR2X1 U16433 ( .IN1(n15201), .IN2(n8472), .Q(g21899) );
  NAND2X0 U16434 ( .IN1(n8906), .IN2(g9019), .QN(n15201) );
  NAND2X0 U16435 ( .IN1(n15202), .IN2(n15203), .QN(g21898) );
  NAND2X0 U16436 ( .IN1(n8472), .IN2(n8908), .QN(n15203) );
  INVX0 U16437 ( .INP(n15204), .ZN(n15202) );
  NOR2X0 U16438 ( .IN1(n8900), .IN2(n8511), .QN(n15204) );
  XOR2X1 U16439 ( .IN1(n15205), .IN2(n8473), .Q(g21897) );
  NAND2X0 U16440 ( .IN1(n8905), .IN2(g8839), .QN(n15205) );
  NAND2X0 U16441 ( .IN1(n15206), .IN2(n15207), .QN(g21896) );
  NAND2X0 U16442 ( .IN1(n8473), .IN2(n8906), .QN(n15207) );
  NAND2X0 U16443 ( .IN1(n9010), .IN2(g4245), .QN(n15206) );
  NAND2X0 U16444 ( .IN1(n15208), .IN2(n15209), .QN(g21895) );
  NAND2X0 U16445 ( .IN1(n15210), .IN2(g4264), .QN(n15209) );
  NAND2X0 U16446 ( .IN1(n15211), .IN2(n8908), .QN(n15210) );
  NAND2X0 U16447 ( .IN1(n5763), .IN2(g4258), .QN(n15211) );
  NAND2X0 U16448 ( .IN1(n15212), .IN2(g4269), .QN(n15208) );
  INVX0 U16449 ( .INP(n14997), .ZN(n15212) );
  NOR2X0 U16450 ( .IN1(g21893), .IN2(n15213), .QN(n14997) );
  NOR2X0 U16451 ( .IN1(g4264), .IN2(n8928), .QN(n15213) );
  NAND2X0 U16452 ( .IN1(n15214), .IN2(n15215), .QN(g21894) );
  NAND2X0 U16453 ( .IN1(n15216), .IN2(g4258), .QN(n15215) );
  NAND2X0 U16454 ( .IN1(n8905), .IN2(g4264), .QN(n15216) );
  NAND2X0 U16455 ( .IN1(g21893), .IN2(g4264), .QN(n15214) );
  NOR2X0 U16456 ( .IN1(g4258), .IN2(n8924), .QN(g21893) );
  NAND2X0 U16457 ( .IN1(n15217), .IN2(n15218), .QN(g21892) );
  NAND2X0 U16458 ( .IN1(n8142), .IN2(n8907), .QN(n15218) );
  NAND2X0 U16459 ( .IN1(n9031), .IN2(g4273), .QN(n15217) );
  NAND2X0 U16460 ( .IN1(n15219), .IN2(n15220), .QN(g21891) );
  NAND2X0 U16461 ( .IN1(n9050), .IN2(g4180), .QN(n15220) );
  NAND2X0 U16462 ( .IN1(n15003), .IN2(n8906), .QN(n15219) );
  NAND2X0 U16463 ( .IN1(n15221), .IN2(n15222), .QN(n15003) );
  NAND2X0 U16464 ( .IN1(n8450), .IN2(g4253), .QN(n15222) );
  NAND2X0 U16465 ( .IN1(n8449), .IN2(n5484), .QN(n15221) );
  NOR2X0 U16466 ( .IN1(n8900), .IN2(DFF_1381_n1), .QN(g21727) );
  NOR2X0 U16467 ( .IN1(n5750), .IN2(n8898), .QN(g18597) );
  INVX0 U16468 ( .INP(g5), .ZN(g12833) );
  NOR2X0 U5116_U2 ( .IN1(g34783), .IN2(n2730), .QN(U5116_n1) );
  INVX0 U5116_U1 ( .INP(U5116_n1), .ZN(g34221) );
  NOR2X0 U5126_U2 ( .IN1(n1376), .IN2(n4896), .QN(U5126_n1) );
  INVX0 U5126_U1 ( .INP(U5126_n1), .ZN(n4895) );
  NOR2X0 U5127_U2 ( .IN1(n4837), .IN2(n4921), .QN(U5127_n1) );
  INVX0 U5127_U1 ( .INP(U5127_n1), .ZN(n4920) );
  NOR2X0 U5128_U2 ( .IN1(n807), .IN2(n1249), .QN(U5128_n1) );
  INVX0 U5128_U1 ( .INP(U5128_n1), .ZN(n5045) );
  NOR2X0 U5129_U2 ( .IN1(g559), .IN2(g9048), .QN(U5129_n1) );
  INVX0 U5129_U1 ( .INP(U5129_n1), .ZN(n4959) );
  INVX0 U5353_U2 ( .INP(n5960), .ZN(U5353_n1) );
  NOR2X0 U5353_U1 ( .IN1(n8575), .IN2(U5353_n1), .QN(n4689) );
  INVX0 U5355_U2 ( .INP(n5961), .ZN(U5355_n1) );
  NOR2X0 U5355_U1 ( .IN1(n8570), .IN2(U5355_n1), .QN(n4708) );
  INVX0 U5961_U2 ( .INP(n3593), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3589), .IN2(U5961_n1), .QN(n3595) );
  INVX0 U5962_U2 ( .INP(n3574), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3570), .IN2(U5962_n1), .QN(n3576) );
  INVX0 U5963_U2 ( .INP(n3517), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3513), .IN2(U5963_n1), .QN(n3519) );
  INVX0 U5964_U2 ( .INP(n3628), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3624), .IN2(U5964_n1), .QN(n3630) );
  INVX0 U5965_U2 ( .INP(n3555), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3551), .IN2(U5965_n1), .QN(n3557) );
  INVX0 U5966_U2 ( .INP(n3646), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3642), .IN2(U5966_n1), .QN(n3648) );
  INVX0 U5967_U2 ( .INP(n3536), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3532), .IN2(U5967_n1), .QN(n3538) );
  INVX0 U5968_U2 ( .INP(n3611), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3607), .IN2(U5968_n1), .QN(n3613) );
  INVX0 U6100_U2 ( .INP(n3635), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n8946), .IN2(U6100_n1), .QN(n4888) );
  INVX0 U6211_U2 ( .INP(n3623), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n1721), .IN2(U6211_n1), .QN(n3622) );
  INVX0 U6212_U2 ( .INP(n3587), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3588), .IN2(U6212_n1), .QN(n3586) );
  INVX0 U6213_U2 ( .INP(n3605), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3606), .IN2(U6213_n1), .QN(n3604) );
  INVX0 U6214_U2 ( .INP(n3568), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3569), .IN2(U6214_n1), .QN(n3567) );
  INVX0 U6215_U2 ( .INP(n3549), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3550), .IN2(U6215_n1), .QN(n3548) );
  INVX0 U6216_U2 ( .INP(n3512), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3006), .IN2(U6216_n1), .QN(n3511) );
  INVX0 U6217_U2 ( .INP(n3531), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3007), .IN2(U6217_n1), .QN(n3530) );
  INVX0 U6218_U2 ( .INP(n3641), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n3003), .IN2(U6218_n1), .QN(n3640) );
  INVX0 U6279_U2 ( .INP(n4537), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5337), .IN2(U6279_n1), .QN(n4201) );
  INVX0 U6280_U2 ( .INP(n4201), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5336), .IN2(U6280_n1), .QN(n3745) );
  INVX0 U6281_U2 ( .INP(n3745), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5294), .IN2(U6281_n1), .QN(n3684) );
  INVX0 U6282_U2 ( .INP(n3684), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5552), .IN2(U6282_n1), .QN(n3274) );
  INVX0 U6283_U2 ( .INP(n3274), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5472), .IN2(U6283_n1), .QN(n2982) );
  INVX0 U6284_U2 ( .INP(n2982), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5476), .IN2(U6284_n1), .QN(n2706) );
  INVX0 U6285_U2 ( .INP(n2706), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5550), .IN2(U6285_n1), .QN(n2649) );
  INVX0 U6286_U2 ( .INP(n2649), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5473), .IN2(U6286_n1), .QN(n2556) );
  INVX0 U6287_U2 ( .INP(n2556), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5475), .IN2(U6287_n1), .QN(n2509) );
  INVX0 U6288_U2 ( .INP(n2509), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5474), .IN2(U6288_n1), .QN(n2487) );
  INVX0 U6289_U2 ( .INP(n2487), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5339), .IN2(U6289_n1), .QN(n2427) );
  INVX0 U6290_U2 ( .INP(n2427), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5672), .IN2(U6290_n1), .QN(n2423) );
  INVX0 U6291_U2 ( .INP(n5), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5335), .IN2(U6291_n1), .QN(n4537) );
  INVX0 U6292_U2 ( .INP(n4959), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n8948), .IN2(U6292_n1), .QN(n2421) );
  INVX0 U6338_U2 ( .INP(n4210), .ZN(U6338_n1) );
  NOR2X1 U6338_U1 ( .IN1(n8944), .IN2(U6338_n1), .QN(n3765) );
  INVX0 U6341_U2 ( .INP(n3765), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n1135), .IN2(U6341_n1), .QN(n3951) );
  INVX0 U6342_U2 ( .INP(n3765), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n750), .IN2(U6342_n1), .QN(n3774) );
  INVX0 U6343_U2 ( .INP(n3765), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n1073), .IN2(U6343_n1), .QN(n3842) );
  INVX0 U6344_U2 ( .INP(n3765), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n1009), .IN2(U6344_n1), .QN(n3808) );
  INVX0 U6345_U2 ( .INP(n3765), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n744), .IN2(U6345_n1), .QN(n3908) );
  INVX0 U6346_U2 ( .INP(n3765), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n99), .IN2(U6346_n1), .QN(n3984) );
  INVX0 U6347_U2 ( .INP(n3765), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n494), .IN2(U6347_n1), .QN(n3875) );
  INVX0 U6348_U2 ( .INP(n3765), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n112), .IN2(U6348_n1), .QN(n4015) );
  INVX0 U6349_U2 ( .INP(n3765), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n746), .IN2(U6349_n1), .QN(n3914) );
  INVX0 U6350_U2 ( .INP(n3765), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n752), .IN2(U6350_n1), .QN(n3780) );
  INVX0 U6351_U2 ( .INP(n3765), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n1136), .IN2(U6351_n1), .QN(n3957) );
  INVX0 U6352_U2 ( .INP(n3765), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n1074), .IN2(U6352_n1), .QN(n3848) );
  INVX0 U6353_U2 ( .INP(n3765), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n100), .IN2(U6353_n1), .QN(n3990) );
  INVX0 U6354_U2 ( .INP(n3765), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n1010), .IN2(U6354_n1), .QN(n3814) );
  INVX0 U6355_U2 ( .INP(n3765), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n496), .IN2(U6355_n1), .QN(n3881) );
  INVX0 U6356_U2 ( .INP(n3765), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n114), .IN2(U6356_n1), .QN(n4022) );
  INVX0 U6357_U2 ( .INP(n3765), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n113), .IN2(U6357_n1), .QN(n4027) );
  INVX0 U6358_U2 ( .INP(n3765), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n751), .IN2(U6358_n1), .QN(n3785) );
  INVX0 U6359_U2 ( .INP(n3765), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n1137), .IN2(U6359_n1), .QN(n3962) );
  INVX0 U6360_U2 ( .INP(n3765), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n1075), .IN2(U6360_n1), .QN(n3853) );
  INVX0 U6361_U2 ( .INP(n3765), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n495), .IN2(U6361_n1), .QN(n3886) );
  INVX0 U6362_U2 ( .INP(n3765), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n1011), .IN2(U6362_n1), .QN(n3819) );
  INVX0 U6363_U2 ( .INP(n3765), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n101), .IN2(U6363_n1), .QN(n3995) );
  INVX0 U6364_U2 ( .INP(n3765), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n745), .IN2(U6364_n1), .QN(n3919) );
  INVX0 U6365_U2 ( .INP(n3682), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5471), .IN2(U6365_n1), .QN(n3272) );
  INVX0 U6366_U2 ( .INP(n3272), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5331), .IN2(U6366_n1), .QN(n2980) );
  INVX0 U6367_U2 ( .INP(n2980), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5332), .IN2(U6367_n1), .QN(n2704) );
  INVX0 U6368_U2 ( .INP(n2704), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5333), .IN2(U6368_n1), .QN(n2647) );
  INVX0 U6369_U2 ( .INP(n2647), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5334), .IN2(U6369_n1), .QN(n2554) );
  INVX0 U6370_U2 ( .INP(n2554), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5330), .IN2(U6370_n1), .QN(n2507) );
  INVX0 U6371_U2 ( .INP(n2507), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5551), .IN2(U6371_n1), .QN(n2485) );
  INVX0 U6372_U2 ( .INP(n2485), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5293), .IN2(U6372_n1), .QN(n2425) );
  INVX0 U6373_U2 ( .INP(n2425), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5292), .IN2(U6373_n1), .QN(n2419) );
  INVX0 U6374_U2 ( .INP(n55), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5470), .IN2(U6374_n1), .QN(n3682) );
  INVX0 U6375_U2 ( .INP(n2419), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5291), .IN2(U6375_n1), .QN(n2405) );
  INVX0 U6417_U2 ( .INP(n4198), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n8947), .IN2(U6417_n1), .QN(n2404) );
  INVX0 U6446_U2 ( .INP(g110), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n1782), .IN2(U6446_n1), .QN(n3524) );
  INVX0 U6465_U2 ( .INP(n3653), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5600), .IN2(U6465_n1), .QN(n4388) );
  INVX0 U6497_U2 ( .INP(n811), .ZN(U6497_n1) );
  NOR2X0 U6497_U1 ( .IN1(n3635), .IN2(U6497_n1), .QN(n3005) );
  INVX0 U6523_U2 ( .INP(n4946), .ZN(U6523_n1) );
  NOR2X0 U6523_U1 ( .IN1(n8947), .IN2(U6523_n1), .QN(n4945) );
  INVX0 U6542_U2 ( .INP(n811), .ZN(U6542_n1) );
  NOR2X0 U6542_U1 ( .IN1(n5300), .IN2(U6542_n1), .QN(n3525) );
  INVX0 U6552_U2 ( .INP(n3281), .ZN(U6552_n1) );
  NOR2X0 U6552_U1 ( .IN1(n5676), .IN2(U6552_n1), .QN(n3277) );
  INVX0 U6553_U2 ( .INP(n3276), .ZN(U6553_n1) );
  NOR2X0 U6553_U1 ( .IN1(n5680), .IN2(U6553_n1), .QN(n2989) );
  INVX0 U6554_U2 ( .INP(n3277), .ZN(U6554_n1) );
  NOR2X0 U6554_U1 ( .IN1(n5677), .IN2(U6554_n1), .QN(n2991) );
  INVX0 U6555_U2 ( .INP(n56), .ZN(U6555_n1) );
  NOR2X0 U6555_U1 ( .IN1(n5561), .IN2(U6555_n1), .QN(n3281) );
  INVX0 U6556_U2 ( .INP(n53), .ZN(U6556_n1) );
  NOR2X0 U6556_U1 ( .IN1(n5679), .IN2(U6556_n1), .QN(n3276) );
  INVX0 U6559_U2 ( .INP(n2991), .ZN(U6559_n1) );
  NOR2X0 U6559_U1 ( .IN1(n5678), .IN2(U6559_n1), .QN(n2710) );
  INVX0 U6560_U2 ( .INP(n2989), .ZN(U6560_n1) );
  NOR2X0 U6560_U1 ( .IN1(n5675), .IN2(U6560_n1), .QN(n2707) );
  INVX0 U6561_U2 ( .INP(n3174), .ZN(U6561_n1) );
  NOR2X0 U6561_U1 ( .IN1(n5327), .IN2(U6561_n1), .QN(n3116) );
  INVX0 U6570_U2 ( .INP(n3362), .ZN(U6570_n1) );
  NOR2X0 U6570_U1 ( .IN1(n5477), .IN2(U6570_n1), .QN(n2527) );
  INVX0 U6911_U2 ( .INP(n3115), .ZN(U6911_n1) );
  NOR2X0 U6911_U1 ( .IN1(n2726), .IN2(U6911_n1), .QN(n3111) );
  INVX0 U6912_U2 ( .INP(n3115), .ZN(U6912_n1) );
  NOR2X0 U6912_U1 ( .IN1(n2727), .IN2(U6912_n1), .QN(n3131) );
  INVX0 U6917_U2 ( .INP(n3933), .ZN(U6917_n1) );
  NOR2X0 U6917_U1 ( .IN1(n5350), .IN2(U6917_n1), .QN(n3799) );
  INVX0 U6926_U2 ( .INP(n3664), .ZN(U6926_n1) );
  NOR2X0 U6926_U1 ( .IN1(n5674), .IN2(U6926_n1), .QN(n3662) );
  INVX0 U6927_U2 ( .INP(n3673), .ZN(U6927_n1) );
  NOR2X0 U6927_U1 ( .IN1(n5673), .IN2(U6927_n1), .QN(n3671) );
  INVX0 U6929_U2 ( .INP(n3505), .ZN(U6929_n1) );
  NOR2X0 U6929_U1 ( .IN1(n3506), .IN2(U6929_n1), .QN(n2790) );
  INVX0 U6931_U2 ( .INP(n4490), .ZN(U6931_n1) );
  NOR2X0 U6931_U1 ( .IN1(n5554), .IN2(U6931_n1), .QN(n4178) );
  INVX0 U6932_U2 ( .INP(n4514), .ZN(U6932_n1) );
  NOR2X0 U6932_U1 ( .IN1(n5555), .IN2(U6932_n1), .QN(n4196) );
  INVX0 U6933_U2 ( .INP(n4178), .ZN(U6933_n1) );
  NOR2X0 U6933_U1 ( .IN1(n5558), .IN2(U6933_n1), .QN(n3736) );
  INVX0 U6934_U2 ( .INP(n4196), .ZN(U6934_n1) );
  NOR2X0 U6934_U1 ( .IN1(n5559), .IN2(U6934_n1), .QN(n3741) );
  INVX0 U6935_U2 ( .INP(n3736), .ZN(U6935_n1) );
  NOR2X0 U6935_U1 ( .IN1(n5553), .IN2(U6935_n1), .QN(n3664) );
  INVX0 U6936_U2 ( .INP(n3741), .ZN(U6936_n1) );
  NOR2X0 U6936_U1 ( .IN1(n5560), .IN2(U6936_n1), .QN(n3673) );
  INVX0 U6937_U2 ( .INP(n2601), .ZN(U6937_n1) );
  NOR2X0 U6937_U1 ( .IN1(n5303), .IN2(U6937_n1), .QN(n2598) );
  INVX0 U6938_U2 ( .INP(n1220), .ZN(U6938_n1) );
  NOR2X0 U6938_U1 ( .IN1(n5556), .IN2(U6938_n1), .QN(n4490) );
  INVX0 U6939_U2 ( .INP(n279), .ZN(U6939_n1) );
  NOR2X0 U6939_U1 ( .IN1(n5557), .IN2(U6939_n1), .QN(n4514) );
  INVX0 U6940_U2 ( .INP(n4814), .ZN(U6940_n1) );
  NOR2X0 U6940_U1 ( .IN1(n5422), .IN2(U6940_n1), .QN(n4519) );
  INVX0 U6941_U2 ( .INP(n2607), .ZN(U6941_n1) );
  NOR2X0 U6941_U1 ( .IN1(n5323), .IN2(U6941_n1), .QN(n2594) );
  INVX0 U6944_U2 ( .INP(n3084), .ZN(U6944_n1) );
  NOR2X0 U6944_U1 ( .IN1(n5348), .IN2(U6944_n1), .QN(n3033) );
  INVX0 U6950_U2 ( .INP(n2598), .ZN(U6950_n1) );
  NOR2X0 U6950_U1 ( .IN1(n5365), .IN2(U6950_n1), .QN(n2590) );
  INVX0 U6954_U2 ( .INP(n3122), .ZN(U6954_n1) );
  NOR2X0 U6954_U1 ( .IN1(n2727), .IN2(U6954_n1), .QN(n3125) );
  INVX0 U6955_U2 ( .INP(n686), .ZN(U6955_n1) );
  NOR2X0 U6955_U1 ( .IN1(n2726), .IN2(U6955_n1), .QN(n3105) );
  INVX0 U6956_U2 ( .INP(n3141), .ZN(U6956_n1) );
  NOR2X0 U6956_U1 ( .IN1(n3146), .IN2(U6956_n1), .QN(n3145) );
  INVX0 U6957_U2 ( .INP(n700), .ZN(U6957_n1) );
  NOR2X0 U6957_U1 ( .IN1(n3165), .IN2(U6957_n1), .QN(n3164) );
  INVX0 U7174_U2 ( .INP(n2423), .ZN(U7174_n1) );
  NOR2X0 U7174_U1 ( .IN1(n5288), .IN2(U7174_n1), .QN(n2422) );
  INVX0 U7248_U2 ( .INP(n4172), .ZN(U7248_n1) );
  NOR2X0 U7248_U1 ( .IN1(g1536), .IN2(U7248_n1), .QN(n4173) );
  INVX0 U7249_U2 ( .INP(n4190), .ZN(U7249_n1) );
  NOR2X0 U7249_U1 ( .IN1(g1193), .IN2(U7249_n1), .QN(n4191) );
  INVX0 U7402_U2 ( .INP(n4034), .ZN(U7402_n1) );
  NOR2X0 U7402_U1 ( .IN1(n528), .IN2(U7402_n1), .QN(n4037) );
  INVX0 U7405_U2 ( .INP(n4034), .ZN(U7405_n1) );
  NOR2X0 U7405_U1 ( .IN1(n527), .IN2(U7405_n1), .QN(n4039) );
  INVX0 U7413_U2 ( .INP(n3969), .ZN(U7413_n1) );
  NOR2X0 U7413_U1 ( .IN1(n826), .IN2(U7413_n1), .QN(n3972) );
  INVX0 U7416_U2 ( .INP(n3926), .ZN(U7416_n1) );
  NOR2X0 U7416_U1 ( .IN1(n205), .IN2(U7416_n1), .QN(n3929) );
  INVX0 U7427_U2 ( .INP(n3860), .ZN(U7427_n1) );
  NOR2X0 U7427_U1 ( .IN1(n712), .IN2(U7427_n1), .QN(n3863) );
  INVX0 U7438_U2 ( .INP(n4002), .ZN(U7438_n1) );
  NOR2X0 U7438_U1 ( .IN1(n429), .IN2(U7438_n1), .QN(n4003) );
  INVX0 U7449_U2 ( .INP(n4034), .ZN(U7449_n1) );
  NOR2X0 U7449_U1 ( .IN1(n530), .IN2(U7449_n1), .QN(n4032) );
  INVX0 U7455_U2 ( .INP(n4034), .ZN(U7455_n1) );
  NOR2X0 U7455_U1 ( .IN1(n526), .IN2(U7455_n1), .QN(n4035) );
  INVX0 U7464_U2 ( .INP(n3792), .ZN(U7464_n1) );
  NOR2X0 U7464_U1 ( .IN1(n1403), .IN2(U7464_n1), .QN(n3797) );
  INVX0 U7467_U2 ( .INP(n3792), .ZN(U7467_n1) );
  NOR2X0 U7467_U1 ( .IN1(n1409), .IN2(U7467_n1), .QN(n3790) );
  INVX0 U7482_U2 ( .INP(n3792), .ZN(U7482_n1) );
  NOR2X0 U7482_U1 ( .IN1(n1405), .IN2(U7482_n1), .QN(n3795) );
  INVX0 U7492_U2 ( .INP(n3893), .ZN(U7492_n1) );
  NOR2X0 U7492_U1 ( .IN1(n939), .IN2(U7492_n1), .QN(n3891) );
  INVX0 U7513_U2 ( .INP(n3826), .ZN(U7513_n1) );
  NOR2X0 U7513_U1 ( .IN1(n46), .IN2(U7513_n1), .QN(n3827) );
  INVX0 U7516_U2 ( .INP(n3893), .ZN(U7516_n1) );
  NOR2X0 U7516_U1 ( .IN1(n937), .IN2(U7516_n1), .QN(n3896) );
  INVX0 U7549_U2 ( .INP(n4002), .ZN(U7549_n1) );
  NOR2X0 U7549_U1 ( .IN1(n431), .IN2(U7549_n1), .QN(n4007) );
  INVX0 U7561_U2 ( .INP(n3926), .ZN(U7561_n1) );
  NOR2X0 U7561_U1 ( .IN1(n207), .IN2(U7561_n1), .QN(n3931) );
  INVX0 U7574_U2 ( .INP(n3792), .ZN(U7574_n1) );
  NOR2X0 U7574_U1 ( .IN1(n1401), .IN2(U7574_n1), .QN(n3793) );
  INVX0 U7577_U2 ( .INP(n3926), .ZN(U7577_n1) );
  NOR2X0 U7577_U1 ( .IN1(n214), .IN2(U7577_n1), .QN(n3924) );
  INVX0 U7585_U2 ( .INP(n3826), .ZN(U7585_n1) );
  NOR2X0 U7585_U1 ( .IN1(n44), .IN2(U7585_n1), .QN(n3831) );
  INVX0 U7595_U2 ( .INP(n3826), .ZN(U7595_n1) );
  NOR2X0 U7595_U1 ( .IN1(n42), .IN2(U7595_n1), .QN(n3829) );
  INVX0 U7614_U2 ( .INP(n3926), .ZN(U7614_n1) );
  NOR2X0 U7614_U1 ( .IN1(n209), .IN2(U7614_n1), .QN(n3927) );
  INVX0 U7621_U2 ( .INP(n3969), .ZN(U7621_n1) );
  NOR2X0 U7621_U1 ( .IN1(n828), .IN2(U7621_n1), .QN(n3974) );
  INVX0 U7629_U2 ( .INP(n3893), .ZN(U7629_n1) );
  NOR2X0 U7629_U1 ( .IN1(n936), .IN2(U7629_n1), .QN(n3898) );
  INVX0 U7636_U2 ( .INP(n3969), .ZN(U7636_n1) );
  NOR2X0 U7636_U1 ( .IN1(n830), .IN2(U7636_n1), .QN(n3970) );
  INVX0 U7639_U2 ( .INP(n4002), .ZN(U7639_n1) );
  NOR2X0 U7639_U1 ( .IN1(n438), .IN2(U7639_n1), .QN(n4000) );
  INVX0 U7649_U2 ( .INP(n3860), .ZN(U7649_n1) );
  NOR2X0 U7649_U1 ( .IN1(n714), .IN2(U7649_n1), .QN(n3865) );
  INVX0 U7652_U2 ( .INP(n3860), .ZN(U7652_n1) );
  NOR2X0 U7652_U1 ( .IN1(n716), .IN2(U7652_n1), .QN(n3861) );
  INVX0 U7668_U2 ( .INP(n3826), .ZN(U7668_n1) );
  NOR2X0 U7668_U1 ( .IN1(n51), .IN2(U7668_n1), .QN(n3824) );
  INVX0 U7673_U2 ( .INP(n3893), .ZN(U7673_n1) );
  NOR2X0 U7673_U1 ( .IN1(n935), .IN2(U7673_n1), .QN(n3894) );
  INVX0 U7690_U2 ( .INP(n3969), .ZN(U7690_n1) );
  NOR2X0 U7690_U1 ( .IN1(n835), .IN2(U7690_n1), .QN(n3967) );
  INVX0 U7707_U2 ( .INP(n3860), .ZN(U7707_n1) );
  NOR2X0 U7707_U1 ( .IN1(n720), .IN2(U7707_n1), .QN(n3858) );
  INVX0 U7712_U2 ( .INP(n4002), .ZN(U7712_n1) );
  NOR2X0 U7712_U1 ( .IN1(n433), .IN2(U7712_n1), .QN(n4005) );
  INVX0 U7792_U2 ( .INP(g952), .ZN(U7792_n1) );
  NOR2X0 U7792_U1 ( .IN1(n8946), .IN2(U7792_n1), .QN(n2505) );
  INVX0 U7794_U2 ( .INP(g1296), .ZN(U7794_n1) );
  NOR2X0 U7794_U1 ( .IN1(n8944), .IN2(U7794_n1), .QN(n2499) );
  INVX0 U7895_U2 ( .INP(n2668), .ZN(U7895_n1) );
  NOR2X0 U7895_U1 ( .IN1(g113), .IN2(U7895_n1), .QN(n2760) );
  INVX0 U7897_U2 ( .INP(g6), .ZN(U7897_n1) );
  NOR2X0 U7897_U1 ( .IN1(g31), .IN2(U7897_n1), .QN(n3395) );
  INVX0 U7977_U2 ( .INP(g661), .ZN(U7977_n1) );
  NOR2X0 U7977_U1 ( .IN1(n8947), .IN2(U7977_n1), .QN(n4956) );
  INVX0 U8034_U2 ( .INP(n1242), .ZN(U8034_n1) );
  NOR2X0 U8034_U1 ( .IN1(n5612), .IN2(U8034_n1), .QN(n5026) );
  INVX0 U8036_U2 ( .INP(n3729), .ZN(U8036_n1) );
  NOR2X0 U8036_U1 ( .IN1(n5340), .IN2(U8036_n1), .QN(n3941) );
  INVX0 U8050_U2 ( .INP(n198), .ZN(U8050_n1) );
  NOR2X0 U8050_U1 ( .IN1(g1367), .IN2(U8050_n1), .QN(n3733) );
  INVX0 U8055_U2 ( .INP(g1345), .ZN(U8055_n1) );
  NOR2X0 U8055_U1 ( .IN1(n8946), .IN2(U8055_n1), .QN(n4798) );
  INVX0 U8060_U2 ( .INP(g1002), .ZN(U8060_n1) );
  NOR2X0 U8060_U1 ( .IN1(n8945), .IN2(U8060_n1), .QN(n4805) );
  INVX0 U8070_U2 ( .INP(n199), .ZN(U8070_n1) );
  NOR2X0 U8070_U1 ( .IN1(g1361), .IN2(U8070_n1), .QN(n4175) );
  INVX0 U8074_U2 ( .INP(n543), .ZN(U8074_n1) );
  NOR2X0 U8074_U1 ( .IN1(g1018), .IN2(U8074_n1), .QN(n4193) );
  INVX0 U8088_U2 ( .INP(n542), .ZN(U8088_n1) );
  NOR2X0 U8088_U1 ( .IN1(g1024), .IN2(U8088_n1), .QN(n3738) );
  INVX0 U8112_U2 ( .INP(n4525), .ZN(U8112_n1) );
  NOR2X0 U8112_U1 ( .IN1(n4523), .IN2(U8112_n1), .QN(n4524) );
  INVX0 U8113_U2 ( .INP(n4526), .ZN(U8113_n1) );
  NOR2X0 U8113_U1 ( .IN1(n5751), .IN2(U8113_n1), .QN(n4523) );
  INVX0 U8147_U2 ( .INP(g4659), .ZN(U8147_n1) );
  NOR2X0 U8147_U1 ( .IN1(n2573), .IN2(U8147_n1), .QN(n2577) );
  INVX0 U8165_U2 ( .INP(g4849), .ZN(U8165_n1) );
  NOR2X0 U8165_U1 ( .IN1(n2563), .IN2(U8165_n1), .QN(n2567) );
  INVX0 U8185_U2 ( .INP(n853), .ZN(U8185_n1) );
  NOR2X0 U8185_U1 ( .IN1(g1046), .IN2(U8185_n1), .QN(n4938) );
  INVX0 U8192_U2 ( .INP(n192), .ZN(U8192_n1) );
  NOR2X0 U8192_U1 ( .IN1(g1389), .IN2(U8192_n1), .QN(n4913) );
  INVX0 U8210_U2 ( .INP(n4722), .ZN(U8210_n1) );
  NOR2X0 U8210_U1 ( .IN1(n1242), .IN2(U8210_n1), .QN(n4714) );
  INVX0 U8223_U2 ( .INP(n4518), .ZN(U8223_n1) );
  NOR2X0 U8223_U1 ( .IN1(n4516), .IN2(U8223_n1), .QN(n4517) );
  INVX0 U8224_U2 ( .INP(n4519), .ZN(U8224_n1) );
  NOR2X0 U8224_U1 ( .IN1(n5728), .IN2(U8224_n1), .QN(n4516) );
  INVX0 U8281_U2 ( .INP(n4819), .ZN(U8281_n1) );
  NOR2X0 U8281_U1 ( .IN1(n8947), .IN2(U8281_n1), .QN(n5111) );
  INVX0 U8307_U2 ( .INP(g29216), .ZN(U8307_n1) );
  NOR2X0 U8307_U1 ( .IN1(n8947), .IN2(U8307_n1), .QN(g26900) );
  INVX0 U8974_U2 ( .INP(n3362), .ZN(U8974_n1) );
  NOR2X0 U8974_U1 ( .IN1(test_so25), .IN2(U8974_n1), .QN(n2552) );
  INVX0 U8975_U2 ( .INP(n3174), .ZN(U8975_n1) );
  NOR2X0 U8975_U1 ( .IN1(g528), .IN2(U8975_n1), .QN(n3195) );
  INVX0 U9065_U2 ( .INP(g4145), .ZN(U9065_n1) );
  NOR2X0 U9065_U1 ( .IN1(n8945), .IN2(U9065_n1), .QN(n4721) );
  INVX0 U9070_U2 ( .INP(g2841), .ZN(U9070_n1) );
  NOR2X0 U9070_U1 ( .IN1(n8945), .IN2(U9070_n1), .QN(n3730) );
  INVX0 U9075_U2 ( .INP(g19), .ZN(U9075_n1) );
  NOR2X0 U9075_U1 ( .IN1(g9), .IN2(U9075_n1), .QN(n3362) );
  INVX0 U9076_U2 ( .INP(g113), .ZN(U9076_n1) );
  NOR2X0 U9076_U1 ( .IN1(n8944), .IN2(U9076_n1), .QN(g25694) );
  INVX0 U9080_U2 ( .INP(n4305), .ZN(U9080_n1) );
  NOR2X0 U9080_U1 ( .IN1(n8946), .IN2(U9080_n1), .QN(g29277) );
  INVX0 U9084_U2 ( .INP(g4423), .ZN(U9084_n1) );
  NOR2X0 U9084_U1 ( .IN1(n8945), .IN2(U9084_n1), .QN(g26953) );
  INVX0 U9085_U2 ( .INP(g64), .ZN(U9085_n1) );
  NOR2X0 U9085_U1 ( .IN1(n8945), .IN2(U9085_n1), .QN(g24212) );
  INVX0 U9086_U2 ( .INP(n4283), .ZN(U9086_n1) );
  NOR2X0 U9086_U1 ( .IN1(n8946), .IN2(U9086_n1), .QN(g29279) );
  INVX0 U9090_U2 ( .INP(g125), .ZN(U9090_n1) );
  NOR2X0 U9090_U1 ( .IN1(n8944), .IN2(U9090_n1), .QN(g25688) );
  INVX0 U9098_U2 ( .INP(g4681), .ZN(U9098_n1) );
  NOR2X0 U9098_U1 ( .IN1(n2774), .IN2(U9098_n1), .QN(g34028) );
  INVX0 U9099_U2 ( .INP(n2595), .ZN(U9099_n1) );
  NOR2X0 U9099_U1 ( .IN1(n2608), .IN2(U9099_n1), .QN(g34449) );
  INVX0 U9101_U2 ( .INP(g6745), .ZN(U9101_n1) );
  NOR2X0 U9101_U1 ( .IN1(n8944), .IN2(U9101_n1), .QN(g26880) );
  INVX0 U9107_U2 ( .INP(n4448), .ZN(U9107_n1) );
  NOR2X0 U9107_U1 ( .IN1(n8579), .IN2(U9107_n1), .QN(n4447) );
  INVX0 U9111_U2 ( .INP(n4403), .ZN(U9111_n1) );
  NOR2X0 U9111_U1 ( .IN1(n8576), .IN2(U9111_n1), .QN(n4402) );
  INVX0 U9116_U2 ( .INP(n1411), .ZN(U9116_n1) );
  NOR2X0 U9116_U1 ( .IN1(n8583), .IN2(U9116_n1), .QN(n4425) );
  INVX0 U9120_U2 ( .INP(n4437), .ZN(U9120_n1) );
  NOR2X0 U9120_U1 ( .IN1(n8573), .IN2(U9120_n1), .QN(n4436) );
  INVX0 U9124_U2 ( .INP(n4392), .ZN(U9124_n1) );
  NOR2X0 U9124_U1 ( .IN1(n8580), .IN2(U9124_n1), .QN(n4391) );
  INVX0 U9128_U2 ( .INP(n4380), .ZN(U9128_n1) );
  NOR2X0 U9128_U1 ( .IN1(n8574), .IN2(U9128_n1), .QN(n4379) );
  INVX0 U9132_U2 ( .INP(n4415), .ZN(U9132_n1) );
  NOR2X0 U9132_U1 ( .IN1(n8581), .IN2(U9132_n1), .QN(n4414) );
  INVX0 U9136_U2 ( .INP(n4459), .ZN(U9136_n1) );
  NOR2X0 U9136_U1 ( .IN1(n8582), .IN2(U9136_n1), .QN(n4458) );
  INVX0 U9315_U2 ( .INP(n5016), .ZN(U9315_n1) );
  NOR2X0 U9315_U1 ( .IN1(n5753), .IN2(U9315_n1), .QN(n5014) );
  INVX0 U9453_U2 ( .INP(n3065), .ZN(U9453_n1) );
  NOR2X0 U9453_U1 ( .IN1(n8577), .IN2(U9453_n1), .QN(n3064) );
  INVX0 U9825_U2 ( .INP(g112), .ZN(U9825_n1) );
  NOR2X0 U9825_U1 ( .IN1(n1782), .IN2(U9825_n1), .QN(n3115) );
  INVX0 U9886_U2 ( .INP(g370), .ZN(U9886_n1) );
  NOR2X0 U9886_U1 ( .IN1(n1161), .IN2(U9886_n1), .QN(n4948) );
  INVX0 U9927_U2 ( .INP(n3933), .ZN(U9927_n1) );
  NOR2X0 U9927_U1 ( .IN1(g4098), .IN2(U9927_n1), .QN(n3833) );
  INVX0 U9953_U2 ( .INP(g671), .ZN(U9953_n1) );
  NOR2X0 U9953_U1 ( .IN1(n8569), .IN2(U9953_n1), .QN(n4526) );
  INVX0 U9957_U2 ( .INP(g4843), .ZN(U9957_n1) );
  NOR2X0 U9957_U1 ( .IN1(n5283), .IN2(U9957_n1), .QN(n2563) );
  INVX0 U9958_U2 ( .INP(test_so19), .ZN(U9958_n1) );
  NOR2X0 U9958_U1 ( .IN1(n5656), .IN2(U9958_n1), .QN(n2573) );
  INVX0 U9968_U2 ( .INP(n3084), .ZN(U9968_n1) );
  NOR2X0 U9968_U1 ( .IN1(g4358), .IN2(U9968_n1), .QN(n3023) );
  INVX0 U9972_U2 ( .INP(g681), .ZN(U9972_n1) );
  NOR2X0 U9972_U1 ( .IN1(n4535), .IN2(U9972_n1), .QN(n5112) );
  INVX0 U9992_U2 ( .INP(n3675), .ZN(U9992_n1) );
  NOR2X0 U9992_U1 ( .IN1(n3676), .IN2(U9992_n1), .QN(n2644) );
  INVX0 U10314_U2 ( .INP(g667), .ZN(U10314_n1) );
  NOR2X0 U10314_U1 ( .IN1(g686), .IN2(U10314_n1), .QN(n4962) );
  INVX0 U10318_U2 ( .INP(g5092), .ZN(U10318_n1) );
  NOR2X0 U10318_U1 ( .IN1(n5681), .IN2(U10318_n1), .QN(n5016) );
endmodule

