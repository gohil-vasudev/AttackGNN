module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;

  XOR2_X1 U537 ( .A(n521), .B(n522), .Z(Result_9_) );
  XOR2_X1 U538 ( .A(n523), .B(n524), .Z(n522) );
  XNOR2_X1 U539 ( .A(n525), .B(n526), .ZN(Result_8_) );
  XNOR2_X1 U540 ( .A(n527), .B(n528), .ZN(n526) );
  XNOR2_X1 U541 ( .A(n529), .B(n530), .ZN(Result_7_) );
  NOR2_X1 U542 ( .A1(n531), .A2(n532), .ZN(Result_6_) );
  NOR2_X1 U543 ( .A1(n533), .A2(n534), .ZN(n532) );
  XOR2_X1 U544 ( .A(n535), .B(n536), .Z(Result_5_) );
  XNOR2_X1 U545 ( .A(n531), .B(n537), .ZN(n536) );
  INV_X1 U546 ( .A(n538), .ZN(n531) );
  XOR2_X1 U547 ( .A(n539), .B(n540), .Z(Result_4_) );
  XOR2_X1 U548 ( .A(n541), .B(n542), .Z(Result_3_) );
  NAND2_X1 U549 ( .A1(n543), .A2(n544), .ZN(n541) );
  NAND2_X1 U550 ( .A1(n545), .A2(n546), .ZN(n544) );
  INV_X1 U551 ( .A(n547), .ZN(n543) );
  XOR2_X1 U552 ( .A(n548), .B(n549), .Z(Result_2_) );
  XNOR2_X1 U553 ( .A(n550), .B(n551), .ZN(Result_1_) );
  NOR2_X1 U554 ( .A1(n552), .A2(n553), .ZN(n551) );
  XOR2_X1 U555 ( .A(n554), .B(n555), .Z(Result_14_) );
  NOR2_X1 U556 ( .A1(n556), .A2(n557), .ZN(n555) );
  XOR2_X1 U557 ( .A(n558), .B(n559), .Z(Result_13_) );
  XOR2_X1 U558 ( .A(n560), .B(n561), .Z(n559) );
  XNOR2_X1 U559 ( .A(n562), .B(n563), .ZN(Result_12_) );
  NAND2_X1 U560 ( .A1(n564), .A2(n565), .ZN(n562) );
  XOR2_X1 U561 ( .A(n566), .B(n567), .Z(Result_11_) );
  XOR2_X1 U562 ( .A(n568), .B(n569), .Z(n567) );
  NOR2_X1 U563 ( .A1(n570), .A2(n557), .ZN(n569) );
  XOR2_X1 U564 ( .A(n571), .B(n572), .Z(Result_10_) );
  XOR2_X1 U565 ( .A(n573), .B(n574), .Z(n571) );
  NOR2_X1 U566 ( .A1(n575), .A2(n557), .ZN(n574) );
  NAND2_X1 U567 ( .A1(n576), .A2(n577), .ZN(Result_0_) );
  NAND2_X1 U568 ( .A1(n578), .A2(n579), .ZN(n577) );
  NOR2_X1 U569 ( .A1(n552), .A2(n580), .ZN(n576) );
  NOR2_X1 U570 ( .A1(n553), .A2(n550), .ZN(n580) );
  NAND2_X1 U571 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U572 ( .A1(n581), .A2(n582), .ZN(n548) );
  NAND2_X1 U573 ( .A1(n583), .A2(n584), .ZN(n582) );
  NOR2_X1 U574 ( .A1(n547), .A2(n585), .ZN(n581) );
  NOR2_X1 U575 ( .A1(n545), .A2(n542), .ZN(n585) );
  NAND2_X1 U576 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U577 ( .A1(n586), .A2(n587), .ZN(n539) );
  NAND2_X1 U578 ( .A1(n537), .A2(n588), .ZN(n586) );
  NAND2_X1 U579 ( .A1(n535), .A2(n538), .ZN(n588) );
  NAND2_X1 U580 ( .A1(n533), .A2(n534), .ZN(n538) );
  XOR2_X1 U581 ( .A(n589), .B(n590), .Z(n534) );
  NOR2_X1 U582 ( .A1(n591), .A2(n530), .ZN(n533) );
  XNOR2_X1 U583 ( .A(n592), .B(n593), .ZN(n530) );
  XOR2_X1 U584 ( .A(n594), .B(n595), .Z(n592) );
  INV_X1 U585 ( .A(n529), .ZN(n591) );
  NAND2_X1 U586 ( .A1(n596), .A2(n597), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n528), .A2(n598), .ZN(n597) );
  INV_X1 U588 ( .A(n599), .ZN(n598) );
  NOR2_X1 U589 ( .A1(n527), .A2(n525), .ZN(n599) );
  NOR2_X1 U590 ( .A1(n557), .A2(n600), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n525), .A2(n527), .ZN(n596) );
  NAND2_X1 U592 ( .A1(n601), .A2(n602), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n524), .A2(n603), .ZN(n602) );
  INV_X1 U594 ( .A(n604), .ZN(n603) );
  NOR2_X1 U595 ( .A1(n523), .A2(n521), .ZN(n604) );
  NOR2_X1 U596 ( .A1(n605), .A2(n557), .ZN(n524) );
  NAND2_X1 U597 ( .A1(n521), .A2(n523), .ZN(n601) );
  NAND2_X1 U598 ( .A1(n606), .A2(n607), .ZN(n523) );
  NAND2_X1 U599 ( .A1(n608), .A2(n609), .ZN(n607) );
  NOR2_X1 U600 ( .A1(n610), .A2(n575), .ZN(n608) );
  NOR2_X1 U601 ( .A1(n572), .A2(n573), .ZN(n610) );
  NAND2_X1 U602 ( .A1(n572), .A2(n573), .ZN(n606) );
  NAND2_X1 U603 ( .A1(n611), .A2(n612), .ZN(n573) );
  NAND2_X1 U604 ( .A1(n613), .A2(n609), .ZN(n612) );
  NOR2_X1 U605 ( .A1(n614), .A2(n570), .ZN(n613) );
  NOR2_X1 U606 ( .A1(n566), .A2(n568), .ZN(n614) );
  NAND2_X1 U607 ( .A1(n566), .A2(n568), .ZN(n611) );
  NAND2_X1 U608 ( .A1(n564), .A2(n615), .ZN(n568) );
  NAND2_X1 U609 ( .A1(n563), .A2(n565), .ZN(n615) );
  NAND2_X1 U610 ( .A1(n616), .A2(n617), .ZN(n565) );
  NAND2_X1 U611 ( .A1(n609), .A2(n618), .ZN(n617) );
  XNOR2_X1 U612 ( .A(n619), .B(n620), .ZN(n563) );
  XNOR2_X1 U613 ( .A(n621), .B(n622), .ZN(n619) );
  INV_X1 U614 ( .A(n623), .ZN(n564) );
  NOR2_X1 U615 ( .A1(n624), .A2(n616), .ZN(n623) );
  NOR2_X1 U616 ( .A1(n625), .A2(n626), .ZN(n616) );
  INV_X1 U617 ( .A(n627), .ZN(n626) );
  NAND2_X1 U618 ( .A1(n561), .A2(n628), .ZN(n627) );
  NAND2_X1 U619 ( .A1(n558), .A2(n560), .ZN(n628) );
  NOR2_X1 U620 ( .A1(n557), .A2(n629), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n560), .A2(n558), .ZN(n625) );
  XNOR2_X1 U622 ( .A(n630), .B(n631), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n632), .A2(n633), .ZN(n631) );
  NAND2_X1 U624 ( .A1(Result_15_), .A2(n630), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n634), .A2(n556), .ZN(n630) );
  NOR2_X1 U626 ( .A1(n557), .A2(n632), .ZN(Result_15_) );
  INV_X1 U627 ( .A(n609), .ZN(n557) );
  NOR2_X1 U628 ( .A1(n635), .A2(n636), .ZN(n609) );
  NOR2_X1 U629 ( .A1(c_7_), .A2(d_7_), .ZN(n636) );
  XNOR2_X1 U630 ( .A(n637), .B(n638), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n639), .B(n640), .ZN(n637) );
  XNOR2_X1 U632 ( .A(n641), .B(n642), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n643), .B(n644), .ZN(n641) );
  XNOR2_X1 U634 ( .A(n645), .B(n646), .ZN(n521) );
  XNOR2_X1 U635 ( .A(n647), .B(n648), .ZN(n645) );
  XNOR2_X1 U636 ( .A(n649), .B(n650), .ZN(n525) );
  XNOR2_X1 U637 ( .A(n651), .B(n652), .ZN(n649) );
  NAND2_X1 U638 ( .A1(n590), .A2(n589), .ZN(n535) );
  NAND2_X1 U639 ( .A1(n653), .A2(n654), .ZN(n589) );
  NAND2_X1 U640 ( .A1(n595), .A2(n655), .ZN(n654) );
  INV_X1 U641 ( .A(n656), .ZN(n655) );
  NOR2_X1 U642 ( .A1(n594), .A2(n593), .ZN(n656) );
  NOR2_X1 U643 ( .A1(n600), .A2(n634), .ZN(n595) );
  NAND2_X1 U644 ( .A1(n593), .A2(n594), .ZN(n653) );
  NAND2_X1 U645 ( .A1(n657), .A2(n658), .ZN(n594) );
  NAND2_X1 U646 ( .A1(n652), .A2(n659), .ZN(n658) );
  NAND2_X1 U647 ( .A1(n650), .A2(n651), .ZN(n659) );
  NOR2_X1 U648 ( .A1(n605), .A2(n634), .ZN(n652) );
  INV_X1 U649 ( .A(n660), .ZN(n657) );
  NOR2_X1 U650 ( .A1(n650), .A2(n651), .ZN(n660) );
  NOR2_X1 U651 ( .A1(n661), .A2(n662), .ZN(n651) );
  INV_X1 U652 ( .A(n663), .ZN(n662) );
  NAND2_X1 U653 ( .A1(n648), .A2(n664), .ZN(n663) );
  NAND2_X1 U654 ( .A1(n646), .A2(n647), .ZN(n664) );
  NOR2_X1 U655 ( .A1(n575), .A2(n634), .ZN(n648) );
  NOR2_X1 U656 ( .A1(n646), .A2(n647), .ZN(n661) );
  NOR2_X1 U657 ( .A1(n665), .A2(n666), .ZN(n647) );
  INV_X1 U658 ( .A(n667), .ZN(n666) );
  NAND2_X1 U659 ( .A1(n644), .A2(n668), .ZN(n667) );
  NAND2_X1 U660 ( .A1(n643), .A2(n642), .ZN(n668) );
  NOR2_X1 U661 ( .A1(n570), .A2(n634), .ZN(n644) );
  NOR2_X1 U662 ( .A1(n642), .A2(n643), .ZN(n665) );
  NOR2_X1 U663 ( .A1(n669), .A2(n670), .ZN(n643) );
  INV_X1 U664 ( .A(n671), .ZN(n670) );
  NAND2_X1 U665 ( .A1(n640), .A2(n672), .ZN(n671) );
  NAND2_X1 U666 ( .A1(n639), .A2(n638), .ZN(n672) );
  NOR2_X1 U667 ( .A1(n624), .A2(n634), .ZN(n640) );
  NOR2_X1 U668 ( .A1(n638), .A2(n639), .ZN(n669) );
  NOR2_X1 U669 ( .A1(n673), .A2(n674), .ZN(n639) );
  INV_X1 U670 ( .A(n675), .ZN(n674) );
  NAND2_X1 U671 ( .A1(n620), .A2(n676), .ZN(n675) );
  NAND2_X1 U672 ( .A1(n621), .A2(n622), .ZN(n676) );
  NOR2_X1 U673 ( .A1(n629), .A2(n634), .ZN(n620) );
  NOR2_X1 U674 ( .A1(n622), .A2(n621), .ZN(n673) );
  NAND2_X1 U675 ( .A1(n677), .A2(n678), .ZN(n621) );
  INV_X1 U676 ( .A(n679), .ZN(n678) );
  NOR2_X1 U677 ( .A1(n680), .A2(n681), .ZN(n679) );
  NAND2_X1 U678 ( .A1(n554), .A2(n681), .ZN(n622) );
  NOR2_X1 U679 ( .A1(n632), .A2(n634), .ZN(n554) );
  XNOR2_X1 U680 ( .A(n635), .B(n682), .ZN(n634) );
  XOR2_X1 U681 ( .A(d_6_), .B(c_6_), .Z(n682) );
  XNOR2_X1 U682 ( .A(n683), .B(n684), .ZN(n638) );
  XOR2_X1 U683 ( .A(n677), .B(n685), .Z(n684) );
  XOR2_X1 U684 ( .A(n686), .B(n687), .Z(n642) );
  XNOR2_X1 U685 ( .A(n688), .B(n689), .ZN(n686) );
  XNOR2_X1 U686 ( .A(n690), .B(n691), .ZN(n646) );
  XOR2_X1 U687 ( .A(n692), .B(n693), .Z(n691) );
  XOR2_X1 U688 ( .A(n694), .B(n695), .Z(n650) );
  XNOR2_X1 U689 ( .A(n696), .B(n697), .ZN(n694) );
  XNOR2_X1 U690 ( .A(n698), .B(n699), .ZN(n593) );
  XNOR2_X1 U691 ( .A(n700), .B(n701), .ZN(n698) );
  XNOR2_X1 U692 ( .A(n702), .B(n703), .ZN(n590) );
  XNOR2_X1 U693 ( .A(n704), .B(n705), .ZN(n702) );
  NOR2_X1 U694 ( .A1(n706), .A2(n707), .ZN(n537) );
  INV_X1 U695 ( .A(n587), .ZN(n707) );
  NAND2_X1 U696 ( .A1(n708), .A2(n709), .ZN(n587) );
  NOR2_X1 U697 ( .A1(n709), .A2(n708), .ZN(n706) );
  XNOR2_X1 U698 ( .A(n710), .B(n711), .ZN(n708) );
  XNOR2_X1 U699 ( .A(n712), .B(n713), .ZN(n711) );
  NAND2_X1 U700 ( .A1(n714), .A2(n715), .ZN(n709) );
  NAND2_X1 U701 ( .A1(n705), .A2(n716), .ZN(n715) );
  NAND2_X1 U702 ( .A1(n703), .A2(n704), .ZN(n716) );
  NOR2_X1 U703 ( .A1(n633), .A2(n600), .ZN(n705) );
  INV_X1 U704 ( .A(n717), .ZN(n714) );
  NOR2_X1 U705 ( .A1(n703), .A2(n704), .ZN(n717) );
  NOR2_X1 U706 ( .A1(n718), .A2(n719), .ZN(n704) );
  INV_X1 U707 ( .A(n720), .ZN(n719) );
  NAND2_X1 U708 ( .A1(n701), .A2(n721), .ZN(n720) );
  NAND2_X1 U709 ( .A1(n699), .A2(n700), .ZN(n721) );
  NOR2_X1 U710 ( .A1(n605), .A2(n633), .ZN(n701) );
  NOR2_X1 U711 ( .A1(n699), .A2(n700), .ZN(n718) );
  NOR2_X1 U712 ( .A1(n722), .A2(n723), .ZN(n700) );
  INV_X1 U713 ( .A(n724), .ZN(n723) );
  NAND2_X1 U714 ( .A1(n697), .A2(n725), .ZN(n724) );
  NAND2_X1 U715 ( .A1(n696), .A2(n695), .ZN(n725) );
  NOR2_X1 U716 ( .A1(n575), .A2(n633), .ZN(n697) );
  NOR2_X1 U717 ( .A1(n695), .A2(n696), .ZN(n722) );
  NOR2_X1 U718 ( .A1(n726), .A2(n727), .ZN(n696) );
  INV_X1 U719 ( .A(n728), .ZN(n727) );
  NAND2_X1 U720 ( .A1(n693), .A2(n729), .ZN(n728) );
  NAND2_X1 U721 ( .A1(n692), .A2(n690), .ZN(n729) );
  NOR2_X1 U722 ( .A1(n570), .A2(n633), .ZN(n693) );
  NOR2_X1 U723 ( .A1(n690), .A2(n692), .ZN(n726) );
  NOR2_X1 U724 ( .A1(n730), .A2(n731), .ZN(n692) );
  INV_X1 U725 ( .A(n732), .ZN(n731) );
  NAND2_X1 U726 ( .A1(n689), .A2(n733), .ZN(n732) );
  NAND2_X1 U727 ( .A1(n688), .A2(n687), .ZN(n733) );
  NOR2_X1 U728 ( .A1(n633), .A2(n624), .ZN(n689) );
  NOR2_X1 U729 ( .A1(n687), .A2(n688), .ZN(n730) );
  NOR2_X1 U730 ( .A1(n734), .A2(n735), .ZN(n688) );
  INV_X1 U731 ( .A(n736), .ZN(n735) );
  NAND2_X1 U732 ( .A1(n683), .A2(n737), .ZN(n736) );
  NAND2_X1 U733 ( .A1(n685), .A2(n677), .ZN(n737) );
  NOR2_X1 U734 ( .A1(n633), .A2(n629), .ZN(n683) );
  NOR2_X1 U735 ( .A1(n677), .A2(n685), .ZN(n734) );
  NAND2_X1 U736 ( .A1(n738), .A2(n739), .ZN(n685) );
  NAND2_X1 U737 ( .A1(n740), .A2(n741), .ZN(n739) );
  NAND2_X1 U738 ( .A1(n742), .A2(n743), .ZN(n741) );
  INV_X1 U739 ( .A(n744), .ZN(n740) );
  NOR2_X1 U740 ( .A1(n745), .A2(n556), .ZN(n744) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n633), .A2(n556), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n746), .B(n747), .ZN(n633) );
  XOR2_X1 U744 ( .A(d_5_), .B(c_5_), .Z(n747) );
  XNOR2_X1 U745 ( .A(n748), .B(n749), .ZN(n687) );
  XOR2_X1 U746 ( .A(n738), .B(n750), .Z(n749) );
  XOR2_X1 U747 ( .A(n751), .B(n752), .Z(n690) );
  XNOR2_X1 U748 ( .A(n753), .B(n754), .ZN(n751) );
  XOR2_X1 U749 ( .A(n755), .B(n756), .Z(n695) );
  XNOR2_X1 U750 ( .A(n757), .B(n758), .ZN(n756) );
  XOR2_X1 U751 ( .A(n759), .B(n760), .Z(n699) );
  XNOR2_X1 U752 ( .A(n761), .B(n762), .ZN(n760) );
  XOR2_X1 U753 ( .A(n763), .B(n764), .Z(n703) );
  XNOR2_X1 U754 ( .A(n765), .B(n766), .ZN(n764) );
  XOR2_X1 U755 ( .A(n767), .B(n768), .Z(n540) );
  NOR2_X1 U756 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U757 ( .A(n583), .B(n584), .ZN(n545) );
  NAND2_X1 U758 ( .A1(n769), .A2(n770), .ZN(n584) );
  NAND2_X1 U759 ( .A1(n771), .A2(n772), .ZN(n770) );
  NAND2_X1 U760 ( .A1(n773), .A2(n774), .ZN(n772) );
  INV_X1 U761 ( .A(n775), .ZN(n769) );
  NOR2_X1 U762 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U763 ( .A(n776), .B(n777), .Z(n583) );
  XOR2_X1 U764 ( .A(n778), .B(n779), .Z(n776) );
  NOR2_X1 U765 ( .A1(n600), .A2(n780), .ZN(n779) );
  NAND2_X1 U766 ( .A1(n768), .A2(n767), .ZN(n546) );
  NAND2_X1 U767 ( .A1(n781), .A2(n782), .ZN(n767) );
  NAND2_X1 U768 ( .A1(n713), .A2(n783), .ZN(n782) );
  INV_X1 U769 ( .A(n784), .ZN(n783) );
  NOR2_X1 U770 ( .A1(n712), .A2(n710), .ZN(n784) );
  NOR2_X1 U771 ( .A1(n745), .A2(n600), .ZN(n713) );
  NAND2_X1 U772 ( .A1(n710), .A2(n712), .ZN(n781) );
  NAND2_X1 U773 ( .A1(n785), .A2(n786), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n766), .A2(n787), .ZN(n786) );
  INV_X1 U775 ( .A(n788), .ZN(n787) );
  NOR2_X1 U776 ( .A1(n765), .A2(n763), .ZN(n788) );
  NOR2_X1 U777 ( .A1(n605), .A2(n745), .ZN(n766) );
  NAND2_X1 U778 ( .A1(n763), .A2(n765), .ZN(n785) );
  NAND2_X1 U779 ( .A1(n789), .A2(n790), .ZN(n765) );
  NAND2_X1 U780 ( .A1(n762), .A2(n791), .ZN(n790) );
  INV_X1 U781 ( .A(n792), .ZN(n791) );
  NOR2_X1 U782 ( .A1(n761), .A2(n759), .ZN(n792) );
  NOR2_X1 U783 ( .A1(n575), .A2(n745), .ZN(n762) );
  NAND2_X1 U784 ( .A1(n759), .A2(n761), .ZN(n789) );
  NAND2_X1 U785 ( .A1(n793), .A2(n794), .ZN(n761) );
  NAND2_X1 U786 ( .A1(n758), .A2(n795), .ZN(n794) );
  INV_X1 U787 ( .A(n796), .ZN(n795) );
  NOR2_X1 U788 ( .A1(n755), .A2(n757), .ZN(n796) );
  NOR2_X1 U789 ( .A1(n570), .A2(n745), .ZN(n758) );
  NAND2_X1 U790 ( .A1(n755), .A2(n757), .ZN(n793) );
  NAND2_X1 U791 ( .A1(n797), .A2(n798), .ZN(n757) );
  NAND2_X1 U792 ( .A1(n754), .A2(n799), .ZN(n798) );
  NAND2_X1 U793 ( .A1(n752), .A2(n753), .ZN(n799) );
  NOR2_X1 U794 ( .A1(n624), .A2(n745), .ZN(n754) );
  INV_X1 U795 ( .A(n800), .ZN(n797) );
  NOR2_X1 U796 ( .A1(n752), .A2(n753), .ZN(n800) );
  NOR2_X1 U797 ( .A1(n801), .A2(n802), .ZN(n753) );
  INV_X1 U798 ( .A(n803), .ZN(n802) );
  NAND2_X1 U799 ( .A1(n748), .A2(n804), .ZN(n803) );
  NAND2_X1 U800 ( .A1(n750), .A2(n738), .ZN(n804) );
  NOR2_X1 U801 ( .A1(n745), .A2(n629), .ZN(n748) );
  NOR2_X1 U802 ( .A1(n738), .A2(n750), .ZN(n801) );
  NAND2_X1 U803 ( .A1(n805), .A2(n806), .ZN(n750) );
  NAND2_X1 U804 ( .A1(n807), .A2(n808), .ZN(n806) );
  NAND2_X1 U805 ( .A1(n680), .A2(n809), .ZN(n738) );
  NOR2_X1 U806 ( .A1(n745), .A2(n632), .ZN(n680) );
  XOR2_X1 U807 ( .A(n810), .B(n811), .Z(n745) );
  XNOR2_X1 U808 ( .A(c_4_), .B(d_4_), .ZN(n810) );
  XOR2_X1 U809 ( .A(n812), .B(n813), .Z(n752) );
  XOR2_X1 U810 ( .A(n814), .B(n805), .Z(n813) );
  XOR2_X1 U811 ( .A(n815), .B(n816), .Z(n755) );
  XOR2_X1 U812 ( .A(n817), .B(n818), .Z(n816) );
  XNOR2_X1 U813 ( .A(n819), .B(n820), .ZN(n759) );
  XNOR2_X1 U814 ( .A(n821), .B(n822), .ZN(n820) );
  XNOR2_X1 U815 ( .A(n823), .B(n824), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n825), .B(n826), .ZN(n824) );
  XNOR2_X1 U817 ( .A(n827), .B(n828), .ZN(n710) );
  XNOR2_X1 U818 ( .A(n829), .B(n830), .ZN(n828) );
  XNOR2_X1 U819 ( .A(n771), .B(n831), .ZN(n768) );
  XNOR2_X1 U820 ( .A(n773), .B(n774), .ZN(n831) );
  NAND2_X1 U821 ( .A1(n742), .A2(n578), .ZN(n774) );
  NOR2_X1 U822 ( .A1(n832), .A2(n833), .ZN(n773) );
  INV_X1 U823 ( .A(n834), .ZN(n833) );
  NAND2_X1 U824 ( .A1(n827), .A2(n835), .ZN(n834) );
  NAND2_X1 U825 ( .A1(n829), .A2(n830), .ZN(n835) );
  XNOR2_X1 U826 ( .A(n836), .B(n837), .ZN(n827) );
  XNOR2_X1 U827 ( .A(n838), .B(n839), .ZN(n837) );
  NOR2_X1 U828 ( .A1(n830), .A2(n829), .ZN(n832) );
  NOR2_X1 U829 ( .A1(n840), .A2(n841), .ZN(n829) );
  INV_X1 U830 ( .A(n842), .ZN(n841) );
  NAND2_X1 U831 ( .A1(n823), .A2(n843), .ZN(n842) );
  NAND2_X1 U832 ( .A1(n825), .A2(n826), .ZN(n843) );
  XOR2_X1 U833 ( .A(n844), .B(n845), .Z(n823) );
  XOR2_X1 U834 ( .A(n846), .B(n847), .Z(n844) );
  NOR2_X1 U835 ( .A1(n826), .A2(n825), .ZN(n840) );
  NOR2_X1 U836 ( .A1(n848), .A2(n849), .ZN(n825) );
  INV_X1 U837 ( .A(n850), .ZN(n849) );
  NAND2_X1 U838 ( .A1(n819), .A2(n851), .ZN(n850) );
  NAND2_X1 U839 ( .A1(n821), .A2(n822), .ZN(n851) );
  XNOR2_X1 U840 ( .A(n852), .B(n853), .ZN(n819) );
  NAND2_X1 U841 ( .A1(n854), .A2(n855), .ZN(n852) );
  NOR2_X1 U842 ( .A1(n822), .A2(n821), .ZN(n848) );
  NOR2_X1 U843 ( .A1(n856), .A2(n857), .ZN(n821) );
  INV_X1 U844 ( .A(n858), .ZN(n857) );
  NAND2_X1 U845 ( .A1(n815), .A2(n859), .ZN(n858) );
  NAND2_X1 U846 ( .A1(n818), .A2(n817), .ZN(n859) );
  XNOR2_X1 U847 ( .A(n860), .B(n861), .ZN(n815) );
  NOR2_X1 U848 ( .A1(n780), .A2(n629), .ZN(n861) );
  XNOR2_X1 U849 ( .A(n862), .B(n863), .ZN(n860) );
  NOR2_X1 U850 ( .A1(n818), .A2(n817), .ZN(n856) );
  NAND2_X1 U851 ( .A1(n864), .A2(n865), .ZN(n817) );
  NAND2_X1 U852 ( .A1(n866), .A2(n814), .ZN(n865) );
  NAND2_X1 U853 ( .A1(n867), .A2(n742), .ZN(n814) );
  INV_X1 U854 ( .A(n868), .ZN(n866) );
  NOR2_X1 U855 ( .A1(n805), .A2(n812), .ZN(n868) );
  NAND2_X1 U856 ( .A1(n812), .A2(n805), .ZN(n864) );
  NAND2_X1 U857 ( .A1(n809), .A2(n869), .ZN(n805) );
  INV_X1 U858 ( .A(n808), .ZN(n809) );
  NAND2_X1 U859 ( .A1(n742), .A2(n870), .ZN(n808) );
  XOR2_X1 U860 ( .A(n871), .B(n872), .Z(n812) );
  NOR2_X1 U861 ( .A1(n556), .A2(n780), .ZN(n872) );
  NAND2_X1 U862 ( .A1(n743), .A2(n873), .ZN(n871) );
  NAND2_X1 U863 ( .A1(n618), .A2(n742), .ZN(n818) );
  NAND2_X1 U864 ( .A1(n874), .A2(n742), .ZN(n822) );
  NAND2_X1 U865 ( .A1(n875), .A2(n742), .ZN(n826) );
  INV_X1 U866 ( .A(n575), .ZN(n875) );
  NAND2_X1 U867 ( .A1(n876), .A2(n742), .ZN(n830) );
  XOR2_X1 U868 ( .A(n877), .B(n878), .Z(n742) );
  XOR2_X1 U869 ( .A(d_3_), .B(c_3_), .Z(n878) );
  XNOR2_X1 U870 ( .A(n879), .B(n880), .ZN(n771) );
  NAND2_X1 U871 ( .A1(n881), .A2(n882), .ZN(n879) );
  XOR2_X1 U872 ( .A(n883), .B(n884), .Z(n549) );
  INV_X1 U873 ( .A(n885), .ZN(n553) );
  NAND2_X1 U874 ( .A1(n886), .A2(n887), .ZN(n885) );
  XOR2_X1 U875 ( .A(n579), .B(n888), .Z(n886) );
  NOR2_X1 U876 ( .A1(n889), .A2(n887), .ZN(n552) );
  NAND2_X1 U877 ( .A1(n884), .A2(n883), .ZN(n887) );
  NAND2_X1 U878 ( .A1(n890), .A2(n891), .ZN(n883) );
  NAND2_X1 U879 ( .A1(n892), .A2(n893), .ZN(n891) );
  NOR2_X1 U880 ( .A1(n894), .A2(n600), .ZN(n892) );
  INV_X1 U881 ( .A(n578), .ZN(n600) );
  NOR2_X1 U882 ( .A1(n777), .A2(n778), .ZN(n894) );
  NAND2_X1 U883 ( .A1(n777), .A2(n778), .ZN(n890) );
  NAND2_X1 U884 ( .A1(n881), .A2(n895), .ZN(n778) );
  NAND2_X1 U885 ( .A1(n880), .A2(n882), .ZN(n895) );
  NAND2_X1 U886 ( .A1(n896), .A2(n897), .ZN(n882) );
  NAND2_X1 U887 ( .A1(n876), .A2(n893), .ZN(n897) );
  INV_X1 U888 ( .A(n898), .ZN(n896) );
  XOR2_X1 U889 ( .A(n899), .B(n900), .Z(n880) );
  XOR2_X1 U890 ( .A(n901), .B(n902), .Z(n899) );
  NAND2_X1 U891 ( .A1(n898), .A2(n876), .ZN(n881) );
  NOR2_X1 U892 ( .A1(n903), .A2(n904), .ZN(n898) );
  NOR2_X1 U893 ( .A1(n905), .A2(n838), .ZN(n904) );
  NOR2_X1 U894 ( .A1(n575), .A2(n780), .ZN(n838) );
  INV_X1 U895 ( .A(n906), .ZN(n905) );
  NAND2_X1 U896 ( .A1(n836), .A2(n839), .ZN(n906) );
  NOR2_X1 U897 ( .A1(n839), .A2(n836), .ZN(n903) );
  XNOR2_X1 U898 ( .A(n907), .B(n908), .ZN(n836) );
  XNOR2_X1 U899 ( .A(n909), .B(n910), .ZN(n908) );
  NAND2_X1 U900 ( .A1(n911), .A2(n912), .ZN(n839) );
  NAND2_X1 U901 ( .A1(n847), .A2(n913), .ZN(n912) );
  INV_X1 U902 ( .A(n914), .ZN(n913) );
  NOR2_X1 U903 ( .A1(n846), .A2(n845), .ZN(n914) );
  NOR2_X1 U904 ( .A1(n570), .A2(n780), .ZN(n847) );
  NAND2_X1 U905 ( .A1(n845), .A2(n846), .ZN(n911) );
  NAND2_X1 U906 ( .A1(n854), .A2(n915), .ZN(n846) );
  NAND2_X1 U907 ( .A1(n853), .A2(n855), .ZN(n915) );
  NAND2_X1 U908 ( .A1(n916), .A2(n917), .ZN(n855) );
  NAND2_X1 U909 ( .A1(n618), .A2(n893), .ZN(n917) );
  INV_X1 U910 ( .A(n918), .ZN(n916) );
  XNOR2_X1 U911 ( .A(n919), .B(n920), .ZN(n853) );
  XNOR2_X1 U912 ( .A(n921), .B(n922), .ZN(n920) );
  NAND2_X1 U913 ( .A1(n923), .A2(n870), .ZN(n919) );
  NAND2_X1 U914 ( .A1(n618), .A2(n918), .ZN(n854) );
  NAND2_X1 U915 ( .A1(n924), .A2(n925), .ZN(n918) );
  NAND2_X1 U916 ( .A1(n926), .A2(n867), .ZN(n925) );
  INV_X1 U917 ( .A(n629), .ZN(n867) );
  NOR2_X1 U918 ( .A1(n927), .A2(n780), .ZN(n926) );
  NOR2_X1 U919 ( .A1(n862), .A2(n863), .ZN(n927) );
  NAND2_X1 U920 ( .A1(n863), .A2(n862), .ZN(n924) );
  NOR2_X1 U921 ( .A1(n928), .A2(n929), .ZN(n862) );
  NOR2_X1 U922 ( .A1(n930), .A2(n931), .ZN(n929) );
  INV_X1 U923 ( .A(n922), .ZN(n928) );
  INV_X1 U924 ( .A(n932), .ZN(n863) );
  NAND2_X1 U925 ( .A1(n931), .A2(n869), .ZN(n932) );
  INV_X1 U926 ( .A(n807), .ZN(n869) );
  NAND2_X1 U927 ( .A1(n743), .A2(n893), .ZN(n807) );
  INV_X1 U928 ( .A(n780), .ZN(n893) );
  XNOR2_X1 U929 ( .A(n933), .B(n934), .ZN(n780) );
  XOR2_X1 U930 ( .A(d_2_), .B(c_2_), .Z(n934) );
  XOR2_X1 U931 ( .A(n935), .B(n936), .Z(n845) );
  XOR2_X1 U932 ( .A(n937), .B(n938), .Z(n935) );
  XNOR2_X1 U933 ( .A(n939), .B(n940), .ZN(n777) );
  XNOR2_X1 U934 ( .A(n941), .B(n942), .ZN(n940) );
  XOR2_X1 U935 ( .A(n943), .B(n944), .Z(n884) );
  XOR2_X1 U936 ( .A(n945), .B(n946), .Z(n943) );
  INV_X1 U937 ( .A(n947), .ZN(n889) );
  NOR2_X1 U938 ( .A1(n579), .A2(n888), .ZN(n947) );
  NAND2_X1 U939 ( .A1(n578), .A2(n923), .ZN(n888) );
  NAND2_X1 U940 ( .A1(n948), .A2(n949), .ZN(n579) );
  NAND2_X1 U941 ( .A1(n944), .A2(n950), .ZN(n949) );
  NAND2_X1 U942 ( .A1(n946), .A2(n945), .ZN(n950) );
  NOR2_X1 U943 ( .A1(n605), .A2(n951), .ZN(n944) );
  INV_X1 U944 ( .A(n952), .ZN(n948) );
  NOR2_X1 U945 ( .A1(n945), .A2(n946), .ZN(n952) );
  NOR2_X1 U946 ( .A1(n953), .A2(n954), .ZN(n946) );
  INV_X1 U947 ( .A(n955), .ZN(n954) );
  NAND2_X1 U948 ( .A1(n939), .A2(n956), .ZN(n955) );
  NAND2_X1 U949 ( .A1(n941), .A2(n942), .ZN(n956) );
  NOR2_X1 U950 ( .A1(n575), .A2(n951), .ZN(n939) );
  NOR2_X1 U951 ( .A1(n942), .A2(n941), .ZN(n953) );
  NOR2_X1 U952 ( .A1(n957), .A2(n958), .ZN(n941) );
  INV_X1 U953 ( .A(n959), .ZN(n958) );
  NAND2_X1 U954 ( .A1(n900), .A2(n960), .ZN(n959) );
  NAND2_X1 U955 ( .A1(n902), .A2(n901), .ZN(n960) );
  NOR2_X1 U956 ( .A1(n575), .A2(n961), .ZN(n900) );
  XNOR2_X1 U957 ( .A(n962), .B(n963), .ZN(n575) );
  XOR2_X1 U958 ( .A(b_2_), .B(a_2_), .Z(n963) );
  NOR2_X1 U959 ( .A1(n901), .A2(n902), .ZN(n957) );
  NOR2_X1 U960 ( .A1(n964), .A2(n965), .ZN(n902) );
  INV_X1 U961 ( .A(n966), .ZN(n965) );
  NAND2_X1 U962 ( .A1(n907), .A2(n967), .ZN(n966) );
  NAND2_X1 U963 ( .A1(n909), .A2(n910), .ZN(n967) );
  NOR2_X1 U964 ( .A1(n624), .A2(n951), .ZN(n907) );
  NOR2_X1 U965 ( .A1(n910), .A2(n909), .ZN(n964) );
  INV_X1 U966 ( .A(n968), .ZN(n909) );
  NAND2_X1 U967 ( .A1(n969), .A2(n970), .ZN(n968) );
  NAND2_X1 U968 ( .A1(n936), .A2(n971), .ZN(n970) );
  INV_X1 U969 ( .A(n972), .ZN(n971) );
  NOR2_X1 U970 ( .A1(n937), .A2(n938), .ZN(n972) );
  NOR2_X1 U971 ( .A1(n629), .A2(n951), .ZN(n936) );
  NAND2_X1 U972 ( .A1(n938), .A2(n937), .ZN(n969) );
  NAND2_X1 U973 ( .A1(n922), .A2(n973), .ZN(n937) );
  NAND2_X1 U974 ( .A1(n974), .A2(n921), .ZN(n973) );
  NOR2_X1 U975 ( .A1(n629), .A2(n961), .ZN(n921) );
  XNOR2_X1 U976 ( .A(n975), .B(n976), .ZN(n629) );
  XOR2_X1 U977 ( .A(b_5_), .B(a_5_), .Z(n976) );
  NOR2_X1 U978 ( .A1(n556), .A2(n951), .ZN(n974) );
  NAND2_X1 U979 ( .A1(n931), .A2(n930), .ZN(n922) );
  NOR2_X1 U980 ( .A1(n632), .A2(n951), .ZN(n930) );
  INV_X1 U981 ( .A(n923), .ZN(n951) );
  INV_X1 U982 ( .A(n743), .ZN(n632) );
  NOR2_X1 U983 ( .A1(n977), .A2(n978), .ZN(n743) );
  NOR2_X1 U984 ( .A1(a_7_), .A2(b_7_), .ZN(n978) );
  NOR2_X1 U985 ( .A1(n961), .A2(n556), .ZN(n931) );
  INV_X1 U986 ( .A(n870), .ZN(n556) );
  XOR2_X1 U987 ( .A(n977), .B(n979), .Z(n870) );
  XNOR2_X1 U988 ( .A(b_6_), .B(n980), .ZN(n979) );
  NOR2_X1 U989 ( .A1(n624), .A2(n961), .ZN(n938) );
  INV_X1 U990 ( .A(n618), .ZN(n624) );
  XNOR2_X1 U991 ( .A(n981), .B(n982), .ZN(n618) );
  XNOR2_X1 U992 ( .A(a_4_), .B(b_4_), .ZN(n981) );
  NAND2_X1 U993 ( .A1(n874), .A2(n873), .ZN(n910) );
  NAND2_X1 U994 ( .A1(n874), .A2(n923), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n983), .B(n984), .ZN(n923) );
  XOR2_X1 U996 ( .A(d_0_), .B(c_0_), .Z(n984) );
  NAND2_X1 U997 ( .A1(n985), .A2(n986), .ZN(n983) );
  NAND2_X1 U998 ( .A1(n987), .A2(n988), .ZN(n986) );
  NAND2_X1 U999 ( .A1(c_1_), .A2(n989), .ZN(n987) );
  INV_X1 U1000 ( .A(n990), .ZN(n985) );
  NOR2_X1 U1001 ( .A1(n989), .A2(c_1_), .ZN(n990) );
  INV_X1 U1002 ( .A(n570), .ZN(n874) );
  XNOR2_X1 U1003 ( .A(n991), .B(n992), .ZN(n570) );
  XOR2_X1 U1004 ( .A(b_3_), .B(a_3_), .Z(n992) );
  NAND2_X1 U1005 ( .A1(n876), .A2(n873), .ZN(n942) );
  INV_X1 U1006 ( .A(n605), .ZN(n876) );
  XNOR2_X1 U1007 ( .A(n993), .B(n994), .ZN(n605) );
  XNOR2_X1 U1008 ( .A(n995), .B(a_1_), .ZN(n994) );
  NAND2_X1 U1009 ( .A1(n873), .A2(n578), .ZN(n945) );
  XNOR2_X1 U1010 ( .A(n996), .B(n997), .ZN(n578) );
  XOR2_X1 U1011 ( .A(b_0_), .B(a_0_), .Z(n997) );
  NAND2_X1 U1012 ( .A1(n998), .A2(n999), .ZN(n996) );
  NAND2_X1 U1013 ( .A1(n1000), .A2(n995), .ZN(n999) );
  INV_X1 U1014 ( .A(b_1_), .ZN(n995) );
  NAND2_X1 U1015 ( .A1(a_1_), .A2(n993), .ZN(n1000) );
  INV_X1 U1016 ( .A(n1001), .ZN(n998) );
  NOR2_X1 U1017 ( .A1(n993), .A2(a_1_), .ZN(n1001) );
  NAND2_X1 U1018 ( .A1(n1002), .A2(n1003), .ZN(n993) );
  NAND2_X1 U1019 ( .A1(b_2_), .A2(n1004), .ZN(n1003) );
  INV_X1 U1020 ( .A(n1005), .ZN(n1004) );
  NOR2_X1 U1021 ( .A1(n962), .A2(a_2_), .ZN(n1005) );
  NAND2_X1 U1022 ( .A1(a_2_), .A2(n962), .ZN(n1002) );
  NAND2_X1 U1023 ( .A1(n1006), .A2(n1007), .ZN(n962) );
  NAND2_X1 U1024 ( .A1(b_3_), .A2(n1008), .ZN(n1007) );
  INV_X1 U1025 ( .A(n1009), .ZN(n1008) );
  NOR2_X1 U1026 ( .A1(n991), .A2(a_3_), .ZN(n1009) );
  NAND2_X1 U1027 ( .A1(a_3_), .A2(n991), .ZN(n1006) );
  NAND2_X1 U1028 ( .A1(n1010), .A2(n1011), .ZN(n991) );
  NAND2_X1 U1029 ( .A1(b_4_), .A2(n1012), .ZN(n1011) );
  INV_X1 U1030 ( .A(n1013), .ZN(n1012) );
  NOR2_X1 U1031 ( .A1(n982), .A2(a_4_), .ZN(n1013) );
  NAND2_X1 U1032 ( .A1(a_4_), .A2(n982), .ZN(n1010) );
  NAND2_X1 U1033 ( .A1(n1014), .A2(n1015), .ZN(n982) );
  NAND2_X1 U1034 ( .A1(b_5_), .A2(n1016), .ZN(n1015) );
  INV_X1 U1035 ( .A(n1017), .ZN(n1016) );
  NOR2_X1 U1036 ( .A1(n975), .A2(a_5_), .ZN(n1017) );
  NAND2_X1 U1037 ( .A1(a_5_), .A2(n975), .ZN(n1014) );
  NAND2_X1 U1038 ( .A1(n1018), .A2(n1019), .ZN(n975) );
  NAND2_X1 U1039 ( .A1(b_6_), .A2(n1020), .ZN(n1019) );
  NAND2_X1 U1040 ( .A1(n980), .A2(n1021), .ZN(n1020) );
  INV_X1 U1041 ( .A(a_6_), .ZN(n980) );
  NAND2_X1 U1042 ( .A1(n977), .A2(a_6_), .ZN(n1018) );
  INV_X1 U1043 ( .A(n1021), .ZN(n977) );
  NAND2_X1 U1044 ( .A1(b_7_), .A2(a_7_), .ZN(n1021) );
  INV_X1 U1045 ( .A(n961), .ZN(n873) );
  XNOR2_X1 U1046 ( .A(n989), .B(n1022), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(n988), .B(c_1_), .ZN(n1022) );
  INV_X1 U1048 ( .A(d_1_), .ZN(n988) );
  NAND2_X1 U1049 ( .A1(n1023), .A2(n1024), .ZN(n989) );
  NAND2_X1 U1050 ( .A1(d_2_), .A2(n1025), .ZN(n1024) );
  INV_X1 U1051 ( .A(n1026), .ZN(n1025) );
  NOR2_X1 U1052 ( .A1(n933), .A2(c_2_), .ZN(n1026) );
  NAND2_X1 U1053 ( .A1(c_2_), .A2(n933), .ZN(n1023) );
  NAND2_X1 U1054 ( .A1(n1027), .A2(n1028), .ZN(n933) );
  NAND2_X1 U1055 ( .A1(d_3_), .A2(n1029), .ZN(n1028) );
  INV_X1 U1056 ( .A(n1030), .ZN(n1029) );
  NOR2_X1 U1057 ( .A1(n877), .A2(c_3_), .ZN(n1030) );
  NAND2_X1 U1058 ( .A1(c_3_), .A2(n877), .ZN(n1027) );
  NAND2_X1 U1059 ( .A1(n1031), .A2(n1032), .ZN(n877) );
  NAND2_X1 U1060 ( .A1(d_4_), .A2(n1033), .ZN(n1032) );
  INV_X1 U1061 ( .A(n1034), .ZN(n1033) );
  NOR2_X1 U1062 ( .A1(n811), .A2(c_4_), .ZN(n1034) );
  NAND2_X1 U1063 ( .A1(c_4_), .A2(n811), .ZN(n1031) );
  NAND2_X1 U1064 ( .A1(n1035), .A2(n1036), .ZN(n811) );
  NAND2_X1 U1065 ( .A1(d_5_), .A2(n1037), .ZN(n1036) );
  INV_X1 U1066 ( .A(n1038), .ZN(n1037) );
  NOR2_X1 U1067 ( .A1(n746), .A2(c_5_), .ZN(n1038) );
  NAND2_X1 U1068 ( .A1(c_5_), .A2(n746), .ZN(n1035) );
  NAND2_X1 U1069 ( .A1(n1039), .A2(n1040), .ZN(n746) );
  NAND2_X1 U1070 ( .A1(d_6_), .A2(n1041), .ZN(n1040) );
  INV_X1 U1071 ( .A(n1042), .ZN(n1041) );
  NOR2_X1 U1072 ( .A1(c_6_), .A2(n635), .ZN(n1042) );
  NAND2_X1 U1073 ( .A1(c_6_), .A2(n635), .ZN(n1039) );
  INV_X1 U1074 ( .A(n1043), .ZN(n635) );
  NAND2_X1 U1075 ( .A1(d_7_), .A2(c_7_), .ZN(n1043) );
endmodule

