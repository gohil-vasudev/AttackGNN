module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n670_, new_n456_, new_n170_, new_n246_, new_n682_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n605_, new_n107_, new_n182_, new_n407_, new_n625_, new_n151_, new_n513_, new_n592_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n563_, new_n148_, new_n662_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n217_, new_n269_, new_n512_, new_n129_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n106_, N69 );
nand g001 ( new_n107_, new_n106_, N65 );
not g002 ( new_n108_, N65 );
nand g003 ( new_n109_, new_n108_, N69 );
not g004 ( new_n110_, N77 );
nand g005 ( new_n111_, new_n110_, N73 );
not g006 ( new_n112_, N73 );
nand g007 ( new_n113_, new_n112_, N77 );
nand g008 ( new_n114_, new_n111_, new_n113_ );
nand g009 ( new_n115_, new_n114_, new_n107_, new_n109_ );
nand g010 ( new_n116_, new_n107_, new_n109_ );
nand g011 ( new_n117_, new_n116_, new_n111_, new_n113_ );
nand g012 ( new_n118_, new_n115_, new_n117_ );
not g013 ( new_n119_, N93 );
nand g014 ( new_n120_, new_n119_, N89 );
not g015 ( new_n121_, N89 );
nand g016 ( new_n122_, new_n121_, N93 );
not g017 ( new_n123_, N85 );
nand g018 ( new_n124_, new_n123_, N81 );
not g019 ( new_n125_, N81 );
nand g020 ( new_n126_, new_n125_, N85 );
nand g021 ( new_n127_, new_n124_, new_n126_ );
nand g022 ( new_n128_, new_n127_, new_n120_, new_n122_ );
nand g023 ( new_n129_, new_n120_, new_n122_ );
nand g024 ( new_n130_, new_n129_, new_n124_, new_n126_ );
nand g025 ( new_n131_, new_n128_, new_n130_ );
not g026 ( new_n132_, new_n131_ );
nand g027 ( new_n133_, new_n132_, new_n118_ );
not g028 ( new_n134_, new_n118_ );
nand g029 ( new_n135_, new_n134_, new_n131_ );
nand g030 ( new_n136_, new_n133_, new_n135_ );
nand g031 ( new_n137_, N129, N137 );
nand g032 ( new_n138_, new_n136_, new_n137_ );
nand g033 ( new_n139_, new_n133_, new_n135_, N129, N137 );
nand g034 ( new_n140_, new_n138_, new_n139_ );
not g035 ( new_n141_, keyIn_0_9 );
not g036 ( new_n142_, N49 );
nand g037 ( new_n143_, new_n142_, N33 );
not g038 ( new_n144_, N33 );
nand g039 ( new_n145_, new_n144_, N49 );
not g040 ( new_n146_, N17 );
nand g041 ( new_n147_, new_n146_, N1 );
not g042 ( new_n148_, N1 );
nand g043 ( new_n149_, new_n148_, N17 );
nand g044 ( new_n150_, new_n147_, new_n149_ );
nand g045 ( new_n151_, new_n150_, new_n143_, new_n145_ );
nand g046 ( new_n152_, new_n143_, new_n145_ );
nand g047 ( new_n153_, new_n152_, new_n147_, new_n149_ );
nand g048 ( new_n154_, new_n151_, new_n153_ );
nand g049 ( new_n155_, new_n154_, new_n141_ );
nand g050 ( new_n156_, new_n151_, new_n153_, keyIn_0_9 );
nand g051 ( new_n157_, new_n155_, new_n156_ );
nand g052 ( new_n158_, new_n140_, new_n157_ );
nand g053 ( new_n159_, new_n138_, new_n139_, new_n155_, new_n156_ );
nand g054 ( new_n160_, new_n158_, new_n159_ );
not g055 ( new_n161_, keyIn_0_24 );
not g056 ( new_n162_, new_n160_ );
not g057 ( new_n163_, N117 );
nand g058 ( new_n164_, new_n163_, N113 );
not g059 ( new_n165_, N113 );
nand g060 ( new_n166_, new_n165_, N117 );
nand g061 ( new_n167_, new_n164_, new_n166_ );
nand g062 ( new_n168_, new_n167_, keyIn_0_4 );
not g063 ( new_n169_, keyIn_0_4 );
nand g064 ( new_n170_, new_n164_, new_n166_, new_n169_ );
nand g065 ( new_n171_, new_n168_, new_n170_ );
not g066 ( new_n172_, N125 );
nand g067 ( new_n173_, new_n172_, N121 );
not g068 ( new_n174_, N121 );
nand g069 ( new_n175_, new_n174_, N125 );
nand g070 ( new_n176_, new_n173_, new_n175_ );
nand g071 ( new_n177_, new_n171_, new_n176_ );
nand g072 ( new_n178_, new_n168_, new_n170_, new_n173_, new_n175_ );
nand g073 ( new_n179_, new_n177_, new_n178_ );
not g074 ( new_n180_, N109 );
nand g075 ( new_n181_, new_n180_, N105 );
not g076 ( new_n182_, N105 );
nand g077 ( new_n183_, new_n182_, N109 );
nand g078 ( new_n184_, new_n181_, new_n183_ );
nand g079 ( new_n185_, new_n184_, keyIn_0_3 );
not g080 ( new_n186_, keyIn_0_3 );
nand g081 ( new_n187_, new_n181_, new_n183_, new_n186_ );
not g082 ( new_n188_, N101 );
nand g083 ( new_n189_, new_n188_, N97 );
not g084 ( new_n190_, N97 );
nand g085 ( new_n191_, new_n190_, N101 );
nand g086 ( new_n192_, new_n189_, new_n191_ );
nand g087 ( new_n193_, new_n185_, new_n187_, new_n192_ );
nand g088 ( new_n194_, new_n185_, new_n187_ );
nand g089 ( new_n195_, new_n194_, new_n189_, new_n191_ );
nand g090 ( new_n196_, new_n195_, new_n193_ );
not g091 ( new_n197_, new_n196_ );
nand g092 ( new_n198_, new_n197_, new_n179_ );
not g093 ( new_n199_, new_n179_ );
nand g094 ( new_n200_, new_n199_, new_n196_ );
nand g095 ( new_n201_, new_n198_, new_n200_ );
nand g096 ( new_n202_, N130, N137 );
nand g097 ( new_n203_, new_n201_, new_n202_ );
nand g098 ( new_n204_, new_n198_, new_n200_, N130, N137 );
not g099 ( new_n205_, N21 );
nand g100 ( new_n206_, new_n205_, N5 );
not g101 ( new_n207_, N5 );
nand g102 ( new_n208_, new_n207_, N21 );
not g103 ( new_n209_, N53 );
nand g104 ( new_n210_, new_n209_, N37 );
not g105 ( new_n211_, N37 );
nand g106 ( new_n212_, new_n211_, N53 );
nand g107 ( new_n213_, new_n210_, new_n212_ );
nand g108 ( new_n214_, new_n213_, new_n206_, new_n208_ );
nand g109 ( new_n215_, new_n206_, new_n208_ );
nand g110 ( new_n216_, new_n215_, new_n210_, new_n212_ );
nand g111 ( new_n217_, new_n214_, new_n216_ );
nand g112 ( new_n218_, new_n203_, new_n204_, new_n217_ );
nand g113 ( new_n219_, new_n203_, new_n204_ );
nand g114 ( new_n220_, new_n219_, new_n214_, new_n216_ );
nand g115 ( new_n221_, new_n220_, new_n218_ );
nand g116 ( new_n222_, new_n196_, new_n134_ );
nand g117 ( new_n223_, new_n197_, new_n118_ );
nand g118 ( new_n224_, new_n223_, new_n222_ );
nand g119 ( new_n225_, N131, N137 );
nand g120 ( new_n226_, new_n224_, new_n225_ );
nand g121 ( new_n227_, new_n223_, N131, N137, new_n222_ );
not g122 ( new_n228_, keyIn_0_6 );
not g123 ( new_n229_, N57 );
nand g124 ( new_n230_, new_n229_, N41 );
not g125 ( new_n231_, N41 );
nand g126 ( new_n232_, new_n231_, N57 );
nand g127 ( new_n233_, new_n230_, new_n232_ );
nand g128 ( new_n234_, new_n233_, new_n228_ );
nand g129 ( new_n235_, new_n230_, new_n232_, keyIn_0_6 );
not g130 ( new_n236_, N9 );
nor g131 ( new_n237_, new_n236_, N25 );
not g132 ( new_n238_, N25 );
nor g133 ( new_n239_, new_n238_, N9 );
nor g134 ( new_n240_, new_n237_, new_n239_ );
nand g135 ( new_n241_, new_n234_, new_n235_, new_n240_ );
nand g136 ( new_n242_, new_n234_, new_n235_ );
not g137 ( new_n243_, new_n240_ );
nand g138 ( new_n244_, new_n242_, new_n243_ );
nand g139 ( new_n245_, new_n244_, new_n241_ );
nand g140 ( new_n246_, new_n226_, new_n227_, new_n245_ );
nand g141 ( new_n247_, new_n226_, new_n227_ );
nand g142 ( new_n248_, new_n247_, new_n241_, new_n244_ );
nand g143 ( new_n249_, new_n248_, new_n246_ );
nand g144 ( new_n250_, new_n221_, new_n249_, keyIn_0_12 );
not g145 ( new_n251_, new_n221_ );
nand g146 ( new_n252_, new_n249_, keyIn_0_12 );
nand g147 ( new_n253_, new_n252_, new_n251_ );
nand g148 ( new_n254_, new_n179_, new_n132_ );
nand g149 ( new_n255_, new_n199_, new_n131_ );
nand g150 ( new_n256_, new_n255_, new_n254_ );
nand g151 ( new_n257_, N132, N137 );
nand g152 ( new_n258_, new_n256_, new_n257_ );
nand g153 ( new_n259_, new_n255_, N132, N137, new_n254_ );
not g154 ( new_n260_, N29 );
nand g155 ( new_n261_, new_n260_, N13 );
not g156 ( new_n262_, N13 );
nand g157 ( new_n263_, new_n262_, N29 );
not g158 ( new_n264_, N61 );
nand g159 ( new_n265_, new_n264_, N45 );
not g160 ( new_n266_, N45 );
nand g161 ( new_n267_, new_n266_, N61 );
nand g162 ( new_n268_, new_n265_, new_n267_ );
nand g163 ( new_n269_, new_n268_, new_n261_, new_n263_ );
nand g164 ( new_n270_, new_n261_, new_n263_ );
nand g165 ( new_n271_, new_n270_, new_n265_, new_n267_ );
nand g166 ( new_n272_, new_n269_, new_n271_ );
nand g167 ( new_n273_, new_n258_, new_n259_, new_n272_ );
nand g168 ( new_n274_, new_n258_, new_n259_ );
nand g169 ( new_n275_, new_n274_, new_n269_, new_n271_ );
nand g170 ( new_n276_, new_n275_, new_n273_ );
not g171 ( new_n277_, new_n276_ );
nand g172 ( new_n278_, new_n253_, new_n162_, new_n250_, new_n277_ );
nor g173 ( new_n279_, new_n277_, new_n249_ );
nand g174 ( new_n280_, new_n160_, keyIn_0_11 );
not g175 ( new_n281_, keyIn_0_11 );
nand g176 ( new_n282_, new_n162_, new_n281_ );
nand g177 ( new_n283_, new_n282_, new_n280_ );
not g178 ( new_n284_, new_n283_ );
nand g179 ( new_n285_, new_n279_, new_n251_, new_n284_ );
nand g180 ( new_n286_, new_n285_, keyIn_0_19 );
not g181 ( new_n287_, keyIn_0_19 );
nand g182 ( new_n288_, new_n279_, new_n284_, new_n287_, new_n251_ );
nand g183 ( new_n289_, new_n286_, new_n288_ );
nand g184 ( new_n290_, new_n221_, keyIn_0_13 );
not g185 ( new_n291_, keyIn_0_13 );
nand g186 ( new_n292_, new_n251_, new_n291_ );
nand g187 ( new_n293_, new_n292_, new_n290_ );
nor g188 ( new_n294_, new_n249_, new_n276_, new_n162_ );
nand g189 ( new_n295_, new_n293_, new_n294_ );
nand g190 ( new_n296_, new_n289_, new_n278_, new_n295_ );
nand g191 ( new_n297_, new_n209_, N49 );
nand g192 ( new_n298_, new_n142_, N53 );
nand g193 ( new_n299_, new_n264_, N57 );
nand g194 ( new_n300_, new_n229_, N61 );
nand g195 ( new_n301_, new_n299_, new_n300_ );
nand g196 ( new_n302_, new_n301_, new_n297_, new_n298_ );
nand g197 ( new_n303_, new_n297_, new_n298_ );
nand g198 ( new_n304_, new_n303_, new_n299_, new_n300_ );
nand g199 ( new_n305_, new_n302_, new_n304_ );
not g200 ( new_n306_, keyIn_0_8 );
nand g201 ( new_n307_, new_n266_, N41 );
nand g202 ( new_n308_, new_n231_, N45 );
nand g203 ( new_n309_, new_n307_, new_n308_ );
nand g204 ( new_n310_, new_n309_, keyIn_0_2 );
not g205 ( new_n311_, keyIn_0_2 );
nand g206 ( new_n312_, new_n307_, new_n308_, new_n311_ );
nand g207 ( new_n313_, new_n310_, new_n312_ );
not g208 ( new_n314_, keyIn_0_1 );
nand g209 ( new_n315_, new_n211_, N33 );
nand g210 ( new_n316_, new_n144_, N37 );
nand g211 ( new_n317_, new_n315_, new_n316_, new_n314_ );
nand g212 ( new_n318_, new_n315_, new_n316_ );
nand g213 ( new_n319_, new_n318_, keyIn_0_1 );
nand g214 ( new_n320_, new_n313_, new_n317_, new_n319_ );
nand g215 ( new_n321_, new_n319_, new_n317_ );
nand g216 ( new_n322_, new_n321_, new_n310_, new_n312_ );
nand g217 ( new_n323_, new_n320_, new_n322_ );
nand g218 ( new_n324_, new_n323_, new_n306_ );
nand g219 ( new_n325_, new_n320_, new_n322_, keyIn_0_8 );
nand g220 ( new_n326_, new_n324_, new_n325_ );
nand g221 ( new_n327_, new_n326_, new_n305_ );
not g222 ( new_n328_, new_n305_ );
nand g223 ( new_n329_, new_n324_, new_n328_, new_n325_ );
nand g224 ( new_n330_, new_n327_, new_n329_ );
nand g225 ( new_n331_, N134, N137 );
nand g226 ( new_n332_, new_n330_, new_n331_ );
nand g227 ( new_n333_, new_n327_, N134, N137, new_n329_ );
nand g228 ( new_n334_, new_n332_, new_n333_ );
nand g229 ( new_n335_, new_n123_, N69 );
nand g230 ( new_n336_, new_n106_, N85 );
nand g231 ( new_n337_, new_n163_, N101 );
nand g232 ( new_n338_, new_n188_, N117 );
nand g233 ( new_n339_, new_n337_, new_n338_ );
nand g234 ( new_n340_, new_n339_, new_n335_, new_n336_ );
nand g235 ( new_n341_, new_n335_, new_n336_ );
nand g236 ( new_n342_, new_n341_, new_n337_, new_n338_ );
nand g237 ( new_n343_, new_n340_, new_n342_ );
not g238 ( new_n344_, new_n343_ );
nand g239 ( new_n345_, new_n334_, new_n344_ );
nand g240 ( new_n346_, new_n332_, new_n333_, new_n343_ );
nand g241 ( new_n347_, new_n345_, new_n346_ );
nand g242 ( new_n348_, new_n347_, keyIn_0_14 );
not g243 ( new_n349_, new_n348_ );
not g244 ( new_n350_, keyIn_0_14 );
not g245 ( new_n351_, new_n347_ );
nand g246 ( new_n352_, new_n351_, new_n350_ );
not g247 ( new_n353_, new_n352_ );
nand g248 ( new_n354_, new_n205_, N17 );
nand g249 ( new_n355_, new_n146_, N21 );
nand g250 ( new_n356_, new_n354_, new_n355_ );
nand g251 ( new_n357_, new_n356_, keyIn_0_0 );
not g252 ( new_n358_, keyIn_0_0 );
nand g253 ( new_n359_, new_n354_, new_n355_, new_n358_ );
nor g254 ( new_n360_, new_n238_, N29 );
nor g255 ( new_n361_, new_n260_, N25 );
nor g256 ( new_n362_, new_n360_, new_n361_ );
not g257 ( new_n363_, new_n362_ );
nand g258 ( new_n364_, new_n363_, new_n357_, new_n359_ );
nand g259 ( new_n365_, new_n357_, new_n359_ );
nand g260 ( new_n366_, new_n365_, new_n362_ );
nand g261 ( new_n367_, new_n366_, new_n364_ );
nand g262 ( new_n368_, new_n207_, N1 );
nand g263 ( new_n369_, new_n148_, N5 );
nand g264 ( new_n370_, new_n262_, N9 );
nand g265 ( new_n371_, new_n236_, N13 );
nand g266 ( new_n372_, new_n370_, new_n371_ );
nand g267 ( new_n373_, new_n372_, new_n368_, new_n369_ );
nand g268 ( new_n374_, new_n368_, new_n369_ );
nand g269 ( new_n375_, new_n374_, new_n370_, new_n371_ );
nand g270 ( new_n376_, new_n373_, new_n375_ );
not g271 ( new_n377_, new_n376_ );
nand g272 ( new_n378_, new_n367_, new_n377_ );
nand g273 ( new_n379_, new_n366_, new_n364_, new_n376_ );
nand g274 ( new_n380_, new_n378_, new_n379_ );
nand g275 ( new_n381_, N133, N137 );
nand g276 ( new_n382_, new_n380_, new_n381_ );
nand g277 ( new_n383_, new_n378_, N133, N137, new_n379_ );
nand g278 ( new_n384_, new_n382_, new_n383_ );
nand g279 ( new_n385_, new_n125_, N65 );
nand g280 ( new_n386_, new_n108_, N81 );
nand g281 ( new_n387_, new_n165_, N97 );
nand g282 ( new_n388_, new_n190_, N113 );
nand g283 ( new_n389_, new_n387_, new_n388_ );
nand g284 ( new_n390_, new_n389_, new_n385_, new_n386_ );
nand g285 ( new_n391_, new_n385_, new_n386_ );
nand g286 ( new_n392_, new_n391_, new_n387_, new_n388_ );
nand g287 ( new_n393_, new_n390_, new_n392_ );
not g288 ( new_n394_, new_n393_ );
nand g289 ( new_n395_, new_n384_, new_n394_ );
nand g290 ( new_n396_, new_n382_, new_n383_, new_n393_ );
nand g291 ( new_n397_, new_n395_, new_n396_ );
not g292 ( new_n398_, new_n397_ );
nor g293 ( new_n399_, new_n353_, new_n349_, new_n398_ );
nand g294 ( new_n400_, new_n366_, new_n305_, new_n364_ );
nand g295 ( new_n401_, new_n367_, new_n328_ );
nand g296 ( new_n402_, new_n401_, N136, N137, new_n400_ );
nand g297 ( new_n403_, new_n401_, new_n400_ );
nand g298 ( new_n404_, N136, N137 );
nand g299 ( new_n405_, new_n403_, new_n404_ );
nand g300 ( new_n406_, new_n405_, keyIn_0_10, new_n402_ );
not g301 ( new_n407_, keyIn_0_10 );
nand g302 ( new_n408_, new_n405_, new_n402_ );
nand g303 ( new_n409_, new_n408_, new_n407_ );
nand g304 ( new_n410_, new_n119_, N77 );
nand g305 ( new_n411_, new_n110_, N93 );
nand g306 ( new_n412_, new_n172_, N109 );
nand g307 ( new_n413_, new_n180_, N125 );
nand g308 ( new_n414_, new_n412_, new_n413_ );
nand g309 ( new_n415_, new_n414_, new_n410_, new_n411_ );
nand g310 ( new_n416_, new_n410_, new_n411_ );
nand g311 ( new_n417_, new_n416_, new_n412_, new_n413_ );
nand g312 ( new_n418_, new_n415_, new_n417_ );
nand g313 ( new_n419_, new_n409_, new_n406_, new_n418_ );
nand g314 ( new_n420_, new_n409_, new_n406_ );
not g315 ( new_n421_, new_n418_ );
nand g316 ( new_n422_, new_n420_, new_n421_ );
nand g317 ( new_n423_, new_n422_, new_n419_ );
not g318 ( new_n424_, new_n423_ );
nand g319 ( new_n425_, new_n424_, keyIn_0_15 );
not g320 ( new_n426_, keyIn_0_15 );
nand g321 ( new_n427_, new_n423_, new_n426_ );
nand g322 ( new_n428_, new_n425_, new_n427_ );
nand g323 ( new_n429_, new_n326_, new_n376_ );
nand g324 ( new_n430_, new_n324_, new_n325_, new_n377_ );
nand g325 ( new_n431_, new_n429_, new_n430_ );
nand g326 ( new_n432_, new_n431_, keyIn_0_5 );
not g327 ( new_n433_, keyIn_0_5 );
nand g328 ( new_n434_, new_n429_, new_n433_, new_n430_ );
nand g329 ( new_n435_, new_n432_, new_n434_ );
nand g330 ( new_n436_, N135, N137 );
nand g331 ( new_n437_, new_n435_, new_n436_ );
nand g332 ( new_n438_, new_n432_, N135, N137, new_n434_ );
not g333 ( new_n439_, keyIn_0_7 );
nand g334 ( new_n440_, new_n174_, N105 );
nand g335 ( new_n441_, new_n182_, N121 );
nand g336 ( new_n442_, new_n440_, new_n441_ );
nand g337 ( new_n443_, new_n442_, new_n439_ );
nand g338 ( new_n444_, new_n440_, new_n441_, keyIn_0_7 );
nand g339 ( new_n445_, new_n443_, new_n444_ );
nor g340 ( new_n446_, new_n112_, N89 );
nor g341 ( new_n447_, new_n121_, N73 );
nor g342 ( new_n448_, new_n446_, new_n447_ );
not g343 ( new_n449_, new_n448_ );
nand g344 ( new_n450_, new_n445_, new_n449_ );
nand g345 ( new_n451_, new_n443_, new_n444_, new_n448_ );
nand g346 ( new_n452_, new_n437_, new_n438_, new_n450_, new_n451_ );
nand g347 ( new_n453_, new_n437_, new_n438_ );
nand g348 ( new_n454_, new_n450_, new_n451_ );
nand g349 ( new_n455_, new_n453_, new_n454_ );
nand g350 ( new_n456_, new_n455_, new_n452_ );
nand g351 ( new_n457_, new_n428_, new_n456_ );
not g352 ( new_n458_, new_n457_ );
nand g353 ( new_n459_, new_n296_, new_n399_, new_n458_ );
nand g354 ( new_n460_, new_n459_, new_n161_ );
nand g355 ( new_n461_, new_n296_, keyIn_0_24, new_n399_, new_n458_ );
nand g356 ( new_n462_, new_n460_, new_n461_ );
not g357 ( new_n463_, new_n462_ );
nand g358 ( new_n464_, new_n463_, new_n160_ );
nand g359 ( new_n465_, new_n464_, N1 );
nand g360 ( new_n466_, new_n463_, new_n148_, new_n160_ );
nand g361 ( N724, new_n465_, new_n466_ );
nand g362 ( new_n468_, new_n463_, new_n221_ );
nand g363 ( new_n469_, new_n468_, N5 );
nand g364 ( new_n470_, new_n463_, new_n207_, new_n221_ );
nand g365 ( N725, new_n469_, new_n470_ );
not g366 ( new_n472_, keyIn_0_30 );
nand g367 ( new_n473_, new_n460_, new_n236_, new_n249_, new_n461_ );
nand g368 ( new_n474_, new_n460_, new_n249_, new_n461_ );
nand g369 ( new_n475_, new_n474_, N9 );
nand g370 ( new_n476_, new_n475_, new_n473_ );
nand g371 ( new_n477_, new_n476_, new_n472_ );
nand g372 ( new_n478_, new_n475_, keyIn_0_30, new_n473_ );
nand g373 ( new_n479_, new_n477_, new_n478_ );
not g374 ( N726, new_n479_ );
nand g375 ( new_n481_, new_n460_, new_n276_, new_n461_ );
nand g376 ( new_n482_, new_n481_, N13 );
nand g377 ( new_n483_, new_n463_, new_n262_, new_n276_ );
nand g378 ( new_n484_, new_n483_, new_n482_ );
nand g379 ( new_n485_, new_n484_, keyIn_0_31 );
not g380 ( new_n486_, keyIn_0_31 );
nand g381 ( new_n487_, new_n483_, new_n486_, new_n482_ );
nand g382 ( N727, new_n485_, new_n487_ );
not g383 ( new_n489_, new_n456_ );
nand g384 ( new_n490_, new_n296_, new_n423_, new_n489_ );
not g385 ( new_n491_, new_n490_ );
nand g386 ( new_n492_, new_n351_, new_n397_ );
not g387 ( new_n493_, new_n492_ );
nand g388 ( new_n494_, new_n491_, new_n493_ );
not g389 ( new_n495_, new_n494_ );
nand g390 ( new_n496_, new_n495_, new_n160_ );
nand g391 ( new_n497_, new_n496_, N17 );
nand g392 ( new_n498_, new_n495_, new_n146_, new_n160_ );
nand g393 ( N728, new_n497_, new_n498_ );
nand g394 ( new_n500_, new_n495_, new_n221_ );
nand g395 ( new_n501_, new_n500_, N21 );
nand g396 ( new_n502_, new_n495_, new_n205_, new_n221_ );
nand g397 ( N729, new_n501_, new_n502_ );
not g398 ( new_n504_, keyIn_0_25 );
nand g399 ( new_n505_, new_n495_, new_n249_ );
nand g400 ( new_n506_, new_n505_, new_n504_ );
nand g401 ( new_n507_, new_n495_, keyIn_0_25, new_n249_ );
nand g402 ( new_n508_, new_n506_, new_n238_, new_n507_ );
nand g403 ( new_n509_, new_n506_, new_n507_ );
nand g404 ( new_n510_, new_n509_, N25 );
nand g405 ( N730, new_n510_, new_n508_ );
nand g406 ( new_n512_, new_n495_, new_n276_ );
nand g407 ( new_n513_, new_n512_, keyIn_0_26 );
not g408 ( new_n514_, keyIn_0_26 );
nand g409 ( new_n515_, new_n495_, new_n514_, new_n276_ );
nand g410 ( new_n516_, new_n513_, new_n515_ );
nand g411 ( new_n517_, new_n516_, N29 );
nand g412 ( new_n518_, new_n513_, new_n260_, new_n515_ );
nand g413 ( N731, new_n517_, new_n518_ );
nand g414 ( new_n520_, new_n398_, keyIn_0_16 );
not g415 ( new_n521_, keyIn_0_16 );
nand g416 ( new_n522_, new_n397_, new_n521_ );
nand g417 ( new_n523_, new_n520_, new_n522_ );
nand g418 ( new_n524_, new_n456_, new_n347_, new_n424_, new_n523_ );
not g419 ( new_n525_, new_n524_ );
nand g420 ( new_n526_, new_n296_, new_n160_, new_n525_ );
nand g421 ( new_n527_, new_n526_, N33 );
nand g422 ( new_n528_, new_n296_, new_n144_, new_n160_, new_n525_ );
nand g423 ( N732, new_n527_, new_n528_ );
nand g424 ( new_n530_, new_n296_, new_n221_, new_n525_ );
nand g425 ( new_n531_, new_n530_, N37 );
nand g426 ( new_n532_, new_n296_, new_n211_, new_n221_, new_n525_ );
nand g427 ( N733, new_n531_, new_n532_ );
nand g428 ( new_n534_, new_n296_, new_n249_, new_n525_ );
nand g429 ( new_n535_, new_n534_, N41 );
nand g430 ( new_n536_, new_n296_, new_n231_, new_n249_, new_n525_ );
nand g431 ( N734, new_n535_, new_n536_ );
nand g432 ( new_n538_, new_n296_, new_n276_, new_n525_ );
nand g433 ( new_n539_, new_n538_, N45 );
nand g434 ( new_n540_, new_n296_, new_n266_, new_n276_, new_n525_ );
nand g435 ( N735, new_n539_, new_n540_ );
nand g436 ( new_n542_, new_n398_, keyIn_0_17 );
not g437 ( new_n543_, keyIn_0_17 );
nand g438 ( new_n544_, new_n397_, new_n543_ );
nand g439 ( new_n545_, new_n491_, new_n347_, new_n542_, new_n544_ );
not g440 ( new_n546_, new_n545_ );
nand g441 ( new_n547_, new_n546_, new_n160_ );
nand g442 ( new_n548_, new_n547_, N49 );
nand g443 ( new_n549_, new_n546_, new_n142_, new_n160_ );
nand g444 ( N736, new_n548_, new_n549_ );
nand g445 ( new_n551_, new_n546_, new_n221_ );
nand g446 ( new_n552_, new_n551_, N53 );
nand g447 ( new_n553_, new_n546_, new_n209_, new_n221_ );
nand g448 ( N737, new_n552_, new_n553_ );
nand g449 ( new_n555_, new_n546_, new_n249_ );
nand g450 ( new_n556_, new_n555_, N57 );
nand g451 ( new_n557_, new_n546_, new_n229_, new_n249_ );
nand g452 ( N738, new_n556_, new_n557_ );
nand g453 ( new_n559_, new_n546_, new_n276_ );
nand g454 ( new_n560_, new_n559_, N61 );
nand g455 ( new_n561_, new_n546_, new_n264_, new_n276_ );
nand g456 ( N739, new_n560_, new_n561_ );
not g457 ( new_n563_, keyIn_0_20 );
nand g458 ( new_n564_, new_n345_, new_n346_, new_n398_ );
not g459 ( new_n565_, new_n564_ );
nand g460 ( new_n566_, new_n489_, new_n563_, new_n423_, new_n565_ );
nand g461 ( new_n567_, new_n565_, new_n455_, new_n423_, new_n452_ );
nand g462 ( new_n568_, new_n567_, keyIn_0_20 );
nand g463 ( new_n569_, new_n566_, new_n568_ );
nand g464 ( new_n570_, new_n456_, new_n424_, new_n565_ );
nand g465 ( new_n571_, new_n570_, keyIn_0_21 );
not g466 ( new_n572_, keyIn_0_21 );
nand g467 ( new_n573_, new_n456_, new_n572_, new_n424_, new_n565_ );
nand g468 ( new_n574_, new_n571_, new_n573_ );
nand g469 ( new_n575_, new_n422_, new_n398_, new_n419_ );
not g470 ( new_n576_, new_n575_ );
nand g471 ( new_n577_, new_n455_, new_n347_, new_n452_, new_n576_ );
nand g472 ( new_n578_, new_n577_, keyIn_0_22 );
not g473 ( new_n579_, keyIn_0_22 );
nor g474 ( new_n580_, new_n351_, new_n575_ );
nand g475 ( new_n581_, new_n580_, new_n579_, new_n452_, new_n455_ );
nand g476 ( new_n582_, new_n578_, new_n581_ );
nand g477 ( new_n583_, new_n456_, keyIn_0_18 );
not g478 ( new_n584_, keyIn_0_18 );
nand g479 ( new_n585_, new_n455_, new_n584_, new_n452_ );
nor g480 ( new_n586_, new_n492_, new_n423_ );
nand g481 ( new_n587_, new_n583_, new_n586_, new_n585_ );
nand g482 ( new_n588_, new_n582_, new_n587_ );
not g483 ( new_n589_, new_n588_ );
nand g484 ( new_n590_, new_n589_, keyIn_0_23, new_n569_, new_n574_ );
not g485 ( new_n591_, keyIn_0_23 );
nand g486 ( new_n592_, new_n574_, new_n569_, new_n582_, new_n587_ );
nand g487 ( new_n593_, new_n592_, new_n591_ );
nand g488 ( new_n594_, new_n593_, new_n590_ );
not g489 ( new_n595_, new_n594_ );
nand g490 ( new_n596_, new_n277_, new_n249_ );
nand g491 ( new_n597_, new_n251_, new_n160_ );
nor g492 ( new_n598_, new_n597_, new_n596_ );
nand g493 ( new_n599_, new_n595_, new_n397_, new_n598_ );
nand g494 ( new_n600_, new_n599_, N65 );
nand g495 ( new_n601_, new_n595_, new_n397_ );
not g496 ( new_n602_, new_n601_ );
nand g497 ( new_n603_, new_n602_, new_n108_, new_n598_ );
nand g498 ( N740, new_n603_, new_n600_ );
nand g499 ( new_n605_, new_n595_, new_n347_, new_n598_ );
nand g500 ( new_n606_, new_n605_, N69 );
nand g501 ( new_n607_, new_n595_, new_n347_ );
not g502 ( new_n608_, new_n607_ );
nand g503 ( new_n609_, new_n608_, new_n106_, new_n598_ );
nand g504 ( N741, new_n609_, new_n606_ );
nand g505 ( new_n611_, new_n595_, new_n456_, new_n598_ );
nand g506 ( new_n612_, new_n611_, N73 );
nand g507 ( new_n613_, new_n595_, new_n456_ );
not g508 ( new_n614_, new_n613_ );
nand g509 ( new_n615_, new_n614_, new_n112_, new_n598_ );
nand g510 ( N742, new_n615_, new_n612_ );
nand g511 ( new_n617_, new_n595_, new_n423_, new_n598_ );
nand g512 ( new_n618_, new_n617_, N77 );
nand g513 ( new_n619_, new_n595_, new_n423_ );
not g514 ( new_n620_, new_n619_ );
nand g515 ( new_n621_, new_n620_, new_n110_, new_n598_ );
nand g516 ( N743, new_n621_, new_n618_ );
not g517 ( new_n623_, new_n279_ );
nor g518 ( new_n624_, new_n623_, new_n597_ );
nand g519 ( new_n625_, new_n595_, new_n397_, new_n624_ );
nand g520 ( new_n626_, new_n625_, N81 );
nand g521 ( new_n627_, new_n602_, new_n125_, new_n624_ );
nand g522 ( N744, new_n627_, new_n626_ );
not g523 ( new_n629_, keyIn_0_27 );
nand g524 ( new_n630_, new_n593_, new_n590_, new_n347_, new_n624_ );
nand g525 ( new_n631_, new_n630_, new_n629_ );
nand g526 ( new_n632_, new_n595_, keyIn_0_27, new_n347_, new_n624_ );
nand g527 ( new_n633_, new_n632_, new_n631_ );
nand g528 ( new_n634_, new_n633_, new_n123_ );
nand g529 ( new_n635_, new_n632_, N85, new_n631_ );
nand g530 ( N745, new_n634_, new_n635_ );
nand g531 ( new_n637_, new_n595_, new_n456_, new_n624_ );
nand g532 ( new_n638_, new_n637_, N89 );
nand g533 ( new_n639_, new_n614_, new_n121_, new_n624_ );
nand g534 ( N746, new_n639_, new_n638_ );
nand g535 ( new_n641_, new_n595_, new_n423_, new_n624_ );
nand g536 ( new_n642_, new_n641_, N93 );
nand g537 ( new_n643_, new_n620_, new_n119_, new_n624_ );
nand g538 ( N747, new_n643_, new_n642_ );
nand g539 ( new_n645_, new_n221_, new_n162_ );
nor g540 ( new_n646_, new_n596_, new_n645_ );
nand g541 ( new_n647_, new_n595_, new_n397_, new_n646_ );
nand g542 ( new_n648_, new_n647_, N97 );
nand g543 ( new_n649_, new_n602_, new_n190_, new_n646_ );
nand g544 ( N748, new_n649_, new_n648_ );
nand g545 ( new_n651_, new_n595_, new_n347_, new_n646_ );
nand g546 ( new_n652_, new_n651_, N101 );
nand g547 ( new_n653_, new_n608_, new_n188_, new_n646_ );
nand g548 ( N749, new_n653_, new_n652_ );
nand g549 ( new_n655_, new_n595_, new_n456_, new_n646_ );
nand g550 ( new_n656_, new_n655_, N105 );
nand g551 ( new_n657_, new_n614_, new_n182_, new_n646_ );
nand g552 ( N750, new_n657_, new_n656_ );
nand g553 ( new_n659_, new_n593_, new_n590_, new_n423_, new_n646_ );
nand g554 ( new_n660_, new_n659_, keyIn_0_28 );
not g555 ( new_n661_, keyIn_0_28 );
nand g556 ( new_n662_, new_n595_, new_n661_, new_n423_, new_n646_ );
nand g557 ( new_n663_, new_n662_, new_n660_ );
nand g558 ( new_n664_, new_n663_, new_n180_ );
nand g559 ( new_n665_, new_n662_, N109, new_n660_ );
nand g560 ( N751, new_n664_, new_n665_ );
nor g561 ( new_n667_, new_n623_, new_n645_ );
nand g562 ( new_n668_, new_n595_, new_n397_, new_n667_ );
nand g563 ( new_n669_, new_n668_, N113 );
nand g564 ( new_n670_, new_n602_, new_n165_, new_n667_ );
nand g565 ( N752, new_n670_, new_n669_ );
nand g566 ( new_n672_, new_n593_, new_n590_, new_n347_, new_n667_ );
nand g567 ( new_n673_, new_n672_, keyIn_0_29 );
not g568 ( new_n674_, keyIn_0_29 );
nand g569 ( new_n675_, new_n595_, new_n674_, new_n347_, new_n667_ );
nand g570 ( new_n676_, new_n675_, new_n673_ );
nand g571 ( new_n677_, new_n676_, N117 );
nand g572 ( new_n678_, new_n675_, new_n163_, new_n673_ );
nand g573 ( N753, new_n677_, new_n678_ );
nand g574 ( new_n680_, new_n595_, new_n456_, new_n667_ );
nand g575 ( new_n681_, new_n680_, N121 );
nand g576 ( new_n682_, new_n614_, new_n174_, new_n667_ );
nand g577 ( N754, new_n682_, new_n681_ );
nand g578 ( new_n684_, new_n595_, new_n423_, new_n667_ );
nand g579 ( new_n685_, new_n684_, N125 );
nand g580 ( new_n686_, new_n620_, new_n172_, new_n667_ );
nand g581 ( N755, new_n686_, new_n685_ );
endmodule