module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n318_, new_n155_, new_n163_, new_n236_, new_n238_, new_n148_, new_n321_, new_n92_, new_n79_, new_n122_, new_n324_, new_n250_, new_n113_, new_n111_, new_n288_, new_n158_, new_n97_, new_n252_, new_n202_, new_n262_, new_n296_, new_n160_, new_n308_, new_n312_, new_n271_, new_n274_, new_n100_, new_n242_, new_n232_, new_n218_, new_n115_, new_n258_, new_n76_, new_n190_, new_n307_, new_n176_, new_n305_, new_n156_, new_n223_, new_n283_, new_n306_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n339_, new_n213_, new_n134_, new_n197_, new_n205_, new_n82_, new_n141_, new_n323_, new_n259_, new_n206_, new_n109_, new_n254_, new_n227_, new_n222_, new_n85_, new_n265_, new_n246_, new_n170_, new_n256_, new_n328_, new_n266_, new_n278_, new_n304_, new_n173_, new_n220_, new_n268_, new_n217_, new_n101_, new_n269_, new_n194_, new_n214_, new_n116_, new_n129_, new_n138_, new_n142_, new_n299_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n139_, new_n240_, new_n314_, new_n352_, new_n118_, new_n165_, new_n123_, new_n127_, new_n211_, new_n126_, new_n342_, new_n327_, new_n216_, new_n177_, new_n77_, new_n196_, new_n280_, new_n264_, new_n319_, new_n235_, new_n273_, new_n224_, new_n301_, new_n169_, new_n338_, new_n317_, new_n210_, new_n102_, new_n343_, new_n143_, new_n344_, new_n207_, new_n125_, new_n145_, new_n267_, new_n287_, new_n253_, new_n140_, new_n247_, new_n90_, new_n237_, new_n330_, new_n234_, new_n149_, new_n294_, new_n187_, new_n260_, new_n86_, new_n311_, new_n251_, new_n189_, new_n300_, new_n84_, new_n292_, new_n195_, new_n106_, new_n263_, new_n215_, new_n331_, new_n334_, new_n152_, new_n341_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n81_, new_n320_, new_n349_, new_n244_, new_n172_, new_n133_, new_n277_, new_n257_, new_n245_, new_n212_, new_n89_, new_n151_, new_n286_, new_n335_, new_n347_, new_n193_, new_n231_, new_n313_, new_n78_, new_n239_, new_n272_, new_n91_, new_n282_, new_n346_, new_n198_, new_n201_, new_n128_, new_n192_, new_n199_, new_n146_, new_n88_, new_n208_, new_n348_, new_n98_, new_n159_, new_n83_, new_n110_, new_n228_, new_n315_, new_n302_, new_n322_, new_n191_, new_n124_, new_n95_, new_n289_, new_n326_, new_n179_, new_n225_, new_n164_, new_n230_, new_n175_, new_n226_, new_n281_, new_n104_, new_n185_, new_n87_, new_n103_, new_n112_, new_n171_, new_n248_, new_n350_, new_n117_, new_n121_, new_n167_, new_n221_, new_n243_, new_n200_, new_n298_, new_n184_, new_n99_, new_n131_, new_n154_, new_n255_, new_n329_, new_n249_, new_n136_, new_n233_, new_n284_, new_n119_, new_n293_, new_n96_, new_n178_, new_n168_, new_n174_, new_n297_, new_n279_, new_n150_, new_n295_, new_n120_, new_n132_, new_n166_, new_n108_, new_n137_, new_n162_, new_n183_, new_n303_, new_n105_, new_n161_, new_n147_, new_n285_, new_n340_, new_n80_, new_n333_, new_n229_, new_n209_, new_n351_, new_n290_, new_n203_, new_n316_, new_n94_, new_n204_, new_n325_, new_n181_, new_n135_, new_n180_, new_n276_, new_n332_;

not g000 ( new_n76_, N17 );
xnor g001 ( new_n77_, keyIn_0_1, N11 );
or g002 ( new_n78_, new_n77_, new_n76_ );
xor g003 ( new_n79_, new_n78_, keyIn_0_10 );
not g004 ( new_n80_, N4 );
xnor g005 ( new_n81_, keyIn_0_0, N1 );
or g006 ( new_n82_, new_n81_, new_n80_ );
xnor g007 ( new_n83_, new_n82_, keyIn_0_9 );
or g008 ( new_n84_, keyIn_0_8, N102 );
and g009 ( new_n85_, keyIn_0_8, N102 );
not g010 ( new_n86_, new_n85_ );
and g011 ( new_n87_, new_n86_, N108 );
and g012 ( new_n88_, new_n87_, new_n84_ );
xnor g013 ( new_n89_, new_n88_, keyIn_0_17 );
and g014 ( new_n90_, new_n89_, new_n83_ );
and g015 ( new_n91_, new_n90_, new_n79_ );
xnor g016 ( new_n92_, keyIn_0_3, N37 );
and g017 ( new_n93_, new_n92_, N43 );
xnor g018 ( new_n94_, new_n93_, keyIn_0_12 );
not g019 ( new_n95_, keyIn_0_2 );
or g020 ( new_n96_, new_n95_, N24 );
not g021 ( new_n97_, N24 );
or g022 ( new_n98_, new_n97_, keyIn_0_2 );
and g023 ( new_n99_, new_n98_, N30 );
and g024 ( new_n100_, new_n99_, new_n96_ );
xnor g025 ( new_n101_, new_n100_, keyIn_0_11 );
and g026 ( new_n102_, new_n101_, new_n94_ );
xnor g027 ( new_n103_, keyIn_0_4, N50 );
and g028 ( new_n104_, new_n103_, N56 );
xnor g029 ( new_n105_, new_n104_, keyIn_0_13 );
not g030 ( new_n106_, keyIn_0_5 );
or g031 ( new_n107_, new_n106_, N63 );
not g032 ( new_n108_, N63 );
or g033 ( new_n109_, new_n108_, keyIn_0_5 );
and g034 ( new_n110_, new_n109_, N69 );
and g035 ( new_n111_, new_n110_, new_n107_ );
xnor g036 ( new_n112_, new_n111_, keyIn_0_14 );
and g037 ( new_n113_, new_n112_, new_n105_ );
xnor g038 ( new_n114_, keyIn_0_7, N89 );
and g039 ( new_n115_, new_n114_, N95 );
xor g040 ( new_n116_, new_n115_, keyIn_0_16 );
not g041 ( new_n117_, keyIn_0_6 );
not g042 ( new_n118_, N76 );
and g043 ( new_n119_, new_n117_, new_n118_ );
not g044 ( new_n120_, N82 );
and g045 ( new_n121_, keyIn_0_6, N76 );
or g046 ( new_n122_, new_n121_, new_n120_ );
or g047 ( new_n123_, new_n122_, new_n119_ );
xnor g048 ( new_n124_, new_n123_, keyIn_0_15 );
and g049 ( new_n125_, new_n124_, new_n116_ );
and g050 ( new_n126_, new_n113_, new_n125_ );
and g051 ( new_n127_, new_n126_, new_n102_ );
and g052 ( new_n128_, new_n127_, new_n91_ );
xnor g053 ( new_n129_, new_n128_, keyIn_0_18 );
not g054 ( N223, new_n129_ );
not g055 ( new_n131_, keyIn_0_26 );
not g056 ( new_n132_, keyIn_0_19 );
xnor g057 ( new_n133_, new_n129_, new_n132_ );
xor g058 ( new_n134_, new_n133_, new_n124_ );
not g059 ( new_n135_, new_n134_ );
and g060 ( new_n136_, new_n135_, new_n131_ );
or g061 ( new_n137_, new_n136_, new_n120_ );
and g062 ( new_n138_, new_n134_, keyIn_0_26 );
or g063 ( new_n139_, new_n138_, N86 );
or g064 ( new_n140_, new_n137_, new_n139_ );
not g065 ( new_n141_, N108 );
xor g066 ( new_n142_, new_n133_, new_n89_ );
not g067 ( new_n143_, new_n142_ );
and g068 ( new_n144_, new_n143_, keyIn_0_28 );
or g069 ( new_n145_, new_n144_, new_n141_ );
not g070 ( new_n146_, keyIn_0_28 );
and g071 ( new_n147_, new_n142_, new_n146_ );
or g072 ( new_n148_, new_n147_, N112 );
or g073 ( new_n149_, new_n145_, new_n148_ );
and g074 ( new_n150_, new_n140_, new_n149_ );
not g075 ( new_n151_, N43 );
xor g076 ( new_n152_, new_n133_, new_n94_ );
not g077 ( new_n153_, new_n152_ );
and g078 ( new_n154_, new_n153_, keyIn_0_23 );
or g079 ( new_n155_, new_n154_, new_n151_ );
not g080 ( new_n156_, keyIn_0_23 );
and g081 ( new_n157_, new_n152_, new_n156_ );
or g082 ( new_n158_, new_n157_, N47 );
or g083 ( new_n159_, new_n155_, new_n158_ );
not g084 ( new_n160_, N30 );
xor g085 ( new_n161_, new_n133_, new_n101_ );
not g086 ( new_n162_, new_n161_ );
and g087 ( new_n163_, new_n162_, keyIn_0_22 );
or g088 ( new_n164_, new_n163_, new_n160_ );
not g089 ( new_n165_, keyIn_0_22 );
and g090 ( new_n166_, new_n161_, new_n165_ );
or g091 ( new_n167_, new_n166_, N34 );
or g092 ( new_n168_, new_n164_, new_n167_ );
and g093 ( new_n169_, new_n159_, new_n168_ );
and g094 ( new_n170_, new_n150_, new_n169_ );
not g095 ( new_n171_, N95 );
xor g096 ( new_n172_, new_n133_, new_n116_ );
xnor g097 ( new_n173_, new_n172_, keyIn_0_27 );
or g098 ( new_n174_, new_n173_, new_n171_ );
or g099 ( new_n175_, new_n174_, N99 );
not g100 ( new_n176_, N56 );
xnor g101 ( new_n177_, new_n133_, new_n105_ );
and g102 ( new_n178_, new_n177_, keyIn_0_24 );
or g103 ( new_n179_, new_n178_, new_n176_ );
not g104 ( new_n180_, keyIn_0_24 );
not g105 ( new_n181_, new_n105_ );
xnor g106 ( new_n182_, new_n133_, new_n181_ );
and g107 ( new_n183_, new_n182_, new_n180_ );
or g108 ( new_n184_, new_n183_, N60 );
or g109 ( new_n185_, new_n179_, new_n184_ );
not g110 ( new_n186_, N69 );
not g111 ( new_n187_, keyIn_0_25 );
xnor g112 ( new_n188_, new_n133_, new_n112_ );
and g113 ( new_n189_, new_n188_, new_n187_ );
or g114 ( new_n190_, new_n189_, new_n186_ );
not g115 ( new_n191_, new_n112_ );
xnor g116 ( new_n192_, new_n133_, new_n191_ );
and g117 ( new_n193_, new_n192_, keyIn_0_25 );
or g118 ( new_n194_, new_n193_, N73 );
or g119 ( new_n195_, new_n190_, new_n194_ );
and g120 ( new_n196_, new_n185_, new_n195_ );
not g121 ( new_n197_, keyIn_0_20 );
xnor g122 ( new_n198_, new_n133_, new_n83_ );
and g123 ( new_n199_, new_n198_, new_n197_ );
or g124 ( new_n200_, new_n199_, new_n80_ );
not g125 ( new_n201_, new_n83_ );
xnor g126 ( new_n202_, new_n133_, new_n201_ );
and g127 ( new_n203_, new_n202_, keyIn_0_20 );
or g128 ( new_n204_, new_n203_, N8 );
or g129 ( new_n205_, new_n200_, new_n204_ );
xnor g130 ( new_n206_, new_n133_, new_n79_ );
and g131 ( new_n207_, new_n206_, keyIn_0_21 );
or g132 ( new_n208_, new_n207_, new_n76_ );
not g133 ( new_n209_, keyIn_0_21 );
not g134 ( new_n210_, new_n79_ );
xnor g135 ( new_n211_, new_n133_, new_n210_ );
and g136 ( new_n212_, new_n211_, new_n209_ );
or g137 ( new_n213_, new_n212_, N21 );
or g138 ( new_n214_, new_n208_, new_n213_ );
and g139 ( new_n215_, new_n205_, new_n214_ );
and g140 ( new_n216_, new_n196_, new_n215_ );
and g141 ( new_n217_, new_n216_, new_n175_ );
and g142 ( new_n218_, new_n217_, new_n170_ );
xnor g143 ( N329, new_n218_, keyIn_0_29 );
not g144 ( new_n220_, keyIn_0_30 );
xnor g145 ( new_n221_, N329, new_n159_ );
or g146 ( new_n222_, new_n157_, N53 );
or g147 ( new_n223_, new_n155_, new_n222_ );
or g148 ( new_n224_, new_n221_, new_n223_ );
xnor g149 ( new_n225_, N329, new_n168_ );
or g150 ( new_n226_, new_n166_, N40 );
or g151 ( new_n227_, new_n164_, new_n226_ );
or g152 ( new_n228_, new_n225_, new_n227_ );
not g153 ( new_n229_, new_n140_ );
or g154 ( new_n230_, N329, new_n229_ );
or g155 ( new_n231_, new_n140_, keyIn_0_29 );
and g156 ( new_n232_, new_n230_, new_n231_ );
or g157 ( new_n233_, new_n138_, N92 );
or g158 ( new_n234_, new_n137_, new_n233_ );
or g159 ( new_n235_, new_n232_, new_n234_ );
and g160 ( new_n236_, new_n235_, new_n228_ );
and g161 ( new_n237_, new_n236_, new_n224_ );
xnor g162 ( new_n238_, N329, new_n205_ );
or g163 ( new_n239_, new_n203_, N14 );
or g164 ( new_n240_, new_n200_, new_n239_ );
or g165 ( new_n241_, new_n238_, new_n240_ );
xnor g166 ( new_n242_, N329, new_n214_ );
or g167 ( new_n243_, new_n212_, N27 );
or g168 ( new_n244_, new_n208_, new_n243_ );
or g169 ( new_n245_, new_n242_, new_n244_ );
and g170 ( new_n246_, new_n241_, new_n245_ );
xnor g171 ( new_n247_, N329, new_n175_ );
or g172 ( new_n248_, new_n174_, N105 );
or g173 ( new_n249_, new_n247_, new_n248_ );
not g174 ( new_n250_, new_n149_ );
or g175 ( new_n251_, N329, new_n250_ );
or g176 ( new_n252_, new_n149_, keyIn_0_29 );
and g177 ( new_n253_, new_n251_, new_n252_ );
or g178 ( new_n254_, new_n147_, N115 );
or g179 ( new_n255_, new_n145_, new_n254_ );
or g180 ( new_n256_, new_n253_, new_n255_ );
and g181 ( new_n257_, new_n256_, new_n249_ );
xnor g182 ( new_n258_, N329, new_n185_ );
or g183 ( new_n259_, new_n183_, N66 );
or g184 ( new_n260_, new_n179_, new_n259_ );
or g185 ( new_n261_, new_n258_, new_n260_ );
xnor g186 ( new_n262_, N329, new_n195_ );
or g187 ( new_n263_, new_n193_, N79 );
or g188 ( new_n264_, new_n190_, new_n263_ );
or g189 ( new_n265_, new_n262_, new_n264_ );
and g190 ( new_n266_, new_n261_, new_n265_ );
and g191 ( new_n267_, new_n257_, new_n266_ );
and g192 ( new_n268_, new_n267_, new_n246_ );
and g193 ( new_n269_, new_n268_, new_n237_ );
xnor g194 ( N370, new_n269_, new_n220_ );
and g195 ( new_n271_, N370, N27 );
and g196 ( new_n272_, N329, N21 );
and g197 ( new_n273_, N223, N11 );
or g198 ( new_n274_, new_n273_, new_n76_ );
or g199 ( new_n275_, new_n272_, new_n274_ );
or g200 ( new_n276_, new_n271_, new_n275_ );
and g201 ( new_n277_, N370, N40 );
and g202 ( new_n278_, N329, N34 );
and g203 ( new_n279_, N223, N24 );
or g204 ( new_n280_, new_n279_, new_n160_ );
or g205 ( new_n281_, new_n278_, new_n280_ );
or g206 ( new_n282_, new_n277_, new_n281_ );
and g207 ( new_n283_, new_n276_, new_n282_ );
and g208 ( new_n284_, N370, N53 );
and g209 ( new_n285_, N329, N47 );
and g210 ( new_n286_, N223, N37 );
or g211 ( new_n287_, new_n286_, new_n151_ );
or g212 ( new_n288_, new_n285_, new_n287_ );
or g213 ( new_n289_, new_n284_, new_n288_ );
and g214 ( new_n290_, N370, N66 );
and g215 ( new_n291_, N329, N60 );
and g216 ( new_n292_, N223, N50 );
or g217 ( new_n293_, new_n292_, new_n176_ );
or g218 ( new_n294_, new_n291_, new_n293_ );
or g219 ( new_n295_, new_n290_, new_n294_ );
and g220 ( new_n296_, new_n289_, new_n295_ );
and g221 ( new_n297_, new_n283_, new_n296_ );
and g222 ( new_n298_, N370, N115 );
and g223 ( new_n299_, N329, N112 );
and g224 ( new_n300_, N223, N102 );
or g225 ( new_n301_, new_n300_, new_n141_ );
or g226 ( new_n302_, new_n299_, new_n301_ );
or g227 ( new_n303_, new_n298_, new_n302_ );
and g228 ( new_n304_, N370, N79 );
and g229 ( new_n305_, N329, N73 );
and g230 ( new_n306_, N223, N63 );
or g231 ( new_n307_, new_n306_, new_n186_ );
or g232 ( new_n308_, new_n305_, new_n307_ );
or g233 ( new_n309_, new_n304_, new_n308_ );
and g234 ( new_n310_, new_n303_, new_n309_ );
and g235 ( new_n311_, N370, N92 );
and g236 ( new_n312_, N329, N86 );
and g237 ( new_n313_, N223, N76 );
or g238 ( new_n314_, new_n313_, new_n120_ );
or g239 ( new_n315_, new_n312_, new_n314_ );
or g240 ( new_n316_, new_n311_, new_n315_ );
and g241 ( new_n317_, N370, N105 );
and g242 ( new_n318_, N329, N99 );
and g243 ( new_n319_, N223, N89 );
or g244 ( new_n320_, new_n319_, new_n171_ );
or g245 ( new_n321_, new_n318_, new_n320_ );
or g246 ( new_n322_, new_n317_, new_n321_ );
and g247 ( new_n323_, new_n316_, new_n322_ );
and g248 ( new_n324_, new_n310_, new_n323_ );
and g249 ( new_n325_, new_n297_, new_n324_ );
and g250 ( new_n326_, new_n325_, keyIn_0_31 );
not g251 ( new_n327_, new_n326_ );
or g252 ( new_n328_, new_n325_, keyIn_0_31 );
and g253 ( new_n329_, N370, N14 );
and g254 ( new_n330_, N329, N8 );
and g255 ( new_n331_, N223, N1 );
or g256 ( new_n332_, new_n331_, new_n80_ );
or g257 ( new_n333_, new_n330_, new_n332_ );
or g258 ( new_n334_, new_n329_, new_n333_ );
and g259 ( new_n335_, new_n328_, new_n334_ );
and g260 ( N421, new_n335_, new_n327_ );
not g261 ( N430, new_n297_ );
not g262 ( new_n338_, new_n309_ );
and g263 ( new_n339_, new_n338_, new_n295_ );
and g264 ( new_n340_, new_n339_, new_n289_ );
not g265 ( new_n341_, new_n283_ );
not g266 ( new_n342_, new_n316_ );
and g267 ( new_n343_, new_n296_, new_n342_ );
or g268 ( new_n344_, new_n343_, new_n341_ );
or g269 ( N431, new_n344_, new_n340_ );
not g270 ( new_n346_, new_n276_ );
not g271 ( new_n347_, new_n322_ );
and g272 ( new_n348_, new_n347_, new_n316_ );
not g273 ( new_n349_, new_n289_ );
or g274 ( new_n350_, new_n339_, new_n349_ );
or g275 ( new_n351_, new_n350_, new_n348_ );
and g276 ( new_n352_, new_n351_, new_n282_ );
or g277 ( N432, new_n352_, new_n346_ );
endmodule