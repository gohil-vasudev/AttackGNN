module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973;

  OR2_X1 U503 ( .A1(n487), .A2(n488), .ZN(Result_9_) );
  AND2_X1 U504 ( .A1(n489), .A2(n490), .ZN(n488) );
  XNOR2_X1 U505 ( .A(n491), .B(n492), .ZN(n489) );
  XOR2_X1 U506 ( .A(n493), .B(n494), .Z(n492) );
  AND2_X1 U507 ( .A1(n495), .A2(n496), .ZN(n487) );
  XOR2_X1 U508 ( .A(n497), .B(n498), .Z(n495) );
  AND2_X1 U509 ( .A1(n499), .A2(n500), .ZN(n498) );
  OR2_X1 U510 ( .A1(n501), .A2(n502), .ZN(Result_8_) );
  AND2_X1 U511 ( .A1(n503), .A2(n490), .ZN(n502) );
  XNOR2_X1 U512 ( .A(n504), .B(n505), .ZN(n503) );
  XOR2_X1 U513 ( .A(n506), .B(n507), .Z(n505) );
  AND2_X1 U514 ( .A1(n508), .A2(n496), .ZN(n501) );
  XOR2_X1 U515 ( .A(n509), .B(n510), .Z(n508) );
  OR2_X1 U516 ( .A1(a_0_), .A2(n511), .ZN(n510) );
  OR2_X1 U517 ( .A1(n512), .A2(n513), .ZN(n509) );
  AND2_X1 U518 ( .A1(n514), .A2(n515), .ZN(n513) );
  AND2_X1 U519 ( .A1(n497), .A2(n516), .ZN(n512) );
  OR2_X1 U520 ( .A1(n517), .A2(n518), .ZN(n497) );
  INV_X1 U521 ( .A(n519), .ZN(n518) );
  AND2_X1 U522 ( .A1(n520), .A2(n521), .ZN(n517) );
  AND2_X1 U523 ( .A1(n490), .A2(n522), .ZN(Result_7_) );
  XOR2_X1 U524 ( .A(n523), .B(n524), .Z(n522) );
  AND3_X1 U525 ( .A1(n525), .A2(n526), .A3(n490), .ZN(Result_6_) );
  OR2_X1 U526 ( .A1(n527), .A2(n528), .ZN(n525) );
  XOR2_X1 U527 ( .A(n529), .B(n530), .Z(n528) );
  INV_X1 U528 ( .A(n531), .ZN(n527) );
  OR2_X1 U529 ( .A1(n523), .A2(n524), .ZN(n531) );
  AND2_X1 U530 ( .A1(n490), .A2(n532), .ZN(Result_5_) );
  XNOR2_X1 U531 ( .A(n533), .B(n534), .ZN(n532) );
  OR2_X1 U532 ( .A1(n535), .A2(n536), .ZN(n533) );
  AND2_X1 U533 ( .A1(n537), .A2(n490), .ZN(Result_4_) );
  XOR2_X1 U534 ( .A(n538), .B(n539), .Z(n537) );
  AND2_X1 U535 ( .A1(n490), .A2(n540), .ZN(Result_3_) );
  XOR2_X1 U536 ( .A(n541), .B(n542), .Z(n540) );
  AND2_X1 U537 ( .A1(n543), .A2(n544), .ZN(n542) );
  OR2_X1 U538 ( .A1(n545), .A2(n546), .ZN(n544) );
  AND2_X1 U539 ( .A1(n547), .A2(n548), .ZN(n546) );
  INV_X1 U540 ( .A(n549), .ZN(n543) );
  AND2_X1 U541 ( .A1(n550), .A2(n490), .ZN(Result_2_) );
  XOR2_X1 U542 ( .A(n551), .B(n552), .Z(n550) );
  AND2_X1 U543 ( .A1(n490), .A2(n553), .ZN(Result_1_) );
  XOR2_X1 U544 ( .A(n554), .B(n555), .Z(n553) );
  AND2_X1 U545 ( .A1(n556), .A2(n557), .ZN(n555) );
  OR2_X1 U546 ( .A1(n558), .A2(n559), .ZN(n557) );
  AND2_X1 U547 ( .A1(n560), .A2(n561), .ZN(n559) );
  INV_X1 U548 ( .A(n562), .ZN(n556) );
  OR2_X1 U549 ( .A1(n563), .A2(n564), .ZN(Result_15_) );
  AND2_X1 U550 ( .A1(n490), .A2(n565), .ZN(n564) );
  AND2_X1 U551 ( .A1(n566), .A2(n496), .ZN(n563) );
  XOR2_X1 U552 ( .A(b_7_), .B(a_7_), .Z(n566) );
  OR2_X1 U553 ( .A1(n567), .A2(n568), .ZN(Result_14_) );
  AND2_X1 U554 ( .A1(n569), .A2(n496), .ZN(n568) );
  XOR2_X1 U555 ( .A(n570), .B(n565), .Z(n569) );
  OR2_X1 U556 ( .A1(n571), .A2(n572), .ZN(n570) );
  AND2_X1 U557 ( .A1(n490), .A2(n573), .ZN(n567) );
  OR2_X1 U558 ( .A1(n574), .A2(n575), .ZN(n573) );
  AND2_X1 U559 ( .A1(a_7_), .A2(n576), .ZN(n575) );
  OR2_X1 U560 ( .A1(n577), .A2(n572), .ZN(n576) );
  INV_X1 U561 ( .A(n578), .ZN(n572) );
  AND2_X1 U562 ( .A1(b_6_), .A2(n579), .ZN(n577) );
  AND3_X1 U563 ( .A1(a_6_), .A2(n580), .A3(b_7_), .ZN(n574) );
  OR2_X1 U564 ( .A1(n581), .A2(n582), .ZN(Result_13_) );
  AND2_X1 U565 ( .A1(n583), .A2(n490), .ZN(n582) );
  XNOR2_X1 U566 ( .A(n584), .B(n585), .ZN(n583) );
  XOR2_X1 U567 ( .A(n586), .B(n587), .Z(n585) );
  AND2_X1 U568 ( .A1(n588), .A2(n496), .ZN(n581) );
  XOR2_X1 U569 ( .A(n589), .B(n590), .Z(n588) );
  OR2_X1 U570 ( .A1(n591), .A2(n592), .ZN(n590) );
  INV_X1 U571 ( .A(n593), .ZN(n592) );
  OR2_X1 U572 ( .A1(n594), .A2(n595), .ZN(Result_12_) );
  AND2_X1 U573 ( .A1(n596), .A2(n490), .ZN(n595) );
  XNOR2_X1 U574 ( .A(n597), .B(n598), .ZN(n596) );
  XOR2_X1 U575 ( .A(n599), .B(n600), .Z(n598) );
  AND2_X1 U576 ( .A1(n601), .A2(n496), .ZN(n594) );
  XOR2_X1 U577 ( .A(n602), .B(n603), .Z(n601) );
  AND2_X1 U578 ( .A1(n604), .A2(n605), .ZN(n603) );
  OR2_X1 U579 ( .A1(n606), .A2(n607), .ZN(Result_11_) );
  AND2_X1 U580 ( .A1(n608), .A2(n490), .ZN(n607) );
  XNOR2_X1 U581 ( .A(n609), .B(n610), .ZN(n608) );
  XOR2_X1 U582 ( .A(n611), .B(n612), .Z(n610) );
  AND2_X1 U583 ( .A1(n613), .A2(n496), .ZN(n606) );
  XNOR2_X1 U584 ( .A(n614), .B(n615), .ZN(n613) );
  OR2_X1 U585 ( .A1(n616), .A2(n617), .ZN(n614) );
  INV_X1 U586 ( .A(n618), .ZN(n617) );
  OR2_X1 U587 ( .A1(n619), .A2(n620), .ZN(Result_10_) );
  AND2_X1 U588 ( .A1(n621), .A2(n490), .ZN(n620) );
  XNOR2_X1 U589 ( .A(n622), .B(n623), .ZN(n621) );
  XOR2_X1 U590 ( .A(n624), .B(n625), .Z(n623) );
  AND2_X1 U591 ( .A1(n626), .A2(n496), .ZN(n619) );
  XNOR2_X1 U592 ( .A(n520), .B(n627), .ZN(n626) );
  AND2_X1 U593 ( .A1(n521), .A2(n519), .ZN(n627) );
  OR2_X1 U594 ( .A1(a_2_), .A2(b_2_), .ZN(n519) );
  OR2_X1 U595 ( .A1(n628), .A2(n629), .ZN(n520) );
  AND2_X1 U596 ( .A1(n630), .A2(n631), .ZN(n629) );
  AND2_X1 U597 ( .A1(n615), .A2(n632), .ZN(n628) );
  OR2_X1 U598 ( .A1(n633), .A2(n634), .ZN(n615) );
  INV_X1 U599 ( .A(n605), .ZN(n634) );
  OR2_X1 U600 ( .A1(a_4_), .A2(b_4_), .ZN(n605) );
  AND2_X1 U601 ( .A1(n635), .A2(n604), .ZN(n633) );
  INV_X1 U602 ( .A(n602), .ZN(n635) );
  AND2_X1 U603 ( .A1(n636), .A2(n637), .ZN(n602) );
  OR2_X1 U604 ( .A1(a_5_), .A2(b_5_), .ZN(n637) );
  OR2_X1 U605 ( .A1(n589), .A2(n638), .ZN(n636) );
  OR2_X1 U606 ( .A1(n639), .A2(n640), .ZN(n589) );
  AND2_X1 U607 ( .A1(n565), .A2(n641), .ZN(n639) );
  OR2_X1 U608 ( .A1(a_6_), .A2(b_6_), .ZN(n641) );
  AND2_X1 U609 ( .A1(n490), .A2(n642), .ZN(Result_0_) );
  OR3_X1 U610 ( .A1(n562), .A2(n643), .A3(n644), .ZN(n642) );
  AND2_X1 U611 ( .A1(n554), .A2(n558), .ZN(n644) );
  AND2_X1 U612 ( .A1(n551), .A2(n552), .ZN(n554) );
  XOR2_X1 U613 ( .A(n561), .B(n560), .Z(n552) );
  OR2_X1 U614 ( .A1(n645), .A2(n646), .ZN(n551) );
  INV_X1 U615 ( .A(n647), .ZN(n646) );
  OR2_X1 U616 ( .A1(n648), .A2(n549), .ZN(n645) );
  AND3_X1 U617 ( .A1(n548), .A2(n547), .A3(n545), .ZN(n549) );
  AND2_X1 U618 ( .A1(n541), .A2(n545), .ZN(n648) );
  AND2_X1 U619 ( .A1(n649), .A2(n647), .ZN(n545) );
  OR2_X1 U620 ( .A1(n650), .A2(n651), .ZN(n647) );
  INV_X1 U621 ( .A(n652), .ZN(n649) );
  AND2_X1 U622 ( .A1(n650), .A2(n651), .ZN(n652) );
  OR2_X1 U623 ( .A1(n653), .A2(n654), .ZN(n651) );
  AND2_X1 U624 ( .A1(n655), .A2(n656), .ZN(n654) );
  AND2_X1 U625 ( .A1(n657), .A2(n658), .ZN(n653) );
  OR2_X1 U626 ( .A1(n656), .A2(n655), .ZN(n658) );
  XNOR2_X1 U627 ( .A(n659), .B(n660), .ZN(n650) );
  XNOR2_X1 U628 ( .A(n661), .B(n662), .ZN(n660) );
  AND2_X1 U629 ( .A1(n538), .A2(n539), .ZN(n541) );
  XOR2_X1 U630 ( .A(n548), .B(n547), .Z(n539) );
  INV_X1 U631 ( .A(n663), .ZN(n547) );
  OR2_X1 U632 ( .A1(n664), .A2(n665), .ZN(n663) );
  AND2_X1 U633 ( .A1(n666), .A2(n667), .ZN(n665) );
  AND2_X1 U634 ( .A1(n668), .A2(n669), .ZN(n664) );
  OR2_X1 U635 ( .A1(n667), .A2(n666), .ZN(n669) );
  XOR2_X1 U636 ( .A(n670), .B(n657), .Z(n548) );
  XOR2_X1 U637 ( .A(n671), .B(n672), .Z(n657) );
  XOR2_X1 U638 ( .A(n673), .B(n674), .Z(n672) );
  XNOR2_X1 U639 ( .A(n656), .B(n655), .ZN(n670) );
  OR2_X1 U640 ( .A1(n675), .A2(n676), .ZN(n655) );
  AND2_X1 U641 ( .A1(n677), .A2(n678), .ZN(n676) );
  AND2_X1 U642 ( .A1(n679), .A2(n680), .ZN(n675) );
  OR2_X1 U643 ( .A1(n678), .A2(n677), .ZN(n680) );
  OR2_X1 U644 ( .A1(n631), .A2(n681), .ZN(n656) );
  OR2_X1 U645 ( .A1(n682), .A2(n683), .ZN(n538) );
  OR2_X1 U646 ( .A1(n684), .A2(n685), .ZN(n682) );
  AND2_X1 U647 ( .A1(n535), .A2(n686), .ZN(n685) );
  AND2_X1 U648 ( .A1(n536), .A2(n686), .ZN(n684) );
  INV_X1 U649 ( .A(n534), .ZN(n686) );
  OR2_X1 U650 ( .A1(n687), .A2(n683), .ZN(n534) );
  INV_X1 U651 ( .A(n688), .ZN(n683) );
  OR2_X1 U652 ( .A1(n689), .A2(n690), .ZN(n688) );
  AND2_X1 U653 ( .A1(n689), .A2(n690), .ZN(n687) );
  OR2_X1 U654 ( .A1(n691), .A2(n692), .ZN(n690) );
  AND2_X1 U655 ( .A1(n693), .A2(n694), .ZN(n692) );
  AND2_X1 U656 ( .A1(n695), .A2(n696), .ZN(n691) );
  OR2_X1 U657 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U658 ( .A(n668), .B(n697), .Z(n689) );
  XOR2_X1 U659 ( .A(n667), .B(n666), .Z(n697) );
  OR2_X1 U660 ( .A1(n698), .A2(n681), .ZN(n666) );
  OR2_X1 U661 ( .A1(n699), .A2(n700), .ZN(n667) );
  AND2_X1 U662 ( .A1(n701), .A2(n702), .ZN(n700) );
  AND2_X1 U663 ( .A1(n703), .A2(n704), .ZN(n699) );
  OR2_X1 U664 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U665 ( .A(n705), .B(n679), .ZN(n668) );
  XNOR2_X1 U666 ( .A(n706), .B(n707), .ZN(n679) );
  XNOR2_X1 U667 ( .A(n521), .B(n708), .ZN(n706) );
  XNOR2_X1 U668 ( .A(n678), .B(n677), .ZN(n705) );
  OR2_X1 U669 ( .A1(n709), .A2(n710), .ZN(n677) );
  AND2_X1 U670 ( .A1(n711), .A2(n712), .ZN(n710) );
  AND2_X1 U671 ( .A1(n713), .A2(n714), .ZN(n709) );
  OR2_X1 U672 ( .A1(n712), .A2(n711), .ZN(n714) );
  OR2_X1 U673 ( .A1(n631), .A2(n514), .ZN(n678) );
  INV_X1 U674 ( .A(n526), .ZN(n536) );
  OR4_X1 U675 ( .A1(n524), .A2(n523), .A3(n535), .A4(n715), .ZN(n526) );
  AND2_X1 U676 ( .A1(n529), .A2(n530), .ZN(n715) );
  INV_X1 U677 ( .A(n716), .ZN(n535) );
  OR2_X1 U678 ( .A1(n529), .A2(n530), .ZN(n716) );
  OR2_X1 U679 ( .A1(n717), .A2(n718), .ZN(n530) );
  AND2_X1 U680 ( .A1(n719), .A2(n720), .ZN(n718) );
  AND2_X1 U681 ( .A1(n721), .A2(n722), .ZN(n717) );
  OR2_X1 U682 ( .A1(n720), .A2(n719), .ZN(n722) );
  XOR2_X1 U683 ( .A(n693), .B(n723), .Z(n529) );
  XOR2_X1 U684 ( .A(n696), .B(n694), .Z(n723) );
  OR2_X1 U685 ( .A1(n724), .A2(n681), .ZN(n694) );
  OR2_X1 U686 ( .A1(n725), .A2(n726), .ZN(n696) );
  AND2_X1 U687 ( .A1(n727), .A2(n728), .ZN(n726) );
  AND2_X1 U688 ( .A1(n729), .A2(n730), .ZN(n725) );
  OR2_X1 U689 ( .A1(n728), .A2(n727), .ZN(n730) );
  XOR2_X1 U690 ( .A(n701), .B(n731), .Z(n693) );
  XOR2_X1 U691 ( .A(n704), .B(n702), .Z(n731) );
  OR2_X1 U692 ( .A1(n698), .A2(n514), .ZN(n702) );
  OR2_X1 U693 ( .A1(n732), .A2(n733), .ZN(n704) );
  AND2_X1 U694 ( .A1(n734), .A2(n735), .ZN(n733) );
  AND2_X1 U695 ( .A1(n736), .A2(n737), .ZN(n732) );
  OR2_X1 U696 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U697 ( .A(n738), .B(n713), .ZN(n701) );
  XNOR2_X1 U698 ( .A(n739), .B(n740), .ZN(n713) );
  XNOR2_X1 U699 ( .A(n741), .B(n742), .ZN(n739) );
  XNOR2_X1 U700 ( .A(n712), .B(n711), .ZN(n738) );
  OR2_X1 U701 ( .A1(n743), .A2(n744), .ZN(n711) );
  AND2_X1 U702 ( .A1(n745), .A2(n632), .ZN(n744) );
  AND2_X1 U703 ( .A1(n746), .A2(n747), .ZN(n743) );
  OR2_X1 U704 ( .A1(n632), .A2(n745), .ZN(n747) );
  OR2_X1 U705 ( .A1(n631), .A2(n748), .ZN(n712) );
  OR2_X1 U706 ( .A1(n749), .A2(n750), .ZN(n523) );
  AND2_X1 U707 ( .A1(n507), .A2(n506), .ZN(n750) );
  AND2_X1 U708 ( .A1(n504), .A2(n751), .ZN(n749) );
  OR2_X1 U709 ( .A1(n506), .A2(n507), .ZN(n751) );
  OR2_X1 U710 ( .A1(n681), .A2(n579), .ZN(n507) );
  OR2_X1 U711 ( .A1(n752), .A2(n753), .ZN(n506) );
  AND2_X1 U712 ( .A1(n494), .A2(n493), .ZN(n753) );
  AND2_X1 U713 ( .A1(n491), .A2(n754), .ZN(n752) );
  OR2_X1 U714 ( .A1(n493), .A2(n494), .ZN(n754) );
  OR2_X1 U715 ( .A1(n514), .A2(n579), .ZN(n494) );
  OR2_X1 U716 ( .A1(n755), .A2(n756), .ZN(n493) );
  AND2_X1 U717 ( .A1(n625), .A2(n624), .ZN(n756) );
  AND2_X1 U718 ( .A1(n622), .A2(n757), .ZN(n755) );
  OR2_X1 U719 ( .A1(n625), .A2(n624), .ZN(n757) );
  OR2_X1 U720 ( .A1(n758), .A2(n759), .ZN(n624) );
  AND2_X1 U721 ( .A1(n612), .A2(n611), .ZN(n759) );
  AND2_X1 U722 ( .A1(n609), .A2(n760), .ZN(n758) );
  OR2_X1 U723 ( .A1(n612), .A2(n611), .ZN(n760) );
  OR2_X1 U724 ( .A1(n761), .A2(n762), .ZN(n611) );
  AND2_X1 U725 ( .A1(n600), .A2(n599), .ZN(n762) );
  AND2_X1 U726 ( .A1(n597), .A2(n763), .ZN(n761) );
  OR2_X1 U727 ( .A1(n600), .A2(n599), .ZN(n763) );
  OR2_X1 U728 ( .A1(n764), .A2(n765), .ZN(n599) );
  AND2_X1 U729 ( .A1(n587), .A2(n586), .ZN(n765) );
  AND2_X1 U730 ( .A1(n584), .A2(n766), .ZN(n764) );
  OR2_X1 U731 ( .A1(n587), .A2(n586), .ZN(n766) );
  INV_X1 U732 ( .A(n767), .ZN(n586) );
  AND2_X1 U733 ( .A1(n640), .A2(n565), .ZN(n767) );
  AND2_X1 U734 ( .A1(a_7_), .A2(b_7_), .ZN(n565) );
  OR2_X1 U735 ( .A1(n768), .A2(n579), .ZN(n587) );
  XOR2_X1 U736 ( .A(n769), .B(n640), .Z(n584) );
  AND2_X1 U737 ( .A1(b_6_), .A2(a_6_), .ZN(n640) );
  OR2_X1 U738 ( .A1(n770), .A2(n579), .ZN(n600) );
  XNOR2_X1 U739 ( .A(n771), .B(n772), .ZN(n597) );
  XNOR2_X1 U740 ( .A(n773), .B(n774), .ZN(n771) );
  OR2_X1 U741 ( .A1(n630), .A2(n579), .ZN(n612) );
  XOR2_X1 U742 ( .A(n775), .B(n776), .Z(n609) );
  XOR2_X1 U743 ( .A(n777), .B(n778), .Z(n776) );
  OR2_X1 U744 ( .A1(n748), .A2(n579), .ZN(n625) );
  XOR2_X1 U745 ( .A(n779), .B(n780), .Z(n622) );
  XOR2_X1 U746 ( .A(n781), .B(n782), .Z(n780) );
  XOR2_X1 U747 ( .A(n783), .B(n784), .Z(n491) );
  XOR2_X1 U748 ( .A(n785), .B(n786), .Z(n784) );
  XOR2_X1 U749 ( .A(n787), .B(n788), .Z(n504) );
  XOR2_X1 U750 ( .A(n789), .B(n790), .Z(n788) );
  XOR2_X1 U751 ( .A(n721), .B(n791), .Z(n524) );
  XOR2_X1 U752 ( .A(n720), .B(n719), .Z(n791) );
  OR2_X1 U753 ( .A1(n792), .A2(n681), .ZN(n719) );
  OR2_X1 U754 ( .A1(n793), .A2(n794), .ZN(n720) );
  AND2_X1 U755 ( .A1(n790), .A2(n789), .ZN(n794) );
  AND2_X1 U756 ( .A1(n787), .A2(n795), .ZN(n793) );
  OR2_X1 U757 ( .A1(n789), .A2(n790), .ZN(n795) );
  OR2_X1 U758 ( .A1(n792), .A2(n514), .ZN(n790) );
  OR2_X1 U759 ( .A1(n796), .A2(n797), .ZN(n789) );
  AND2_X1 U760 ( .A1(n786), .A2(n785), .ZN(n797) );
  AND2_X1 U761 ( .A1(n783), .A2(n798), .ZN(n796) );
  OR2_X1 U762 ( .A1(n785), .A2(n786), .ZN(n798) );
  OR2_X1 U763 ( .A1(n792), .A2(n748), .ZN(n786) );
  OR2_X1 U764 ( .A1(n799), .A2(n800), .ZN(n785) );
  AND2_X1 U765 ( .A1(n782), .A2(n781), .ZN(n800) );
  AND2_X1 U766 ( .A1(n779), .A2(n801), .ZN(n799) );
  OR2_X1 U767 ( .A1(n782), .A2(n781), .ZN(n801) );
  OR2_X1 U768 ( .A1(n802), .A2(n803), .ZN(n781) );
  AND2_X1 U769 ( .A1(n778), .A2(n777), .ZN(n803) );
  AND2_X1 U770 ( .A1(n775), .A2(n804), .ZN(n802) );
  OR2_X1 U771 ( .A1(n778), .A2(n777), .ZN(n804) );
  OR2_X1 U772 ( .A1(n805), .A2(n806), .ZN(n777) );
  AND2_X1 U773 ( .A1(n773), .A2(n774), .ZN(n806) );
  AND2_X1 U774 ( .A1(n772), .A2(n807), .ZN(n805) );
  OR2_X1 U775 ( .A1(n773), .A2(n774), .ZN(n807) );
  OR2_X1 U776 ( .A1(n580), .A2(n808), .ZN(n774) );
  OR2_X1 U777 ( .A1(n792), .A2(n809), .ZN(n580) );
  OR2_X1 U778 ( .A1(n768), .A2(n792), .ZN(n773) );
  XNOR2_X1 U779 ( .A(n810), .B(n808), .ZN(n772) );
  OR2_X1 U780 ( .A1(n724), .A2(n811), .ZN(n808) );
  OR2_X1 U781 ( .A1(n698), .A2(n809), .ZN(n810) );
  OR2_X1 U782 ( .A1(n792), .A2(n770), .ZN(n778) );
  XNOR2_X1 U783 ( .A(n812), .B(n813), .ZN(n775) );
  XOR2_X1 U784 ( .A(n814), .B(n638), .Z(n812) );
  INV_X1 U785 ( .A(n815), .ZN(n638) );
  OR2_X1 U786 ( .A1(n630), .A2(n792), .ZN(n782) );
  XOR2_X1 U787 ( .A(n816), .B(n817), .Z(n779) );
  XOR2_X1 U788 ( .A(n818), .B(n819), .Z(n817) );
  XOR2_X1 U789 ( .A(n820), .B(n821), .Z(n783) );
  XOR2_X1 U790 ( .A(n822), .B(n823), .Z(n821) );
  XOR2_X1 U791 ( .A(n824), .B(n825), .Z(n787) );
  XOR2_X1 U792 ( .A(n826), .B(n827), .Z(n825) );
  XOR2_X1 U793 ( .A(n729), .B(n828), .Z(n721) );
  XOR2_X1 U794 ( .A(n728), .B(n727), .Z(n828) );
  OR2_X1 U795 ( .A1(n724), .A2(n514), .ZN(n727) );
  OR2_X1 U796 ( .A1(n829), .A2(n830), .ZN(n728) );
  AND2_X1 U797 ( .A1(n827), .A2(n826), .ZN(n830) );
  AND2_X1 U798 ( .A1(n824), .A2(n831), .ZN(n829) );
  OR2_X1 U799 ( .A1(n826), .A2(n827), .ZN(n831) );
  OR2_X1 U800 ( .A1(n724), .A2(n748), .ZN(n827) );
  OR2_X1 U801 ( .A1(n832), .A2(n833), .ZN(n826) );
  AND2_X1 U802 ( .A1(n823), .A2(n822), .ZN(n833) );
  AND2_X1 U803 ( .A1(n820), .A2(n834), .ZN(n832) );
  OR2_X1 U804 ( .A1(n822), .A2(n823), .ZN(n834) );
  OR2_X1 U805 ( .A1(n630), .A2(n724), .ZN(n823) );
  OR2_X1 U806 ( .A1(n835), .A2(n836), .ZN(n822) );
  AND2_X1 U807 ( .A1(n819), .A2(n818), .ZN(n836) );
  AND2_X1 U808 ( .A1(n816), .A2(n837), .ZN(n835) );
  OR2_X1 U809 ( .A1(n819), .A2(n818), .ZN(n837) );
  OR2_X1 U810 ( .A1(n838), .A2(n839), .ZN(n818) );
  AND2_X1 U811 ( .A1(n813), .A2(n815), .ZN(n839) );
  AND2_X1 U812 ( .A1(n840), .A2(n814), .ZN(n838) );
  OR2_X1 U813 ( .A1(n841), .A2(n842), .ZN(n814) );
  AND2_X1 U814 ( .A1(n843), .A2(n844), .ZN(n841) );
  OR2_X1 U815 ( .A1(n813), .A2(n815), .ZN(n840) );
  OR2_X1 U816 ( .A1(n768), .A2(n724), .ZN(n815) );
  OR2_X1 U817 ( .A1(n843), .A2(n769), .ZN(n813) );
  OR2_X1 U818 ( .A1(n724), .A2(n809), .ZN(n769) );
  OR2_X1 U819 ( .A1(n724), .A2(n770), .ZN(n819) );
  XNOR2_X1 U820 ( .A(n845), .B(n846), .ZN(n816) );
  XOR2_X1 U821 ( .A(n847), .B(n842), .Z(n845) );
  INV_X1 U822 ( .A(n848), .ZN(n842) );
  XNOR2_X1 U823 ( .A(n849), .B(n850), .ZN(n820) );
  XNOR2_X1 U824 ( .A(n604), .B(n851), .ZN(n849) );
  XOR2_X1 U825 ( .A(n852), .B(n853), .Z(n824) );
  XOR2_X1 U826 ( .A(n854), .B(n855), .Z(n853) );
  XOR2_X1 U827 ( .A(n736), .B(n856), .Z(n729) );
  XOR2_X1 U828 ( .A(n735), .B(n734), .Z(n856) );
  OR2_X1 U829 ( .A1(n698), .A2(n748), .ZN(n734) );
  OR2_X1 U830 ( .A1(n857), .A2(n858), .ZN(n735) );
  AND2_X1 U831 ( .A1(n855), .A2(n854), .ZN(n858) );
  AND2_X1 U832 ( .A1(n852), .A2(n859), .ZN(n857) );
  OR2_X1 U833 ( .A1(n854), .A2(n855), .ZN(n859) );
  OR2_X1 U834 ( .A1(n630), .A2(n698), .ZN(n855) );
  OR2_X1 U835 ( .A1(n860), .A2(n861), .ZN(n854) );
  AND2_X1 U836 ( .A1(n851), .A2(n604), .ZN(n861) );
  AND2_X1 U837 ( .A1(n850), .A2(n862), .ZN(n860) );
  OR2_X1 U838 ( .A1(n604), .A2(n851), .ZN(n862) );
  OR2_X1 U839 ( .A1(n863), .A2(n864), .ZN(n851) );
  AND2_X1 U840 ( .A1(n846), .A2(n848), .ZN(n864) );
  AND2_X1 U841 ( .A1(n865), .A2(n847), .ZN(n863) );
  OR2_X1 U842 ( .A1(n866), .A2(n867), .ZN(n847) );
  INV_X1 U843 ( .A(n868), .ZN(n867) );
  AND2_X1 U844 ( .A1(n869), .A2(n870), .ZN(n866) );
  OR2_X1 U845 ( .A1(n809), .A2(n871), .ZN(n870) );
  OR2_X1 U846 ( .A1(n631), .A2(n811), .ZN(n869) );
  OR2_X1 U847 ( .A1(n846), .A2(n848), .ZN(n865) );
  OR2_X1 U848 ( .A1(n844), .A2(n843), .ZN(n848) );
  OR2_X1 U849 ( .A1(n698), .A2(n811), .ZN(n843) );
  OR2_X1 U850 ( .A1(n698), .A2(n768), .ZN(n846) );
  OR2_X1 U851 ( .A1(n698), .A2(n770), .ZN(n604) );
  XNOR2_X1 U852 ( .A(n872), .B(n868), .ZN(n850) );
  XNOR2_X1 U853 ( .A(n873), .B(n874), .ZN(n872) );
  XNOR2_X1 U854 ( .A(n875), .B(n876), .ZN(n852) );
  XNOR2_X1 U855 ( .A(n877), .B(n878), .ZN(n875) );
  XNOR2_X1 U856 ( .A(n879), .B(n746), .ZN(n736) );
  XNOR2_X1 U857 ( .A(n880), .B(n881), .ZN(n746) );
  XNOR2_X1 U858 ( .A(n882), .B(n883), .ZN(n880) );
  XNOR2_X1 U859 ( .A(n632), .B(n745), .ZN(n879) );
  OR2_X1 U860 ( .A1(n884), .A2(n885), .ZN(n745) );
  AND2_X1 U861 ( .A1(n878), .A2(n877), .ZN(n885) );
  AND2_X1 U862 ( .A1(n876), .A2(n886), .ZN(n884) );
  OR2_X1 U863 ( .A1(n877), .A2(n878), .ZN(n886) );
  OR2_X1 U864 ( .A1(n887), .A2(n888), .ZN(n878) );
  AND2_X1 U865 ( .A1(n868), .A2(n874), .ZN(n888) );
  AND2_X1 U866 ( .A1(n889), .A2(n873), .ZN(n887) );
  OR2_X1 U867 ( .A1(n890), .A2(n891), .ZN(n873) );
  AND2_X1 U868 ( .A1(n892), .A2(n893), .ZN(n890) );
  OR2_X1 U869 ( .A1(n874), .A2(n868), .ZN(n889) );
  OR2_X1 U870 ( .A1(n844), .A2(n893), .ZN(n868) );
  OR2_X1 U871 ( .A1(n631), .A2(n809), .ZN(n844) );
  OR2_X1 U872 ( .A1(n631), .A2(n768), .ZN(n874) );
  OR2_X1 U873 ( .A1(n631), .A2(n770), .ZN(n877) );
  XNOR2_X1 U874 ( .A(n894), .B(n895), .ZN(n876) );
  XOR2_X1 U875 ( .A(n896), .B(n891), .Z(n894) );
  INV_X1 U876 ( .A(n897), .ZN(n891) );
  OR2_X1 U877 ( .A1(n630), .A2(n631), .ZN(n632) );
  AND2_X1 U878 ( .A1(n898), .A2(b_0_), .ZN(n643) );
  AND3_X1 U879 ( .A1(n561), .A2(n560), .A3(n558), .ZN(n562) );
  AND2_X1 U880 ( .A1(n899), .A2(b_0_), .ZN(n558) );
  INV_X1 U881 ( .A(n898), .ZN(n899) );
  OR3_X1 U882 ( .A1(n900), .A2(n901), .A3(n902), .ZN(n560) );
  XOR2_X1 U883 ( .A(n898), .B(n903), .Z(n902) );
  AND2_X1 U884 ( .A1(b_0_), .A2(a_1_), .ZN(n903) );
  AND2_X1 U885 ( .A1(b_1_), .A2(a_0_), .ZN(n898) );
  OR2_X1 U886 ( .A1(n904), .A2(n905), .ZN(n561) );
  AND2_X1 U887 ( .A1(n662), .A2(n659), .ZN(n905) );
  XNOR2_X1 U888 ( .A(n906), .B(n901), .ZN(n659) );
  INV_X1 U889 ( .A(n907), .ZN(n901) );
  OR2_X1 U890 ( .A1(n908), .A2(n909), .ZN(n907) );
  AND2_X1 U891 ( .A1(n910), .A2(n911), .ZN(n909) );
  AND2_X1 U892 ( .A1(n912), .A2(n913), .ZN(n908) );
  OR2_X1 U893 ( .A1(n911), .A2(n910), .ZN(n912) );
  OR2_X1 U894 ( .A1(n914), .A2(n900), .ZN(n906) );
  INV_X1 U895 ( .A(n915), .ZN(n900) );
  OR3_X1 U896 ( .A1(n748), .A2(n511), .A3(n516), .ZN(n915) );
  AND2_X1 U897 ( .A1(n916), .A2(n516), .ZN(n914) );
  OR2_X1 U898 ( .A1(n515), .A2(n514), .ZN(n516) );
  OR2_X1 U899 ( .A1(n748), .A2(n511), .ZN(n916) );
  AND2_X1 U900 ( .A1(b_2_), .A2(a_0_), .ZN(n662) );
  INV_X1 U901 ( .A(n661), .ZN(n904) );
  OR2_X1 U902 ( .A1(n917), .A2(n918), .ZN(n661) );
  AND2_X1 U903 ( .A1(n674), .A2(n673), .ZN(n918) );
  AND2_X1 U904 ( .A1(n671), .A2(n919), .ZN(n917) );
  OR2_X1 U905 ( .A1(n673), .A2(n674), .ZN(n919) );
  OR2_X1 U906 ( .A1(n871), .A2(n514), .ZN(n674) );
  OR2_X1 U907 ( .A1(n920), .A2(n921), .ZN(n673) );
  AND2_X1 U908 ( .A1(n708), .A2(n521), .ZN(n921) );
  AND2_X1 U909 ( .A1(n707), .A2(n922), .ZN(n920) );
  OR2_X1 U910 ( .A1(n521), .A2(n708), .ZN(n922) );
  OR2_X1 U911 ( .A1(n923), .A2(n924), .ZN(n708) );
  AND2_X1 U912 ( .A1(n741), .A2(n742), .ZN(n924) );
  AND2_X1 U913 ( .A1(n740), .A2(n925), .ZN(n923) );
  OR2_X1 U914 ( .A1(n742), .A2(n741), .ZN(n925) );
  OR2_X1 U915 ( .A1(n926), .A2(n927), .ZN(n741) );
  AND2_X1 U916 ( .A1(n883), .A2(n882), .ZN(n927) );
  AND2_X1 U917 ( .A1(n881), .A2(n928), .ZN(n926) );
  OR2_X1 U918 ( .A1(n882), .A2(n883), .ZN(n928) );
  OR2_X1 U919 ( .A1(n770), .A2(n871), .ZN(n883) );
  OR2_X1 U920 ( .A1(n929), .A2(n930), .ZN(n882) );
  AND2_X1 U921 ( .A1(n895), .A2(n897), .ZN(n930) );
  AND2_X1 U922 ( .A1(n931), .A2(n896), .ZN(n929) );
  OR2_X1 U923 ( .A1(n932), .A2(n933), .ZN(n896) );
  AND2_X1 U924 ( .A1(n934), .A2(n935), .ZN(n932) );
  OR2_X1 U925 ( .A1(n809), .A2(n511), .ZN(n934) );
  OR2_X1 U926 ( .A1(n897), .A2(n895), .ZN(n931) );
  OR2_X1 U927 ( .A1(n768), .A2(n871), .ZN(n895) );
  OR2_X1 U928 ( .A1(n893), .A2(n892), .ZN(n897) );
  OR2_X1 U929 ( .A1(n515), .A2(n809), .ZN(n892) );
  OR2_X1 U930 ( .A1(n811), .A2(n871), .ZN(n893) );
  XOR2_X1 U931 ( .A(n936), .B(n933), .Z(n881) );
  INV_X1 U932 ( .A(n937), .ZN(n933) );
  OR2_X1 U933 ( .A1(n938), .A2(n939), .ZN(n936) );
  INV_X1 U934 ( .A(n940), .ZN(n939) );
  AND2_X1 U935 ( .A1(n941), .A2(n942), .ZN(n938) );
  OR2_X1 U936 ( .A1(n811), .A2(n511), .ZN(n941) );
  OR2_X1 U937 ( .A1(n630), .A2(n871), .ZN(n742) );
  XOR2_X1 U938 ( .A(n943), .B(n944), .Z(n740) );
  XOR2_X1 U939 ( .A(n945), .B(n946), .Z(n943) );
  OR2_X1 U940 ( .A1(n748), .A2(n871), .ZN(n521) );
  XOR2_X1 U941 ( .A(n947), .B(n948), .Z(n707) );
  XOR2_X1 U942 ( .A(n949), .B(n950), .Z(n948) );
  XOR2_X1 U943 ( .A(n910), .B(n951), .Z(n671) );
  XOR2_X1 U944 ( .A(n911), .B(n913), .Z(n951) );
  OR2_X1 U945 ( .A1(n630), .A2(n511), .ZN(n913) );
  OR2_X1 U946 ( .A1(n952), .A2(n953), .ZN(n911) );
  AND2_X1 U947 ( .A1(n947), .A2(n949), .ZN(n953) );
  AND2_X1 U948 ( .A1(n954), .A2(n950), .ZN(n952) );
  OR2_X1 U949 ( .A1(n515), .A2(n630), .ZN(n950) );
  INV_X1 U950 ( .A(a_3_), .ZN(n630) );
  OR2_X1 U951 ( .A1(n949), .A2(n947), .ZN(n954) );
  OR2_X1 U952 ( .A1(n770), .A2(n511), .ZN(n947) );
  OR2_X1 U953 ( .A1(n955), .A2(n956), .ZN(n949) );
  AND2_X1 U954 ( .A1(n944), .A2(n946), .ZN(n956) );
  AND2_X1 U955 ( .A1(n945), .A2(n957), .ZN(n955) );
  OR2_X1 U956 ( .A1(n946), .A2(n944), .ZN(n957) );
  OR2_X1 U957 ( .A1(n768), .A2(n511), .ZN(n944) );
  OR2_X1 U958 ( .A1(n515), .A2(n770), .ZN(n946) );
  INV_X1 U959 ( .A(a_4_), .ZN(n770) );
  AND2_X1 U960 ( .A1(n940), .A2(n937), .ZN(n945) );
  OR3_X1 U961 ( .A1(n809), .A2(n511), .A3(n935), .ZN(n937) );
  OR2_X1 U962 ( .A1(n515), .A2(n811), .ZN(n935) );
  INV_X1 U963 ( .A(a_7_), .ZN(n809) );
  OR3_X1 U964 ( .A1(n811), .A2(n511), .A3(n942), .ZN(n940) );
  OR2_X1 U965 ( .A1(n515), .A2(n768), .ZN(n942) );
  INV_X1 U966 ( .A(a_5_), .ZN(n768) );
  INV_X1 U967 ( .A(b_0_), .ZN(n511) );
  INV_X1 U968 ( .A(a_6_), .ZN(n811) );
  OR2_X1 U969 ( .A1(n515), .A2(n748), .ZN(n910) );
  INV_X1 U970 ( .A(a_2_), .ZN(n748) );
  INV_X1 U971 ( .A(n496), .ZN(n490) );
  OR2_X1 U972 ( .A1(n958), .A2(n959), .ZN(n496) );
  AND2_X1 U973 ( .A1(n960), .A2(n681), .ZN(n959) );
  AND2_X1 U974 ( .A1(b_0_), .A2(n961), .ZN(n958) );
  OR2_X1 U975 ( .A1(n960), .A2(n681), .ZN(n961) );
  INV_X1 U976 ( .A(a_0_), .ZN(n681) );
  AND2_X1 U977 ( .A1(n962), .A2(n500), .ZN(n960) );
  OR2_X1 U978 ( .A1(b_1_), .A2(n514), .ZN(n500) );
  INV_X1 U979 ( .A(a_1_), .ZN(n514) );
  INV_X1 U980 ( .A(n963), .ZN(n962) );
  AND3_X1 U981 ( .A1(n964), .A2(n499), .A3(n965), .ZN(n963) );
  OR2_X1 U982 ( .A1(a_2_), .A2(n871), .ZN(n965) );
  OR2_X1 U983 ( .A1(a_1_), .A2(n515), .ZN(n499) );
  INV_X1 U984 ( .A(b_1_), .ZN(n515) );
  OR3_X1 U985 ( .A1(n616), .A2(n966), .A3(n967), .ZN(n964) );
  AND2_X1 U986 ( .A1(a_2_), .A2(n871), .ZN(n967) );
  INV_X1 U987 ( .A(b_2_), .ZN(n871) );
  AND3_X1 U988 ( .A1(n618), .A2(n968), .A3(n969), .ZN(n966) );
  OR3_X1 U989 ( .A1(n591), .A2(n970), .A3(n971), .ZN(n969) );
  AND2_X1 U990 ( .A1(a_4_), .A2(n698), .ZN(n971) );
  AND3_X1 U991 ( .A1(n593), .A2(n578), .A3(n972), .ZN(n970) );
  OR2_X1 U992 ( .A1(n973), .A2(n571), .ZN(n972) );
  AND2_X1 U993 ( .A1(n792), .A2(a_6_), .ZN(n571) );
  AND2_X1 U994 ( .A1(a_7_), .A2(n579), .ZN(n973) );
  INV_X1 U995 ( .A(b_7_), .ZN(n579) );
  OR2_X1 U996 ( .A1(a_6_), .A2(n792), .ZN(n578) );
  INV_X1 U997 ( .A(b_6_), .ZN(n792) );
  OR2_X1 U998 ( .A1(a_5_), .A2(n724), .ZN(n593) );
  AND2_X1 U999 ( .A1(n724), .A2(a_5_), .ZN(n591) );
  INV_X1 U1000 ( .A(b_5_), .ZN(n724) );
  OR2_X1 U1001 ( .A1(a_4_), .A2(n698), .ZN(n968) );
  INV_X1 U1002 ( .A(b_4_), .ZN(n698) );
  OR2_X1 U1003 ( .A1(a_3_), .A2(n631), .ZN(n618) );
  AND2_X1 U1004 ( .A1(n631), .A2(a_3_), .ZN(n616) );
  INV_X1 U1005 ( .A(b_3_), .ZN(n631) );
endmodule

