module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n642_, new_n211_, new_n552_, new_n342_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n318_, new_n622_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n179_, new_n572_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n598_, new_n570_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n563_, new_n148_, new_n662_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n138_, keyIn_0_41 );
xnor g001 ( new_n139_, N81, N85 );
xnor g002 ( new_n140_, N89, N93 );
xnor g003 ( new_n141_, new_n139_, new_n140_ );
not g004 ( new_n142_, new_n141_ );
xor g005 ( new_n143_, N65, N69 );
xnor g006 ( new_n144_, N73, N77 );
nand g007 ( new_n145_, new_n144_, keyIn_0_6 );
not g008 ( new_n146_, keyIn_0_6 );
not g009 ( new_n147_, N73 );
not g010 ( new_n148_, N77 );
nand g011 ( new_n149_, new_n147_, new_n148_ );
nand g012 ( new_n150_, N73, N77 );
nand g013 ( new_n151_, new_n149_, new_n146_, new_n150_ );
nand g014 ( new_n152_, new_n145_, new_n151_ );
nand g015 ( new_n153_, new_n152_, keyIn_0_5 );
not g016 ( new_n154_, keyIn_0_5 );
nand g017 ( new_n155_, new_n145_, new_n154_, new_n151_ );
nand g018 ( new_n156_, new_n153_, new_n143_, new_n155_ );
not g019 ( new_n157_, new_n143_ );
nand g020 ( new_n158_, new_n153_, new_n155_ );
nand g021 ( new_n159_, new_n158_, new_n157_ );
nand g022 ( new_n160_, new_n159_, new_n156_ );
nand g023 ( new_n161_, new_n160_, new_n142_ );
nand g024 ( new_n162_, new_n159_, new_n141_, new_n156_ );
nand g025 ( new_n163_, new_n161_, new_n162_ );
nand g026 ( new_n164_, N129, N137 );
nand g027 ( new_n165_, new_n163_, new_n164_ );
nand g028 ( new_n166_, new_n161_, N129, N137, new_n162_ );
nand g029 ( new_n167_, new_n165_, new_n166_ );
xnor g030 ( new_n168_, N1, N17 );
xnor g031 ( new_n169_, N33, N49 );
xnor g032 ( new_n170_, new_n168_, new_n169_ );
xnor g033 ( new_n171_, new_n167_, new_n170_ );
xnor g034 ( new_n172_, N97, N101 );
xnor g035 ( new_n173_, N105, N109 );
xnor g036 ( new_n174_, new_n172_, new_n173_ );
xnor g037 ( new_n175_, new_n174_, keyIn_0_18 );
nand g038 ( new_n176_, new_n160_, new_n175_ );
not g039 ( new_n177_, keyIn_0_18 );
xnor g040 ( new_n178_, new_n174_, new_n177_ );
nand g041 ( new_n179_, new_n178_, new_n156_, new_n159_ );
nand g042 ( new_n180_, new_n176_, new_n179_ );
nand g043 ( new_n181_, N131, N137 );
nand g044 ( new_n182_, new_n180_, new_n181_ );
nand g045 ( new_n183_, new_n176_, N131, new_n179_, N137 );
nand g046 ( new_n184_, new_n182_, new_n183_ );
xnor g047 ( new_n185_, N9, N25 );
xnor g048 ( new_n186_, N41, N57 );
xnor g049 ( new_n187_, new_n185_, new_n186_ );
nand g050 ( new_n188_, new_n184_, new_n187_ );
not g051 ( new_n189_, new_n187_ );
nand g052 ( new_n190_, new_n182_, new_n183_, new_n189_ );
nand g053 ( new_n191_, new_n188_, new_n190_ );
nand g054 ( new_n192_, new_n191_, keyIn_0_24 );
not g055 ( new_n193_, keyIn_0_24 );
nand g056 ( new_n194_, new_n188_, new_n193_, new_n190_ );
nand g057 ( new_n195_, new_n192_, new_n194_ );
nand g058 ( new_n196_, new_n195_, keyIn_0_26 );
not g059 ( new_n197_, keyIn_0_23 );
not g060 ( new_n198_, N121 );
not g061 ( new_n199_, N125 );
nand g062 ( new_n200_, new_n198_, new_n199_ );
nand g063 ( new_n201_, N121, N125 );
nand g064 ( new_n202_, new_n200_, new_n201_ );
nand g065 ( new_n203_, new_n202_, keyIn_0_7 );
not g066 ( new_n204_, keyIn_0_7 );
nand g067 ( new_n205_, new_n200_, new_n204_, new_n201_ );
xnor g068 ( new_n206_, N113, N117 );
nand g069 ( new_n207_, new_n203_, new_n205_, new_n206_ );
nand g070 ( new_n208_, new_n203_, new_n205_ );
not g071 ( new_n209_, new_n206_ );
nand g072 ( new_n210_, new_n208_, new_n209_ );
nand g073 ( new_n211_, new_n210_, new_n207_ );
nand g074 ( new_n212_, new_n211_, keyIn_0_19 );
not g075 ( new_n213_, keyIn_0_19 );
nand g076 ( new_n214_, new_n210_, new_n213_, new_n207_ );
nand g077 ( new_n215_, new_n212_, new_n214_ );
nand g078 ( new_n216_, new_n215_, new_n141_ );
nand g079 ( new_n217_, new_n212_, new_n142_, new_n214_ );
nand g080 ( new_n218_, new_n216_, new_n217_ );
nand g081 ( new_n219_, N132, N137 );
xnor g082 ( new_n220_, new_n219_, keyIn_0_9 );
not g083 ( new_n221_, new_n220_ );
nand g084 ( new_n222_, new_n218_, new_n221_ );
nand g085 ( new_n223_, new_n216_, new_n217_, new_n220_ );
nand g086 ( new_n224_, new_n222_, new_n223_ );
nand g087 ( new_n225_, new_n224_, new_n197_ );
nand g088 ( new_n226_, new_n222_, keyIn_0_23, new_n223_ );
nand g089 ( new_n227_, new_n225_, new_n226_ );
xor g090 ( new_n228_, N13, N29 );
xnor g091 ( new_n229_, new_n228_, keyIn_0_14 );
xnor g092 ( new_n230_, N45, N61 );
xnor g093 ( new_n231_, new_n229_, new_n230_ );
xnor g094 ( new_n232_, new_n227_, new_n231_ );
not g095 ( new_n233_, keyIn_0_26 );
nand g096 ( new_n234_, new_n192_, new_n233_, new_n194_ );
not g097 ( new_n235_, new_n234_ );
nand g098 ( new_n236_, new_n215_, new_n178_ );
nand g099 ( new_n237_, new_n175_, new_n212_, new_n214_ );
nand g100 ( new_n238_, new_n236_, new_n237_ );
nand g101 ( new_n239_, new_n238_, keyIn_0_22 );
not g102 ( new_n240_, keyIn_0_22 );
nand g103 ( new_n241_, new_n236_, new_n237_, new_n240_ );
nand g104 ( new_n242_, new_n239_, new_n241_ );
nand g105 ( new_n243_, N130, N137 );
xor g106 ( new_n244_, new_n243_, keyIn_0_8 );
not g107 ( new_n245_, new_n244_ );
nand g108 ( new_n246_, new_n242_, new_n245_ );
nand g109 ( new_n247_, new_n239_, new_n241_, new_n244_ );
nand g110 ( new_n248_, new_n246_, new_n247_ );
xor g111 ( new_n249_, N5, N21 );
xnor g112 ( new_n250_, new_n249_, keyIn_0_12 );
xor g113 ( new_n251_, N37, N53 );
xnor g114 ( new_n252_, new_n251_, keyIn_0_13 );
xnor g115 ( new_n253_, new_n250_, new_n252_ );
nand g116 ( new_n254_, new_n248_, new_n253_ );
not g117 ( new_n255_, new_n253_ );
nand g118 ( new_n256_, new_n246_, new_n247_, new_n255_ );
nand g119 ( new_n257_, new_n254_, new_n171_, new_n256_ );
nor g120 ( new_n258_, new_n235_, new_n257_ );
nand g121 ( new_n259_, new_n258_, keyIn_0_36, new_n196_, new_n232_ );
not g122 ( new_n260_, keyIn_0_36 );
not g123 ( new_n261_, new_n257_ );
nand g124 ( new_n262_, new_n261_, new_n196_, new_n232_, new_n234_ );
nand g125 ( new_n263_, new_n262_, new_n260_ );
nand g126 ( new_n264_, new_n259_, new_n263_ );
not g127 ( new_n265_, new_n171_ );
nand g128 ( new_n266_, new_n254_, new_n256_ );
nand g129 ( new_n267_, new_n266_, new_n195_, new_n265_ );
not g130 ( new_n268_, new_n195_ );
not g131 ( new_n269_, new_n266_ );
xnor g132 ( new_n270_, new_n171_, keyIn_0_25 );
nand g133 ( new_n271_, new_n270_, new_n268_, new_n269_ );
nand g134 ( new_n272_, new_n271_, new_n267_ );
nand g135 ( new_n273_, new_n272_, new_n232_ );
not g136 ( new_n274_, new_n232_ );
nand g137 ( new_n275_, new_n274_, new_n265_, new_n195_, new_n269_ );
nand g138 ( new_n276_, new_n264_, new_n273_, new_n275_ );
not g139 ( new_n277_, new_n276_ );
not g140 ( new_n278_, keyIn_0_21 );
not g141 ( new_n279_, N37 );
not g142 ( new_n280_, N33 );
nand g143 ( new_n281_, new_n280_, keyIn_0_2 );
not g144 ( new_n282_, keyIn_0_2 );
nand g145 ( new_n283_, new_n282_, N33 );
nand g146 ( new_n284_, new_n281_, new_n283_ );
nand g147 ( new_n285_, new_n284_, new_n279_ );
nand g148 ( new_n286_, new_n281_, new_n283_, N37 );
xnor g149 ( new_n287_, N41, N45 );
nand g150 ( new_n288_, new_n287_, keyIn_0_3 );
not g151 ( new_n289_, keyIn_0_3 );
not g152 ( new_n290_, N41 );
not g153 ( new_n291_, N45 );
nand g154 ( new_n292_, new_n290_, new_n291_ );
nand g155 ( new_n293_, N41, N45 );
nand g156 ( new_n294_, new_n292_, new_n289_, new_n293_ );
nand g157 ( new_n295_, new_n285_, new_n288_, new_n286_, new_n294_ );
nand g158 ( new_n296_, new_n285_, new_n286_ );
nand g159 ( new_n297_, new_n288_, new_n294_ );
nand g160 ( new_n298_, new_n296_, new_n297_ );
nand g161 ( new_n299_, new_n298_, keyIn_0_17, new_n295_ );
not g162 ( new_n300_, keyIn_0_17 );
nand g163 ( new_n301_, new_n298_, new_n295_ );
nand g164 ( new_n302_, new_n301_, new_n300_ );
nand g165 ( new_n303_, new_n302_, new_n299_ );
not g166 ( new_n304_, N5 );
nand g167 ( new_n305_, new_n304_, N1 );
not g168 ( new_n306_, N1 );
nand g169 ( new_n307_, new_n306_, N5 );
not g170 ( new_n308_, N9 );
not g171 ( new_n309_, N13 );
nand g172 ( new_n310_, new_n308_, new_n309_ );
nand g173 ( new_n311_, N9, N13 );
nand g174 ( new_n312_, new_n310_, new_n305_, new_n307_, new_n311_ );
nand g175 ( new_n313_, new_n305_, new_n307_ );
nand g176 ( new_n314_, new_n310_, new_n311_ );
nand g177 ( new_n315_, new_n313_, new_n314_ );
nand g178 ( new_n316_, new_n315_, new_n312_ );
nand g179 ( new_n317_, new_n316_, keyIn_0_16 );
not g180 ( new_n318_, keyIn_0_16 );
nand g181 ( new_n319_, new_n315_, new_n318_, new_n312_ );
nand g182 ( new_n320_, new_n317_, new_n319_ );
not g183 ( new_n321_, new_n320_ );
nand g184 ( new_n322_, new_n303_, new_n321_ );
nand g185 ( new_n323_, new_n302_, new_n299_, new_n320_ );
nand g186 ( new_n324_, new_n322_, new_n323_ );
nand g187 ( new_n325_, new_n324_, new_n278_ );
nand g188 ( new_n326_, new_n322_, keyIn_0_21, new_n323_ );
nand g189 ( new_n327_, new_n325_, new_n326_ );
nand g190 ( new_n328_, N135, N137 );
xor g191 ( new_n329_, new_n328_, keyIn_0_10 );
not g192 ( new_n330_, new_n329_ );
nand g193 ( new_n331_, new_n327_, new_n330_ );
nand g194 ( new_n332_, new_n325_, new_n326_, new_n329_ );
nand g195 ( new_n333_, new_n331_, new_n332_ );
xor g196 ( new_n334_, N73, N89 );
xnor g197 ( new_n335_, N105, N121 );
xnor g198 ( new_n336_, new_n334_, new_n335_ );
xnor g199 ( new_n337_, new_n336_, keyIn_0_20 );
not g200 ( new_n338_, new_n337_ );
nand g201 ( new_n339_, new_n333_, new_n338_ );
nand g202 ( new_n340_, new_n331_, new_n332_, new_n337_ );
nand g203 ( new_n341_, new_n339_, new_n340_ );
not g204 ( new_n342_, new_n341_ );
nor g205 ( new_n343_, new_n277_, new_n342_ );
not g206 ( new_n344_, keyIn_0_4 );
xnor g207 ( new_n345_, N57, N61 );
xnor g208 ( new_n346_, new_n345_, new_n344_ );
xor g209 ( new_n347_, N49, N53 );
xnor g210 ( new_n348_, new_n346_, new_n347_ );
nand g211 ( new_n349_, new_n303_, new_n348_ );
not g212 ( new_n350_, new_n347_ );
nand g213 ( new_n351_, new_n346_, new_n350_ );
xnor g214 ( new_n352_, new_n345_, keyIn_0_4 );
nand g215 ( new_n353_, new_n352_, new_n347_ );
nand g216 ( new_n354_, new_n351_, new_n353_ );
nand g217 ( new_n355_, new_n302_, new_n299_, new_n354_ );
nand g218 ( new_n356_, new_n349_, new_n355_ );
nand g219 ( new_n357_, N134, N137 );
nand g220 ( new_n358_, new_n356_, new_n357_ );
nand g221 ( new_n359_, new_n349_, N134, N137, new_n355_ );
xnor g222 ( new_n360_, N69, N85 );
xnor g223 ( new_n361_, N101, N117 );
xnor g224 ( new_n362_, new_n360_, new_n361_ );
not g225 ( new_n363_, new_n362_ );
nand g226 ( new_n364_, new_n358_, new_n359_, new_n363_ );
nand g227 ( new_n365_, new_n358_, new_n359_ );
nand g228 ( new_n366_, new_n365_, new_n362_ );
nand g229 ( new_n367_, new_n366_, new_n364_ );
not g230 ( new_n368_, new_n367_ );
not g231 ( new_n369_, N17 );
not g232 ( new_n370_, N21 );
nand g233 ( new_n371_, new_n369_, new_n370_ );
nand g234 ( new_n372_, N17, N21 );
nand g235 ( new_n373_, new_n371_, new_n372_ );
nand g236 ( new_n374_, new_n373_, keyIn_0_0 );
not g237 ( new_n375_, keyIn_0_0 );
nand g238 ( new_n376_, new_n371_, new_n375_, new_n372_ );
nand g239 ( new_n377_, new_n374_, new_n376_ );
not g240 ( new_n378_, N25 );
not g241 ( new_n379_, N29 );
nand g242 ( new_n380_, new_n378_, new_n379_ );
nand g243 ( new_n381_, N25, N29 );
nand g244 ( new_n382_, new_n380_, new_n381_ );
nand g245 ( new_n383_, new_n382_, keyIn_0_1 );
not g246 ( new_n384_, keyIn_0_1 );
nand g247 ( new_n385_, new_n380_, new_n384_, new_n381_ );
nand g248 ( new_n386_, new_n383_, new_n385_ );
nand g249 ( new_n387_, new_n377_, new_n386_ );
nand g250 ( new_n388_, new_n374_, new_n383_, new_n376_, new_n385_ );
nand g251 ( new_n389_, new_n387_, new_n388_ );
nand g252 ( new_n390_, new_n389_, new_n317_, new_n319_ );
nand g253 ( new_n391_, new_n320_, new_n387_, new_n388_ );
nand g254 ( new_n392_, new_n390_, new_n391_ );
nand g255 ( new_n393_, N133, N137 );
nand g256 ( new_n394_, new_n392_, new_n393_ );
nand g257 ( new_n395_, new_n390_, new_n391_, N133, N137 );
nand g258 ( new_n396_, new_n394_, new_n395_ );
xnor g259 ( new_n397_, N97, N113 );
xnor g260 ( new_n398_, new_n397_, keyIn_0_15 );
xor g261 ( new_n399_, N65, N81 );
xnor g262 ( new_n400_, new_n398_, new_n399_ );
not g263 ( new_n401_, new_n400_ );
nand g264 ( new_n402_, new_n396_, new_n401_ );
nand g265 ( new_n403_, new_n394_, new_n395_, new_n400_ );
nand g266 ( new_n404_, new_n402_, new_n403_ );
nand g267 ( new_n405_, new_n348_, new_n389_ );
nand g268 ( new_n406_, new_n354_, new_n387_, new_n388_ );
nand g269 ( new_n407_, N136, N137 );
xnor g270 ( new_n408_, new_n407_, keyIn_0_11 );
nand g271 ( new_n409_, new_n405_, new_n406_, new_n408_ );
nand g272 ( new_n410_, new_n405_, new_n406_ );
not g273 ( new_n411_, new_n408_ );
nand g274 ( new_n412_, new_n410_, new_n411_ );
nand g275 ( new_n413_, new_n412_, new_n409_ );
xnor g276 ( new_n414_, N77, N93 );
xnor g277 ( new_n415_, N109, N125 );
xnor g278 ( new_n416_, new_n414_, new_n415_ );
nand g279 ( new_n417_, new_n413_, new_n416_ );
not g280 ( new_n418_, new_n416_ );
nand g281 ( new_n419_, new_n412_, new_n409_, new_n418_ );
nand g282 ( new_n420_, new_n417_, new_n419_ );
not g283 ( new_n421_, new_n420_ );
nand g284 ( new_n422_, new_n368_, new_n404_, new_n421_ );
not g285 ( new_n423_, new_n422_ );
nand g286 ( new_n424_, new_n343_, new_n171_, new_n423_ );
xnor g287 ( new_n425_, new_n424_, new_n138_ );
nand g288 ( new_n426_, new_n425_, N1 );
xnor g289 ( new_n427_, new_n424_, keyIn_0_41 );
nand g290 ( new_n428_, new_n427_, new_n306_ );
nand g291 ( N724, new_n426_, new_n428_ );
not g292 ( new_n430_, keyIn_0_42 );
nand g293 ( new_n431_, new_n343_, new_n266_, new_n423_ );
xnor g294 ( new_n432_, new_n431_, new_n430_ );
nand g295 ( new_n433_, new_n432_, new_n304_ );
xnor g296 ( new_n434_, new_n431_, keyIn_0_42 );
nand g297 ( new_n435_, new_n434_, N5 );
nand g298 ( N725, new_n433_, new_n435_ );
nand g299 ( new_n437_, new_n343_, new_n423_ );
not g300 ( new_n438_, new_n437_ );
nand g301 ( new_n439_, new_n438_, new_n268_ );
xnor g302 ( N726, new_n439_, N9 );
nand g303 ( new_n441_, new_n438_, new_n274_ );
xnor g304 ( N727, new_n441_, N13 );
nand g305 ( new_n443_, new_n368_, new_n404_, new_n420_ );
nor g306 ( new_n444_, new_n277_, new_n341_, new_n443_ );
nand g307 ( new_n445_, new_n444_, new_n171_ );
xnor g308 ( new_n446_, new_n445_, N17 );
nand g309 ( new_n447_, new_n446_, keyIn_0_54 );
not g310 ( new_n448_, keyIn_0_54 );
xnor g311 ( new_n449_, new_n445_, new_n369_ );
nand g312 ( new_n450_, new_n449_, new_n448_ );
nand g313 ( N728, new_n447_, new_n450_ );
nand g314 ( new_n452_, new_n444_, new_n266_ );
xnor g315 ( new_n453_, new_n452_, N21 );
nand g316 ( new_n454_, new_n453_, keyIn_0_55 );
not g317 ( new_n455_, keyIn_0_55 );
xnor g318 ( new_n456_, new_n452_, new_n370_ );
nand g319 ( new_n457_, new_n456_, new_n455_ );
nand g320 ( N729, new_n454_, new_n457_ );
nand g321 ( new_n459_, new_n444_, new_n268_ );
xnor g322 ( N730, new_n459_, N25 );
not g323 ( new_n461_, keyIn_0_43 );
nand g324 ( new_n462_, new_n444_, new_n274_ );
xnor g325 ( new_n463_, new_n462_, new_n461_ );
nand g326 ( new_n464_, new_n463_, N29 );
xnor g327 ( new_n465_, new_n462_, keyIn_0_43 );
nand g328 ( new_n466_, new_n465_, new_n379_ );
nand g329 ( N731, new_n464_, new_n466_ );
not g330 ( new_n468_, new_n404_ );
nand g331 ( new_n469_, new_n367_, new_n421_, new_n468_ );
not g332 ( new_n470_, new_n469_ );
nand g333 ( new_n471_, new_n343_, new_n171_, new_n470_ );
xnor g334 ( new_n472_, new_n471_, N33 );
nand g335 ( new_n473_, new_n472_, keyIn_0_56 );
not g336 ( new_n474_, keyIn_0_56 );
xnor g337 ( new_n475_, new_n471_, new_n280_ );
nand g338 ( new_n476_, new_n475_, new_n474_ );
nand g339 ( N732, new_n473_, new_n476_ );
nand g340 ( new_n478_, new_n343_, new_n266_, new_n470_ );
xnor g341 ( new_n479_, new_n478_, new_n279_ );
nand g342 ( new_n480_, new_n479_, keyIn_0_57 );
not g343 ( new_n481_, keyIn_0_57 );
xnor g344 ( new_n482_, new_n478_, N37 );
nand g345 ( new_n483_, new_n482_, new_n481_ );
nand g346 ( N733, new_n480_, new_n483_ );
not g347 ( new_n485_, keyIn_0_44 );
nand g348 ( new_n486_, new_n343_, new_n268_, new_n470_ );
xnor g349 ( new_n487_, new_n486_, new_n485_ );
nand g350 ( new_n488_, new_n487_, N41 );
xnor g351 ( new_n489_, new_n486_, keyIn_0_44 );
nand g352 ( new_n490_, new_n489_, new_n290_ );
nand g353 ( N734, new_n488_, new_n490_ );
nand g354 ( new_n492_, new_n276_, new_n274_, new_n341_, new_n470_ );
xnor g355 ( new_n493_, new_n492_, keyIn_0_45 );
nand g356 ( new_n494_, new_n493_, new_n291_ );
not g357 ( new_n495_, keyIn_0_45 );
xnor g358 ( new_n496_, new_n492_, new_n495_ );
nand g359 ( new_n497_, new_n496_, N45 );
nand g360 ( new_n498_, new_n494_, new_n497_ );
nand g361 ( new_n499_, new_n498_, keyIn_0_58 );
not g362 ( new_n500_, keyIn_0_58 );
nand g363 ( new_n501_, new_n494_, new_n497_, new_n500_ );
nand g364 ( N735, new_n499_, new_n501_ );
not g365 ( new_n503_, N49 );
not g366 ( new_n504_, keyIn_0_39 );
xnor g367 ( new_n505_, new_n341_, keyIn_0_27 );
nand g368 ( new_n506_, new_n505_, new_n367_, new_n468_, new_n420_ );
not g369 ( new_n507_, new_n506_ );
nand g370 ( new_n508_, new_n276_, new_n507_ );
nand g371 ( new_n509_, new_n508_, new_n504_ );
nand g372 ( new_n510_, new_n276_, keyIn_0_39, new_n507_ );
nand g373 ( new_n511_, new_n509_, new_n510_ );
nand g374 ( new_n512_, new_n511_, new_n503_, new_n171_ );
nand g375 ( new_n513_, new_n511_, new_n171_ );
nand g376 ( new_n514_, new_n513_, N49 );
nand g377 ( new_n515_, new_n514_, new_n512_ );
nand g378 ( new_n516_, new_n515_, keyIn_0_59 );
not g379 ( new_n517_, keyIn_0_59 );
nand g380 ( new_n518_, new_n514_, new_n517_, new_n512_ );
nand g381 ( N736, new_n516_, new_n518_ );
not g382 ( new_n520_, keyIn_0_46 );
nand g383 ( new_n521_, new_n511_, new_n520_, new_n266_ );
nand g384 ( new_n522_, new_n511_, new_n266_ );
nand g385 ( new_n523_, new_n522_, keyIn_0_46 );
nand g386 ( new_n524_, new_n523_, new_n521_ );
nand g387 ( new_n525_, new_n524_, N53 );
not g388 ( new_n526_, N53 );
nand g389 ( new_n527_, new_n523_, new_n526_, new_n521_ );
nand g390 ( N737, new_n525_, new_n527_ );
nand g391 ( new_n529_, new_n511_, new_n268_ );
xnor g392 ( N738, new_n529_, N57 );
nand g393 ( new_n531_, new_n511_, new_n274_ );
xnor g394 ( N739, new_n531_, N61 );
not g395 ( new_n533_, N65 );
not g396 ( new_n534_, keyIn_0_40 );
not g397 ( new_n535_, keyIn_0_37 );
not g398 ( new_n536_, keyIn_0_31 );
nand g399 ( new_n537_, new_n339_, new_n536_, new_n340_ );
nand g400 ( new_n538_, new_n341_, keyIn_0_31 );
nand g401 ( new_n539_, new_n538_, new_n535_, new_n470_, new_n537_ );
nand g402 ( new_n540_, new_n538_, new_n470_, new_n537_ );
nand g403 ( new_n541_, new_n540_, keyIn_0_37 );
not g404 ( new_n542_, keyIn_0_32 );
nand g405 ( new_n543_, new_n339_, new_n542_, new_n340_ );
nand g406 ( new_n544_, new_n341_, keyIn_0_32 );
not g407 ( new_n545_, keyIn_0_33 );
nand g408 ( new_n546_, new_n420_, new_n545_ );
nand g409 ( new_n547_, new_n417_, keyIn_0_33, new_n419_ );
nand g410 ( new_n548_, new_n546_, new_n547_ );
nor g411 ( new_n549_, new_n548_, new_n367_, new_n468_ );
nand g412 ( new_n550_, new_n544_, new_n543_, new_n549_ );
nand g413 ( new_n551_, new_n367_, keyIn_0_28 );
not g414 ( new_n552_, keyIn_0_28 );
nand g415 ( new_n553_, new_n366_, new_n552_, new_n364_ );
nand g416 ( new_n554_, new_n551_, new_n553_ );
nor g417 ( new_n555_, new_n421_, new_n404_ );
nand g418 ( new_n556_, new_n554_, new_n339_, new_n340_, new_n555_ );
not g419 ( new_n557_, keyIn_0_30 );
xnor g420 ( new_n558_, new_n420_, new_n557_ );
not g421 ( new_n559_, keyIn_0_29 );
nand g422 ( new_n560_, new_n402_, new_n559_, new_n403_ );
nand g423 ( new_n561_, new_n404_, keyIn_0_29 );
nand g424 ( new_n562_, new_n561_, new_n560_ );
nor g425 ( new_n563_, new_n562_, new_n367_ );
nand g426 ( new_n564_, new_n341_, new_n558_, new_n563_ );
nand g427 ( new_n565_, new_n556_, new_n564_ );
not g428 ( new_n566_, new_n565_ );
nand g429 ( new_n567_, new_n541_, new_n566_, new_n539_, new_n550_ );
nand g430 ( new_n568_, new_n567_, keyIn_0_38 );
not g431 ( new_n569_, keyIn_0_38 );
not g432 ( new_n570_, new_n550_ );
nor g433 ( new_n571_, new_n570_, new_n565_ );
nand g434 ( new_n572_, new_n571_, new_n569_, new_n539_, new_n541_ );
nand g435 ( new_n573_, new_n268_, new_n232_ );
nor g436 ( new_n574_, new_n573_, new_n257_ );
nand g437 ( new_n575_, new_n568_, new_n572_, new_n534_, new_n574_ );
nand g438 ( new_n576_, new_n568_, new_n572_, new_n574_ );
nand g439 ( new_n577_, new_n576_, keyIn_0_40 );
nand g440 ( new_n578_, new_n577_, new_n575_ );
nand g441 ( new_n579_, new_n578_, new_n404_ );
nand g442 ( new_n580_, new_n579_, keyIn_0_47 );
not g443 ( new_n581_, keyIn_0_47 );
nand g444 ( new_n582_, new_n578_, new_n581_, new_n404_ );
nand g445 ( new_n583_, new_n580_, new_n582_ );
nand g446 ( new_n584_, new_n583_, new_n533_ );
nand g447 ( new_n585_, new_n580_, N65, new_n582_ );
nand g448 ( N740, new_n584_, new_n585_ );
not g449 ( new_n587_, N69 );
nand g450 ( new_n588_, new_n578_, new_n367_ );
nand g451 ( new_n589_, new_n588_, keyIn_0_48 );
not g452 ( new_n590_, keyIn_0_48 );
nand g453 ( new_n591_, new_n578_, new_n590_, new_n367_ );
nand g454 ( new_n592_, new_n589_, new_n591_ );
nand g455 ( new_n593_, new_n592_, new_n587_ );
nand g456 ( new_n594_, new_n589_, N69, new_n591_ );
nand g457 ( N741, new_n593_, new_n594_ );
nand g458 ( new_n596_, new_n578_, new_n341_ );
xnor g459 ( N742, new_n596_, N73 );
nand g460 ( new_n598_, new_n578_, new_n420_ );
nand g461 ( new_n599_, new_n598_, N77 );
nand g462 ( new_n600_, new_n578_, new_n148_, new_n420_ );
nand g463 ( new_n601_, new_n599_, new_n600_ );
nand g464 ( new_n602_, new_n601_, keyIn_0_60 );
not g465 ( new_n603_, keyIn_0_60 );
nand g466 ( new_n604_, new_n599_, new_n603_, new_n600_ );
nand g467 ( N743, new_n602_, new_n604_ );
xnor g468 ( new_n606_, new_n567_, new_n569_ );
xnor g469 ( new_n607_, new_n266_, keyIn_0_34 );
nor g470 ( new_n608_, new_n607_, new_n265_, new_n268_, new_n232_ );
nand g471 ( new_n609_, new_n606_, new_n608_ );
not g472 ( new_n610_, new_n609_ );
nand g473 ( new_n611_, new_n610_, new_n404_ );
xnor g474 ( N744, new_n611_, N81 );
nand g475 ( new_n613_, new_n606_, new_n367_, new_n608_ );
xnor g476 ( new_n614_, new_n613_, keyIn_0_49 );
xnor g477 ( N745, new_n614_, N85 );
nand g478 ( new_n616_, new_n606_, new_n341_, new_n608_ );
xnor g479 ( new_n617_, new_n616_, N89 );
xnor g480 ( N746, new_n617_, keyIn_0_61 );
nand g481 ( new_n619_, new_n610_, new_n420_ );
xnor g482 ( N747, new_n619_, N93 );
xor g483 ( new_n621_, new_n171_, keyIn_0_35 );
nor g484 ( new_n622_, new_n573_, new_n621_, new_n269_ );
nand g485 ( new_n623_, new_n606_, new_n622_ );
not g486 ( new_n624_, new_n623_ );
nand g487 ( new_n625_, new_n624_, new_n404_ );
xnor g488 ( N748, new_n625_, N97 );
nand g489 ( new_n627_, new_n606_, new_n367_, new_n622_ );
xnor g490 ( new_n628_, new_n627_, keyIn_0_50 );
xnor g491 ( N749, new_n628_, N101 );
nand g492 ( new_n630_, new_n624_, new_n341_ );
xnor g493 ( N750, new_n630_, N105 );
nand g494 ( new_n632_, new_n624_, new_n420_ );
xnor g495 ( N751, new_n632_, N109 );
nand g496 ( new_n634_, new_n274_, new_n265_, new_n195_, new_n266_ );
not g497 ( new_n635_, new_n634_ );
nand g498 ( new_n636_, new_n606_, new_n404_, new_n635_ );
xnor g499 ( N752, new_n636_, N113 );
not g500 ( new_n638_, N117 );
nand g501 ( new_n639_, new_n606_, new_n367_, new_n635_ );
xnor g502 ( new_n640_, new_n639_, keyIn_0_51 );
xnor g503 ( N753, new_n640_, new_n638_ );
not g504 ( new_n642_, keyIn_0_62 );
nand g505 ( new_n643_, new_n568_, new_n572_, new_n341_, new_n635_ );
xnor g506 ( new_n644_, new_n643_, keyIn_0_52 );
nand g507 ( new_n645_, new_n644_, new_n198_ );
not g508 ( new_n646_, keyIn_0_52 );
xnor g509 ( new_n647_, new_n643_, new_n646_ );
nand g510 ( new_n648_, new_n647_, N121 );
nand g511 ( new_n649_, new_n645_, new_n648_ );
nand g512 ( new_n650_, new_n649_, new_n642_ );
nand g513 ( new_n651_, new_n645_, new_n648_, keyIn_0_62 );
nand g514 ( N754, new_n650_, new_n651_ );
not g515 ( new_n653_, keyIn_0_63 );
nand g516 ( new_n654_, new_n568_, new_n572_, new_n420_, new_n635_ );
xnor g517 ( new_n655_, new_n654_, keyIn_0_53 );
nand g518 ( new_n656_, new_n655_, N125 );
not g519 ( new_n657_, keyIn_0_53 );
xnor g520 ( new_n658_, new_n654_, new_n657_ );
nand g521 ( new_n659_, new_n658_, new_n199_ );
nand g522 ( new_n660_, new_n656_, new_n659_ );
nand g523 ( new_n661_, new_n660_, new_n653_ );
nand g524 ( new_n662_, new_n656_, new_n659_, keyIn_0_63 );
nand g525 ( N755, new_n661_, new_n662_ );
endmodule