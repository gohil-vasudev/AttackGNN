module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n170_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n121_, new_n415_, new_n537_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n108_, keyIn_0_26 );
and g001 ( new_n109_, keyIn_0_14, N89 );
not g002 ( new_n110_, keyIn_0_14 );
not g003 ( new_n111_, N89 );
and g004 ( new_n112_, new_n110_, new_n111_ );
or g005 ( new_n113_, new_n112_, new_n109_ );
and g006 ( new_n114_, new_n113_, new_n108_, N95 );
not g007 ( new_n115_, N95 );
not g008 ( new_n116_, new_n109_ );
or g009 ( new_n117_, keyIn_0_14, N89 );
and g010 ( new_n118_, new_n116_, new_n117_ );
or g011 ( new_n119_, new_n118_, new_n115_ );
and g012 ( new_n120_, new_n119_, keyIn_0_26 );
or g013 ( new_n121_, new_n120_, new_n114_ );
not g014 ( new_n122_, keyIn_0_25 );
and g015 ( new_n123_, keyIn_0_12, N76 );
not g016 ( new_n124_, new_n123_ );
or g017 ( new_n125_, keyIn_0_12, N76 );
and g018 ( new_n126_, new_n124_, new_n125_ );
not g019 ( new_n127_, new_n126_ );
and g020 ( new_n128_, new_n127_, new_n122_, N82 );
not g021 ( new_n129_, N82 );
or g022 ( new_n130_, new_n126_, new_n129_ );
and g023 ( new_n131_, new_n130_, keyIn_0_25 );
or g024 ( new_n132_, new_n131_, new_n128_ );
not g025 ( new_n133_, keyIn_0_27 );
or g026 ( new_n134_, keyIn_0_16, N102 );
and g027 ( new_n135_, keyIn_0_16, N102 );
not g028 ( new_n136_, new_n135_ );
and g029 ( new_n137_, new_n136_, N108, new_n134_ );
not g030 ( new_n138_, new_n137_ );
or g031 ( new_n139_, new_n138_, new_n133_ );
or g032 ( new_n140_, new_n137_, keyIn_0_27 );
and g033 ( new_n141_, new_n139_, new_n140_ );
and g034 ( new_n142_, new_n121_, new_n132_, new_n141_ );
not g035 ( new_n143_, keyIn_0_23 );
not g036 ( new_n144_, N56 );
not g037 ( new_n145_, keyIn_0_8 );
or g038 ( new_n146_, new_n145_, N50 );
not g039 ( new_n147_, N50 );
or g040 ( new_n148_, new_n147_, keyIn_0_8 );
and g041 ( new_n149_, new_n146_, new_n148_ );
or g042 ( new_n150_, new_n149_, new_n144_ );
and g043 ( new_n151_, new_n150_, new_n143_ );
not g044 ( new_n152_, new_n149_ );
and g045 ( new_n153_, new_n152_, keyIn_0_23, N56 );
or g046 ( new_n154_, new_n151_, new_n153_ );
not g047 ( new_n155_, keyIn_0_24 );
not g048 ( new_n156_, keyIn_0_10 );
not g049 ( new_n157_, N63 );
and g050 ( new_n158_, new_n156_, new_n157_ );
and g051 ( new_n159_, keyIn_0_10, N63 );
or g052 ( new_n160_, new_n158_, new_n159_ );
and g053 ( new_n161_, new_n160_, N69 );
or g054 ( new_n162_, new_n161_, new_n155_ );
not g055 ( new_n163_, N69 );
not g056 ( new_n164_, new_n160_ );
or g057 ( new_n165_, new_n164_, keyIn_0_24, new_n163_ );
and g058 ( new_n166_, new_n162_, new_n165_ );
and g059 ( new_n167_, new_n154_, new_n166_ );
not g060 ( new_n168_, keyIn_0_4 );
not g061 ( new_n169_, N24 );
and g062 ( new_n170_, new_n168_, new_n169_ );
and g063 ( new_n171_, keyIn_0_4, N24 );
or g064 ( new_n172_, new_n170_, new_n171_ );
and g065 ( new_n173_, new_n172_, N30 );
or g066 ( new_n174_, new_n173_, keyIn_0_21 );
not g067 ( new_n175_, keyIn_0_21 );
not g068 ( new_n176_, N30 );
not g069 ( new_n177_, new_n172_ );
or g070 ( new_n178_, new_n177_, new_n175_, new_n176_ );
and g071 ( new_n179_, new_n174_, new_n178_ );
not g072 ( new_n180_, keyIn_0_6 );
not g073 ( new_n181_, N37 );
and g074 ( new_n182_, new_n180_, new_n181_ );
and g075 ( new_n183_, keyIn_0_6, N37 );
or g076 ( new_n184_, new_n182_, new_n183_ );
and g077 ( new_n185_, new_n184_, N43 );
or g078 ( new_n186_, new_n185_, keyIn_0_22 );
not g079 ( new_n187_, keyIn_0_22 );
not g080 ( new_n188_, N43 );
not g081 ( new_n189_, new_n184_ );
or g082 ( new_n190_, new_n189_, new_n187_, new_n188_ );
and g083 ( new_n191_, new_n186_, new_n190_ );
not g084 ( new_n192_, keyIn_0_18 );
not g085 ( new_n193_, keyIn_0_0 );
or g086 ( new_n194_, new_n193_, N1 );
not g087 ( new_n195_, N1 );
or g088 ( new_n196_, new_n195_, keyIn_0_0 );
and g089 ( new_n197_, new_n194_, new_n196_ );
not g090 ( new_n198_, new_n197_ );
and g091 ( new_n199_, new_n198_, new_n192_, N4 );
not g092 ( new_n200_, N4 );
or g093 ( new_n201_, new_n197_, new_n200_ );
and g094 ( new_n202_, new_n201_, keyIn_0_18 );
or g095 ( new_n203_, new_n202_, new_n199_ );
not g096 ( new_n204_, N17 );
or g097 ( new_n205_, keyIn_0_2, N11 );
not g098 ( new_n206_, new_n205_ );
and g099 ( new_n207_, keyIn_0_2, N11 );
or g100 ( new_n208_, new_n206_, new_n204_, new_n207_ );
and g101 ( new_n209_, new_n208_, keyIn_0_20 );
not g102 ( new_n210_, keyIn_0_20 );
not g103 ( new_n211_, new_n207_ );
and g104 ( new_n212_, new_n211_, new_n210_, N17, new_n205_ );
or g105 ( new_n213_, new_n209_, new_n212_ );
and g106 ( new_n214_, new_n203_, new_n179_, new_n191_, new_n213_ );
and g107 ( new_n215_, new_n214_, keyIn_0_36, new_n142_, new_n167_ );
not g108 ( new_n216_, new_n215_ );
and g109 ( new_n217_, new_n179_, new_n191_ );
and g110 ( new_n218_, new_n203_, new_n213_ );
and g111 ( new_n219_, new_n142_, new_n167_, new_n218_, new_n217_ );
or g112 ( new_n220_, new_n219_, keyIn_0_36 );
and g113 ( N223, new_n220_, new_n216_ );
not g114 ( new_n222_, keyIn_0_60 );
not g115 ( new_n223_, new_n132_ );
or g116 ( new_n224_, N223, keyIn_0_37 );
and g117 ( new_n225_, new_n220_, keyIn_0_37, new_n216_ );
not g118 ( new_n226_, new_n225_ );
and g119 ( new_n227_, new_n224_, new_n226_ );
or g120 ( new_n228_, new_n227_, new_n223_ );
and g121 ( new_n229_, new_n227_, new_n223_ );
not g122 ( new_n230_, new_n229_ );
and g123 ( new_n231_, new_n230_, new_n228_ );
or g124 ( new_n232_, new_n231_, keyIn_0_44 );
and g125 ( new_n233_, new_n231_, keyIn_0_44 );
not g126 ( new_n234_, new_n233_ );
and g127 ( new_n235_, new_n234_, new_n232_ );
not g128 ( new_n236_, keyIn_0_33 );
and g129 ( new_n237_, keyIn_0_13, N82 );
or g130 ( new_n238_, keyIn_0_13, N82 );
not g131 ( new_n239_, new_n238_ );
or g132 ( new_n240_, new_n239_, N86, new_n237_ );
and g133 ( new_n241_, new_n240_, new_n236_ );
not g134 ( new_n242_, new_n241_ );
or g135 ( new_n243_, new_n240_, new_n236_ );
and g136 ( new_n244_, new_n242_, new_n243_ );
or g137 ( new_n245_, new_n235_, new_n244_ );
or g138 ( new_n246_, new_n245_, keyIn_0_53 );
not g139 ( new_n247_, keyIn_0_53 );
not g140 ( new_n248_, new_n232_ );
or g141 ( new_n249_, new_n248_, new_n233_ );
not g142 ( new_n250_, new_n244_ );
and g143 ( new_n251_, new_n249_, new_n250_ );
or g144 ( new_n252_, new_n251_, new_n247_ );
not g145 ( new_n253_, new_n141_ );
or g146 ( new_n254_, new_n227_, new_n253_ );
and g147 ( new_n255_, new_n224_, new_n253_, new_n226_ );
not g148 ( new_n256_, new_n255_ );
and g149 ( new_n257_, new_n254_, new_n256_ );
or g150 ( new_n258_, new_n257_, keyIn_0_46 );
and g151 ( new_n259_, new_n254_, keyIn_0_46, new_n256_ );
not g152 ( new_n260_, new_n259_ );
and g153 ( new_n261_, new_n258_, new_n260_ );
not g154 ( new_n262_, new_n261_ );
not g155 ( new_n263_, keyIn_0_35 );
not g156 ( new_n264_, N108 );
and g157 ( new_n265_, new_n264_, keyIn_0_17 );
not g158 ( new_n266_, new_n265_ );
or g159 ( new_n267_, new_n264_, keyIn_0_17 );
and g160 ( new_n268_, new_n266_, new_n267_ );
not g161 ( new_n269_, new_n268_ );
or g162 ( new_n270_, new_n269_, N112 );
and g163 ( new_n271_, new_n270_, new_n263_ );
not g164 ( new_n272_, new_n271_ );
or g165 ( new_n273_, new_n270_, new_n263_ );
and g166 ( new_n274_, new_n272_, new_n273_ );
and g167 ( new_n275_, new_n262_, keyIn_0_55, new_n274_ );
not g168 ( new_n276_, keyIn_0_55 );
not g169 ( new_n277_, new_n274_ );
or g170 ( new_n278_, new_n261_, new_n277_ );
and g171 ( new_n279_, new_n278_, new_n276_ );
or g172 ( new_n280_, new_n279_, new_n275_ );
not g173 ( new_n281_, keyIn_0_54 );
not g174 ( new_n282_, new_n121_ );
or g175 ( new_n283_, new_n227_, new_n282_ );
and g176 ( new_n284_, new_n224_, new_n282_, new_n226_ );
not g177 ( new_n285_, new_n284_ );
and g178 ( new_n286_, new_n283_, new_n285_ );
or g179 ( new_n287_, new_n286_, keyIn_0_45 );
and g180 ( new_n288_, new_n283_, keyIn_0_45, new_n285_ );
not g181 ( new_n289_, new_n288_ );
and g182 ( new_n290_, new_n287_, new_n289_ );
not g183 ( new_n291_, new_n290_ );
and g184 ( new_n292_, new_n115_, keyIn_0_15 );
not g185 ( new_n293_, new_n292_ );
or g186 ( new_n294_, new_n115_, keyIn_0_15 );
and g187 ( new_n295_, new_n293_, new_n294_ );
not g188 ( new_n296_, new_n295_ );
or g189 ( new_n297_, new_n296_, N99 );
and g190 ( new_n298_, new_n297_, keyIn_0_34 );
not g191 ( new_n299_, new_n298_ );
or g192 ( new_n300_, new_n297_, keyIn_0_34 );
and g193 ( new_n301_, new_n299_, new_n300_ );
and g194 ( new_n302_, new_n291_, new_n281_, new_n301_ );
not g195 ( new_n303_, new_n301_ );
or g196 ( new_n304_, new_n290_, new_n303_ );
and g197 ( new_n305_, new_n304_, keyIn_0_54 );
or g198 ( new_n306_, new_n305_, new_n302_ );
and g199 ( new_n307_, new_n280_, new_n306_, new_n246_, new_n252_ );
not g200 ( new_n308_, keyIn_0_51 );
not g201 ( new_n309_, new_n154_ );
or g202 ( new_n310_, new_n227_, new_n309_ );
and g203 ( new_n311_, new_n227_, new_n309_ );
not g204 ( new_n312_, new_n311_ );
and g205 ( new_n313_, new_n312_, new_n310_ );
or g206 ( new_n314_, new_n313_, keyIn_0_42 );
and g207 ( new_n315_, new_n312_, keyIn_0_42, new_n310_ );
not g208 ( new_n316_, new_n315_ );
not g209 ( new_n317_, N60 );
and g210 ( new_n318_, keyIn_0_9, N56 );
not g211 ( new_n319_, new_n318_ );
or g212 ( new_n320_, keyIn_0_9, N56 );
and g213 ( new_n321_, new_n319_, new_n320_ );
and g214 ( new_n322_, new_n321_, new_n317_ );
or g215 ( new_n323_, new_n322_, keyIn_0_31 );
not g216 ( new_n324_, keyIn_0_31 );
not g217 ( new_n325_, new_n322_ );
or g218 ( new_n326_, new_n325_, new_n324_ );
and g219 ( new_n327_, new_n326_, new_n323_ );
and g220 ( new_n328_, new_n314_, new_n316_, new_n327_ );
not g221 ( new_n329_, new_n328_ );
and g222 ( new_n330_, new_n329_, new_n308_ );
and g223 ( new_n331_, new_n328_, keyIn_0_51 );
or g224 ( new_n332_, new_n330_, new_n331_ );
not g225 ( new_n333_, new_n166_ );
or g226 ( new_n334_, new_n227_, new_n333_ );
and g227 ( new_n335_, new_n227_, new_n333_ );
not g228 ( new_n336_, new_n335_ );
and g229 ( new_n337_, new_n336_, new_n334_ );
or g230 ( new_n338_, new_n337_, keyIn_0_43 );
and g231 ( new_n339_, new_n336_, keyIn_0_43, new_n334_ );
not g232 ( new_n340_, new_n339_ );
not g233 ( new_n341_, keyIn_0_32 );
and g234 ( new_n342_, new_n163_, keyIn_0_11 );
not g235 ( new_n343_, new_n342_ );
or g236 ( new_n344_, new_n163_, keyIn_0_11 );
and g237 ( new_n345_, new_n343_, new_n344_ );
or g238 ( new_n346_, new_n345_, N73 );
not g239 ( new_n347_, new_n346_ );
or g240 ( new_n348_, new_n347_, new_n341_ );
or g241 ( new_n349_, new_n346_, keyIn_0_32 );
and g242 ( new_n350_, new_n348_, new_n349_ );
and g243 ( new_n351_, new_n338_, new_n340_, new_n350_ );
not g244 ( new_n352_, new_n351_ );
and g245 ( new_n353_, new_n352_, keyIn_0_52 );
not g246 ( new_n354_, keyIn_0_52 );
and g247 ( new_n355_, new_n351_, new_n354_ );
or g248 ( new_n356_, new_n353_, new_n355_ );
and g249 ( new_n357_, new_n332_, new_n356_ );
not g250 ( new_n358_, keyIn_0_38 );
not g251 ( new_n359_, new_n203_ );
or g252 ( new_n360_, new_n227_, new_n359_ );
and g253 ( new_n361_, new_n227_, new_n359_ );
not g254 ( new_n362_, new_n361_ );
and g255 ( new_n363_, new_n362_, new_n360_ );
or g256 ( new_n364_, new_n363_, new_n358_ );
and g257 ( new_n365_, new_n363_, new_n358_ );
not g258 ( new_n366_, new_n365_ );
not g259 ( new_n367_, keyIn_0_19 );
and g260 ( new_n368_, keyIn_0_1, N4 );
not g261 ( new_n369_, new_n368_ );
or g262 ( new_n370_, keyIn_0_1, N4 );
and g263 ( new_n371_, new_n369_, new_n370_ );
or g264 ( new_n372_, new_n371_, N8 );
and g265 ( new_n373_, new_n372_, new_n367_ );
not g266 ( new_n374_, new_n372_ );
and g267 ( new_n375_, new_n374_, keyIn_0_19 );
or g268 ( new_n376_, new_n375_, new_n373_ );
and g269 ( new_n377_, new_n366_, keyIn_0_47, new_n364_, new_n376_ );
not g270 ( new_n378_, new_n377_ );
and g271 ( new_n379_, new_n366_, new_n364_, new_n376_ );
or g272 ( new_n380_, new_n379_, keyIn_0_47 );
and g273 ( new_n381_, new_n380_, new_n378_ );
not g274 ( new_n382_, keyIn_0_48 );
not g275 ( new_n383_, keyIn_0_39 );
not g276 ( new_n384_, new_n213_ );
or g277 ( new_n385_, new_n227_, new_n384_ );
and g278 ( new_n386_, new_n227_, new_n384_ );
not g279 ( new_n387_, new_n386_ );
and g280 ( new_n388_, new_n387_, new_n385_ );
and g281 ( new_n389_, new_n388_, new_n383_ );
not g282 ( new_n390_, new_n388_ );
and g283 ( new_n391_, new_n390_, keyIn_0_39 );
or g284 ( new_n392_, new_n391_, new_n389_ );
not g285 ( new_n393_, new_n392_ );
and g286 ( new_n394_, new_n204_, keyIn_0_3 );
not g287 ( new_n395_, new_n394_ );
or g288 ( new_n396_, new_n204_, keyIn_0_3 );
and g289 ( new_n397_, new_n395_, new_n396_ );
or g290 ( new_n398_, new_n397_, N21 );
and g291 ( new_n399_, new_n398_, keyIn_0_28 );
not g292 ( new_n400_, new_n399_ );
or g293 ( new_n401_, new_n398_, keyIn_0_28 );
and g294 ( new_n402_, new_n400_, new_n401_ );
not g295 ( new_n403_, new_n402_ );
or g296 ( new_n404_, new_n393_, new_n382_, new_n403_ );
and g297 ( new_n405_, new_n392_, new_n402_ );
or g298 ( new_n406_, new_n405_, keyIn_0_48 );
and g299 ( new_n407_, new_n381_, new_n406_, new_n404_ );
not g300 ( new_n408_, keyIn_0_49 );
not g301 ( new_n409_, new_n179_ );
or g302 ( new_n410_, new_n227_, new_n409_ );
and g303 ( new_n411_, new_n227_, new_n409_ );
not g304 ( new_n412_, new_n411_ );
and g305 ( new_n413_, new_n412_, new_n410_ );
and g306 ( new_n414_, new_n413_, keyIn_0_40 );
not g307 ( new_n415_, new_n414_ );
or g308 ( new_n416_, new_n413_, keyIn_0_40 );
not g309 ( new_n417_, N34 );
and g310 ( new_n418_, keyIn_0_5, N30 );
not g311 ( new_n419_, new_n418_ );
or g312 ( new_n420_, keyIn_0_5, N30 );
and g313 ( new_n421_, new_n419_, new_n420_ );
and g314 ( new_n422_, new_n421_, new_n417_ );
not g315 ( new_n423_, new_n422_ );
and g316 ( new_n424_, new_n423_, keyIn_0_29 );
not g317 ( new_n425_, keyIn_0_29 );
and g318 ( new_n426_, new_n422_, new_n425_ );
or g319 ( new_n427_, new_n424_, new_n426_ );
and g320 ( new_n428_, new_n415_, new_n408_, new_n416_, new_n427_ );
not g321 ( new_n429_, new_n428_ );
and g322 ( new_n430_, new_n415_, new_n416_, new_n427_ );
or g323 ( new_n431_, new_n430_, new_n408_ );
and g324 ( new_n432_, new_n431_, new_n429_ );
not g325 ( new_n433_, new_n191_ );
or g326 ( new_n434_, new_n227_, new_n433_ );
not g327 ( new_n435_, new_n434_ );
and g328 ( new_n436_, new_n227_, new_n433_ );
or g329 ( new_n437_, new_n435_, new_n436_ );
and g330 ( new_n438_, new_n437_, keyIn_0_41 );
not g331 ( new_n439_, keyIn_0_41 );
not g332 ( new_n440_, new_n436_ );
and g333 ( new_n441_, new_n440_, new_n434_ );
and g334 ( new_n442_, new_n441_, new_n439_ );
or g335 ( new_n443_, new_n438_, new_n442_ );
not g336 ( new_n444_, keyIn_0_30 );
and g337 ( new_n445_, new_n188_, keyIn_0_7 );
not g338 ( new_n446_, new_n445_ );
or g339 ( new_n447_, new_n188_, keyIn_0_7 );
and g340 ( new_n448_, new_n446_, new_n447_ );
not g341 ( new_n449_, new_n448_ );
or g342 ( new_n450_, new_n449_, N47 );
and g343 ( new_n451_, new_n450_, new_n444_ );
not g344 ( new_n452_, new_n451_ );
or g345 ( new_n453_, new_n450_, new_n444_ );
and g346 ( new_n454_, new_n452_, new_n453_ );
and g347 ( new_n455_, new_n443_, new_n454_ );
or g348 ( new_n456_, new_n455_, keyIn_0_50 );
not g349 ( new_n457_, keyIn_0_50 );
not g350 ( new_n458_, new_n443_ );
not g351 ( new_n459_, new_n454_ );
or g352 ( new_n460_, new_n458_, new_n457_, new_n459_ );
and g353 ( new_n461_, new_n432_, new_n456_, new_n460_ );
and g354 ( new_n462_, new_n407_, new_n461_ );
and g355 ( new_n463_, new_n462_, new_n222_, new_n307_, new_n357_ );
not g356 ( new_n464_, new_n463_ );
and g357 ( new_n465_, new_n307_, new_n357_, new_n407_, new_n461_ );
or g358 ( new_n466_, new_n465_, new_n222_ );
and g359 ( N329, new_n466_, new_n464_ );
not g360 ( new_n468_, keyIn_0_62 );
and g361 ( new_n469_, new_n406_, new_n404_ );
not g362 ( new_n470_, new_n469_ );
not g363 ( new_n471_, keyIn_0_61 );
or g364 ( new_n472_, N329, new_n471_ );
and g365 ( new_n473_, new_n466_, new_n464_, new_n471_ );
not g366 ( new_n474_, new_n473_ );
and g367 ( new_n475_, new_n472_, new_n470_, new_n474_ );
not g368 ( new_n476_, new_n475_ );
and g369 ( new_n477_, new_n472_, new_n474_ );
or g370 ( new_n478_, new_n477_, new_n470_ );
and g371 ( new_n479_, new_n478_, new_n476_ );
or g372 ( new_n480_, new_n393_, N27, new_n397_ );
or g373 ( new_n481_, new_n479_, new_n480_ );
not g374 ( new_n482_, new_n356_ );
and g375 ( new_n483_, new_n472_, new_n482_, new_n474_ );
not g376 ( new_n484_, new_n483_ );
or g377 ( new_n485_, new_n477_, new_n482_ );
and g378 ( new_n486_, new_n485_, new_n484_ );
not g379 ( new_n487_, N79 );
not g380 ( new_n488_, new_n345_ );
and g381 ( new_n489_, new_n338_, new_n487_, new_n340_, new_n488_ );
and g382 ( new_n490_, new_n489_, keyIn_0_56 );
not g383 ( new_n491_, new_n490_ );
or g384 ( new_n492_, new_n489_, keyIn_0_56 );
and g385 ( new_n493_, new_n491_, new_n492_ );
or g386 ( new_n494_, new_n486_, new_n493_ );
not g387 ( new_n495_, new_n381_ );
and g388 ( new_n496_, new_n472_, new_n495_, new_n474_ );
not g389 ( new_n497_, new_n496_ );
or g390 ( new_n498_, new_n477_, new_n495_ );
and g391 ( new_n499_, new_n498_, new_n497_ );
not g392 ( new_n500_, N14 );
not g393 ( new_n501_, new_n371_ );
and g394 ( new_n502_, new_n366_, new_n500_, new_n364_, new_n501_ );
not g395 ( new_n503_, new_n502_ );
or g396 ( new_n504_, new_n499_, new_n503_ );
and g397 ( new_n505_, new_n481_, new_n494_, new_n504_ );
and g398 ( new_n506_, new_n456_, new_n460_ );
not g399 ( new_n507_, new_n506_ );
and g400 ( new_n508_, new_n472_, new_n507_, new_n474_ );
not g401 ( new_n509_, new_n508_ );
or g402 ( new_n510_, new_n477_, new_n507_ );
and g403 ( new_n511_, new_n510_, new_n509_ );
or g404 ( new_n512_, new_n458_, N53, new_n449_ );
or g405 ( new_n513_, new_n511_, new_n512_ );
not g406 ( new_n514_, new_n332_ );
and g407 ( new_n515_, new_n472_, new_n514_, new_n474_ );
not g408 ( new_n516_, new_n515_ );
or g409 ( new_n517_, new_n477_, new_n514_ );
and g410 ( new_n518_, new_n517_, new_n516_ );
not g411 ( new_n519_, N66 );
and g412 ( new_n520_, new_n314_, new_n519_, new_n316_, new_n321_ );
not g413 ( new_n521_, new_n520_ );
or g414 ( new_n522_, new_n518_, new_n521_ );
and g415 ( new_n523_, new_n513_, new_n522_ );
not g416 ( new_n524_, new_n306_ );
and g417 ( new_n525_, new_n472_, new_n524_, new_n474_ );
not g418 ( new_n526_, new_n525_ );
or g419 ( new_n527_, new_n477_, new_n524_ );
and g420 ( new_n528_, new_n527_, new_n526_ );
not g421 ( new_n529_, keyIn_0_58 );
or g422 ( new_n530_, new_n290_, N105, new_n296_ );
and g423 ( new_n531_, new_n530_, new_n529_ );
not g424 ( new_n532_, new_n530_ );
and g425 ( new_n533_, new_n532_, keyIn_0_58 );
or g426 ( new_n534_, new_n533_, new_n531_ );
or g427 ( new_n535_, new_n528_, new_n534_ );
not g428 ( new_n536_, new_n280_ );
and g429 ( new_n537_, new_n472_, new_n536_, new_n474_ );
not g430 ( new_n538_, new_n537_ );
or g431 ( new_n539_, new_n477_, new_n536_ );
and g432 ( new_n540_, new_n539_, new_n538_ );
not g433 ( new_n541_, keyIn_0_59 );
or g434 ( new_n542_, new_n261_, N115, new_n269_ );
not g435 ( new_n543_, new_n542_ );
and g436 ( new_n544_, new_n543_, new_n541_ );
and g437 ( new_n545_, new_n542_, keyIn_0_59 );
or g438 ( new_n546_, new_n544_, new_n545_ );
or g439 ( new_n547_, new_n540_, new_n546_ );
not g440 ( new_n548_, new_n246_ );
not g441 ( new_n549_, new_n252_ );
or g442 ( new_n550_, new_n549_, new_n548_ );
and g443 ( new_n551_, new_n472_, new_n550_, new_n474_ );
not g444 ( new_n552_, new_n551_ );
or g445 ( new_n553_, new_n477_, new_n550_ );
and g446 ( new_n554_, new_n553_, new_n552_ );
or g447 ( new_n555_, new_n235_, N92, new_n237_, new_n239_ );
and g448 ( new_n556_, new_n555_, keyIn_0_57 );
not g449 ( new_n557_, keyIn_0_57 );
not g450 ( new_n558_, new_n555_ );
and g451 ( new_n559_, new_n558_, new_n557_ );
or g452 ( new_n560_, new_n559_, new_n556_ );
or g453 ( new_n561_, new_n554_, new_n560_ );
not g454 ( new_n562_, new_n432_ );
and g455 ( new_n563_, new_n472_, new_n562_, new_n474_ );
not g456 ( new_n564_, new_n563_ );
or g457 ( new_n565_, new_n477_, new_n562_ );
and g458 ( new_n566_, new_n565_, new_n564_ );
not g459 ( new_n567_, N40 );
and g460 ( new_n568_, new_n415_, new_n567_, new_n416_, new_n421_ );
not g461 ( new_n569_, new_n568_ );
or g462 ( new_n570_, new_n566_, new_n569_ );
and g463 ( new_n571_, new_n535_, new_n547_, new_n561_, new_n570_ );
and g464 ( new_n572_, new_n571_, new_n468_, new_n505_, new_n523_ );
not g465 ( new_n573_, new_n572_ );
and g466 ( new_n574_, new_n535_, new_n547_ );
and g467 ( new_n575_, new_n561_, new_n570_ );
and g468 ( new_n576_, new_n505_, new_n523_, new_n574_, new_n575_ );
or g469 ( new_n577_, new_n576_, new_n468_ );
and g470 ( N370, new_n577_, new_n573_ );
and g471 ( new_n579_, new_n577_, N27, new_n573_ );
and g472 ( new_n580_, N329, N21 );
and g473 ( new_n581_, N223, N11 );
or g474 ( new_n582_, new_n580_, new_n204_, new_n581_ );
or g475 ( new_n583_, new_n579_, new_n582_ );
and g476 ( new_n584_, new_n577_, N40, new_n573_ );
and g477 ( new_n585_, N329, N34 );
and g478 ( new_n586_, N223, N24 );
or g479 ( new_n587_, new_n585_, new_n176_, new_n586_ );
or g480 ( new_n588_, new_n584_, new_n587_ );
and g481 ( new_n589_, new_n583_, new_n588_ );
and g482 ( new_n590_, new_n577_, N53, new_n573_ );
and g483 ( new_n591_, N329, N47 );
and g484 ( new_n592_, N223, N37 );
or g485 ( new_n593_, new_n591_, new_n188_, new_n592_ );
or g486 ( new_n594_, new_n590_, new_n593_ );
and g487 ( new_n595_, new_n577_, N66, new_n573_ );
and g488 ( new_n596_, N329, N60 );
and g489 ( new_n597_, N223, N50 );
or g490 ( new_n598_, new_n596_, new_n144_, new_n597_ );
or g491 ( new_n599_, new_n595_, new_n598_ );
and g492 ( new_n600_, new_n594_, new_n599_ );
and g493 ( new_n601_, new_n577_, N79, new_n573_ );
and g494 ( new_n602_, N329, N73 );
and g495 ( new_n603_, N223, N63 );
or g496 ( new_n604_, new_n602_, new_n163_, new_n603_ );
or g497 ( new_n605_, new_n601_, new_n604_ );
and g498 ( new_n606_, new_n577_, N92, new_n573_ );
and g499 ( new_n607_, N329, N86 );
and g500 ( new_n608_, N223, N76 );
or g501 ( new_n609_, new_n607_, new_n129_, new_n608_ );
or g502 ( new_n610_, new_n606_, new_n609_ );
and g503 ( new_n611_, new_n605_, new_n610_ );
and g504 ( new_n612_, new_n577_, N115, new_n573_ );
and g505 ( new_n613_, N329, N112 );
and g506 ( new_n614_, N223, N102 );
or g507 ( new_n615_, new_n613_, new_n264_, new_n614_ );
or g508 ( new_n616_, new_n612_, new_n615_ );
and g509 ( new_n617_, new_n577_, N105, new_n573_ );
and g510 ( new_n618_, N329, N99 );
and g511 ( new_n619_, N223, N89 );
or g512 ( new_n620_, new_n618_, new_n115_, new_n619_ );
or g513 ( new_n621_, new_n617_, new_n620_ );
and g514 ( new_n622_, new_n616_, new_n621_ );
and g515 ( new_n623_, new_n589_, new_n600_, new_n611_, new_n622_ );
not g516 ( new_n624_, new_n623_ );
and g517 ( new_n625_, new_n624_, keyIn_0_63 );
not g518 ( new_n626_, keyIn_0_63 );
and g519 ( new_n627_, new_n623_, new_n626_ );
or g520 ( new_n628_, new_n625_, new_n627_ );
and g521 ( new_n629_, N370, N14 );
and g522 ( new_n630_, N329, N8 );
and g523 ( new_n631_, N223, N1 );
or g524 ( new_n632_, new_n629_, new_n200_, new_n630_, new_n631_ );
and g525 ( N421, new_n628_, new_n632_ );
and g526 ( new_n634_, new_n589_, new_n600_ );
not g527 ( N430, new_n634_ );
not g528 ( new_n636_, new_n589_ );
not g529 ( new_n637_, new_n611_ );
and g530 ( new_n638_, new_n637_, new_n600_ );
or g531 ( N431, new_n638_, new_n636_ );
not g532 ( new_n640_, new_n583_ );
not g533 ( new_n641_, new_n594_ );
not g534 ( new_n642_, new_n617_ );
not g535 ( new_n643_, new_n620_ );
and g536 ( new_n644_, new_n610_, new_n642_, new_n643_ );
not g537 ( new_n645_, new_n601_ );
not g538 ( new_n646_, new_n604_ );
and g539 ( new_n647_, new_n599_, new_n645_, new_n646_ );
or g540 ( new_n648_, new_n644_, new_n647_, new_n641_ );
and g541 ( new_n649_, new_n648_, new_n588_ );
or g542 ( N432, new_n649_, new_n640_ );
endmodule