module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n92_, new_n79_, new_n250_, new_n113_, new_n288_, new_n371_, new_n97_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n173_, new_n220_, new_n130_, new_n419_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n214_, new_n451_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n352_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n317_, new_n102_, new_n344_, new_n143_, new_n287_, new_n125_, new_n145_, new_n253_, new_n403_, new_n90_, new_n237_, new_n234_, new_n149_, new_n472_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n133_, new_n257_, new_n212_, new_n151_, new_n364_, new_n449_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n382_, new_n272_, new_n282_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n88_, new_n360_, new_n98_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n87_, new_n387_, new_n103_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n221_, new_n385_, new_n450_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n461_, new_n459_, new_n174_, new_n297_, new_n361_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n105_, new_n340_, new_n147_, new_n285_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n325_, new_n417_, new_n180_, new_n332_, new_n318_, new_n453_, new_n163_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n111_, new_n158_, new_n252_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n274_, new_n372_, new_n100_, new_n242_, new_n218_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n470_, new_n423_, new_n205_, new_n213_, new_n134_, new_n141_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n432_, new_n265_, new_n370_, new_n256_, new_n278_, new_n304_, new_n381_, new_n388_, new_n217_, new_n101_, new_n269_, new_n194_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n327_, new_n216_, new_n431_, new_n77_, new_n196_, new_n280_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n338_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n465_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n277_, new_n245_, new_n402_, new_n474_, new_n89_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n289_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n96_, new_n178_, new_n437_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n406_, new_n356_, new_n333_, new_n229_, new_n290_, new_n464_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n76_, N17 );
or g001 ( new_n77_, keyIn_0_0, N11 );
and g002 ( new_n78_, keyIn_0_0, N11 );
not g003 ( new_n79_, new_n78_ );
and g004 ( new_n80_, new_n79_, new_n77_ );
or g005 ( new_n81_, new_n80_, new_n76_ );
and g006 ( new_n82_, new_n81_, keyIn_0_3 );
not g007 ( new_n83_, keyIn_0_3 );
not g008 ( new_n84_, new_n77_ );
or g009 ( new_n85_, new_n84_, new_n78_ );
and g010 ( new_n86_, new_n85_, new_n83_, N17 );
or g011 ( new_n87_, new_n82_, new_n86_ );
not g012 ( new_n88_, N82 );
or g013 ( new_n89_, new_n88_, N76 );
not g014 ( new_n90_, N30 );
or g015 ( new_n91_, new_n90_, N24 );
and g016 ( new_n92_, new_n89_, new_n91_ );
not g017 ( new_n93_, N1 );
and g018 ( new_n94_, new_n93_, N4 );
not g019 ( new_n95_, new_n94_ );
not g020 ( new_n96_, N50 );
and g021 ( new_n97_, new_n96_, N56 );
not g022 ( new_n98_, new_n97_ );
not g023 ( new_n99_, N43 );
or g024 ( new_n100_, new_n99_, N37 );
not g025 ( new_n101_, N108 );
or g026 ( new_n102_, new_n101_, N102 );
and g027 ( new_n103_, new_n100_, new_n102_ );
and g028 ( new_n104_, new_n92_, new_n103_, new_n95_, new_n98_ );
not g029 ( new_n105_, N89 );
or g030 ( new_n106_, new_n105_, keyIn_0_2 );
not g031 ( new_n107_, keyIn_0_2 );
or g032 ( new_n108_, new_n107_, N89 );
and g033 ( new_n109_, new_n106_, new_n108_, N95 );
or g034 ( new_n110_, new_n109_, keyIn_0_5 );
not g035 ( new_n111_, keyIn_0_5 );
not g036 ( new_n112_, N95 );
not g037 ( new_n113_, new_n106_ );
and g038 ( new_n114_, new_n105_, keyIn_0_2 );
or g039 ( new_n115_, new_n113_, new_n114_, new_n111_, new_n112_ );
and g040 ( new_n116_, new_n110_, new_n115_ );
not g041 ( new_n117_, new_n116_ );
not g042 ( new_n118_, keyIn_0_1 );
not g043 ( new_n119_, N63 );
and g044 ( new_n120_, new_n118_, new_n119_ );
and g045 ( new_n121_, keyIn_0_1, N63 );
or g046 ( new_n122_, new_n120_, new_n121_ );
and g047 ( new_n123_, new_n122_, N69 );
or g048 ( new_n124_, new_n123_, keyIn_0_4 );
not g049 ( new_n125_, keyIn_0_4 );
not g050 ( new_n126_, N69 );
or g051 ( new_n127_, keyIn_0_1, N63 );
not g052 ( new_n128_, new_n121_ );
and g053 ( new_n129_, new_n128_, new_n127_ );
or g054 ( new_n130_, new_n129_, new_n125_, new_n126_ );
and g055 ( new_n131_, new_n124_, new_n130_ );
and g056 ( new_n132_, new_n87_, new_n131_, new_n104_, new_n117_ );
or g057 ( new_n133_, new_n132_, keyIn_0_6 );
not g058 ( new_n134_, keyIn_0_6 );
and g059 ( new_n135_, new_n85_, N17 );
or g060 ( new_n136_, new_n135_, new_n83_ );
not g061 ( new_n137_, new_n86_ );
and g062 ( new_n138_, new_n136_, new_n137_ );
not g063 ( new_n139_, new_n104_ );
or g064 ( new_n140_, new_n129_, new_n126_ );
and g065 ( new_n141_, new_n140_, new_n125_ );
not g066 ( new_n142_, new_n130_ );
or g067 ( new_n143_, new_n116_, new_n141_, new_n142_ );
or g068 ( new_n144_, new_n143_, new_n138_, new_n134_, new_n139_ );
and g069 ( new_n145_, new_n133_, new_n144_ );
not g070 ( N223, new_n145_ );
not g071 ( new_n147_, keyIn_0_12 );
or g072 ( new_n148_, new_n145_, keyIn_0_7 );
and g073 ( new_n149_, new_n133_, keyIn_0_7, new_n144_ );
not g074 ( new_n150_, new_n149_ );
and g075 ( new_n151_, new_n148_, new_n150_ );
or g076 ( new_n152_, new_n151_, new_n116_ );
and g077 ( new_n153_, new_n148_, new_n116_, new_n150_ );
not g078 ( new_n154_, new_n153_ );
and g079 ( new_n155_, new_n152_, new_n154_ );
or g080 ( new_n156_, new_n155_, keyIn_0_10 );
and g081 ( new_n157_, new_n152_, keyIn_0_10, new_n154_ );
not g082 ( new_n158_, new_n157_ );
and g083 ( new_n159_, new_n156_, new_n158_ );
or g084 ( new_n160_, new_n159_, new_n112_, N99 );
and g085 ( new_n161_, new_n160_, new_n147_ );
not g086 ( new_n162_, new_n161_ );
not g087 ( new_n163_, N99 );
not g088 ( new_n164_, new_n159_ );
and g089 ( new_n165_, new_n164_, keyIn_0_12, N95, new_n163_ );
not g090 ( new_n166_, new_n165_ );
not g091 ( new_n167_, keyIn_0_11 );
or g092 ( new_n168_, new_n151_, new_n94_ );
and g093 ( new_n169_, new_n148_, new_n94_, new_n150_ );
not g094 ( new_n170_, new_n169_ );
and g095 ( new_n171_, new_n168_, new_n170_ );
or g096 ( new_n172_, new_n171_, keyIn_0_8 );
and g097 ( new_n173_, new_n168_, keyIn_0_8, new_n170_ );
not g098 ( new_n174_, new_n173_ );
and g099 ( new_n175_, new_n172_, new_n174_ );
not g100 ( new_n176_, N4 );
or g101 ( new_n177_, new_n176_, N8 );
or g102 ( new_n178_, new_n175_, new_n177_ );
and g103 ( new_n179_, new_n178_, new_n167_ );
not g104 ( new_n180_, N8 );
not g105 ( new_n181_, new_n175_ );
and g106 ( new_n182_, new_n181_, keyIn_0_11, N4, new_n180_ );
or g107 ( new_n183_, new_n179_, new_n182_ );
not g108 ( new_n184_, N21 );
or g109 ( new_n185_, new_n151_, new_n138_ );
and g110 ( new_n186_, new_n151_, new_n138_ );
not g111 ( new_n187_, new_n186_ );
and g112 ( new_n188_, new_n187_, keyIn_0_9, new_n185_ );
not g113 ( new_n189_, new_n188_ );
and g114 ( new_n190_, new_n187_, new_n185_ );
or g115 ( new_n191_, new_n190_, keyIn_0_9 );
and g116 ( new_n192_, new_n191_, N17, new_n184_, new_n189_ );
not g117 ( new_n193_, new_n192_ );
not g118 ( new_n194_, new_n91_ );
or g119 ( new_n195_, new_n151_, new_n194_ );
and g120 ( new_n196_, new_n151_, new_n194_ );
not g121 ( new_n197_, new_n196_ );
and g122 ( new_n198_, new_n197_, new_n195_ );
or g123 ( new_n199_, new_n198_, new_n90_ );
or g124 ( new_n200_, new_n199_, N34 );
not g125 ( new_n201_, new_n100_ );
or g126 ( new_n202_, new_n151_, new_n201_ );
and g127 ( new_n203_, new_n151_, new_n201_ );
not g128 ( new_n204_, new_n203_ );
and g129 ( new_n205_, new_n204_, new_n202_ );
or g130 ( new_n206_, new_n205_, new_n99_ );
or g131 ( new_n207_, new_n206_, N47 );
and g132 ( new_n208_, new_n200_, new_n207_ );
not g133 ( new_n209_, new_n89_ );
or g134 ( new_n210_, new_n151_, new_n209_ );
and g135 ( new_n211_, new_n151_, new_n209_ );
not g136 ( new_n212_, new_n211_ );
and g137 ( new_n213_, new_n212_, new_n210_ );
or g138 ( new_n214_, new_n213_, new_n88_, N86 );
not g139 ( new_n215_, N56 );
or g140 ( new_n216_, new_n151_, new_n97_ );
and g141 ( new_n217_, new_n151_, new_n97_ );
not g142 ( new_n218_, new_n217_ );
and g143 ( new_n219_, new_n218_, new_n216_ );
or g144 ( new_n220_, new_n219_, new_n215_, N60 );
not g145 ( new_n221_, new_n131_ );
or g146 ( new_n222_, new_n151_, new_n221_ );
and g147 ( new_n223_, new_n151_, new_n221_ );
not g148 ( new_n224_, new_n223_ );
and g149 ( new_n225_, new_n224_, new_n222_ );
or g150 ( new_n226_, new_n225_, new_n126_, N73 );
not g151 ( new_n227_, new_n102_ );
or g152 ( new_n228_, new_n151_, new_n227_ );
and g153 ( new_n229_, new_n151_, new_n227_ );
not g154 ( new_n230_, new_n229_ );
and g155 ( new_n231_, new_n230_, new_n228_ );
or g156 ( new_n232_, new_n231_, new_n101_, N112 );
and g157 ( new_n233_, new_n214_, new_n220_, new_n232_, new_n226_ );
and g158 ( new_n234_, new_n208_, new_n193_, new_n233_ );
and g159 ( new_n235_, new_n183_, new_n162_, new_n166_, new_n234_ );
or g160 ( new_n236_, new_n235_, keyIn_0_13 );
not g161 ( new_n237_, keyIn_0_13 );
or g162 ( new_n238_, new_n161_, new_n165_ );
not g163 ( new_n239_, new_n183_ );
not g164 ( new_n240_, new_n234_ );
or g165 ( new_n241_, new_n239_, new_n238_, new_n237_, new_n240_ );
and g166 ( new_n242_, new_n236_, new_n241_ );
not g167 ( N329, new_n242_ );
not g168 ( new_n244_, keyIn_0_19 );
not g169 ( new_n245_, new_n220_ );
not g170 ( new_n246_, keyIn_0_15 );
or g171 ( new_n247_, new_n242_, new_n246_ );
and g172 ( new_n248_, new_n236_, new_n246_, new_n241_ );
not g173 ( new_n249_, new_n248_ );
and g174 ( new_n250_, new_n247_, new_n249_ );
or g175 ( new_n251_, new_n250_, new_n245_ );
and g176 ( new_n252_, new_n247_, new_n245_, new_n249_ );
not g177 ( new_n253_, new_n252_ );
and g178 ( new_n254_, new_n251_, new_n253_ );
or g179 ( new_n255_, new_n254_, keyIn_0_17 );
and g180 ( new_n256_, new_n251_, keyIn_0_17, new_n253_ );
not g181 ( new_n257_, new_n256_ );
and g182 ( new_n258_, new_n255_, new_n257_ );
or g183 ( new_n259_, new_n219_, new_n215_ );
or g184 ( new_n260_, new_n259_, N66 );
or g185 ( new_n261_, new_n258_, new_n260_ );
and g186 ( new_n262_, new_n261_, new_n244_ );
not g187 ( new_n263_, new_n258_ );
not g188 ( new_n264_, new_n260_ );
and g189 ( new_n265_, new_n263_, keyIn_0_19, new_n264_ );
or g190 ( new_n266_, new_n262_, new_n265_ );
not g191 ( new_n267_, keyIn_0_16 );
or g192 ( new_n268_, new_n250_, new_n239_ );
and g193 ( new_n269_, new_n247_, new_n239_, new_n249_ );
not g194 ( new_n270_, new_n269_ );
and g195 ( new_n271_, new_n268_, new_n267_, new_n270_ );
not g196 ( new_n272_, new_n271_ );
not g197 ( new_n273_, keyIn_0_14 );
or g198 ( new_n274_, new_n175_, new_n176_, N14 );
and g199 ( new_n275_, new_n274_, new_n273_ );
not g200 ( new_n276_, new_n274_ );
and g201 ( new_n277_, new_n276_, keyIn_0_14 );
or g202 ( new_n278_, new_n277_, new_n275_ );
and g203 ( new_n279_, new_n268_, new_n270_ );
or g204 ( new_n280_, new_n279_, new_n267_ );
and g205 ( new_n281_, new_n280_, new_n272_, new_n278_ );
or g206 ( new_n282_, new_n281_, keyIn_0_18 );
and g207 ( new_n283_, new_n280_, keyIn_0_18, new_n272_, new_n278_ );
not g208 ( new_n284_, new_n283_ );
and g209 ( new_n285_, new_n282_, new_n284_ );
not g210 ( new_n286_, new_n285_ );
or g211 ( new_n287_, new_n213_, new_n88_ );
not g212 ( new_n288_, new_n214_ );
or g213 ( new_n289_, new_n250_, new_n288_ );
and g214 ( new_n290_, new_n250_, new_n288_ );
not g215 ( new_n291_, new_n290_ );
and g216 ( new_n292_, new_n291_, new_n289_ );
or g217 ( new_n293_, new_n292_, N92, new_n287_ );
and g218 ( new_n294_, new_n191_, N17, new_n189_ );
not g219 ( new_n295_, new_n294_ );
or g220 ( new_n296_, new_n250_, new_n192_ );
and g221 ( new_n297_, new_n250_, new_n192_ );
not g222 ( new_n298_, new_n297_ );
and g223 ( new_n299_, new_n298_, new_n296_ );
or g224 ( new_n300_, new_n299_, N27, new_n295_ );
not g225 ( new_n301_, new_n200_ );
or g226 ( new_n302_, new_n250_, new_n301_ );
and g227 ( new_n303_, new_n250_, new_n301_ );
not g228 ( new_n304_, new_n303_ );
and g229 ( new_n305_, new_n304_, new_n302_ );
or g230 ( new_n306_, new_n305_, N40, new_n199_ );
and g231 ( new_n307_, new_n293_, new_n306_, new_n300_ );
not g232 ( new_n308_, new_n232_ );
or g233 ( new_n309_, new_n250_, new_n308_ );
and g234 ( new_n310_, new_n250_, new_n308_ );
not g235 ( new_n311_, new_n310_ );
and g236 ( new_n312_, new_n311_, new_n309_ );
or g237 ( new_n313_, new_n312_, new_n101_, N115, new_n231_ );
or g238 ( new_n314_, new_n225_, new_n126_ );
not g239 ( new_n315_, new_n226_ );
or g240 ( new_n316_, new_n250_, new_n315_ );
and g241 ( new_n317_, new_n250_, new_n315_ );
not g242 ( new_n318_, new_n317_ );
and g243 ( new_n319_, new_n318_, new_n316_ );
or g244 ( new_n320_, new_n319_, N79, new_n314_ );
and g245 ( new_n321_, new_n313_, new_n320_ );
not g246 ( new_n322_, new_n207_ );
or g247 ( new_n323_, new_n250_, new_n322_ );
and g248 ( new_n324_, new_n250_, new_n322_ );
not g249 ( new_n325_, new_n324_ );
and g250 ( new_n326_, new_n325_, new_n323_ );
or g251 ( new_n327_, new_n326_, N53, new_n206_ );
or g252 ( new_n328_, new_n159_, new_n112_ );
or g253 ( new_n329_, new_n250_, new_n238_ );
and g254 ( new_n330_, new_n250_, new_n238_ );
not g255 ( new_n331_, new_n330_ );
and g256 ( new_n332_, new_n331_, new_n329_ );
or g257 ( new_n333_, new_n332_, N105, new_n328_ );
and g258 ( new_n334_, new_n327_, new_n333_ );
and g259 ( new_n335_, new_n321_, new_n307_, new_n334_ );
and g260 ( new_n336_, new_n266_, new_n286_, new_n335_ );
or g261 ( new_n337_, new_n336_, keyIn_0_20 );
not g262 ( new_n338_, keyIn_0_20 );
not g263 ( new_n339_, new_n262_ );
not g264 ( new_n340_, new_n265_ );
and g265 ( new_n341_, new_n339_, new_n340_ );
not g266 ( new_n342_, new_n335_ );
or g267 ( new_n343_, new_n341_, new_n338_, new_n285_, new_n342_ );
and g268 ( new_n344_, new_n337_, new_n343_ );
not g269 ( N370, new_n344_ );
not g270 ( new_n346_, keyIn_0_25 );
or g271 ( new_n347_, new_n344_, keyIn_0_21 );
not g272 ( new_n348_, keyIn_0_21 );
not g273 ( new_n349_, new_n336_ );
and g274 ( new_n350_, new_n349_, new_n338_ );
not g275 ( new_n351_, new_n343_ );
or g276 ( new_n352_, new_n350_, new_n351_, new_n348_ );
and g277 ( new_n353_, new_n347_, new_n352_ );
not g278 ( new_n354_, new_n353_ );
and g279 ( new_n355_, new_n354_, keyIn_0_23, N53 );
not g280 ( new_n356_, keyIn_0_23 );
not g281 ( new_n357_, N53 );
or g282 ( new_n358_, new_n353_, new_n357_ );
and g283 ( new_n359_, new_n358_, new_n356_ );
and g284 ( new_n360_, N329, N47 );
and g285 ( new_n361_, N223, N37 );
or g286 ( new_n362_, new_n360_, new_n99_, new_n361_ );
or g287 ( new_n363_, new_n359_, new_n355_, new_n362_ );
and g288 ( new_n364_, new_n363_, new_n346_ );
not g289 ( new_n365_, new_n355_ );
not g290 ( new_n366_, new_n359_ );
not g291 ( new_n367_, new_n362_ );
and g292 ( new_n368_, new_n366_, keyIn_0_25, new_n365_, new_n367_ );
or g293 ( new_n369_, new_n364_, new_n368_ );
and g294 ( new_n370_, new_n354_, N66 );
and g295 ( new_n371_, N329, N60 );
and g296 ( new_n372_, N223, N50 );
or g297 ( new_n373_, new_n370_, new_n215_, new_n371_, new_n372_ );
and g298 ( new_n374_, new_n369_, new_n373_ );
not g299 ( new_n375_, keyIn_0_22 );
not g300 ( new_n376_, N40 );
or g301 ( new_n377_, new_n353_, new_n376_ );
or g302 ( new_n378_, new_n377_, new_n375_ );
and g303 ( new_n379_, new_n377_, new_n375_ );
not g304 ( new_n380_, new_n379_ );
and g305 ( new_n381_, N329, N34 );
and g306 ( new_n382_, N223, N24 );
or g307 ( new_n383_, new_n381_, new_n90_, new_n382_ );
not g308 ( new_n384_, new_n383_ );
and g309 ( new_n385_, new_n380_, new_n378_, new_n384_ );
or g310 ( new_n386_, new_n385_, keyIn_0_24 );
not g311 ( new_n387_, keyIn_0_24 );
and g312 ( new_n388_, new_n354_, N40 );
and g313 ( new_n389_, new_n388_, keyIn_0_22 );
or g314 ( new_n390_, new_n389_, new_n379_, new_n387_, new_n383_ );
and g315 ( new_n391_, new_n386_, new_n390_ );
not g316 ( new_n392_, new_n391_ );
and g317 ( new_n393_, new_n354_, N27 );
and g318 ( new_n394_, N329, N21 );
and g319 ( new_n395_, N223, N11 );
or g320 ( new_n396_, new_n393_, new_n76_, new_n394_, new_n395_ );
not g321 ( new_n397_, new_n396_ );
or g322 ( new_n398_, new_n392_, new_n397_ );
not g323 ( new_n399_, new_n398_ );
and g324 ( new_n400_, new_n354_, N92 );
and g325 ( new_n401_, N329, N86 );
and g326 ( new_n402_, N223, N76 );
or g327 ( new_n403_, new_n400_, new_n88_, new_n401_, new_n402_ );
and g328 ( new_n404_, new_n354_, N115 );
and g329 ( new_n405_, N329, N112 );
and g330 ( new_n406_, N223, N102 );
or g331 ( new_n407_, new_n404_, new_n101_, new_n405_, new_n406_ );
and g332 ( new_n408_, new_n354_, N105 );
and g333 ( new_n409_, N329, N99 );
and g334 ( new_n410_, N223, N89 );
or g335 ( new_n411_, new_n408_, new_n112_, new_n409_, new_n410_ );
and g336 ( new_n412_, new_n354_, N79 );
not g337 ( new_n413_, new_n412_ );
and g338 ( new_n414_, N329, N73 );
not g339 ( new_n415_, new_n414_ );
and g340 ( new_n416_, N223, N63 );
not g341 ( new_n417_, new_n416_ );
and g342 ( new_n418_, new_n413_, N69, new_n415_, new_n417_ );
not g343 ( new_n419_, new_n418_ );
and g344 ( new_n420_, new_n419_, new_n403_, new_n407_, new_n411_ );
and g345 ( new_n421_, new_n399_, new_n374_, new_n420_ );
not g346 ( new_n422_, new_n421_ );
and g347 ( new_n423_, new_n354_, N14 );
and g348 ( new_n424_, N329, N8 );
and g349 ( new_n425_, N223, N1 );
or g350 ( new_n426_, new_n423_, new_n176_, new_n424_, new_n425_ );
and g351 ( N421, new_n422_, new_n426_ );
not g352 ( new_n428_, keyIn_0_30 );
not g353 ( new_n429_, keyIn_0_26 );
and g354 ( new_n430_, new_n366_, new_n365_, new_n367_ );
or g355 ( new_n431_, new_n430_, keyIn_0_25 );
not g356 ( new_n432_, new_n368_ );
and g357 ( new_n433_, new_n431_, new_n432_ );
or g358 ( new_n434_, new_n433_, new_n429_ );
and g359 ( new_n435_, new_n431_, new_n429_, new_n432_ );
not g360 ( new_n436_, new_n435_ );
and g361 ( new_n437_, new_n434_, new_n436_ );
or g362 ( new_n438_, new_n437_, keyIn_0_27, new_n392_ );
not g363 ( new_n439_, new_n438_ );
or g364 ( new_n440_, new_n437_, new_n392_ );
and g365 ( new_n441_, new_n440_, keyIn_0_27 );
and g366 ( new_n442_, new_n399_, new_n373_ );
not g367 ( new_n443_, new_n442_ );
or g368 ( new_n444_, new_n441_, new_n439_, new_n443_ );
and g369 ( new_n445_, new_n444_, new_n428_ );
not g370 ( new_n446_, keyIn_0_27 );
and g371 ( new_n447_, new_n369_, keyIn_0_26 );
or g372 ( new_n448_, new_n447_, new_n435_ );
and g373 ( new_n449_, new_n448_, new_n391_ );
or g374 ( new_n450_, new_n449_, new_n446_ );
and g375 ( new_n451_, new_n450_, keyIn_0_30, new_n438_, new_n442_ );
or g376 ( N430, new_n445_, new_n451_ );
not g377 ( new_n453_, keyIn_0_28 );
and g378 ( new_n454_, new_n391_, new_n369_, new_n373_, new_n418_ );
or g379 ( new_n455_, new_n454_, new_n453_ );
and g380 ( new_n456_, new_n454_, new_n453_ );
not g381 ( new_n457_, new_n456_ );
and g382 ( new_n458_, new_n457_, new_n455_ );
not g383 ( new_n459_, new_n458_ );
not g384 ( new_n460_, new_n403_ );
and g385 ( new_n461_, new_n374_, new_n460_ );
or g386 ( N431, new_n459_, new_n398_, new_n461_ );
not g387 ( new_n463_, keyIn_0_29 );
not g388 ( new_n464_, new_n411_ );
and g389 ( new_n465_, new_n464_, new_n403_ );
and g390 ( new_n466_, new_n391_, new_n463_, new_n369_, new_n465_ );
not g391 ( new_n467_, new_n466_ );
and g392 ( new_n468_, new_n391_, new_n369_, new_n465_ );
or g393 ( new_n469_, new_n468_, new_n463_ );
and g394 ( new_n470_, new_n469_, new_n396_, new_n467_ );
and g395 ( new_n471_, new_n450_, new_n438_, new_n458_, new_n470_ );
or g396 ( new_n472_, new_n471_, keyIn_0_31 );
and g397 ( new_n473_, new_n471_, keyIn_0_31 );
not g398 ( new_n474_, new_n473_ );
and g399 ( N432, new_n474_, new_n472_ );
endmodule