module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g4556, g1289, g8943, g1882, n1663, g255,
         g312, g11257, g452, g7032, g123, g6830, g207, g8920, g713, g4340,
         g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695, g11372, g461,
         n1594, g8260, g940, n1712, g11391, g976, g8432, g709, g6088, g1092,
         g6478, g1574, g6795, g1864, g11320, g369, g6500, g1580, g5392, g1736,
         n1637, g10782, n3065, g6216, g1424, g1737, g10858, g1672, g5914,
         g1077, g7590, g1231, g6656, g4, g6728, g5126, g1104, n1658, g7290,
         g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064, g8019, g6545,
         g1543, g256, g315, g6533, g1534, g8820, g622, n1713, g8941, g1927,
         g10859, g1660, g6922, g278, g8772, g1436, g8433, g718, g6526, n1669,
         g10793, g554, g11333, g496, g11392, g981, n1720, g794, g829, n1651,
         g6093, g1095, g8889, g704, g7302, g1265, g6525, g1786, g8429, g682,
         g7292, g1296, g6621, n1668, g7134, n3062, g260, g327, g6333, g1389,
         n1603, g6826, g1371, g1955, g1956, g10860, g1675, g11483, g354, g6392,
         g113, g7626, g639, n1692, g10866, g1684, g8193, g1639, g6983, g1791,
         n1702, g6839, g248, n1598, g4076, g1707, g4293, g1759, g11482, g351,
         g6507, g1604, g6096, g1098, g8250, g932, n1591, g8282, g1896, g8435,
         g736, g6924, g1019, g6819, n3061, g746, g745, g6244, g1419, n1602,
         g6627, n1667, g32, n1865, g6071, g1086, g8046, g1486, g10707, g1730,
         g6198, g1504, g8051, g1470, g8024, g822, g10862, g1678, g8050, g174,
         g7133, g1766, g7930, g1801, g6832, g186, g11308, g959, g6918, g8769,
         g1407, g6909, g1868, g4940, g5404, g1718, n1611, g11265, g396, g6930,
         g1015, g10726, n1650, g4891, n3059, g6224, g1415, g7586, g1227,
         g10770, g1721, n3058, DFF_121_n1, n3057, g6934, g284, g11256, g426,
         g6824, g219, g1360, n3056, DFF_126_n1, g6126, g806, g8767, g1428,
         g6546, g1564, g4238, g1741, g6823, g225, g6928, g281, g11602, g1308,
         g9721, g611, n1609, g4890, n3055, DFF_136_n1, n1586, g1217, g6524,
         g1589, g8045, g1466, g6469, g1571, g6471, g1861, g6821, n3054, g11514,
         g1448, g4480, g1133, n1706, g11610, g1333, g7843, g153, g11310, g962,
         g5536, g11331, g486, n1621, g11380, g471, n1606, g6838, g1397, n1711,
         g8288, g1950, g755, g756, g4892, n3053, DFF_157_n1, g10855, g1101,
         g549, g10898, g105, g10865, g1669, g6822, g6528, g1531, g6180, g1458,
         n1703, g10718, g572, g6912, g1011, n3051, g6234, g1411, g6099, g1074,
         g11259, g444, g8039, g1474, g6059, g1080, g5396, g1713, n1610, g262,
         g333, g6906, g269, g11266, g401, g11294, g1857, n1682, g5421, g9,
         g8649, g664, g11312, g965, g6840, g1400, n1629, g254, g309, g7202,
         g814, g6834, g231, g10795, g557, g875, g869, g6831, g1383, g8060,
         g158, g4893, g627, n1701, g7244, g1023, g6026, g259, n3050,
         DFF_194_n1, g11608, g1327, g7660, g654, g6911, g293, g11640, g1346,
         g8777, g1633, g4274, g1753, g1508, n1707, g7297, g1240, g11326, g538,
         g11269, g416, g11325, g542, g10864, g1681, g11290, g374, g10798, g563,
         g8284, g1914, g11328, g530, g10800, g575, g8944, g1936, n1694, g7183,
         n1674, g4465, g1356, g1317, g11484, g357, g11263, g386, g6501, g1601,
         g6757, g166, g11334, g501, n1690, g6042, g8384, g1840, g6653, n1666,
         g257, g318, g5763, g5849, n3048, g6929, g302, g11488, g342, g7299,
         g1250, g4330, g1163, g1958, n3047, g7257, g1032, g8775, g1432, g5770,
         g1453, n1628, g11486, g363, g261, g330, g4338, g1157, g4500, n3046,
         n3045, DFF_242_n1, g8147, g928, n1604, g6038, g11337, g516, n1620,
         g6045, g7191, g826, g861, g8774, g1627, g7293, g1292, g6907, g290,
         g4903, n3044, g6123, g6506, g1583, g11376, g466, n1646, g6542, g1561,
         g6551, g1546, g6901, g287, g10797, g560, g8505, g617, n1645, n1631,
         g11647, g336, g11340, g456, n1641, g253, g305, n1681, g11625, g345,
         g636, g8, g6502, N599, g6049, g8945, g1945, n1697, g4231, g1738,
         g8040, g1478, n3042, DFF_275_n1, g6155, g1690, n1653, g8043, g1482,
         g5173, g1110, n1677, g6916, g296, g10861, g1663, g8431, g700, g4309,
         g1762, g11485, g360, g6334, g192, g10767, g1657, g8923, g722, n1693,
         g7189, n1673, g10799, g566, g6747, n3041, g6080, g1089, g3381, g5910,
         g1071, g11393, g986, n1722, g11349, g971, g6439, g143, g9266, g1814,
         n1608, g1212, g8940, g1918, g7705, g9269, g1822, n1643, g6820, g237,
         g8042, g1462, g6759, g178, g11487, g366, g802, g837, g9124, g599,
         n1644, g11293, g1854, g11298, g944, g8287, g1941, g8047, g170, g6205,
         g1520, n1710, g8885, g686, n1676, g11305, g953, g5556, n3040, g2478,
         g1765, g10711, g1733, g7303, g5194, g1610, g7541, g1796, n1626,
         g11607, g1324, g6541, g1540, g6827, n3038, g11332, g491, n1691, g4902,
         n3037, DFF_330_n1, g6828, g213, g6516, g1781, n1659, g8938, g1900,
         n1675, g7298, g1245, n3036, g6672, n3035, DFF_336_n1, g8048, g148,
         g798, g833, g8285, g1923, g8254, g936, n1630, g11604, g1314, g849,
         g11636, g1336, g6910, g272, g8173, g1806, g8245, n1716, g8281, g1887,
         n3034, g11314, g968, g4905, n3033, g4484, g1137, n1597, g8937, g1891,
         n1657, g7300, g1255, g6002, n1588, g874, g9110, g591, n1607, g8926,
         g731, n1696, g8631, g7632, g1218, g9150, g605, n1593, g6531, n1665,
         g6786, g182, g11303, g950, g4477, g1129, n1705, g857, g11258, g448,
         g9272, g1828, n1605, g10773, g1727, g6470, g1592, g5083, g1703, g8286,
         g1932, g8773, g1624, g6054, g11260, g440, g11338, g476, n1599, g5918,
         g119, n1613, g8922, g668, n1662, g8049, g139, g4342, g1149, n1685,
         n3031, g6755, n3030, DFF_385_n1, g6897, g263, g7709, g818, g4255,
         g1747, g5543, n1622, g6915, g275, g6513, g1524, g6480, g1577, g6733,
         g810, g11264, g391, g8973, g658, n1615, g6833, g1386, g5996, n1587,
         g4473, g1125, n1708, g5755, g201, n1619, g7295, g1280, n1862, g6068,
         g1083, g7137, g650, g8779, g1636, g853, g11270, g421, g5529, g11306,
         g956, g11291, g378, g4283, g1756, g841, g6894, g1027, g6902, g1003,
         g8765, g1403, g4498, g1145, n1617, g5148, g1107, n1614, g7581, g1223,
         g11267, g406, g10936, g1811, g10784, n3029, g10765, g1654, g6332,
         g197, n1678, g6479, g1595, g6537, g1537, g8434, g727, g6908, g6243,
         n1717, g11324, g481, g3462, n1647, g11609, g1330, g845, g8244, g8194,
         g1512, n3027, DFF_436_n1, g8052, g1490, g4325, g1166, g11481, g348,
         n3026, DFF_441_n1, g7301, g1260, g6035, g8059, g131, n3025, g6015,
         g258, g11330, g521, n1698, g11605, g1318, g8921, g1872, n1616, g8883,
         g677, n1656, n3024, DFF_452_n1, g6523, g1549, g11300, g947, g9555,
         g1834, n1655, g6481, g1598, g4471, g1121, n1618, g11606, g1321,
         g11335, g506, n1600, g10791, g546, g8939, g1909, g6529, g1552, g10776,
         g1687, g6514, g1586, g324, g4490, g1141, n1660, g11639, g1341, g4089,
         g1710, g10785, n3023, g6179, n3022, g8053, g135, g11329, g525, n1695,
         g6515, g1607, g321, g7204, n1672, g11443, g1275, g11603, g8770, g1615,
         g11292, g382, n3020, g6900, g266, g7294, g1284, n1864, g6829, n3019,
         g8428, g673, g4904, n3018, DFF_489_n1, g8054, g162, g11268, g411,
         g11262, g431, n1876, g8283, g1905, g6193, g1515, n1627, g8776, g1630,
         g7143, n1671, g6898, g991, n1871, g7291, g1300, g11478, g339, g6000,
         g4264, g1750, g8768, g1440, g10863, g1666, g6522, g1528, g11641,
         g1351, n1721, g10780, n3017, g8044, g127, n1704, g11579, g1618, g7296,
         g1235, g6923, g299, g11261, g435, n1878, g6638, n1664, g6534, g1555,
         g6895, g995, g8771, g1621, g4506, n3016, g7441, g643, n1612, g8055,
         g1494, g6468, g1567, g8430, g691, g11327, g534, g6508, g1776, n1715,
         g10717, g569, g4334, g1160, n1585, g6679, g1, g11336, g511, g10771,
         g1724, g5445, g12, g8559, g1878, g7219, g5390, n1654, n1512, n1574,
         n1486, n1485, n1544, n1545, n1548, n1530, n1420, n1855, n1472, n1566,
         n1567, n1479, n1858, n1546, n1478, n968, n1137, n1195, n1404, n1229,
         n1262, n1227, n1450, n916, n822, n958, n918, n1054, n1159, n812,
         n1057, n1056, n817, n929, n837, n804, n1016, n1380, n926, n1391,
         n1564, n1231, n1226, n1232, n1260, n1132, n1107, n1154, n1155, n1093,
         n1214, n931, n962, n902, n1193, n1153, n1125, n1099, n917, n857, n806,
         n808, n1097, n1123, n1151, n1090, n1161, n1162, n967, n921, n898,
         n1055, n938, n1150, n1096, n1098, n1213, n1152, n836, n838, Tg1_OUT1,
         Tg1_OUT2, Tg1_OUT3, Tg1_OUT4, Tg1_OUT5, Tg1_OUT6, Tg1_OUT7, Tg1_OUT8,
         Tg2_OUT1, Tg2_OUT2, Tg2_OUT3, Tg2_OUT4, Tg2_OUT5, Tg2_OUT6, Tg2_OUT7,
         Tg2_OUT8, test_se_NOT, Trigger_select, n2, n11, n14, n16, n17, n19,
         n22, n25, n32, n33, n38, n39, n40, n42, n44, n68, n114, n177, n263,
         n280, n367, n374, n382, n387, n2071, n2072, n2073, n2074, n2079,
         n2085, n2094, n2095, n2102, n2103, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2125, n2129, n2130, n2132, n2133, n2134, n2137,
         n2139, n2141, n2143, n2144, n2147, n2154, n2160, n2175, n2195, n2196,
         n2201, n2203, n2221, n2222, n2225, n2226, n2227, n2228, n2229, n2232,
         n2233, n2237, n2240, n2241, n2242, n2243, n2246, n2247, n2248, n2249,
         n2250, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2300, n2301, n2302, n2304, n2306, n2308, n2309, n2310,
         n2311, n2314, n2315, n2316, n2317, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2334, n2336, n2337, n2338, n2339, n2340, n2341,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3021, n3028, n3032, n3039, n3043, n3049, n3052,
         n3060, n3063, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         U1586_n1, U1754_n1, U1798_n1, U1839_n1, U1843_n1, U1877_n1, U1908_n1,
         U1909_n1, U1987_n1, U2031_n1, U2035_n1, U2418_n1, U2468_n1, U2478_n1,
         U2488_n1, U2533_n1, U2534_n1, U2639_n1, U2641_n1, U2654_n1, U2658_n1,
         U2683_n1, U2699_n1, U2846_n1, U2847_n1, U2848_n1, U2859_n1, U2860_n1,
         U2861_n1, U2867_n1, U2879_n1, U2881_n1, U2882_n1, U2883_n1, U2884_n1,
         U2885_n1, U2886_n1, U2887_n1, U2888_n1, U2889_n1, U2890_n1, U2891_n1,
         U2892_n1, U2893_n1, U2894_n1, U2895_n1, U2896_n1, U2897_n1, U2898_n1,
         U2899_n1, U2900_n1, U2901_n1, U2902_n1, U3090_n1, U3092_n1, U3094_n1,
         U3096_n1, U3098_n1, U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(g4556), .SI(test_si1), .SE(n2451), .CLK(n2491), .Q(
        g1289), .QN(n2348) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n2432), .CLK(n2500), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n2427), .CLK(n2502), .Q(g312), 
        .QN(n2289) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n2424), .CLK(n2504), .Q(g452) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n2397), .CLK(n2517), .Q(g123)
         );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n2397), .CLK(n2518), .Q(g207), 
        .QN(n2122) );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n2447), .CLK(n2493), .Q(g713), 
        .QN(n2125) );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n2447), .CLK(n2493), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n2389), .CLK(n2522), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n2375), .CLK(n2528), .Q(
        g1558) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n2420), .CLK(n2506), .Q(
        g695), .QN(n2317) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n2420), .CLK(n2506), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n2429), .CLK(n2502), .Q(g940), .QN(n1712) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n2428), .CLK(n2502), .Q(
        g976), .QN(n2314) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n2370), .CLK(n2531), .Q(g709) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n2412), .CLK(n2510), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n2405), .CLK(n2513), .Q(
        g1574) );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(n2405), .CLK(n2513), .Q(
        g1864), .QN(n2336) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n2383), .CLK(n2524), .Q(
        g369), .QN(n2226) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n2411), .CLK(n2511), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n2410), .CLK(n2511), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(n44), .SI(g1736), .SE(n2410), .CLK(n2511), .Q(n1637), .QN(n4116) );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(n2410), .CLK(n2511), .Q(
        n3065), .QN(n4117) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n2410), .CLK(n2511), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n2410), .CLK(n2511), .Q(
        g1737) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n2394), .CLK(n2519), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n2444), .CLK(n2494), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n2407), .CLK(n2512), .Q(
        g1231), .QN(n2117) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n2446), .CLK(n2493), .Q(g4)
         );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(n2428), .CLK(n2502), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n2381), .CLK(n2525), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n2437), .CLK(n2498), .Q(
        g1304), .QN(n2247) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n2398), .CLK(n2517), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n2446), .CLK(n2493), .Q(
        g1499), .QN(n2281) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n2417), .CLK(n2508), .Q(
        g1444), .QN(n2328) );
  SDFFX1 DFF_37_Q_reg ( .D(n11), .SI(g1444), .SE(n2417), .CLK(n2508), .Q(n3064) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n2403), .CLK(n2515), .Q(
        g4180), .QN(n2134) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n2414), .CLK(n2509), .Q(
        g1543) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n2414), .CLK(n2509), .Q(g315), .QN(n2308) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n2434), .CLK(n2499), .Q(
        g1534) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n2433), .CLK(n2499), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n2366), .CLK(n2533), .Q(
        g1927), .QN(n2237) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n2366), .CLK(n2533), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n2435), .CLK(n2498), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n2435), .CLK(n2498), .Q(
        g1436), .QN(n2325) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n2372), .CLK(n2530), .Q(
        g718) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n2372), .CLK(n2530), .Q(
        g8985), .QN(n1669) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n2372), .CLK(n2530), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n2406), .CLK(n2513), .Q(
        g496) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n2428), .CLK(n2502), .Q(
        g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n33), .SI(g981), .SE(n2428), .CLK(n2502), .Q(g3007)
         );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n2428), .CLK(n2502), .Q(
        test_so1) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n2426), .CLK(n2503), .Q(
        g829), .QN(n1651) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n2393), .CLK(n2519), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n2367), .CLK(n2532), .Q(
        g704), .QN(n2288) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n2437), .CLK(n2497), .Q(
        g1265), .QN(n2243) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n2389), .CLK(n2522), .Q(
        g1786), .QN(n2341) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n2420), .CLK(n2506), .Q(
        g682), .QN(n2221) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n2437), .CLK(n2498), .Q(
        g1296) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n2436), .CLK(n2498), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n2418), .CLK(n2507), .Q(
        g8977), .QN(n1668) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n2382), .CLK(n2525), .Q(
        n3062), .QN(n4111) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n2382), .CLK(n2525), .Q(g327), .QN(n2273) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n2382), .CLK(n2525), .Q(
        g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n2382), .CLK(n2525), .Q(
        g1371) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n2378), .CLK(n2527), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n2378), .CLK(n2527), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n2442), .CLK(n2495), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n2429), .CLK(n2502), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n2373), .CLK(n2530), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n2434), .CLK(n2499), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n2434), .CLK(n2499), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n2388), .CLK(n2522), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n2377), .CLK(n2527), .Q(
        g248), .QN(n1598) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n2377), .CLK(n2527), .Q(
        g1707) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n2377), .CLK(n2527), .Q(
        g1759) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n2377), .CLK(n2528), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n2377), .CLK(n2528), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n2377), .CLK(n2528), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n2419), .CLK(n2506), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n2419), .CLK(n2506), .Q(
        g932), .QN(n1591) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n2421), .CLK(n2505), .Q(
        g1896), .QN(n2222) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n2421), .CLK(n2506), .Q(
        g736), .QN(n2300) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n2419), .CLK(n2506), .Q(
        g1019), .QN(n2229) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n2419), .CLK(n2507), .Q(
        n3061), .QN(n4127) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n2418), .CLK(n2507), .Q(g745) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n2411), .CLK(n2510), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n2411), .CLK(n2511), .Q(
        g8979), .QN(n1667) );
  SDFFX1 DFF_92_Q_reg ( .D(n17), .SI(g8979), .SE(n2445), .CLK(n2493), .Q(g32), 
        .QN(n4113) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n2445), .CLK(n2493), .Q(n1865), .QN(n2094) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n2442), .CLK(n2495), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n2416), .CLK(n2508), .Q(
        g1486), .QN(n2256) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n2415), .CLK(n2508), .Q(
        g1730) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n2415), .CLK(n2508), .Q(
        g1504), .QN(n2139) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n2402), .CLK(n2515), .Q(
        g1470), .QN(n2295) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n2399), .CLK(n2517), .Q(
        g822), .QN(n2344) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n2399), .CLK(n2517), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n2394), .CLK(n2519), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n2390), .CLK(n2521), .Q(
        g174), .QN(n2345) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n2390), .CLK(n2521), .Q(
        g1766), .QN(n2334) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n2388), .CLK(n2522), .Q(
        g1801), .QN(n2339) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n2388), .CLK(n2522), .Q(
        g186), .QN(n2121) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n2387), .CLK(n2522), .Q(
        g959) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n2387), .CLK(n2522), .Q(
        test_so2) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n2369), .CLK(n2532), 
        .Q(g1407) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n2445), .CLK(n2494), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n2444), .CLK(n2494), .Q(
        g4173) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n2413), .CLK(n2509), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n2425), .CLK(n2503), .Q(
        g396) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n2409), .CLK(n2512), .Q(
        g1015), .QN(n2228) );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(n2409), .CLK(n2512), .Q(
        n1650) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n2408), .CLK(n2512), .Q(
        n3059) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n2391), .CLK(n2521), .Q(
        g1415), .QN(n2137) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n2450), .CLK(n2491), .Q(
        g1227), .QN(n2118) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n2450), .CLK(n2491), .Q(
        g1721) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n2429), .CLK(n2502), .Q(
        n3058), .QN(DFF_121_n1) );
  SDFFX1 DFF_122_Q_reg ( .D(n2358), .SI(n3058), .SE(n2401), .CLK(n2515), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(n2448), .CLK(n2492), .Q(
        g284), .QN(n2175) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n2446), .CLK(n2493), .Q(
        g426) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n2382), .CLK(n2525), .Q(
        g219) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n2381), .CLK(n2525), .Q(
        n3056), .QN(DFF_126_n1) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n2381), .CLK(n2525), .Q(
        g806), .QN(n2332) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n2397), .CLK(n2518), .Q(
        g1428), .QN(n2327) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n2397), .CLK(n2518), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n2396), .CLK(n2518), .Q(
        g1564) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n2396), .CLK(n2518), .Q(
        g1741) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n2396), .CLK(n2518), .Q(
        g225), .QN(n2282) );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(n2374), .CLK(n2529), .Q(
        g281) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n2374), .CLK(n2529), .Q(
        g1308) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n2448), .CLK(n2492), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n2408), .CLK(n2512), .Q(
        n3055), .QN(DFF_136_n1) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n2407), .CLK(n2512), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n2369), .CLK(n2532), .Q(
        g1589) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n2416), .CLK(n2508), .Q(
        g1466), .QN(n2260) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n2393), .CLK(n2520), .Q(
        g1571), .QN(n2154) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n2392), .CLK(n2520), .Q(
        g1861), .QN(n2338) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n2392), .CLK(n2520), .Q(
        n3054), .QN(n4118) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n2443), .CLK(n2495), .Q(
        g1448), .QN(n2262) );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(n2442), .CLK(n2495), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n2443), .CLK(n2494), .Q(
        g1333) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n2443), .CLK(n2494), .Q(
        g153), .QN(n2278) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n2368), .CLK(n2532), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(n2444), .CLK(n2494), .Q(
        g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n2444), .CLK(n2494), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n2444), .CLK(n2494), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n2409), .CLK(n2511), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n2378), .CLK(n2527), .Q(
        g1397), .QN(n1711) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n2378), .CLK(n2527), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n2422), .CLK(n2505), .Q(
        g1950), .QN(n2302) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n2422), .CLK(n2505), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(g4892), .SI(g756), .SE(n2408), .CLK(n2512), .Q(
        n3053), .QN(DFF_157_n1) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n2376), .CLK(n2528), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n2449), .CLK(n2491), .Q(
        g105), .QN(n2095) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n2449), .CLK(n2491), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n2449), .CLK(n2492), .Q(
        test_so3), .QN(n4112) );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(n2405), .CLK(n2514), 
        .Q(g1531) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n2446), .CLK(n2493), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n2441), .CLK(n2496), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n2412), .CLK(n2510), .Q(
        g1011), .QN(n2267) );
  SDFFX1 DFF_168_Q_reg ( .D(n16), .SI(g1011), .SE(n2411), .CLK(n2510), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n2411), .CLK(n2510), .Q(
        g1411), .QN(n2160) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n2409), .CLK(n2512), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n2424), .CLK(n2504), .Q(
        g444), .QN(n2250) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n2402), .CLK(n2515), .Q(
        g1474), .QN(n2294) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n2414), .CLK(n2509), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n2413), .CLK(n2509), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n2398), .CLK(n2517), .Q(
        g333), .QN(n2291) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n2385), .CLK(n2524), .Q(
        g269) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n2425), .CLK(n2504), .Q(
        g401), .QN(n2274) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n2433), .CLK(n2500), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n2432), .CLK(n2500), .Q(g9), .QN(n2233) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n2421), .CLK(n2506), .Q(g664)
         );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n2400), .CLK(n2516), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n2399), .CLK(n2516), .Q(
        g1400), .QN(n1629) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n2399), .CLK(n2516), .Q(
        g309), .QN(n2072) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n2399), .CLK(n2516), .Q(
        g814), .QN(n2343) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n2392), .CLK(n2520), .Q(
        g231), .QN(n2283) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n2392), .CLK(n2520), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n2392), .CLK(n2520), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n2386), .CLK(n2523), .Q(
        g869), .QN(n2116) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n2386), .CLK(n2523), .Q(
        g1383) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n2386), .CLK(n2523), .Q(
        g158), .QN(n2259) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n2408), .CLK(n2512), .Q(
        g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n2427), .CLK(n2503), .Q(
        g1023), .QN(n2203) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n2426), .CLK(n2503), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n2426), .CLK(n2503), .Q(
        n3050), .QN(DFF_194_n1) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n2383), .CLK(n2525), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(n2382), .CLK(n2525), .Q(
        g654) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n2403), .CLK(n2515), .Q(
        g293) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n2402), .CLK(n2515), .Q(
        g1346) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n2402), .CLK(n2515), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n2388), .CLK(n2522), .Q(
        g1753) );
  SDFFX1 DFF_201_Q_reg ( .D(n2354), .SI(g1753), .SE(n2388), .CLK(n2522), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n2438), .CLK(n2497), .Q(
        g1240) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n2404), .CLK(n2514), .Q(
        g538) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n2424), .CLK(n2504), .Q(
        g416), .QN(n2248) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n2404), .CLK(n2514), .Q(
        g542) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n2394), .CLK(n2519), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n2383), .CLK(n2524), .Q(
        g374), .QN(n2227) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n2383), .CLK(n2524), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n2423), .CLK(n2505), .Q(
        g1914) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n2404), .CLK(n2514), .Q(
        g530), .QN(n2296) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n2403), .CLK(n2514), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n2366), .CLK(n2533), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n2366), .CLK(n2533), .Q(
        g8978), .QN(n1674) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n2366), .CLK(n2533), .Q(
        test_so4), .QN(n2360) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n2367), .CLK(n2533), 
        .Q(g1317) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n2430), .CLK(n2501), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n2429), .CLK(n2501), .Q(
        g386), .QN(n2272) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n2371), .CLK(n2531), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n2371), .CLK(n2531), .Q(
        g166), .QN(n2257) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n2406), .CLK(n2513), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n2398), .CLK(n2517), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n2398), .CLK(n2517), .Q(
        g1840), .QN(n2301) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n2398), .CLK(n2517), .Q(
        g8983), .QN(n1666) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n2391), .CLK(n2520), .Q(
        g318), .QN(n2271) );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(n2426), .CLK(n2503), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n2426), .CLK(n2503), .Q(
        g794), .QN(n2242) );
  SDFFX1 DFF_228_Q_reg ( .D(n25), .SI(g794), .SE(n2426), .CLK(n2503), .Q(n3048) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n2443), .CLK(n2495), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n2409), .CLK(n2511), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n2438), .CLK(n2497), .Q(
        g1250), .QN(n2268) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n2438), .CLK(n2497), .Q(
        g1163) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n2413), .CLK(n2510), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n2443), .CLK(n2494), .Q(
        g1032), .QN(n2201) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n2379), .CLK(n2527), .Q(
        g1432), .QN(n2263) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n2446), .CLK(n2493), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n2393), .CLK(n2519), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n2395), .CLK(n2519), .Q(g330), .QN(n2071) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n2395), .CLK(n2519), .Q(
        g1157), .QN(n4132) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n2395), .CLK(n2519), .Q(
        n3046), .QN(n4130) );
  SDFFX1 DFF_242_Q_reg ( .D(n38), .SI(n3046), .SE(n2394), .CLK(n2519), .Q(
        n3045), .QN(DFF_242_n1) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n2394), .CLK(n2519), .Q(
        g928), .QN(n1604) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n2395), .CLK(n2518), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n2405), .CLK(n2514), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n2403), .CLK(n2514), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n2403), .CLK(n2514), .Q(
        g4178), .QN(n2133) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n2398), .CLK(n2517), .Q(
        g861) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n2380), .CLK(n2526), .Q(
        g1627) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n2436), .CLK(n2498), .Q(
        g1292) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n2436), .CLK(n2498), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n2436), .CLK(n2498), .Q(
        n3044) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n2428), .CLK(n2502), .Q(
        g4176), .QN(n2132) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n2410), .CLK(n2511), .Q(
        g1583) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n2409), .CLK(n2511), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n2405), .CLK(n2514), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n2379), .CLK(n2527), .Q(
        g1546) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n2374), .CLK(n2529), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n2374), .CLK(n2529), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n2374), .CLK(n2529), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n2356), .SI(g617), .SE(n2373), .CLK(n2530), .Q(
        n1631), .QN(n4114) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n2450), .CLK(n2491), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n2391), .CLK(n2521), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n2387), .CLK(n2523), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n2444), .CLK(n2494), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n2433), .CLK(n2499), .Q(g8)
         );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n2433), .CLK(n2500), .Q(
        test_so5) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n2427), .CLK(n2502), .Q(
        g2648) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n2427), .CLK(n2502), .Q(
        g255) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n2432), .CLK(n2500), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n2390), .CLK(n2521), .Q(
        g1738) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n2379), .CLK(n2526), .Q(
        g1478), .QN(n2331) );
  SDFFX1 DFF_275_Q_reg ( .D(n374), .SI(g1478), .SE(n2379), .CLK(n2526), .Q(
        n3042), .QN(DFF_275_n1) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n2376), .CLK(n2528), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n2414), .CLK(n2509), .Q(
        g1482), .QN(n2261) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n2381), .CLK(n2526), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n2370), .CLK(n2531), .Q(
        g296) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n2370), .CLK(n2531), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n2370), .CLK(n2531), .Q(
        g700) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n2412), .CLK(n2510), .Q(
        g1762) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n2412), .CLK(n2510), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n2378), .CLK(n2527), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n2448), .CLK(n2492), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n2448), .CLK(n2492), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n2417), .CLK(n2507), .Q(
        g8980), .QN(n1673) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n2380), .CLK(n2526), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n2449), .CLK(n2492), .Q(
        n3041), .QN(n4129) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n2429), .CLK(n2501), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n2429), .CLK(n2501), .Q(
        g2986) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n2427), .CLK(n2503), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n2446), .CLK(n2493), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n2385), .CLK(n2523), .Q(
        g971), .QN(n2315) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n2385), .CLK(n2523), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n2443), .CLK(n2495), .Q(
        g143), .QN(n2279) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n2431), .CLK(n2500), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n2407), .CLK(n2512), .Q(
        g1212), .QN(n2347) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n2432), .CLK(n2500), .Q(
        g1918), .QN(n2287) );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(n2432), .CLK(n2500), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n2431), .CLK(n2500), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n2419), .CLK(n2507), .Q(
        g237), .QN(n2284) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n2419), .CLK(n2507), .Q(g746), .QN(n2337) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n2376), .CLK(n2528), .Q(
        g1462), .QN(n2330) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n2376), .CLK(n2528), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n2420), .CLK(n2506), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n2400), .CLK(n2516), .Q(g837) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n2373), .CLK(n2530), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n2450), .CLK(n2491), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n2450), .CLK(n2491), .Q(
        g944) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n2422), .CLK(n2505), .Q(
        g1941) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n2393), .CLK(n2520), .Q(
        g170), .QN(n2346) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n2393), .CLK(n2520), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n2420), .CLK(n2506), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n2375), .CLK(n2529), .Q(
        g953) );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(n2413), .CLK(n2510), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(n114), .SI(g1958), .SE(n2413), .CLK(n2510), .Q(
        n3040), .QN(n4115) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n2412), .CLK(n2510), .Q(
        g1765) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n2412), .CLK(n2510), .Q(
        g1733) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n2437), .CLK(n2497), .Q(
        test_so6) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n2441), .CLK(n2496), 
        .Q(g1610) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n2383), .CLK(n2525), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n2383), .CLK(n2525), .Q(
        g1324) );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(n2415), .CLK(n2508), .Q(
        g1540) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n2415), .CLK(n2509), .Q(
        n3038), .QN(n4126) );
  SDFFX1 DFF_328_Q_reg ( .D(n2357), .SI(n3038), .SE(n2407), .CLK(n2513), .Q(
        g3069) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n2406), .CLK(n2513), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n2368), .CLK(n2532), .Q(
        n3037), .QN(DFF_330_n1) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n2415), .CLK(n2509), .Q(
        g213), .QN(n2123) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n2389), .CLK(n2522), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n2367), .CLK(n2533), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n2438), .CLK(n2497), .Q(
        g1245), .QN(n2265) );
  SDFFX1 DFF_335_Q_reg ( .D(n2), .SI(g1245), .SE(n2438), .CLK(n2497), .Q(n3036), .QN(n4131) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(n2408), .CLK(n2512), .Q(
        n3035), .QN(DFF_336_n1) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n2385), .CLK(n2524), .Q(
        g148), .QN(n2280) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n2385), .CLK(n2524), .Q(g833), .QN(n2074) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n2423), .CLK(n2505), .Q(
        g1923) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n2422), .CLK(n2505), .Q(
        g936), .QN(n1630) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n2390), .CLK(n2521), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n2390), .CLK(n2521), .Q(
        g849), .QN(n2102) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n2389), .CLK(n2521), .Q(
        g1336) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n2389), .CLK(n2521), .Q(
        g272) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n2413), .CLK(n2509), .Q(
        g1806), .QN(n2340) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n2399), .CLK(n2517), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n2421), .CLK(n2505), .Q(
        g1887), .QN(n2196) );
  SDFFX1 DFF_350_Q_reg ( .D(n42), .SI(g1887), .SE(n2421), .CLK(n2505), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n2445), .CLK(n2493), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n2445), .CLK(n2494), .Q(
        n3033), .QN(n4128) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(n2445), .CLK(n2494), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n2432), .CLK(n2500), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n2438), .CLK(n2497), .Q(
        g1255) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n2392), .CLK(n2520), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n2391), .CLK(n2520), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n2374), .CLK(n2529), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n2367), .CLK(n2532), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n2433), .CLK(n2499), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n2451), .CLK(n2491), .Q(
        g1218), .QN(n2119) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n2373), .CLK(n2529), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n2373), .CLK(n2529), .Q(
        g8986), .QN(n1665) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n2373), .CLK(n2529), .Q(
        g182), .QN(n2277) );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(n2400), .CLK(n2516), .Q(
        g950) );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(n2400), .CLK(n2516), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n2400), .CLK(n2516), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n2424), .CLK(n2504), .Q(
        g448) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n2431), .CLK(n2500), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n2440), .CLK(n2496), .Q(
        g1727) );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(n2441), .CLK(n2495), .Q(
        g1592) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n2441), .CLK(n2496), .Q(
        g1703), .QN(n2349) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n2422), .CLK(n2505), .Q(
        g1932) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n2414), .CLK(n2509), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n2450), .CLK(n2491), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n2451), .CLK(n2491), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n2423), .CLK(n2504), .Q(
        g440), .QN(n2249) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n2404), .CLK(n2514), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n2404), .CLK(n2514), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n2447), .CLK(n2492), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n2371), .CLK(n2531), .Q(
        g139), .QN(n2254) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n2370), .CLK(n2531), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(n32), .SI(g1149), .SE(n2370), .CLK(n2531), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n2401), .CLK(n2515), .Q(
        n3030), .QN(DFF_385_n1) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n2401), .CLK(n2516), .Q(
        g263) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n2401), .CLK(n2516), .Q(
        g818) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n2401), .CLK(n2516), .Q(
        g1747) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n2400), .CLK(n2516), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n2386), .CLK(n2523), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n2386), .CLK(n2523), .Q(
        g1524) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n2386), .CLK(n2523), .Q(
        g1577), .QN(n2147) );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(n2425), .CLK(n2503), .Q(
        g810) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n2425), .CLK(n2503), .Q(
        g391), .QN(n2309) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n2448), .CLK(n2492), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n2387), .CLK(n2522), .Q(
        g1386), .QN(n2276) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n2387), .CLK(n2523), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n2387), .CLK(n2523), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(n2385), .CLK(n2523), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n2440), .CLK(n2496), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n2439), .CLK(n2497), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n2376), .CLK(n2528), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n2375), .CLK(n2528), .Q(
        g650) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n2417), .CLK(n2508), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n2368), .CLK(n2532), .Q(
        g853), .QN(n2079) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n2424), .CLK(n2504), .Q(
        g421), .QN(n2290) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n2424), .CLK(n2504), .Q(
        g4174), .QN(n2130) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n2384), .CLK(n2524), .Q(
        g956), .QN(n2085) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n2384), .CLK(n2524), .Q(
        g378), .QN(n2225) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n2375), .CLK(n2528), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n2375), .CLK(n2529), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n2375), .CLK(n2529), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n2449), .CLK(n2491), .Q(
        g1027), .QN(n2350) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n2442), .CLK(n2495), .Q(
        g1003), .QN(n2306) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n2441), .CLK(n2495), .Q(
        g1403), .QN(n2264) );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(n2441), .CLK(n2495), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n2381), .CLK(n2526), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n2381), .CLK(n2526), .Q(
        g1223), .QN(n2120) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n2425), .CLK(n2504), .Q(
        g406), .QN(n2241) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n2440), .CLK(n2496), .Q(
        g1811) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(n2440), .CLK(n2496), .Q(
        n3029), .QN(n4119) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n2440), .CLK(n2496), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(n2440), .CLK(n2496), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n2378), .CLK(n2527), .Q(
        g1595) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n2434), .CLK(n2499), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n2369), .CLK(n2531), .Q(
        g727) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n2366), .CLK(n2533), .Q(
        test_so8) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n2418), .CLK(n2507), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n2418), .CLK(n2507), .Q(
        g481) );
  SDFFX1 DFF_431_Q_reg ( .D(g3462), .SI(g481), .SE(n2418), .CLK(n2507), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n2384), .CLK(n2524), .Q(
        g1330) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n2384), .CLK(n2524), .Q(
        g845), .QN(n2103) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n2384), .CLK(n2524), .Q(
        g4181), .QN(n2129) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n2380), .CLK(n2526), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n2380), .CLK(n2526), .Q(
        n3027), .QN(DFF_436_n1) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n2435), .CLK(n2499), .Q(
        g1490), .QN(n2329) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n2434), .CLK(n2499), .Q(
        g1166), .QN(n2275) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n2414), .CLK(n2509), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n2391), .CLK(n2520), .Q(
        n3026), .QN(DFF_441_n1) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n2437), .CLK(n2497), .Q(
        g1260), .QN(n2240) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n2380), .CLK(n2526), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n2397), .CLK(n2517), .Q(
        g131), .QN(n2253) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n2397), .CLK(n2517), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n2369), .CLK(n2531), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n2368), .CLK(n2532), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n2367), .CLK(n2532), .Q(
        g1318) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n2367), .CLK(n2533), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n2447), .CLK(n2492), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n2447), .CLK(n2492), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n2352), .SI(g2608), .SE(n2449), .CLK(n2492), .Q(
        n3024), .QN(DFF_452_n1) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n2402), .CLK(n2515), .Q(
        g1549) );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(n2402), .CLK(n2515), .Q(
        g947), .QN(n2073) );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(n2401), .CLK(n2515), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n2435), .CLK(n2498), .Q(
        g1598), .QN(n2144) );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(n2435), .CLK(n2499), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n2388), .CLK(n2522), .Q(
        g1321) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n2406), .CLK(n2513), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n2394), .CLK(n2519), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n2431), .CLK(n2501), .Q(
        g1909), .QN(n2316) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n2431), .CLK(n2501), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n2431), .CLK(n2501), .Q(
        g1552), .QN(n2143) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n2430), .CLK(n2501), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n2430), .CLK(n2501), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(n2430), .CLK(n2501), .Q(
        g1586), .QN(n2141) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n2430), .CLK(n2501), .Q(
        g324), .QN(n2269) );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(n2430), .CLK(n2501), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n2389), .CLK(n2521), .Q(
        g1341), .QN(n2311) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n2379), .CLK(n2526), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(n2379), .CLK(n2527), .Q(
        n3023), .QN(n4120) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(n2448), .CLK(n2492), .Q(
        n3022), .QN(n4121) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n2403), .CLK(n2515), .Q(
        g135), .QN(n2255) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n2368), .CLK(n2532), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n2368), .CLK(n2532), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n2442), .CLK(n2495), .Q(
        g1607) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n2442), .CLK(n2495), .Q(
        g321), .QN(n2310) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n2417), .CLK(n2507), .Q(
        g8982), .QN(n1672) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n2439), .CLK(n2497), .Q(
        g1275) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n2433), .CLK(n2500), .Q(
        test_so9) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n2435), .CLK(n2499), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n2384), .CLK(n2524), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(n280), .SI(g382), .SE(n2439), .CLK(n2496), .Q(
        n3020), .QN(n4122) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n2439), .CLK(n2496), .Q(
        g266) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n2439), .CLK(n2496), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n2415), .CLK(n2509), .Q(
        n3019), .QN(n4125) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n2421), .CLK(n2506), .Q(
        g673), .QN(n2195) );
  SDFFX1 DFF_489_Q_reg ( .D(g4904), .SI(g673), .SE(n2436), .CLK(n2498), .Q(
        n3018), .QN(DFF_489_n1) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n2436), .CLK(n2498), .Q(
        g162), .QN(n2258) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n2425), .CLK(n2504), .Q(
        g411), .QN(n2292) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n2423), .CLK(n2504), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n2423), .CLK(n2505), .Q(
        g1905) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n2411), .CLK(n2511), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n2396), .CLK(n2518), .Q(
        g1630) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n2396), .CLK(n2518), .Q(
        g8976), .QN(n1671) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n2376), .CLK(n2528), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n2437), .CLK(n2498), .Q(
        g1300), .QN(n2246) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n2427), .CLK(n2503), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n2372), .CLK(n2530), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n2372), .CLK(n2530), .Q(
        g1750) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n2372), .CLK(n2530), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n2371), .CLK(n2530), .Q(
        g1440), .QN(n2326) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n2371), .CLK(n2530), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(n2371), .CLK(n2530), .Q(
        g1528) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n2407), .CLK(n2513), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(n2407), .CLK(n2513), .Q(
        n3017), .QN(n4123) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n2393), .CLK(n2519), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n2447), .CLK(n2493), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n2439), .CLK(n2497), .Q(
        g1235), .QN(n2266) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n2369), .CLK(n2531), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n2423), .CLK(n2504), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n2418), .CLK(n2507), .Q(
        g8981), .QN(n1664) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(n2416), .CLK(n2508), .Q(
        g1555) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n2416), .CLK(n2508), .Q(
        g995), .QN(n2304) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n2416), .CLK(n2508), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n2416), .CLK(n2508), .Q(
        n3016), .QN(n4124) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(n2408), .CLK(n2512), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n2434), .CLK(n2499), .Q(
        g1494), .QN(n2293) );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(n2391), .CLK(n2521), .Q(
        g1567) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n2420), .CLK(n2506), .Q(
        g691) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n2404), .CLK(n2514), .Q(
        g534) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n2390), .CLK(n2521), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n2396), .CLK(n2518), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n2395), .CLK(n2518), .Q(
        g1160) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n2395), .CLK(n2518), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n2369), .CLK(n2532), .Q(g1) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n2406), .CLK(n2513), .Q(g511) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n2406), .CLK(n2513), .Q(
        g1724) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n2405), .CLK(n2513), .Q(
        g12), .QN(n2232) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n2422), .CLK(n2505), .Q(
        g1878) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n2417), .CLK(n2507), .Q(
        test_so10), .QN(n2361) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n2380), .CLK(n2526), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(g6179), .IN2(n2352), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n19), .IN2(n1132), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n1226), .IN2(n1858), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(g5556), .IN2(n898), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n857), .IN2(n902), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n14), .IN2(n14), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n938), .IN2(n2351), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n2351), .IN2(n2351), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n2351), .IN2(n2351), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n2351), .IN2(n2351), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n68), .IN2(n1162), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n1155), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n929), .IN2(n2355), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n2451), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n968), .S(Trigger_select), .Q(
        g4207) );
  INVX0 U2387 ( .INP(g109), .ZN(n2362) );
  INVX0 U2388 ( .INP(g109), .ZN(n2363) );
  INVX0 U2389 ( .INP(g109), .ZN(n2364) );
  INVX0 U2390 ( .INP(g109), .ZN(n2365) );
  INVX2 U2391 ( .INP(n2351), .ZN(n14) );
  NBUFFX2 U2392 ( .INP(n2542), .Z(n2492) );
  NBUFFX2 U2393 ( .INP(n2542), .Z(n2493) );
  NBUFFX2 U2394 ( .INP(n2542), .Z(n2491) );
  NBUFFX2 U2395 ( .INP(n2535), .Z(n2526) );
  NBUFFX2 U2396 ( .INP(n2540), .Z(n2501) );
  NBUFFX2 U2397 ( .INP(n2536), .Z(n2523) );
  NBUFFX2 U2398 ( .INP(n2537), .Z(n2516) );
  NBUFFX2 U2399 ( .INP(n2541), .Z(n2496) );
  NBUFFX2 U2400 ( .INP(n2537), .Z(n2514) );
  NBUFFX2 U2401 ( .INP(n2536), .Z(n2520) );
  NBUFFX2 U2402 ( .INP(n2534), .Z(n2529) );
  NBUFFX2 U2403 ( .INP(n2536), .Z(n2521) );
  NBUFFX2 U2404 ( .INP(n2539), .Z(n2505) );
  NBUFFX2 U2405 ( .INP(n2541), .Z(n2495) );
  NBUFFX2 U2406 ( .INP(n2535), .Z(n2527) );
  NBUFFX2 U2407 ( .INP(n2539), .Z(n2507) );
  NBUFFX2 U2408 ( .INP(n2541), .Z(n2497) );
  NBUFFX2 U2409 ( .INP(n2534), .Z(n2532) );
  NBUFFX2 U2410 ( .INP(n2540), .Z(n2503) );
  NBUFFX2 U2411 ( .INP(n2534), .Z(n2530) );
  NBUFFX2 U2412 ( .INP(n2540), .Z(n2499) );
  NBUFFX2 U2413 ( .INP(n2538), .Z(n2509) );
  NBUFFX2 U2414 ( .INP(n2537), .Z(n2515) );
  NBUFFX2 U2415 ( .INP(n2539), .Z(n2508) );
  NBUFFX2 U2416 ( .INP(n2541), .Z(n2498) );
  NBUFFX2 U2417 ( .INP(n2535), .Z(n2525) );
  NBUFFX2 U2419 ( .INP(n2538), .Z(n2512) );
  NBUFFX2 U2420 ( .INP(n2541), .Z(n2494) );
  NBUFFX2 U2421 ( .INP(n2536), .Z(n2519) );
  NBUFFX2 U2422 ( .INP(n2538), .Z(n2511) );
  NBUFFX2 U2423 ( .INP(n2535), .Z(n2524) );
  NBUFFX2 U2424 ( .INP(n2538), .Z(n2513) );
  NBUFFX2 U2425 ( .INP(n2538), .Z(n2510) );
  NBUFFX2 U2426 ( .INP(n2534), .Z(n2531) );
  NBUFFX2 U2427 ( .INP(n2539), .Z(n2506) );
  NBUFFX2 U2428 ( .INP(n2535), .Z(n2528) );
  NBUFFX2 U2429 ( .INP(n2536), .Z(n2522) );
  NBUFFX2 U2430 ( .INP(n2537), .Z(n2518) );
  NBUFFX2 U2431 ( .INP(n2537), .Z(n2517) );
  NBUFFX2 U2432 ( .INP(n2539), .Z(n2504) );
  NBUFFX2 U2433 ( .INP(n2540), .Z(n2502) );
  NBUFFX2 U2434 ( .INP(n2540), .Z(n2500) );
  NBUFFX2 U2435 ( .INP(n2534), .Z(n2533) );
  NBUFFX2 U2436 ( .INP(n2480), .Z(n2366) );
  NBUFFX2 U2437 ( .INP(n2480), .Z(n2367) );
  NBUFFX2 U2438 ( .INP(n2479), .Z(n2368) );
  NBUFFX2 U2439 ( .INP(n2479), .Z(n2369) );
  NBUFFX2 U2440 ( .INP(n2479), .Z(n2370) );
  NBUFFX2 U2441 ( .INP(n2478), .Z(n2371) );
  NBUFFX2 U2442 ( .INP(n2478), .Z(n2372) );
  NBUFFX2 U2443 ( .INP(n2478), .Z(n2373) );
  NBUFFX2 U2444 ( .INP(n2477), .Z(n2374) );
  NBUFFX2 U2445 ( .INP(n2477), .Z(n2375) );
  NBUFFX2 U2446 ( .INP(n2477), .Z(n2376) );
  NBUFFX2 U2447 ( .INP(n2476), .Z(n2377) );
  NBUFFX2 U2448 ( .INP(n2476), .Z(n2378) );
  NBUFFX2 U2449 ( .INP(n2476), .Z(n2379) );
  NBUFFX2 U2450 ( .INP(n2475), .Z(n2380) );
  NBUFFX2 U2451 ( .INP(n2475), .Z(n2381) );
  NBUFFX2 U2452 ( .INP(n2475), .Z(n2382) );
  NBUFFX2 U2453 ( .INP(n2474), .Z(n2383) );
  NBUFFX2 U2454 ( .INP(n2474), .Z(n2384) );
  NBUFFX2 U2455 ( .INP(n2474), .Z(n2385) );
  NBUFFX2 U2456 ( .INP(n2473), .Z(n2386) );
  NBUFFX2 U2457 ( .INP(n2473), .Z(n2387) );
  NBUFFX2 U2458 ( .INP(n2473), .Z(n2388) );
  NBUFFX2 U2459 ( .INP(n2472), .Z(n2389) );
  NBUFFX2 U2460 ( .INP(n2472), .Z(n2390) );
  NBUFFX2 U2461 ( .INP(n2472), .Z(n2391) );
  NBUFFX2 U2462 ( .INP(n2471), .Z(n2392) );
  NBUFFX2 U2463 ( .INP(n2471), .Z(n2393) );
  NBUFFX2 U2464 ( .INP(n2471), .Z(n2394) );
  NBUFFX2 U2465 ( .INP(n2470), .Z(n2395) );
  NBUFFX2 U2466 ( .INP(n2470), .Z(n2396) );
  NBUFFX2 U2467 ( .INP(n2470), .Z(n2397) );
  NBUFFX2 U2469 ( .INP(n2469), .Z(n2398) );
  NBUFFX2 U2470 ( .INP(n2469), .Z(n2399) );
  NBUFFX2 U2471 ( .INP(n2469), .Z(n2400) );
  NBUFFX2 U2472 ( .INP(n2468), .Z(n2401) );
  NBUFFX2 U2473 ( .INP(n2468), .Z(n2402) );
  NBUFFX2 U2474 ( .INP(n2468), .Z(n2403) );
  NBUFFX2 U2475 ( .INP(n2467), .Z(n2404) );
  NBUFFX2 U2476 ( .INP(n2467), .Z(n2405) );
  NBUFFX2 U2477 ( .INP(n2467), .Z(n2406) );
  NBUFFX2 U2479 ( .INP(n2466), .Z(n2407) );
  NBUFFX2 U2480 ( .INP(n2466), .Z(n2408) );
  NBUFFX2 U2481 ( .INP(n2466), .Z(n2409) );
  NBUFFX2 U2482 ( .INP(n2465), .Z(n2410) );
  NBUFFX2 U2483 ( .INP(n2465), .Z(n2411) );
  NBUFFX2 U2484 ( .INP(n2465), .Z(n2412) );
  NBUFFX2 U2485 ( .INP(n2464), .Z(n2413) );
  NBUFFX2 U2486 ( .INP(n2464), .Z(n2414) );
  NBUFFX2 U2487 ( .INP(n2464), .Z(n2415) );
  NBUFFX2 U2489 ( .INP(n2463), .Z(n2416) );
  NBUFFX2 U2490 ( .INP(n2463), .Z(n2417) );
  NBUFFX2 U2491 ( .INP(n2463), .Z(n2418) );
  NBUFFX2 U2492 ( .INP(n2462), .Z(n2419) );
  NBUFFX2 U2493 ( .INP(n2462), .Z(n2420) );
  NBUFFX2 U2494 ( .INP(n2462), .Z(n2421) );
  NBUFFX2 U2495 ( .INP(n2461), .Z(n2422) );
  NBUFFX2 U2496 ( .INP(n2461), .Z(n2423) );
  NBUFFX2 U2497 ( .INP(n2461), .Z(n2424) );
  NBUFFX2 U2498 ( .INP(n2460), .Z(n2425) );
  NBUFFX2 U2499 ( .INP(n2460), .Z(n2426) );
  NBUFFX2 U2500 ( .INP(n2460), .Z(n2427) );
  NBUFFX2 U2501 ( .INP(n2459), .Z(n2428) );
  NBUFFX2 U2502 ( .INP(n2459), .Z(n2429) );
  NBUFFX2 U2503 ( .INP(n2459), .Z(n2430) );
  NBUFFX2 U2504 ( .INP(n2458), .Z(n2431) );
  NBUFFX2 U2505 ( .INP(n2458), .Z(n2432) );
  NBUFFX2 U2506 ( .INP(n2458), .Z(n2433) );
  NBUFFX2 U2507 ( .INP(n2457), .Z(n2434) );
  NBUFFX2 U2508 ( .INP(n2457), .Z(n2435) );
  NBUFFX2 U2509 ( .INP(n2457), .Z(n2436) );
  NBUFFX2 U2510 ( .INP(n2456), .Z(n2437) );
  NBUFFX2 U2511 ( .INP(n2456), .Z(n2438) );
  NBUFFX2 U2512 ( .INP(n2456), .Z(n2439) );
  NBUFFX2 U2513 ( .INP(n2455), .Z(n2440) );
  NBUFFX2 U2514 ( .INP(n2455), .Z(n2441) );
  NBUFFX2 U2515 ( .INP(n2455), .Z(n2442) );
  NBUFFX2 U2516 ( .INP(n2454), .Z(n2443) );
  NBUFFX2 U2517 ( .INP(n2454), .Z(n2444) );
  NBUFFX2 U2518 ( .INP(n2454), .Z(n2445) );
  NBUFFX2 U2519 ( .INP(n2453), .Z(n2446) );
  NBUFFX2 U2520 ( .INP(n2453), .Z(n2447) );
  NBUFFX2 U2521 ( .INP(n2453), .Z(n2448) );
  NBUFFX2 U2522 ( .INP(n2452), .Z(n2449) );
  NBUFFX2 U2523 ( .INP(n2452), .Z(n2450) );
  NBUFFX2 U2524 ( .INP(n2452), .Z(n2451) );
  NBUFFX2 U2525 ( .INP(n2490), .Z(n2452) );
  NBUFFX2 U2526 ( .INP(n2490), .Z(n2453) );
  NBUFFX2 U2527 ( .INP(n2489), .Z(n2454) );
  NBUFFX2 U2528 ( .INP(n2489), .Z(n2455) );
  NBUFFX2 U2529 ( .INP(n2489), .Z(n2456) );
  NBUFFX2 U2530 ( .INP(n2488), .Z(n2457) );
  NBUFFX2 U2531 ( .INP(n2488), .Z(n2458) );
  NBUFFX2 U2532 ( .INP(n2488), .Z(n2459) );
  NBUFFX2 U2535 ( .INP(n2487), .Z(n2460) );
  NBUFFX2 U2536 ( .INP(n2487), .Z(n2461) );
  NBUFFX2 U2537 ( .INP(n2487), .Z(n2462) );
  NBUFFX2 U2538 ( .INP(n2486), .Z(n2463) );
  NBUFFX2 U2539 ( .INP(n2486), .Z(n2464) );
  NBUFFX2 U2540 ( .INP(n2486), .Z(n2465) );
  NBUFFX2 U2541 ( .INP(n2485), .Z(n2466) );
  NBUFFX2 U2542 ( .INP(n2485), .Z(n2467) );
  NBUFFX2 U2543 ( .INP(n2485), .Z(n2468) );
  NBUFFX2 U2544 ( .INP(n2484), .Z(n2469) );
  NBUFFX2 U2545 ( .INP(n2484), .Z(n2470) );
  NBUFFX2 U2546 ( .INP(n2484), .Z(n2471) );
  NBUFFX2 U2547 ( .INP(n2483), .Z(n2472) );
  NBUFFX2 U2548 ( .INP(n2483), .Z(n2473) );
  NBUFFX2 U2549 ( .INP(n2483), .Z(n2474) );
  NBUFFX2 U2550 ( .INP(n2482), .Z(n2475) );
  NBUFFX2 U2551 ( .INP(n2482), .Z(n2476) );
  NBUFFX2 U2552 ( .INP(n2482), .Z(n2477) );
  NBUFFX2 U2553 ( .INP(n2481), .Z(n2478) );
  NBUFFX2 U2554 ( .INP(n2481), .Z(n2479) );
  NBUFFX2 U2555 ( .INP(n2481), .Z(n2480) );
  NBUFFX2 U2556 ( .INP(test_se), .Z(n2481) );
  NBUFFX2 U2557 ( .INP(n2486), .Z(n2482) );
  NBUFFX2 U2558 ( .INP(n2463), .Z(n2483) );
  NBUFFX2 U2559 ( .INP(n2464), .Z(n2484) );
  NBUFFX2 U2560 ( .INP(n2465), .Z(n2485) );
  NBUFFX2 U2561 ( .INP(test_se), .Z(n2486) );
  NBUFFX2 U2562 ( .INP(test_se), .Z(n2487) );
  NBUFFX2 U2563 ( .INP(n2480), .Z(n2488) );
  NBUFFX2 U2564 ( .INP(test_se), .Z(n2489) );
  NBUFFX2 U2565 ( .INP(n2481), .Z(n2490) );
  NBUFFX2 U2566 ( .INP(CK), .Z(n2534) );
  NBUFFX2 U2567 ( .INP(CK), .Z(n2535) );
  NBUFFX2 U2568 ( .INP(CK), .Z(n2536) );
  NBUFFX2 U2569 ( .INP(CK), .Z(n2537) );
  NBUFFX2 U2570 ( .INP(CK), .Z(n2538) );
  NBUFFX2 U2571 ( .INP(CK), .Z(n2539) );
  NBUFFX2 U2572 ( .INP(CK), .Z(n2540) );
  NBUFFX2 U2573 ( .INP(CK), .Z(n2541) );
  NBUFFX2 U2574 ( .INP(CK), .Z(n2542) );
  NAND2X0 U2576 ( .IN1(n2543), .IN2(n2544), .QN(n962) );
  OR2X1 U2577 ( .IN1(n902), .IN2(n1696), .Q(n2544) );
  NAND2X0 U2578 ( .IN1(n2545), .IN2(n1696), .QN(n2543) );
  INVX0 U2579 ( .INP(n2546), .ZN(n2545) );
  NAND2X0 U2580 ( .IN1(n2547), .IN2(n2548), .QN(n917) );
  OR2X1 U2581 ( .IN1(n857), .IN2(n1697), .Q(n2548) );
  NAND2X0 U2582 ( .IN1(n2549), .IN2(n1697), .QN(n2547) );
  INVX0 U2583 ( .INP(n2550), .ZN(n2549) );
  NOR2X0 U2584 ( .IN1(n2551), .IN2(n2552), .QN(n838) );
  INVX0 U2585 ( .INP(n2553), .ZN(n387) );
  NOR2X0 U2586 ( .IN1(n2365), .IN2(n2554), .QN(n2353) );
  NOR2X0 U2587 ( .IN1(n2555), .IN2(n3064), .QN(n2554) );
  INVX0 U2588 ( .INP(n2556), .ZN(n2352) );
  INVX0 U2589 ( .INP(n2557), .ZN(n22) );
  INVX0 U2590 ( .INP(n2558), .ZN(n19) );
  INVX0 U2591 ( .INP(n2559), .ZN(n177) );
  NAND4X0 U2592 ( .IN1(n2560), .IN2(g46), .IN3(n2561), .IN4(n2562), .QN(n1588)
         );
  NAND2X0 U2593 ( .IN1(n2563), .IN2(g46), .QN(n1587) );
  NAND2X0 U2594 ( .IN1(n2564), .IN2(g42), .QN(n1586) );
  NAND2X0 U2595 ( .IN1(n2564), .IN2(n2561), .QN(n1585) );
  AND3X1 U2596 ( .IN1(g47), .IN2(n2565), .IN3(n2560), .Q(n2564) );
  INVX0 U2597 ( .INP(n2566), .ZN(n1229) );
  NAND2X0 U2598 ( .IN1(g4173), .IN2(g4174), .QN(n1214) );
  NAND2X0 U2599 ( .IN1(n1193), .IN2(g4176), .QN(n1153) );
  NAND2X0 U2600 ( .IN1(n2567), .IN2(g806), .QN(n1151) );
  NAND2X0 U2601 ( .IN1(n1125), .IN2(g4178), .QN(n1099) );
  NAND2X0 U2602 ( .IN1(n1123), .IN2(g814), .QN(n1097) );
  NOR2X0 U2603 ( .IN1(n2568), .IN2(n2569), .QN(g9721) );
  XOR2X1 U2604 ( .IN1(g611), .IN2(n2570), .Q(n2568) );
  NOR2X0 U2605 ( .IN1(n2571), .IN2(n2572), .QN(n2570) );
  NOR2X0 U2606 ( .IN1(n2573), .IN2(n2574), .QN(n2572) );
  NOR2X0 U2607 ( .IN1(n2575), .IN2(g617), .QN(n2573) );
  NOR2X0 U2608 ( .IN1(n804), .IN2(n2576), .QN(n2575) );
  INVX0 U2609 ( .INP(n2577), .ZN(n2571) );
  NOR3X0 U2610 ( .IN1(n2569), .IN2(n2578), .IN3(n2579), .QN(g9555) );
  AND3X1 U2611 ( .IN1(g1834), .IN2(n808), .IN3(n926), .Q(n2579) );
  NAND2X0 U2612 ( .IN1(n2301), .IN2(n2580), .QN(n808) );
  OR2X1 U2613 ( .IN1(n2559), .IN2(n812), .Q(n2580) );
  NOR2X0 U2614 ( .IN1(n806), .IN2(g1834), .QN(n2578) );
  NAND3X0 U2615 ( .IN1(n2581), .IN2(n2582), .IN3(n2583), .QN(g9451) );
  AND3X1 U2616 ( .IN1(n2584), .IN2(n2585), .IN3(g18), .Q(g9272) );
  OR2X1 U2617 ( .IN1(n2586), .IN2(n1605), .Q(n2585) );
  NAND3X0 U2618 ( .IN1(n2586), .IN2(n2587), .IN3(n1605), .QN(n2584) );
  NAND2X0 U2619 ( .IN1(n812), .IN2(n2588), .QN(n2586) );
  NAND3X0 U2620 ( .IN1(n2589), .IN2(n2590), .IN3(n2591), .QN(n2588) );
  NAND3X0 U2621 ( .IN1(g1814), .IN2(g1822), .IN3(g1828), .QN(n2590) );
  NOR2X0 U2622 ( .IN1(n2569), .IN2(n2592), .QN(g9269) );
  XOR2X1 U2623 ( .IN1(g1822), .IN2(n2593), .Q(n2592) );
  NAND2X0 U2624 ( .IN1(n812), .IN2(n2594), .QN(n2593) );
  NAND3X0 U2625 ( .IN1(n822), .IN2(n2591), .IN3(n2595), .QN(n2594) );
  NAND2X0 U2626 ( .IN1(n1643), .IN2(n2596), .QN(n2595) );
  NOR2X0 U2627 ( .IN1(n2597), .IN2(n2569), .QN(g9266) );
  XOR2X1 U2628 ( .IN1(n2598), .IN2(n1608), .Q(n2597) );
  NAND2X0 U2629 ( .IN1(n2599), .IN2(n2600), .QN(n2598) );
  NAND3X0 U2630 ( .IN1(n1643), .IN2(n2596), .IN3(n812), .QN(n2600) );
  INVX0 U2631 ( .INP(n817), .ZN(n2596) );
  NAND2X0 U2632 ( .IN1(n812), .IN2(n2601), .QN(n2599) );
  NAND2X0 U2633 ( .IN1(n2602), .IN2(n2559), .QN(n2601) );
  AND3X1 U2634 ( .IN1(n2603), .IN2(n2604), .IN3(g18), .Q(g9150) );
  NAND2X0 U2635 ( .IN1(n2605), .IN2(g605), .QN(n2604) );
  OR3X1 U2636 ( .IN1(n2605), .IN2(n2606), .IN3(g605), .Q(n2603) );
  NAND2X0 U2637 ( .IN1(n2577), .IN2(n2607), .QN(n2605) );
  NAND2X0 U2638 ( .IN1(n804), .IN2(n2608), .QN(n2607) );
  NAND2X0 U2640 ( .IN1(n2609), .IN2(n2610), .QN(n2608) );
  NAND2X0 U2642 ( .IN1(n2611), .IN2(g599), .QN(n2610) );
  NOR2X0 U2643 ( .IN1(n2612), .IN2(n2569), .QN(g9124) );
  XOR2X1 U2644 ( .IN1(g599), .IN2(n836), .Q(n2612) );
  NOR2X0 U2645 ( .IN1(n2613), .IN2(n2569), .QN(g9110) );
  XOR2X1 U2646 ( .IN1(g591), .IN2(n2614), .Q(n2613) );
  NOR2X0 U2647 ( .IN1(n2615), .IN2(n2616), .QN(n2614) );
  NOR2X0 U2648 ( .IN1(n2617), .IN2(n2552), .QN(n2616) );
  NOR2X0 U2649 ( .IN1(n2618), .IN2(n2619), .QN(n2617) );
  INVX0 U2650 ( .INP(n837), .ZN(n2615) );
  NAND3X0 U2651 ( .IN1(n804), .IN2(n1644), .IN3(n2611), .QN(n837) );
  INVX0 U2652 ( .INP(n2620), .ZN(n2611) );
  NAND2X0 U2653 ( .IN1(n2621), .IN2(n2622), .QN(g8973) );
  NAND2X0 U2655 ( .IN1(n2623), .IN2(n2624), .QN(n2622) );
  XNOR2X1 U2656 ( .IN1(n1615), .IN2(n2625), .Q(n2623) );
  NOR2X0 U2657 ( .IN1(n2626), .IN2(n2627), .QN(n2625) );
  INVX0 U2659 ( .INP(n2628), .ZN(n2627) );
  NOR2X0 U2660 ( .IN1(n2629), .IN2(g664), .QN(n2626) );
  NAND2X0 U2661 ( .IN1(n2630), .IN2(n2631), .QN(g8945) );
  NAND2X0 U2662 ( .IN1(n2632), .IN2(n2633), .QN(n2631) );
  XOR2X1 U2663 ( .IN1(n2634), .IN2(n1697), .Q(n2632) );
  NAND3X0 U2664 ( .IN1(n2635), .IN2(n2636), .IN3(n2637), .QN(n2634) );
  NAND2X0 U2665 ( .IN1(n2302), .IN2(n2638), .QN(n2636) );
  NAND3X0 U2666 ( .IN1(n2550), .IN2(n857), .IN3(n2639), .QN(n2635) );
  NAND4X0 U2667 ( .IN1(n2640), .IN2(n2641), .IN3(n921), .IN4(n2642), .QN(n857)
         );
  NOR3X0 U2668 ( .IN1(n1616), .IN2(n1694), .IN3(n1663), .QN(n2642) );
  NAND4X0 U2669 ( .IN1(n1675), .IN2(n2643), .IN3(n1694), .IN4(n2644), .QN(
        n2550) );
  AND3X1 U2670 ( .IN1(n2287), .IN2(n2237), .IN3(n2316), .Q(n2644) );
  NAND2X0 U2671 ( .IN1(n2630), .IN2(n2645), .QN(g8944) );
  NAND2X0 U2672 ( .IN1(n2646), .IN2(n2633), .QN(n2645) );
  XOR2X1 U2673 ( .IN1(n2647), .IN2(n1694), .Q(n2646) );
  NAND2X0 U2674 ( .IN1(n2637), .IN2(n2648), .QN(n2647) );
  NAND3X0 U2675 ( .IN1(n2649), .IN2(n2650), .IN3(n2651), .QN(n2648) );
  NAND2X0 U2676 ( .IN1(n2638), .IN2(g1941), .QN(n2651) );
  NAND3X0 U2677 ( .IN1(n921), .IN2(n2640), .IN3(n2652), .QN(n2650) );
  INVX0 U2678 ( .INP(n2653), .ZN(n2652) );
  NAND3X0 U2679 ( .IN1(n2287), .IN2(n2237), .IN3(n2654), .QN(n2649) );
  NAND2X0 U2680 ( .IN1(n2630), .IN2(n2655), .QN(g8943) );
  NAND2X0 U2681 ( .IN1(n2656), .IN2(n2633), .QN(n2655) );
  XOR2X1 U2682 ( .IN1(n2657), .IN2(n1663), .Q(n2656) );
  NAND3X0 U2684 ( .IN1(n2658), .IN2(n2659), .IN3(n2660), .QN(n2657) );
  NAND2X0 U2685 ( .IN1(n2661), .IN2(n2662), .QN(n2659) );
  NAND2X0 U2686 ( .IN1(n2196), .IN2(n2638), .QN(n2658) );
  NAND2X0 U2687 ( .IN1(n2630), .IN2(n2663), .QN(g8941) );
  NAND2X0 U2688 ( .IN1(n2664), .IN2(n2633), .QN(n2663) );
  XOR2X1 U2689 ( .IN1(n2665), .IN2(n2237), .Q(n2664) );
  NAND2X0 U2690 ( .IN1(n2637), .IN2(n2666), .QN(n2665) );
  NAND3X0 U2691 ( .IN1(n2667), .IN2(n2668), .IN3(n2669), .QN(n2666) );
  NAND2X0 U2692 ( .IN1(n2638), .IN2(g1932), .QN(n2669) );
  NAND2X0 U2693 ( .IN1(n2670), .IN2(n2640), .QN(n2668) );
  NOR3X0 U2694 ( .IN1(n2287), .IN2(n2316), .IN3(n1675), .QN(n2640) );
  NAND2X0 U2695 ( .IN1(n2654), .IN2(n2287), .QN(n2667) );
  INVX0 U2696 ( .INP(n2671), .ZN(n2654) );
  NAND2X0 U2697 ( .IN1(n2630), .IN2(n2672), .QN(g8940) );
  NAND2X0 U2698 ( .IN1(n2673), .IN2(n2633), .QN(n2672) );
  XOR2X1 U2700 ( .IN1(n2674), .IN2(n2287), .Q(n2673) );
  NAND2X0 U2701 ( .IN1(n2637), .IN2(n2675), .QN(n2674) );
  NAND3X0 U2702 ( .IN1(n2676), .IN2(n2671), .IN3(n2677), .QN(n2675) );
  NAND2X0 U2703 ( .IN1(n2638), .IN2(g1923), .QN(n2677) );
  NAND3X0 U2704 ( .IN1(n2316), .IN2(n1675), .IN3(n2678), .QN(n2671) );
  OR3X1 U2705 ( .IN1(n1675), .IN2(n2316), .IN3(n2679), .Q(n2676) );
  NAND2X0 U2706 ( .IN1(n2630), .IN2(n2680), .QN(g8939) );
  NAND2X0 U2707 ( .IN1(n2681), .IN2(n2633), .QN(n2680) );
  XOR2X1 U2708 ( .IN1(n2682), .IN2(n2316), .Q(n2681) );
  NAND2X0 U2709 ( .IN1(n2683), .IN2(n2637), .QN(n2682) );
  NAND3X0 U2710 ( .IN1(n2684), .IN2(n2685), .IN3(n2686), .QN(n2683) );
  NAND2X0 U2711 ( .IN1(n2638), .IN2(g1914), .QN(n2686) );
  OR2X1 U2712 ( .IN1(n2679), .IN2(n1675), .Q(n2685) );
  NAND2X0 U2713 ( .IN1(n2678), .IN2(n1675), .QN(n2684) );
  INVX0 U2714 ( .INP(n2687), .ZN(n2678) );
  NAND2X0 U2715 ( .IN1(n2630), .IN2(n2688), .QN(g8938) );
  NAND2X0 U2716 ( .IN1(n2689), .IN2(n2633), .QN(n2688) );
  XOR2X1 U2717 ( .IN1(n2690), .IN2(n1675), .Q(n2689) );
  NAND2X0 U2718 ( .IN1(n2637), .IN2(n2691), .QN(n2690) );
  NAND3X0 U2719 ( .IN1(n2687), .IN2(n2679), .IN3(n2692), .QN(n2691) );
  NAND2X0 U2720 ( .IN1(g1905), .IN2(n2638), .QN(n2692) );
  INVX0 U2721 ( .INP(n2670), .ZN(n2679) );
  NOR2X0 U2722 ( .IN1(n2653), .IN2(n1657), .QN(n2670) );
  NAND3X0 U2723 ( .IN1(n2641), .IN2(g1882), .IN3(n2661), .QN(n2653) );
  NAND2X0 U2724 ( .IN1(n2639), .IN2(n2643), .QN(n2687) );
  AND4X1 U2725 ( .IN1(n1663), .IN2(n1657), .IN3(n1616), .IN4(n2662), .Q(n2643)
         );
  NAND2X0 U2726 ( .IN1(n2630), .IN2(n2693), .QN(g8937) );
  NAND2X0 U2727 ( .IN1(n2694), .IN2(n2633), .QN(n2693) );
  XOR2X1 U2728 ( .IN1(n2695), .IN2(n1657), .Q(n2694) );
  NAND4X0 U2729 ( .IN1(n2660), .IN2(n2696), .IN3(n2697), .IN4(n2698), .QN(
        n2695) );
  NAND3X0 U2730 ( .IN1(n2639), .IN2(n2662), .IN3(g1882), .QN(n2698) );
  INVX0 U2731 ( .INP(n2641), .ZN(n2662) );
  NAND2X0 U2732 ( .IN1(n2661), .IN2(n1663), .QN(n2697) );
  NOR2X0 U2733 ( .IN1(n2638), .IN2(n1616), .QN(n2661) );
  NAND2X0 U2734 ( .IN1(n2222), .IN2(n2638), .QN(n2696) );
  AND2X1 U2735 ( .IN1(n2637), .IN2(n2699), .Q(n2660) );
  NAND3X0 U2736 ( .IN1(n1616), .IN2(n2641), .IN3(n2639), .QN(n2699) );
  NAND3X0 U2737 ( .IN1(n2589), .IN2(n2591), .IN3(n2700), .QN(n2641) );
  NAND2X0 U2738 ( .IN1(n1643), .IN2(g1814), .QN(n2700) );
  NAND2X0 U2739 ( .IN1(n2701), .IN2(n1605), .QN(n2589) );
  INVX0 U2740 ( .INP(n2602), .ZN(n2701) );
  NAND2X0 U2741 ( .IN1(n2621), .IN2(n2702), .QN(g8926) );
  NAND2X0 U2742 ( .IN1(n2703), .IN2(n2624), .QN(n2702) );
  XNOR2X1 U2743 ( .IN1(n898), .IN2(n1696), .Q(n2703) );
  AND3X1 U2744 ( .IN1(n2704), .IN2(n2705), .IN3(n2628), .Q(n898) );
  NAND2X0 U2745 ( .IN1(n2300), .IN2(n2706), .QN(n2705) );
  NAND3X0 U2746 ( .IN1(n2546), .IN2(n902), .IN3(n2629), .QN(n2704) );
  NAND4X0 U2747 ( .IN1(n2707), .IN2(n2708), .IN3(n967), .IN4(n2709), .QN(n902)
         );
  NOR3X0 U2748 ( .IN1(n1615), .IN2(n1693), .IN3(n1662), .QN(n2709) );
  NAND4X0 U2749 ( .IN1(n1676), .IN2(n2710), .IN3(n1693), .IN4(n2711), .QN(
        n2546) );
  AND3X1 U2750 ( .IN1(n2288), .IN2(n2125), .IN3(n2317), .Q(n2711) );
  NAND2X0 U2751 ( .IN1(n2621), .IN2(n2712), .QN(g8923) );
  NAND2X0 U2752 ( .IN1(n2713), .IN2(n2624), .QN(n2712) );
  XOR2X1 U2753 ( .IN1(n2714), .IN2(n1693), .Q(n2713) );
  NAND2X0 U2754 ( .IN1(n2628), .IN2(n2715), .QN(n2714) );
  NAND3X0 U2755 ( .IN1(n2716), .IN2(n2717), .IN3(n2718), .QN(n2715) );
  NAND2X0 U2756 ( .IN1(n2706), .IN2(g727), .QN(n2718) );
  NAND3X0 U2757 ( .IN1(n967), .IN2(n2707), .IN3(n2719), .QN(n2717) );
  INVX0 U2758 ( .INP(n2720), .ZN(n2719) );
  NAND3X0 U2759 ( .IN1(n2288), .IN2(n2125), .IN3(n2721), .QN(n2716) );
  NAND2X0 U2760 ( .IN1(n2621), .IN2(n2722), .QN(g8922) );
  NAND2X0 U2761 ( .IN1(n2723), .IN2(n2624), .QN(n2722) );
  XOR2X1 U2762 ( .IN1(n2724), .IN2(n1662), .Q(n2723) );
  NAND3X0 U2763 ( .IN1(n2725), .IN2(n2726), .IN3(n2727), .QN(n2724) );
  NAND2X0 U2764 ( .IN1(n2728), .IN2(n2729), .QN(n2726) );
  NAND2X0 U2765 ( .IN1(n2195), .IN2(n2706), .QN(n2725) );
  NAND2X0 U2766 ( .IN1(n2630), .IN2(n2730), .QN(g8921) );
  NAND2X0 U2767 ( .IN1(n2731), .IN2(n2633), .QN(n2730) );
  XNOR2X1 U2768 ( .IN1(n1616), .IN2(n2732), .Q(n2731) );
  NOR2X0 U2769 ( .IN1(n2733), .IN2(n2734), .QN(n2732) );
  INVX0 U2770 ( .INP(n2637), .ZN(n2734) );
  NAND2X0 U2771 ( .IN1(n2639), .IN2(n918), .QN(n2637) );
  NAND2X0 U2772 ( .IN1(n2735), .IN2(n926), .QN(n918) );
  NAND2X0 U2773 ( .IN1(n2736), .IN2(n2559), .QN(n2735) );
  NAND3X0 U2774 ( .IN1(g1814), .IN2(g1834), .IN3(n2301), .QN(n2559) );
  NAND2X0 U2775 ( .IN1(g1857), .IN2(n2737), .QN(n2736) );
  NAND2X0 U2776 ( .IN1(n1643), .IN2(n1605), .QN(n2737) );
  NOR2X0 U2777 ( .IN1(n2639), .IN2(g1878), .QN(n2733) );
  INVX0 U2778 ( .INP(n2638), .ZN(n2639) );
  NAND2X0 U2779 ( .IN1(n2738), .IN2(n2739), .QN(n2638) );
  NAND2X0 U2780 ( .IN1(n926), .IN2(g1840), .QN(n2738) );
  NAND4X0 U2781 ( .IN1(n916), .IN2(n2740), .IN3(n2587), .IN4(n2591), .QN(n2630) );
  INVX0 U2782 ( .INP(n2633), .ZN(n2740) );
  NOR2X0 U2783 ( .IN1(n812), .IN2(n2741), .QN(n2633) );
  NAND2X0 U2784 ( .IN1(n2621), .IN2(n2742), .QN(g8920) );
  NAND2X0 U2785 ( .IN1(n2743), .IN2(n2624), .QN(n2742) );
  XOR2X1 U2786 ( .IN1(n931), .IN2(n2125), .Q(n2743) );
  NAND2X0 U2787 ( .IN1(n2628), .IN2(n2744), .QN(n931) );
  NAND3X0 U2788 ( .IN1(n2745), .IN2(n2746), .IN3(n2747), .QN(n2744) );
  NAND2X0 U2789 ( .IN1(n2706), .IN2(g718), .QN(n2747) );
  NAND2X0 U2790 ( .IN1(n2748), .IN2(n2707), .QN(n2746) );
  NOR3X0 U2791 ( .IN1(n2288), .IN2(n2317), .IN3(n1676), .QN(n2707) );
  NAND2X0 U2792 ( .IN1(n2721), .IN2(n2288), .QN(n2745) );
  INVX0 U2793 ( .INP(n2749), .ZN(n2721) );
  NAND2X0 U2794 ( .IN1(n2621), .IN2(n2750), .QN(g8889) );
  NAND2X0 U2795 ( .IN1(n2751), .IN2(n2624), .QN(n2750) );
  XNOR2X1 U2796 ( .IN1(n938), .IN2(n2288), .Q(n2751) );
  AND2X1 U2797 ( .IN1(n2752), .IN2(n2628), .Q(n938) );
  NAND3X0 U2798 ( .IN1(n2753), .IN2(n2749), .IN3(n2754), .QN(n2752) );
  NAND2X0 U2799 ( .IN1(n2706), .IN2(g709), .QN(n2754) );
  NAND3X0 U2800 ( .IN1(n2317), .IN2(n1676), .IN3(n2755), .QN(n2749) );
  OR3X1 U2801 ( .IN1(n1676), .IN2(n2317), .IN3(n2756), .Q(n2753) );
  NAND2X0 U2802 ( .IN1(n2621), .IN2(n2757), .QN(g8887) );
  NAND2X0 U2803 ( .IN1(n2758), .IN2(n2624), .QN(n2757) );
  XOR2X1 U2804 ( .IN1(n2759), .IN2(n2317), .Q(n2758) );
  NAND2X0 U2805 ( .IN1(n2760), .IN2(n2628), .QN(n2759) );
  NAND3X0 U2806 ( .IN1(n2761), .IN2(n2762), .IN3(n2763), .QN(n2760) );
  NAND2X0 U2807 ( .IN1(n2706), .IN2(g700), .QN(n2763) );
  OR2X1 U2808 ( .IN1(n2756), .IN2(n1676), .Q(n2762) );
  NAND2X0 U2809 ( .IN1(n2755), .IN2(n1676), .QN(n2761) );
  INVX0 U2810 ( .INP(n2764), .ZN(n2755) );
  NAND2X0 U2811 ( .IN1(n2621), .IN2(n2765), .QN(g8885) );
  NAND2X0 U2812 ( .IN1(n2766), .IN2(n2624), .QN(n2765) );
  XOR2X1 U2813 ( .IN1(n2767), .IN2(n1676), .Q(n2766) );
  NAND2X0 U2814 ( .IN1(n2628), .IN2(n2768), .QN(n2767) );
  NAND3X0 U2815 ( .IN1(n2764), .IN2(n2756), .IN3(n2769), .QN(n2768) );
  NAND2X0 U2816 ( .IN1(g691), .IN2(n2706), .QN(n2769) );
  INVX0 U2817 ( .INP(n2748), .ZN(n2756) );
  NOR2X0 U2818 ( .IN1(n2720), .IN2(n1656), .QN(n2748) );
  NAND3X0 U2819 ( .IN1(n2708), .IN2(g668), .IN3(n2728), .QN(n2720) );
  NAND2X0 U2820 ( .IN1(n2629), .IN2(n2710), .QN(n2764) );
  AND4X1 U2821 ( .IN1(n1662), .IN2(n1656), .IN3(n1615), .IN4(n2729), .Q(n2710)
         );
  NAND2X0 U2822 ( .IN1(n2621), .IN2(n2770), .QN(g8883) );
  NAND2X0 U2823 ( .IN1(n2771), .IN2(n2624), .QN(n2770) );
  INVX0 U2824 ( .INP(n2772), .ZN(n2624) );
  XOR2X1 U2825 ( .IN1(n2773), .IN2(n1656), .Q(n2771) );
  NAND4X0 U2826 ( .IN1(n2727), .IN2(n2774), .IN3(n2775), .IN4(n2776), .QN(
        n2773) );
  NAND3X0 U2827 ( .IN1(n2629), .IN2(n2729), .IN3(g668), .QN(n2776) );
  INVX0 U2828 ( .INP(n2708), .ZN(n2729) );
  NAND2X0 U2829 ( .IN1(n2728), .IN2(n1662), .QN(n2775) );
  NOR2X0 U2830 ( .IN1(n2706), .IN2(n1615), .QN(n2728) );
  NAND2X0 U2831 ( .IN1(n2221), .IN2(n2706), .QN(n2774) );
  AND2X1 U2832 ( .IN1(n2628), .IN2(n2777), .Q(n2727) );
  NAND3X0 U2833 ( .IN1(n1615), .IN2(n2708), .IN3(n2629), .QN(n2777) );
  NAND2X0 U2834 ( .IN1(n2609), .IN2(n2778), .QN(n2708) );
  NAND2X0 U2835 ( .IN1(n1644), .IN2(g591), .QN(n2778) );
  AND2X1 U2836 ( .IN1(n2779), .IN2(n2780), .Q(n2609) );
  NAND2X0 U2837 ( .IN1(n1593), .IN2(n2618), .QN(n2780) );
  INVX0 U2838 ( .INP(n2781), .ZN(n2618) );
  NAND2X0 U2839 ( .IN1(n2629), .IN2(n958), .QN(n2628) );
  NAND2X0 U2840 ( .IN1(n2782), .IN2(n2783), .QN(n958) );
  NAND2X0 U2841 ( .IN1(n2784), .IN2(n2576), .QN(n2783) );
  NAND2X0 U2842 ( .IN1(g639), .IN2(n2785), .QN(n2784) );
  NAND2X0 U2843 ( .IN1(n1644), .IN2(n1593), .QN(n2785) );
  INVX0 U2844 ( .INP(n2706), .ZN(n2629) );
  NAND2X0 U2845 ( .IN1(n2786), .IN2(n2787), .QN(n2706) );
  NAND2X0 U2849 ( .IN1(n2782), .IN2(g617), .QN(n2787) );
  NAND4X0 U2850 ( .IN1(n2551), .IN2(n2772), .IN3(n2788), .IN4(n2576), .QN(
        n2621) );
  NAND2X0 U2851 ( .IN1(n2577), .IN2(n2789), .QN(g8820) );
  NAND2X0 U2852 ( .IN1(n2790), .IN2(g622), .QN(n2789) );
  NAND2X0 U2853 ( .IN1(n2772), .IN2(n2791), .QN(n2790) );
  NAND2X0 U2854 ( .IN1(n2788), .IN2(n2576), .QN(n2791) );
  NAND2X0 U2855 ( .IN1(n2552), .IN2(n2788), .QN(n2772) );
  INVX0 U2856 ( .INP(n804), .ZN(n2552) );
  NAND3X0 U2857 ( .IN1(n2619), .IN2(n804), .IN3(n1713), .QN(n2577) );
  INVX0 U2858 ( .INP(n2576), .ZN(n2619) );
  NAND3X0 U2862 ( .IN1(g591), .IN2(g611), .IN3(n1645), .QN(n2576) );
  NAND2X0 U2863 ( .IN1(n2792), .IN2(n2793), .QN(g8779) );
  NAND2X0 U2864 ( .IN1(n968), .IN2(g1636), .QN(n2793) );
  NAND2X0 U2865 ( .IN1(n2794), .IN2(n2795), .QN(n2792) );
  NAND2X0 U2866 ( .IN1(n2796), .IN2(n2797), .QN(g8777) );
  NAND2X0 U2868 ( .IN1(n968), .IN2(g1633), .QN(n2797) );
  NAND2X0 U2869 ( .IN1(n2798), .IN2(n2795), .QN(n2796) );
  NAND2X0 U2870 ( .IN1(n2799), .IN2(n2800), .QN(g8776) );
  NAND2X0 U2871 ( .IN1(n968), .IN2(g1630), .QN(n2800) );
  NAND2X0 U2872 ( .IN1(n2801), .IN2(n2795), .QN(n2799) );
  NOR2X0 U2873 ( .IN1(n2363), .IN2(n2802), .QN(g8775) );
  XOR2X1 U2874 ( .IN1(n2803), .IN2(n2325), .Q(n2802) );
  NAND2X0 U2875 ( .IN1(n2804), .IN2(n2805), .QN(g8774) );
  NAND2X0 U2876 ( .IN1(n968), .IN2(g1627), .QN(n2805) );
  NAND2X0 U2877 ( .IN1(n2803), .IN2(n2795), .QN(n2804) );
  NAND2X0 U2878 ( .IN1(n2806), .IN2(n2807), .QN(n2803) );
  NAND2X0 U2880 ( .IN1(n2808), .IN2(n2569), .QN(n2807) );
  XOR2X1 U2903 ( .IN1(n2809), .IN2(n1706), .Q(n2808) );
  NAND3X0 U2904 ( .IN1(n1654), .IN2(g1107), .IN3(n2810), .QN(n2809) );
  NAND2X0 U2905 ( .IN1(n2811), .IN2(n2812), .QN(g8773) );
  NAND2X0 U2906 ( .IN1(n968), .IN2(g1624), .QN(n2812) );
  NAND2X0 U2907 ( .IN1(n2813), .IN2(n2795), .QN(n2811) );
  NOR2X0 U2908 ( .IN1(n2364), .IN2(n2814), .QN(g8772) );
  XOR2X1 U2909 ( .IN1(n2801), .IN2(n2326), .Q(n2814) );
  NAND2X0 U2910 ( .IN1(n2815), .IN2(n2816), .QN(n2801) );
  NAND2X0 U2911 ( .IN1(n2817), .IN2(n2569), .QN(n2816) );
  XOR2X1 U2912 ( .IN1(n2818), .IN2(n1597), .Q(n2817) );
  NAND3X0 U2913 ( .IN1(g1107), .IN2(g1101), .IN3(n2810), .QN(n2818) );
  NAND2X0 U2914 ( .IN1(n2819), .IN2(n2820), .QN(g8771) );
  NAND2X0 U2915 ( .IN1(n968), .IN2(g1621), .QN(n2820) );
  NAND2X0 U2916 ( .IN1(n2821), .IN2(n2795), .QN(n2819) );
  NAND2X0 U2917 ( .IN1(n2822), .IN2(n2823), .QN(g8770) );
  NAND2X0 U2918 ( .IN1(n968), .IN2(g1615), .QN(n2823) );
  NAND2X0 U2919 ( .IN1(n2824), .IN2(n2795), .QN(n2822) );
  NOR2X0 U2920 ( .IN1(n2362), .IN2(n2825), .QN(g8769) );
  XOR2X1 U2921 ( .IN1(n2824), .IN2(n2327), .Q(n2825) );
  NAND2X0 U2922 ( .IN1(n2826), .IN2(n2827), .QN(n2824) );
  NAND2X0 U2923 ( .IN1(n2828), .IN2(n2569), .QN(n2827) );
  XOR2X1 U2924 ( .IN1(n2829), .IN2(n1618), .Q(n2828) );
  NAND2X0 U2925 ( .IN1(n2810), .IN2(n2830), .QN(n2829) );
  NOR2X0 U2926 ( .IN1(n2365), .IN2(n2831), .QN(g8768) );
  XOR2X1 U2927 ( .IN1(n2798), .IN2(n2328), .Q(n2831) );
  NAND2X0 U2928 ( .IN1(n2832), .IN2(n2833), .QN(n2798) );
  NAND2X0 U2929 ( .IN1(n2834), .IN2(n2569), .QN(n2833) );
  XNOR2X1 U2930 ( .IN1(n1660), .IN2(n2835), .Q(n2834) );
  NOR2X0 U2931 ( .IN1(n2836), .IN2(g1101), .QN(n2835) );
  NOR2X0 U2932 ( .IN1(n2363), .IN2(n2837), .QN(g8767) );
  XOR2X1 U2933 ( .IN1(n2821), .IN2(n2264), .Q(n2837) );
  NAND2X0 U2934 ( .IN1(n2838), .IN2(n2839), .QN(n2821) );
  NAND2X0 U2935 ( .IN1(n2840), .IN2(n2569), .QN(n2839) );
  XNOR2X1 U2936 ( .IN1(n1708), .IN2(n2841), .Q(n2840) );
  NOR2X0 U2937 ( .IN1(g1101), .IN2(n2842), .QN(n2841) );
  NOR2X0 U2938 ( .IN1(n2364), .IN2(n2843), .QN(g8766) );
  XOR2X1 U2939 ( .IN1(n2794), .IN2(n2262), .Q(n2843) );
  NAND2X0 U2940 ( .IN1(n2844), .IN2(n2845), .QN(n2794) );
  NAND2X0 U2941 ( .IN1(n2846), .IN2(n2569), .QN(n2845) );
  XNOR2X1 U2942 ( .IN1(n1617), .IN2(n2847), .Q(n2846) );
  NOR2X0 U2943 ( .IN1(n1654), .IN2(n2836), .QN(n2847) );
  NAND3X0 U2944 ( .IN1(n1614), .IN2(g1110), .IN3(n1658), .QN(n2836) );
  NOR2X0 U2945 ( .IN1(n2362), .IN2(n2848), .QN(g8765) );
  XOR2X1 U2946 ( .IN1(n2813), .IN2(n2263), .Q(n2848) );
  NAND2X0 U2947 ( .IN1(n2849), .IN2(n2850), .QN(n2813) );
  NAND2X0 U2948 ( .IN1(n2851), .IN2(n2569), .QN(n2850) );
  XNOR2X1 U2949 ( .IN1(n1705), .IN2(n2852), .Q(n2851) );
  NOR2X0 U2950 ( .IN1(n1654), .IN2(n2842), .QN(n2852) );
  NAND3X0 U2951 ( .IN1(n1658), .IN2(g1107), .IN3(n1677), .QN(n2842) );
  NAND3X0 U2952 ( .IN1(n2853), .IN2(n2854), .IN3(n2788), .QN(g8649) );
  NAND2X0 U2953 ( .IN1(n2855), .IN2(g736), .QN(n2854) );
  NAND2X0 U2954 ( .IN1(n1016), .IN2(g664), .QN(n2853) );
  NAND2X0 U2955 ( .IN1(n2856), .IN2(n2857), .QN(g8631) );
  NAND2X0 U2956 ( .IN1(n2606), .IN2(n2858), .QN(n2857) );
  NAND3X0 U2957 ( .IN1(n2859), .IN2(g826), .IN3(n2860), .QN(n2858) );
  NAND2X0 U2958 ( .IN1(n2861), .IN2(n2862), .QN(n2860) );
  OR2X1 U2959 ( .IN1(n2332), .IN2(n1622), .Q(n2862) );
  OR2X1 U2960 ( .IN1(n2242), .IN2(n1717), .Q(n2861) );
  NAND2X0 U2961 ( .IN1(n2863), .IN2(n2864), .QN(n2859) );
  NAND2X0 U2962 ( .IN1(g810), .IN2(g814), .QN(n2864) );
  NAND2X0 U2963 ( .IN1(g818), .IN2(g822), .QN(n2863) );
  NAND2X0 U2964 ( .IN1(n2865), .IN2(n2788), .QN(n2856) );
  NAND2X0 U2965 ( .IN1(n2866), .IN2(n2867), .QN(n2865) );
  NAND2X0 U2966 ( .IN1(n2868), .IN2(g636), .QN(n2867) );
  NAND3X0 U2967 ( .IN1(g4892), .IN2(n2869), .IN3(n2870), .QN(n2868) );
  XOR2X1 U2968 ( .IN1(n2871), .IN2(n2872), .Q(n2870) );
  NAND2X0 U2969 ( .IN1(n2873), .IN2(n2874), .QN(n2872) );
  NAND2X0 U2970 ( .IN1(n2781), .IN2(g639), .QN(n2874) );
  NAND3X0 U2971 ( .IN1(n1609), .IN2(n2620), .IN3(n1692), .QN(n2873) );
  NAND2X0 U2972 ( .IN1(g255), .IN2(g622), .QN(n2871) );
  NAND3X0 U2973 ( .IN1(n1644), .IN2(n2875), .IN3(n1609), .QN(n2869) );
  NAND2X0 U2974 ( .IN1(g591), .IN2(n2876), .QN(n2875) );
  NAND2X0 U2975 ( .IN1(n1593), .IN2(g617), .QN(n2876) );
  OR2X1 U2976 ( .IN1(n2779), .IN2(g622), .Q(n2866) );
  NAND2X0 U2977 ( .IN1(n2877), .IN2(n2878), .QN(g8566) );
  NAND2X0 U2978 ( .IN1(n1653), .IN2(g1669), .QN(n2878) );
  NAND2X0 U2979 ( .IN1(g1690), .IN2(g1687), .QN(n2877) );
  NAND2X0 U2980 ( .IN1(n2879), .IN2(n2880), .QN(g8565) );
  NAND2X0 U2981 ( .IN1(n1653), .IN2(g1666), .QN(n2880) );
  NAND2X0 U2982 ( .IN1(g1690), .IN2(g1684), .QN(n2879) );
  NAND2X0 U2983 ( .IN1(n2881), .IN2(n2882), .QN(g8564) );
  NAND2X0 U2984 ( .IN1(n1653), .IN2(g1663), .QN(n2882) );
  NAND2X0 U2985 ( .IN1(g1690), .IN2(g1681), .QN(n2881) );
  NAND2X0 U2986 ( .IN1(n2883), .IN2(n2884), .QN(g8563) );
  NAND2X0 U2987 ( .IN1(n1653), .IN2(g1660), .QN(n2884) );
  NAND2X0 U2988 ( .IN1(g1690), .IN2(g1678), .QN(n2883) );
  NAND2X0 U2989 ( .IN1(n2885), .IN2(n2886), .QN(g8562) );
  NAND2X0 U2990 ( .IN1(n1653), .IN2(g1657), .QN(n2886) );
  NAND2X0 U2991 ( .IN1(g1690), .IN2(g1675), .QN(n2885) );
  NAND2X0 U2992 ( .IN1(n2887), .IN2(n2888), .QN(g8561) );
  NAND2X0 U2993 ( .IN1(n1653), .IN2(g1654), .QN(n2888) );
  NAND2X0 U2994 ( .IN1(g1690), .IN2(g1672), .QN(n2887) );
  NAND3X0 U2995 ( .IN1(n2889), .IN2(n2587), .IN3(n2890), .QN(g8559) );
  NAND2X0 U2996 ( .IN1(n2891), .IN2(g1878), .QN(n2890) );
  NOR2X0 U2997 ( .IN1(n2892), .IN2(n2569), .QN(g8505) );
  XOR2X1 U2998 ( .IN1(g617), .IN2(n2893), .Q(n2892) );
  NOR2X0 U2999 ( .IN1(n2894), .IN2(n2895), .QN(n2893) );
  NOR2X0 U3000 ( .IN1(n2300), .IN2(n1016), .QN(n2895) );
  NOR2X0 U3001 ( .IN1(g617), .IN2(n2786), .QN(n2894) );
  NAND4X0 U3002 ( .IN1(n1609), .IN2(n2782), .IN3(n2896), .IN4(n1644), .QN(
        n2786) );
  NOR2X0 U3003 ( .IN1(n1607), .IN2(g605), .QN(n2896) );
  NAND2X0 U3004 ( .IN1(n2897), .IN2(n2898), .QN(g8435) );
  NAND2X0 U3005 ( .IN1(n2899), .IN2(g736), .QN(n2898) );
  NAND2X0 U3006 ( .IN1(n2855), .IN2(g727), .QN(n2897) );
  NAND2X0 U3007 ( .IN1(n2900), .IN2(n2901), .QN(g8434) );
  NAND2X0 U3008 ( .IN1(n2899), .IN2(g727), .QN(n2901) );
  NAND2X0 U3009 ( .IN1(n2855), .IN2(g718), .QN(n2900) );
  NAND2X0 U3010 ( .IN1(n2902), .IN2(n2903), .QN(g8433) );
  NAND2X0 U3011 ( .IN1(n2899), .IN2(g718), .QN(n2903) );
  NAND2X0 U3012 ( .IN1(n2855), .IN2(g709), .QN(n2902) );
  NAND2X0 U3013 ( .IN1(n2904), .IN2(n2905), .QN(g8432) );
  NAND2X0 U3014 ( .IN1(n2899), .IN2(g709), .QN(n2905) );
  NAND2X0 U3015 ( .IN1(n2855), .IN2(g700), .QN(n2904) );
  NAND2X0 U3016 ( .IN1(n2906), .IN2(n2907), .QN(g8431) );
  NAND2X0 U3017 ( .IN1(n2899), .IN2(g700), .QN(n2907) );
  NAND2X0 U3018 ( .IN1(n2855), .IN2(g691), .QN(n2906) );
  NAND2X0 U3019 ( .IN1(n2908), .IN2(n2909), .QN(g8430) );
  NAND2X0 U3020 ( .IN1(n2899), .IN2(g691), .QN(n2909) );
  NAND2X0 U3021 ( .IN1(n2855), .IN2(g682), .QN(n2908) );
  NAND2X0 U3022 ( .IN1(n2910), .IN2(n2911), .QN(g8429) );
  NAND2X0 U3023 ( .IN1(n2899), .IN2(g682), .QN(n2911) );
  NAND2X0 U3024 ( .IN1(n2855), .IN2(g673), .QN(n2910) );
  NAND2X0 U3025 ( .IN1(n2912), .IN2(n2913), .QN(g8428) );
  NAND2X0 U3026 ( .IN1(n2899), .IN2(g673), .QN(n2913) );
  NOR2X0 U3027 ( .IN1(n2855), .IN2(n2606), .QN(n2899) );
  INVX0 U3028 ( .INP(n2788), .ZN(n2606) );
  NAND2X0 U3029 ( .IN1(n2855), .IN2(g664), .QN(n2912) );
  INVX0 U3030 ( .INP(n1016), .ZN(n2855) );
  NAND3X0 U3031 ( .IN1(n2782), .IN2(g617), .IN3(n1609), .QN(n1016) );
  NOR2X0 U3032 ( .IN1(n2914), .IN2(n2569), .QN(g8384) );
  XOR2X1 U3033 ( .IN1(n2915), .IN2(n2301), .Q(n2914) );
  NAND2X0 U3034 ( .IN1(n2739), .IN2(n2889), .QN(n2915) );
  NAND2X0 U3035 ( .IN1(n2916), .IN2(g1950), .QN(n2889) );
  INVX0 U3036 ( .INP(n929), .ZN(n2739) );
  NOR3X0 U3037 ( .IN1(n2917), .IN2(n367), .IN3(g1822), .QN(n929) );
  NAND2X0 U3038 ( .IN1(n1665), .IN2(n2918), .QN(g8352) );
  NAND2X0 U3039 ( .IN1(n1669), .IN2(n2918), .QN(g8349) );
  NAND2X0 U3040 ( .IN1(n1671), .IN2(n2918), .QN(g8347) );
  NAND2X0 U3041 ( .IN1(n2361), .IN2(n2918), .QN(g8340) );
  NAND2X0 U3042 ( .IN1(n1666), .IN2(n2918), .QN(g8335) );
  NAND2X0 U3043 ( .IN1(n1672), .IN2(n2918), .QN(g8331) );
  NAND2X0 U3044 ( .IN1(n1664), .IN2(n2918), .QN(g8328) );
  NAND2X0 U3045 ( .IN1(n1673), .IN2(n2918), .QN(g8323) );
  NAND2X0 U3046 ( .IN1(n1667), .IN2(n2918), .QN(g8318) );
  NAND2X0 U3047 ( .IN1(n1674), .IN2(n2918), .QN(g8316) );
  NAND2X0 U3048 ( .IN1(n1668), .IN2(n2918), .QN(g8313) );
  INVX0 U3049 ( .INP(g82), .ZN(n2918) );
  NAND2X0 U3050 ( .IN1(n2919), .IN2(n2920), .QN(g8288) );
  NAND2X0 U3051 ( .IN1(n2921), .IN2(g1950), .QN(n2920) );
  NAND2X0 U3052 ( .IN1(n2916), .IN2(g1941), .QN(n2919) );
  NAND2X0 U3053 ( .IN1(n2922), .IN2(n2923), .QN(g8287) );
  NAND2X0 U3054 ( .IN1(n2921), .IN2(g1941), .QN(n2923) );
  NAND2X0 U3055 ( .IN1(n2916), .IN2(g1932), .QN(n2922) );
  NAND2X0 U3056 ( .IN1(n2924), .IN2(n2925), .QN(g8286) );
  NAND2X0 U3057 ( .IN1(n2921), .IN2(g1932), .QN(n2925) );
  NAND2X0 U3058 ( .IN1(n2916), .IN2(g1923), .QN(n2924) );
  NAND2X0 U3059 ( .IN1(n2926), .IN2(n2927), .QN(g8285) );
  NAND2X0 U3060 ( .IN1(n2921), .IN2(g1923), .QN(n2927) );
  NAND2X0 U3061 ( .IN1(n2916), .IN2(g1914), .QN(n2926) );
  NAND2X0 U3062 ( .IN1(n2928), .IN2(n2929), .QN(g8284) );
  NAND2X0 U3063 ( .IN1(n2921), .IN2(g1914), .QN(n2929) );
  NAND2X0 U3064 ( .IN1(n2916), .IN2(g1905), .QN(n2928) );
  NAND2X0 U3065 ( .IN1(n2930), .IN2(n2931), .QN(g8283) );
  NAND2X0 U3066 ( .IN1(n2921), .IN2(g1905), .QN(n2931) );
  NAND2X0 U3067 ( .IN1(n2916), .IN2(g1896), .QN(n2930) );
  NAND2X0 U3068 ( .IN1(n2932), .IN2(n2933), .QN(g8282) );
  NAND2X0 U3069 ( .IN1(n2921), .IN2(g1896), .QN(n2933) );
  NAND2X0 U3070 ( .IN1(n2916), .IN2(g1887), .QN(n2932) );
  NAND2X0 U3071 ( .IN1(n2934), .IN2(n2935), .QN(g8281) );
  NAND2X0 U3072 ( .IN1(n2921), .IN2(g1887), .QN(n2935) );
  NOR2X0 U3073 ( .IN1(n2741), .IN2(n2916), .QN(n2921) );
  NAND2X0 U3074 ( .IN1(n2916), .IN2(g1878), .QN(n2934) );
  INVX0 U3075 ( .INP(n2891), .ZN(n2916) );
  NAND3X0 U3076 ( .IN1(n926), .IN2(g1840), .IN3(n1655), .QN(n2891) );
  NOR2X0 U3077 ( .IN1(n1712), .IN2(n2936), .QN(g8260) );
  NOR2X0 U3078 ( .IN1(n1630), .IN2(n2936), .QN(g8254) );
  NOR2X0 U3079 ( .IN1(n1591), .IN2(n2936), .QN(g8250) );
  NOR2X0 U3080 ( .IN1(n2937), .IN2(n2938), .QN(g8245) );
  XOR2X1 U3081 ( .IN1(n1716), .IN2(n2939), .Q(n2938) );
  AND2X1 U3082 ( .IN1(g822), .IN2(n1090), .Q(n2939) );
  NOR3X0 U3083 ( .IN1(n2940), .IN2(n2941), .IN3(n2942), .QN(g8244) );
  NOR2X0 U3084 ( .IN1(n2943), .IN2(g4181), .QN(n2942) );
  NOR2X0 U3085 ( .IN1(n2134), .IN2(n2944), .QN(n2943) );
  NAND2X0 U3086 ( .IN1(n2945), .IN2(n2946), .QN(g8194) );
  NAND2X0 U3087 ( .IN1(n968), .IN2(g1512), .QN(n2946) );
  NAND2X0 U3088 ( .IN1(n2947), .IN2(n2795), .QN(n2945) );
  XOR2X1 U3089 ( .IN1(n2948), .IN2(n4124), .Q(n2947) );
  OR3X1 U3091 ( .IN1(n1658), .IN2(n1677), .IN3(n2949), .Q(n2948) );
  NAND2X0 U3093 ( .IN1(n2950), .IN2(n2951), .QN(g8193) );
  NAND2X0 U3095 ( .IN1(n968), .IN2(g1639), .QN(n2951) );
  NAND2X0 U3097 ( .IN1(n2952), .IN2(n2795), .QN(n2950) );
  XOR2X1 U3099 ( .IN1(test_so4), .IN2(n2953), .Q(n2952) );
  NOR2X0 U3100 ( .IN1(n2954), .IN2(n2949), .QN(n2953) );
  NAND2X0 U3101 ( .IN1(n1654), .IN2(n1614), .QN(n2949) );
  INVX0 U3102 ( .INP(n2810), .ZN(n2954) );
  NOR2X0 U3103 ( .IN1(g1110), .IN2(n1658), .QN(n2810) );
  NOR2X0 U3104 ( .IN1(n2955), .IN2(g1713), .QN(g8173) );
  NOR2X0 U3105 ( .IN1(n2956), .IN2(n2957), .QN(n2955) );
  NOR2X0 U3106 ( .IN1(n2340), .IN2(n2958), .QN(n2957) );
  NOR2X0 U3107 ( .IN1(n1055), .IN2(n1054), .QN(n2958) );
  AND3X1 U3108 ( .IN1(n1056), .IN2(g1801), .IN3(n1055), .Q(n2956) );
  NAND3X0 U3109 ( .IN1(g1801), .IN2(g1806), .IN3(n1057), .QN(n1055) );
  AND2X1 U3110 ( .IN1(n2959), .IN2(g1796), .Q(n1057) );
  NOR2X0 U3111 ( .IN1(n1604), .IN2(n2936), .QN(g8147) );
  NAND2X0 U3112 ( .IN1(n2960), .IN2(g109), .QN(n2936) );
  NAND3X0 U3113 ( .IN1(n2961), .IN2(DFF_436_n1), .IN3(n2962), .QN(n2960) );
  NOR2X0 U3114 ( .IN1(n2365), .IN2(n2963), .QN(g8060) );
  XOR2X1 U3115 ( .IN1(g6002), .IN2(n2258), .Q(n2963) );
  NOR2X0 U3116 ( .IN1(n2363), .IN2(n2964), .QN(g8059) );
  XOR2X1 U3117 ( .IN1(g6042), .IN2(n2255), .Q(n2964) );
  NOR2X0 U3118 ( .IN1(n2364), .IN2(n2965), .QN(g8055) );
  XNOR2X1 U3119 ( .IN1(n2966), .IN2(n2329), .Q(n2965) );
  NOR2X0 U3120 ( .IN1(n2362), .IN2(n2967), .QN(g8054) );
  XOR2X1 U3121 ( .IN1(g6015), .IN2(n2345), .Q(n2967) );
  NOR2X0 U3122 ( .IN1(n2365), .IN2(n2968), .QN(g8053) );
  XOR2X1 U3123 ( .IN1(g6045), .IN2(n2254), .Q(n2968) );
  NOR2X0 U3125 ( .IN1(n2363), .IN2(n2969), .QN(g8052) );
  XOR2X1 U3126 ( .IN1(n2970), .IN2(n2256), .Q(n2969) );
  NOR2X0 U3127 ( .IN1(n2364), .IN2(n2971), .QN(g8051) );
  XOR2X1 U3128 ( .IN1(n2972), .IN2(n2260), .Q(n2971) );
  NOR2X0 U3129 ( .IN1(n2362), .IN2(n2973), .QN(g8050) );
  XOR2X1 U3130 ( .IN1(g6026), .IN2(n2346), .Q(n2973) );
  NOR2X0 U3131 ( .IN1(n2365), .IN2(n2974), .QN(g8049) );
  XOR2X1 U3132 ( .IN1(g6049), .IN2(n2257), .Q(n2974) );
  NOR2X0 U3133 ( .IN1(n2363), .IN2(n2975), .QN(g8048) );
  XOR2X1 U3134 ( .IN1(g5996), .IN2(n2278), .Q(n2975) );
  NOR2X0 U3135 ( .IN1(n2364), .IN2(n2976), .QN(g8047) );
  XOR2X1 U3136 ( .IN1(g6035), .IN2(n1704), .Q(n2976) );
  NOR2X0 U3137 ( .IN1(n2362), .IN2(n2977), .QN(g8046) );
  XOR2X1 U3138 ( .IN1(n2978), .IN2(n2261), .Q(n2977) );
  NOR2X0 U3139 ( .IN1(n2365), .IN2(n2979), .QN(g8045) );
  XOR2X1 U3140 ( .IN1(n2980), .IN2(n2330), .Q(n2979) );
  NOR2X0 U3141 ( .IN1(n2363), .IN2(n2981), .QN(g8044) );
  XOR2X1 U3142 ( .IN1(g6038), .IN2(n2253), .Q(n2981) );
  NOR2X0 U3143 ( .IN1(n2364), .IN2(n2982), .QN(g8043) );
  XOR2X1 U3144 ( .IN1(n2983), .IN2(n2331), .Q(n2982) );
  NOR2X0 U3145 ( .IN1(n2362), .IN2(n2984), .QN(g8042) );
  XOR2X1 U3146 ( .IN1(n2985), .IN2(n1703), .Q(n2984) );
  NOR2X0 U3147 ( .IN1(n2365), .IN2(n2986), .QN(g8041) );
  XOR2X1 U3148 ( .IN1(n2987), .IN2(n2293), .Q(n2986) );
  NOR2X0 U3149 ( .IN1(n2363), .IN2(n2988), .QN(g8040) );
  XOR2X1 U3150 ( .IN1(n2989), .IN2(n2294), .Q(n2988) );
  NOR2X0 U3151 ( .IN1(n2364), .IN2(n2990), .QN(g8039) );
  XOR2X1 U3152 ( .IN1(n2991), .IN2(n2295), .Q(n2990) );
  NOR2X0 U3153 ( .IN1(n2937), .IN2(n2992), .QN(g8024) );
  XOR2X1 U3154 ( .IN1(n2344), .IN2(n1090), .Q(n2992) );
  NOR2X0 U3155 ( .IN1(n2940), .IN2(n2993), .QN(g8019) );
  XOR2X1 U3156 ( .IN1(n2134), .IN2(n1093), .Q(n2993) );
  NOR2X0 U3157 ( .IN1(g1713), .IN2(n2994), .QN(g7930) );
  XOR2X1 U3158 ( .IN1(n2339), .IN2(n1056), .Q(n2994) );
  NOR2X0 U3159 ( .IN1(n2362), .IN2(n2995), .QN(g7843) );
  XOR2X1 U3160 ( .IN1(g6000), .IN2(n2259), .Q(n2995) );
  NOR3X0 U3161 ( .IN1(n2937), .IN2(n1096), .IN3(n1090), .QN(g7709) );
  NOR3X0 U3162 ( .IN1(n2940), .IN2(n1098), .IN3(n1093), .QN(g7705) );
  NAND3X0 U3163 ( .IN1(n2788), .IN2(n2574), .IN3(n2996), .QN(g7660) );
  NAND2X0 U3164 ( .IN1(n2997), .IN2(g654), .QN(n2996) );
  NOR3X0 U3165 ( .IN1(n2998), .IN2(n2999), .IN3(n3000), .QN(g7632) );
  AND2X1 U3166 ( .IN1(n3001), .IN2(n2119), .Q(n3000) );
  NAND3X0 U3167 ( .IN1(n3002), .IN2(n3003), .IN3(n2788), .QN(g7626) );
  NAND2X0 U3168 ( .IN1(n2574), .IN2(g639), .QN(n3003) );
  NAND3X0 U3169 ( .IN1(n2782), .IN2(n3004), .IN3(n1692), .QN(n3002) );
  NAND3X0 U3170 ( .IN1(n2620), .IN2(n2781), .IN3(n2551), .QN(n3004) );
  AND2X1 U3172 ( .IN1(n2779), .IN2(n3005), .Q(n2551) );
  NAND2X0 U3173 ( .IN1(n1593), .IN2(g599), .QN(n3005) );
  NAND3X0 U3174 ( .IN1(n1607), .IN2(g605), .IN3(n1644), .QN(n2779) );
  NAND2X0 U3175 ( .IN1(n1607), .IN2(g599), .QN(n2781) );
  NAND2X0 U3176 ( .IN1(g591), .IN2(g605), .QN(n2620) );
  NOR2X0 U3177 ( .IN1(n3006), .IN2(n2998), .QN(g7590) );
  NOR2X0 U3178 ( .IN1(n3007), .IN2(g1231), .QN(n3006) );
  NOR2X0 U3179 ( .IN1(n3008), .IN2(n2998), .QN(g7586) );
  NOR2X0 U3180 ( .IN1(n3009), .IN2(n1107), .QN(n3008) );
  AND3X1 U3181 ( .IN1(n3010), .IN2(g1223), .IN3(n2999), .Q(n1107) );
  NOR2X0 U3182 ( .IN1(n2118), .IN2(n3007), .QN(n3009) );
  NOR2X0 U3183 ( .IN1(n3010), .IN2(n3001), .QN(n3007) );
  NOR2X0 U3184 ( .IN1(n2998), .IN2(n3011), .QN(g7581) );
  XOR2X1 U3185 ( .IN1(n2120), .IN2(n2999), .Q(n3011) );
  NOR2X0 U3186 ( .IN1(n3001), .IN2(n2119), .QN(n2999) );
  NAND2X0 U3187 ( .IN1(n3012), .IN2(n3013), .QN(n3001) );
  INVX0 U3188 ( .INP(n3014), .ZN(n3013) );
  NAND2X0 U3189 ( .IN1(n2347), .IN2(g109), .QN(n2998) );
  NOR3X0 U3190 ( .IN1(g1713), .IN2(n3015), .IN3(n3021), .QN(g7541) );
  NOR2X0 U3191 ( .IN1(n68), .IN2(g1796), .QN(n3021) );
  AND2X1 U3192 ( .IN1(g1796), .IN2(n1056), .Q(n3015) );
  NAND2X0 U3193 ( .IN1(n3028), .IN2(n2788), .QN(g7441) );
  XOR2X1 U3194 ( .IN1(n1612), .IN2(g627), .Q(n3028) );
  NAND2X0 U3195 ( .IN1(n3032), .IN2(n3039), .QN(g7303) );
  NAND2X0 U3196 ( .IN1(n3043), .IN2(test_so6), .QN(n3039) );
  NAND2X0 U3197 ( .IN1(n3012), .IN2(g1265), .QN(n3032) );
  NAND2X0 U3198 ( .IN1(n3049), .IN2(n3052), .QN(g7302) );
  NAND2X0 U3199 ( .IN1(n3043), .IN2(g1265), .QN(n3052) );
  NAND2X0 U3200 ( .IN1(n3012), .IN2(g1260), .QN(n3049) );
  NAND2X0 U3201 ( .IN1(n3060), .IN2(n3063), .QN(g7301) );
  NAND2X0 U3202 ( .IN1(n3043), .IN2(g1260), .QN(n3063) );
  NAND2X0 U3203 ( .IN1(n3012), .IN2(g1255), .QN(n3060) );
  NAND2X0 U3204 ( .IN1(n3066), .IN2(n3067), .QN(g7300) );
  NAND2X0 U3205 ( .IN1(n3043), .IN2(g1255), .QN(n3067) );
  NAND2X0 U3206 ( .IN1(n3012), .IN2(g1250), .QN(n3066) );
  NAND2X0 U3207 ( .IN1(n3068), .IN2(n3069), .QN(g7299) );
  NAND2X0 U3208 ( .IN1(n3043), .IN2(g1250), .QN(n3069) );
  NAND2X0 U3209 ( .IN1(n3012), .IN2(g1245), .QN(n3068) );
  NAND2X0 U3210 ( .IN1(n3070), .IN2(n3071), .QN(g7298) );
  NAND2X0 U3211 ( .IN1(n3043), .IN2(g1245), .QN(n3071) );
  NAND2X0 U3212 ( .IN1(n3012), .IN2(g1240), .QN(n3070) );
  NAND2X0 U3213 ( .IN1(n3072), .IN2(n3073), .QN(g7297) );
  NAND2X0 U3214 ( .IN1(n3043), .IN2(g1240), .QN(n3073) );
  NAND2X0 U3215 ( .IN1(n3012), .IN2(g1235), .QN(n3072) );
  NAND2X0 U3216 ( .IN1(n3074), .IN2(n3075), .QN(g7296) );
  NAND2X0 U3217 ( .IN1(n3043), .IN2(g1235), .QN(n3075) );
  NAND2X0 U3218 ( .IN1(n3012), .IN2(g1275), .QN(n3074) );
  NAND2X0 U3219 ( .IN1(n3076), .IN2(n3077), .QN(g7295) );
  NAND2X0 U3220 ( .IN1(n3043), .IN2(g1280), .QN(n3077) );
  NAND2X0 U3221 ( .IN1(n3012), .IN2(g1284), .QN(n3076) );
  NAND2X0 U3222 ( .IN1(n3078), .IN2(n3079), .QN(g7294) );
  NAND2X0 U3223 ( .IN1(n3043), .IN2(g1284), .QN(n3079) );
  NAND2X0 U3224 ( .IN1(n3012), .IN2(g1292), .QN(n3078) );
  NAND2X0 U3225 ( .IN1(n3080), .IN2(n3081), .QN(g7293) );
  NAND2X0 U3226 ( .IN1(n3043), .IN2(g1292), .QN(n3081) );
  NAND2X0 U3227 ( .IN1(n3012), .IN2(g1296), .QN(n3080) );
  NAND2X0 U3228 ( .IN1(n3082), .IN2(n3083), .QN(g7292) );
  NAND2X0 U3229 ( .IN1(n3043), .IN2(g1296), .QN(n3083) );
  NAND2X0 U3230 ( .IN1(n3012), .IN2(g1300), .QN(n3082) );
  NAND2X0 U3231 ( .IN1(n3084), .IN2(n3085), .QN(g7291) );
  NAND2X0 U3232 ( .IN1(n3043), .IN2(g1300), .QN(n3085) );
  NAND2X0 U3233 ( .IN1(n3012), .IN2(g1304), .QN(n3084) );
  NAND2X0 U3234 ( .IN1(n3086), .IN2(n3087), .QN(g7290) );
  NAND2X0 U3235 ( .IN1(n3043), .IN2(g1304), .QN(n3087) );
  NAND2X0 U3236 ( .IN1(n3012), .IN2(test_so6), .QN(n3086) );
  NAND2X0 U3237 ( .IN1(n3088), .IN2(n3089), .QN(g7257) );
  NAND2X0 U3238 ( .IN1(n2795), .IN2(g1077), .QN(n3089) );
  OR2X1 U3239 ( .IN1(n2795), .IN2(n2201), .Q(n3088) );
  NAND2X0 U3240 ( .IN1(n3090), .IN2(n3091), .QN(g7244) );
  NAND2X0 U3241 ( .IN1(n2795), .IN2(g1071), .QN(n3091) );
  OR2X1 U3242 ( .IN1(n2795), .IN2(n2203), .Q(n3090) );
  NAND2X0 U3243 ( .IN1(n2361), .IN2(n3092), .QN(g7219) );
  NAND2X0 U3244 ( .IN1(n1672), .IN2(n3092), .QN(g7204) );
  NOR2X0 U3245 ( .IN1(n2937), .IN2(n3093), .QN(g7202) );
  XOR2X1 U3246 ( .IN1(n2343), .IN2(n1123), .Q(n3093) );
  NOR2X0 U3247 ( .IN1(n2940), .IN2(n3094), .QN(g7191) );
  XOR2X1 U3248 ( .IN1(n2133), .IN2(n1125), .Q(n3094) );
  NAND2X0 U3249 ( .IN1(n1673), .IN2(n3092), .QN(g7189) );
  NAND2X0 U3250 ( .IN1(n1674), .IN2(n3092), .QN(g7183) );
  NAND2X0 U3251 ( .IN1(n1671), .IN2(n3092), .QN(g7143) );
  AND3X1 U3252 ( .IN1(n2788), .IN2(n2574), .IN3(n3095), .Q(g7137) );
  NAND2X0 U3253 ( .IN1(n2997), .IN2(n3096), .QN(n3095) );
  NAND2X0 U3254 ( .IN1(n3097), .IN2(g650), .QN(n3096) );
  AND3X1 U3255 ( .IN1(n2788), .IN2(n2574), .IN3(n3098), .Q(g7134) );
  NAND2X0 U3256 ( .IN1(n3097), .IN2(n3099), .QN(n3098) );
  NAND2X0 U3257 ( .IN1(n3100), .IN2(n3062), .QN(n3099) );
  NAND2X0 U3258 ( .IN1(n1612), .IN2(g627), .QN(n3100) );
  INVX0 U3259 ( .INP(n2782), .ZN(n2574) );
  NOR2X0 U3260 ( .IN1(g654), .IN2(n2997), .QN(n2782) );
  OR2X1 U3261 ( .IN1(g650), .IN2(n3097), .Q(n2997) );
  NAND3X0 U3262 ( .IN1(n1612), .IN2(g627), .IN3(n4111), .QN(n3097) );
  NAND2X0 U3263 ( .IN1(n1610), .IN2(n3101), .QN(g7133) );
  XOR2X1 U3264 ( .IN1(g1766), .IN2(n1054), .Q(n3101) );
  NAND2X0 U3265 ( .IN1(n3102), .IN2(n3103), .QN(g7032) );
  NAND2X0 U3266 ( .IN1(g109), .IN2(g123), .QN(n3103) );
  INVX0 U3267 ( .INP(n1132), .ZN(n3102) );
  NOR4X0 U3268 ( .IN1(n3104), .IN2(n3105), .IN3(n3106), .IN4(n3107), .QN(n1132) );
  NAND4X0 U3269 ( .IN1(n1704), .IN2(n1613), .IN3(g6786), .IN4(n1137), .QN(
        n3107) );
  NAND4X0 U3270 ( .IN1(g166), .IN2(g182), .IN3(g174), .IN4(g170), .QN(n3106)
         );
  NAND4X0 U3271 ( .IN1(n2280), .IN2(n2279), .IN3(n2278), .IN4(n2259), .QN(
        n3105) );
  NAND4X0 U3272 ( .IN1(n2258), .IN2(n2255), .IN3(n2254), .IN4(n2253), .QN(
        n3104) );
  NOR2X0 U3273 ( .IN1(n3108), .IN2(g1713), .QN(g6983) );
  NOR2X0 U3274 ( .IN1(n3109), .IN2(n3110), .QN(n3108) );
  NOR2X0 U3275 ( .IN1(n1702), .IN2(n68), .QN(n3110) );
  AND2X1 U3276 ( .IN1(n2959), .IN2(n263), .Q(n68) );
  NOR3X0 U3277 ( .IN1(n3111), .IN2(n2341), .IN3(n2959), .QN(n3109) );
  NOR3X0 U3278 ( .IN1(n3112), .IN2(n1659), .IN3(n3113), .QN(n2959) );
  NAND2X0 U3279 ( .IN1(n3114), .IN2(n3115), .QN(g6934) );
  OR2X1 U3280 ( .IN1(n3116), .IN2(n2175), .Q(n3115) );
  NAND2X0 U3281 ( .IN1(n3116), .IN2(g170), .QN(n3114) );
  NAND2X0 U3282 ( .IN1(n3117), .IN2(n3118), .QN(g6930) );
  NAND2X0 U3283 ( .IN1(n2795), .IN2(g1074), .QN(n3118) );
  OR2X1 U3284 ( .IN1(n2795), .IN2(n2228), .Q(n3117) );
  NAND2X0 U3285 ( .IN1(n3119), .IN2(n3120), .QN(g6929) );
  NAND2X0 U3286 ( .IN1(n3121), .IN2(g302), .QN(n3120) );
  OR2X1 U3287 ( .IN1(n3121), .IN2(n2279), .Q(n3119) );
  NAND2X0 U3288 ( .IN1(n3122), .IN2(n3123), .QN(g6928) );
  NAND2X0 U3289 ( .IN1(n3121), .IN2(g281), .QN(n3123) );
  NAND2X0 U3290 ( .IN1(n3116), .IN2(g174), .QN(n3122) );
  NAND2X0 U3291 ( .IN1(n3124), .IN2(n3125), .QN(g6924) );
  NAND2X0 U3292 ( .IN1(n2795), .IN2(g1098), .QN(n3125) );
  OR2X1 U3293 ( .IN1(n2795), .IN2(n2229), .Q(n3124) );
  NAND2X0 U3294 ( .IN1(n3126), .IN2(n3127), .QN(g6923) );
  NAND2X0 U3295 ( .IN1(n3121), .IN2(g299), .QN(n3127) );
  NAND2X0 U3296 ( .IN1(n3116), .IN2(g166), .QN(n3126) );
  NAND2X0 U3297 ( .IN1(n3128), .IN2(n3129), .QN(g6922) );
  NAND2X0 U3298 ( .IN1(n3121), .IN2(g278), .QN(n3129) );
  OR2X1 U3299 ( .IN1(n3121), .IN2(n2258), .Q(n3128) );
  NAND2X0 U3300 ( .IN1(n3130), .IN2(n3131), .QN(g6918) );
  NAND2X0 U3301 ( .IN1(n2795), .IN2(g1095), .QN(n3131) );
  NAND2X0 U3302 ( .IN1(test_so2), .IN2(n968), .QN(n3130) );
  NAND2X0 U3303 ( .IN1(n3132), .IN2(n3133), .QN(g6916) );
  NAND2X0 U3304 ( .IN1(n3121), .IN2(g296), .QN(n3133) );
  OR2X1 U3305 ( .IN1(n3121), .IN2(n2254), .Q(n3132) );
  NAND2X0 U3306 ( .IN1(n3134), .IN2(n3135), .QN(g6915) );
  NAND2X0 U3307 ( .IN1(n3121), .IN2(g275), .QN(n3135) );
  OR2X1 U3308 ( .IN1(n3121), .IN2(n2259), .Q(n3134) );
  NAND2X0 U3309 ( .IN1(n3136), .IN2(n3137), .QN(g6912) );
  NAND2X0 U3310 ( .IN1(n2795), .IN2(g1092), .QN(n3137) );
  OR2X1 U3311 ( .IN1(n2795), .IN2(n2267), .Q(n3136) );
  NAND2X0 U3312 ( .IN1(n3138), .IN2(n3139), .QN(g6911) );
  NAND2X0 U3313 ( .IN1(n3121), .IN2(g293), .QN(n3139) );
  OR2X1 U3314 ( .IN1(n3121), .IN2(n2255), .Q(n3138) );
  NAND2X0 U3315 ( .IN1(n3140), .IN2(n3141), .QN(g6910) );
  NAND2X0 U3316 ( .IN1(n3121), .IN2(g272), .QN(n3141) );
  NAND2X0 U3317 ( .IN1(n3116), .IN2(g153), .QN(n3140) );
  NAND2X0 U3318 ( .IN1(n3142), .IN2(n3143), .QN(g6909) );
  NAND2X0 U3319 ( .IN1(n3144), .IN2(g1868), .QN(n3143) );
  NAND2X0 U3320 ( .IN1(n3145), .IN2(n3146), .QN(g6908) );
  NAND2X0 U3321 ( .IN1(n2795), .IN2(g1089), .QN(n3146) );
  NAND2X0 U3322 ( .IN1(test_so8), .IN2(n968), .QN(n3145) );
  NAND2X0 U3323 ( .IN1(n3147), .IN2(n3148), .QN(g6907) );
  NAND2X0 U3324 ( .IN1(n3121), .IN2(g290), .QN(n3148) );
  OR2X1 U3325 ( .IN1(n3121), .IN2(n2253), .Q(n3147) );
  NAND2X0 U3326 ( .IN1(n3149), .IN2(n3150), .QN(g6906) );
  NAND2X0 U3327 ( .IN1(n3121), .IN2(g269), .QN(n3150) );
  OR2X1 U3328 ( .IN1(n3121), .IN2(n2280), .Q(n3149) );
  NAND2X0 U3329 ( .IN1(n3151), .IN2(n3152), .QN(g6902) );
  NAND2X0 U3330 ( .IN1(n2795), .IN2(g1086), .QN(n3152) );
  OR2X1 U3331 ( .IN1(n2795), .IN2(n2306), .Q(n3151) );
  NAND2X0 U3332 ( .IN1(n3153), .IN2(n3154), .QN(g6901) );
  NAND2X0 U3333 ( .IN1(n3121), .IN2(g287), .QN(n3154) );
  OR2X1 U3334 ( .IN1(n3121), .IN2(n1704), .Q(n3153) );
  NAND2X0 U3335 ( .IN1(n3155), .IN2(n3156), .QN(g6900) );
  NAND2X0 U3336 ( .IN1(n3121), .IN2(g266), .QN(n3156) );
  NAND2X0 U3337 ( .IN1(n3116), .IN2(g178), .QN(n3155) );
  NAND2X0 U3338 ( .IN1(n3157), .IN2(n3158), .QN(g6898) );
  NAND2X0 U3339 ( .IN1(n2795), .IN2(g1083), .QN(n3158) );
  OR2X1 U3340 ( .IN1(n2795), .IN2(n1871), .Q(n3157) );
  NAND2X0 U3341 ( .IN1(n3159), .IN2(n3160), .QN(g6897) );
  NAND2X0 U3342 ( .IN1(n3121), .IN2(g263), .QN(n3160) );
  INVX0 U3343 ( .INP(n3116), .ZN(n3121) );
  NAND2X0 U3344 ( .IN1(n3116), .IN2(g182), .QN(n3159) );
  NAND2X0 U3345 ( .IN1(n3161), .IN2(g109), .QN(n3116) );
  NAND2X0 U3346 ( .IN1(n1613), .IN2(n1137), .QN(n3161) );
  NOR2X0 U3347 ( .IN1(n2569), .IN2(n4121), .QN(n1137) );
  NAND2X0 U3348 ( .IN1(n3162), .IN2(n3163), .QN(g6895) );
  NAND2X0 U3349 ( .IN1(n2795), .IN2(g1080), .QN(n3163) );
  OR2X1 U3350 ( .IN1(n2795), .IN2(n2304), .Q(n3162) );
  NAND2X0 U3351 ( .IN1(n3164), .IN2(n3165), .QN(g6894) );
  NAND2X0 U3352 ( .IN1(test_so7), .IN2(n2795), .QN(n3165) );
  OR2X1 U3353 ( .IN1(n2795), .IN2(n2350), .Q(n3164) );
  NOR2X0 U3354 ( .IN1(g1696), .IN2(g4089), .QN(g6842) );
  NOR2X0 U3355 ( .IN1(n1629), .IN2(n2362), .QN(g6841) );
  NOR2X0 U3356 ( .IN1(n1598), .IN2(n2363), .QN(g6840) );
  NOR2X0 U3357 ( .IN1(n1711), .IN2(n2364), .QN(g6839) );
  NOR2X0 U3358 ( .IN1(n4118), .IN2(n2362), .QN(g6834) );
  NOR2X0 U3359 ( .IN1(n4125), .IN2(n2365), .QN(g6830) );
  NOR2X0 U3360 ( .IN1(n4126), .IN2(n2363), .QN(g6828) );
  NOR2X0 U3361 ( .IN1(n4127), .IN2(n2364), .QN(g6820) );
  NOR2X0 U3362 ( .IN1(n3166), .IN2(n3167), .QN(g6795) );
  NOR2X0 U3363 ( .IN1(n3168), .IN2(n39), .QN(n3166) );
  INVX0 U3364 ( .INP(n3144), .ZN(n39) );
  NAND2X0 U3365 ( .IN1(n2336), .IN2(n3169), .QN(n3144) );
  NOR2X0 U3366 ( .IN1(n2336), .IN2(n3169), .QN(n3168) );
  NAND2X0 U3367 ( .IN1(n4128), .IN2(n3170), .QN(g6755) );
  AND3X1 U3368 ( .IN1(n3171), .IN2(g109), .IN3(n4121), .Q(g6747) );
  NAND2X0 U3369 ( .IN1(n4129), .IN2(DFF_452_n1), .QN(n3171) );
  NOR3X0 U3370 ( .IN1(n2937), .IN2(n1150), .IN3(n1123), .QN(g6733) );
  NOR3X0 U3371 ( .IN1(n2940), .IN2(n1152), .IN3(n1125), .QN(g6728) );
  NAND2X0 U3372 ( .IN1(n3172), .IN2(n3173), .QN(g6679) );
  NAND2X0 U3373 ( .IN1(n1155), .IN2(n1154), .QN(n3173) );
  AND4X1 U3374 ( .IN1(n1159), .IN2(g1419), .IN3(g6234), .IN4(n3174), .Q(n1154)
         );
  NOR4X0 U3375 ( .IN1(n2263), .IN2(n2262), .IN3(n1710), .IN4(n1627), .QN(n3174) );
  AND4X1 U3376 ( .IN1(n2264), .IN2(n2160), .IN3(n3175), .IN4(n3176), .Q(n1155)
         );
  NOR4X0 U3377 ( .IN1(n2328), .IN2(n2327), .IN3(n2326), .IN4(n2325), .QN(n3176) );
  NOR2X0 U3378 ( .IN1(g1415), .IN2(g1407), .QN(n3175) );
  NAND2X0 U3379 ( .IN1(g109), .IN2(g1), .QN(n3172) );
  NAND2X0 U3380 ( .IN1(n1701), .IN2(n3177), .QN(g6672) );
  NAND2X0 U3381 ( .IN1(n3178), .IN2(n3179), .QN(g6656) );
  NAND2X0 U3382 ( .IN1(n1162), .IN2(n1161), .QN(n3179) );
  AND4X1 U3383 ( .IN1(n2354), .IN2(g1453), .IN3(n1159), .IN4(n3180), .Q(n1161)
         );
  NOR4X0 U3384 ( .IN1(n2295), .IN2(n2294), .IN3(n2293), .IN4(n1707), .QN(n3180) );
  NOR2X0 U3385 ( .IN1(n2365), .IN2(n2139), .QN(n2354) );
  AND4X1 U3386 ( .IN1(n2281), .IN2(n2261), .IN3(n3181), .IN4(n3182), .Q(n1162)
         );
  NOR4X0 U3387 ( .IN1(n2331), .IN2(n2330), .IN3(n2329), .IN4(g1458), .QN(n3182) );
  NOR2X0 U3388 ( .IN1(g1486), .IN2(g1466), .QN(n3181) );
  NAND2X0 U3389 ( .IN1(g109), .IN2(g4), .QN(n3178) );
  NOR2X0 U3390 ( .IN1(n1666), .IN2(n3183), .QN(g6653) );
  NOR2X0 U3391 ( .IN1(n1664), .IN2(n3183), .QN(g6638) );
  NOR2X0 U3392 ( .IN1(n1667), .IN2(n3183), .QN(g6627) );
  NOR2X0 U3393 ( .IN1(n1668), .IN2(n3183), .QN(g6621) );
  NAND2X0 U3394 ( .IN1(n3184), .IN2(n3185), .QN(g6551) );
  NAND2X0 U3395 ( .IN1(n3186), .IN2(g1546), .QN(n3185) );
  OR2X1 U3396 ( .IN1(n3186), .IN2(n2331), .Q(n3184) );
  NAND2X0 U3397 ( .IN1(n3187), .IN2(n3188), .QN(g6546) );
  NAND2X0 U3398 ( .IN1(n3186), .IN2(g1564), .QN(n3188) );
  NAND2X0 U3399 ( .IN1(n3189), .IN2(g1453), .QN(n3187) );
  NAND2X0 U3400 ( .IN1(n3190), .IN2(n3191), .QN(g6545) );
  NAND2X0 U3401 ( .IN1(n3186), .IN2(g1543), .QN(n3191) );
  OR2X1 U3402 ( .IN1(n3186), .IN2(n2261), .Q(n3190) );
  NAND2X0 U3403 ( .IN1(n3192), .IN2(n3193), .QN(g6542) );
  NAND2X0 U3404 ( .IN1(n3186), .IN2(g1561), .QN(n3193) );
  NAND2X0 U3405 ( .IN1(n3189), .IN2(g1458), .QN(n3192) );
  NAND2X0 U3406 ( .IN1(n3194), .IN2(n3195), .QN(g6541) );
  NAND2X0 U3407 ( .IN1(n3186), .IN2(g1540), .QN(n3195) );
  NAND2X0 U3408 ( .IN1(n3189), .IN2(g1486), .QN(n3194) );
  NAND2X0 U3409 ( .IN1(n3196), .IN2(n3197), .QN(g6538) );
  NAND2X0 U3410 ( .IN1(n3186), .IN2(g1558), .QN(n3197) );
  OR2X1 U3411 ( .IN1(n3186), .IN2(n2330), .Q(n3196) );
  NAND2X0 U3412 ( .IN1(n3198), .IN2(n3199), .QN(g6537) );
  NAND2X0 U3413 ( .IN1(n3186), .IN2(g1537), .QN(n3199) );
  OR2X1 U3414 ( .IN1(n3186), .IN2(n2329), .Q(n3198) );
  NAND2X0 U3415 ( .IN1(n3200), .IN2(n3201), .QN(g6534) );
  NAND2X0 U3416 ( .IN1(n3186), .IN2(g1555), .QN(n3201) );
  NAND2X0 U3417 ( .IN1(n3189), .IN2(g1466), .QN(n3200) );
  NAND2X0 U3418 ( .IN1(n3202), .IN2(n3203), .QN(g6533) );
  NAND2X0 U3419 ( .IN1(n3186), .IN2(g1534), .QN(n3203) );
  NAND2X0 U3420 ( .IN1(n3189), .IN2(g1494), .QN(n3202) );
  NOR2X0 U3421 ( .IN1(n1665), .IN2(n3183), .QN(g6531) );
  NAND2X0 U3422 ( .IN1(n3204), .IN2(n3205), .QN(g6529) );
  OR2X1 U3423 ( .IN1(n3189), .IN2(n2143), .Q(n3205) );
  OR2X1 U3424 ( .IN1(n3186), .IN2(n2295), .Q(n3204) );
  NAND2X0 U3425 ( .IN1(n3206), .IN2(n3207), .QN(g6528) );
  NAND2X0 U3426 ( .IN1(n3186), .IN2(g1531), .QN(n3207) );
  OR2X1 U3427 ( .IN1(n3186), .IN2(n2281), .Q(n3206) );
  NOR2X0 U3428 ( .IN1(n1669), .IN2(n3183), .QN(g6526) );
  NOR2X0 U3429 ( .IN1(g1713), .IN2(n3208), .QN(g6525) );
  XOR2X1 U3430 ( .IN1(g1786), .IN2(n3111), .Q(n3208) );
  NAND2X0 U3431 ( .IN1(n3209), .IN2(n3210), .QN(g6524) );
  NAND2X0 U3432 ( .IN1(n3186), .IN2(g1589), .QN(n3210) );
  OR2X1 U3433 ( .IN1(n3186), .IN2(n2327), .Q(n3209) );
  NAND2X0 U3434 ( .IN1(n3211), .IN2(n3212), .QN(g6523) );
  NAND2X0 U3435 ( .IN1(n3186), .IN2(g1549), .QN(n3212) );
  OR2X1 U3436 ( .IN1(n3186), .IN2(n2294), .Q(n3211) );
  NAND2X0 U3437 ( .IN1(n3213), .IN2(n3214), .QN(g6522) );
  NAND2X0 U3438 ( .IN1(n3186), .IN2(g1528), .QN(n3214) );
  OR2X1 U3439 ( .IN1(n3186), .IN2(n2139), .Q(n3213) );
  NOR3X0 U3440 ( .IN1(g1713), .IN2(n2355), .IN3(n3215), .QN(g6516) );
  NOR2X0 U3441 ( .IN1(n3216), .IN2(g1781), .QN(n3215) );
  INVX0 U3442 ( .INP(n3111), .ZN(n2355) );
  NAND2X0 U3443 ( .IN1(n3216), .IN2(g1781), .QN(n3111) );
  NAND2X0 U3444 ( .IN1(n3217), .IN2(n3218), .QN(g6515) );
  NAND2X0 U3445 ( .IN1(n3186), .IN2(g1607), .QN(n3218) );
  NAND2X0 U3446 ( .IN1(n3189), .IN2(g1448), .QN(n3217) );
  NAND2X0 U3447 ( .IN1(n3219), .IN2(n3220), .QN(g6514) );
  OR2X1 U3448 ( .IN1(n3189), .IN2(n2141), .Q(n3220) );
  NAND2X0 U3449 ( .IN1(n3189), .IN2(g1407), .QN(n3219) );
  NAND2X0 U3450 ( .IN1(n3221), .IN2(n3222), .QN(g6513) );
  NAND2X0 U3451 ( .IN1(n3186), .IN2(g1524), .QN(n3222) );
  OR2X1 U3452 ( .IN1(n3186), .IN2(n1707), .Q(n3221) );
  NOR2X0 U3453 ( .IN1(n3223), .IN2(g1713), .QN(g6508) );
  NOR2X0 U3454 ( .IN1(n3224), .IN2(n3225), .QN(n3223) );
  NOR2X0 U3455 ( .IN1(n1715), .IN2(n3216), .QN(n3225) );
  NOR2X0 U3456 ( .IN1(n3113), .IN2(n1054), .QN(n3216) );
  AND3X1 U3457 ( .IN1(n3226), .IN2(n3113), .IN3(test_so5), .Q(n3224) );
  NAND2X0 U3458 ( .IN1(n3227), .IN2(n3228), .QN(g6507) );
  NAND2X0 U3459 ( .IN1(n3186), .IN2(g1604), .QN(n3228) );
  OR2X1 U3460 ( .IN1(n3186), .IN2(n2328), .Q(n3227) );
  NAND2X0 U3461 ( .IN1(n3229), .IN2(n3230), .QN(g6506) );
  NAND2X0 U3462 ( .IN1(n3186), .IN2(g1583), .QN(n3230) );
  NAND2X0 U3463 ( .IN1(n3189), .IN2(g1424), .QN(n3229) );
  NOR2X0 U3464 ( .IN1(n3231), .IN2(g1713), .QN(g6502) );
  XNOR2X1 U3465 ( .IN1(test_so5), .IN2(n3226), .Q(n3231) );
  NOR2X0 U3466 ( .IN1(n1054), .IN2(n2334), .QN(n3226) );
  NAND2X0 U3467 ( .IN1(n3232), .IN2(n3233), .QN(g6501) );
  NAND2X0 U3468 ( .IN1(n3186), .IN2(g1601), .QN(n3233) );
  OR2X1 U3469 ( .IN1(n3186), .IN2(n2326), .Q(n3232) );
  NAND2X0 U3470 ( .IN1(n3234), .IN2(n3235), .QN(g6500) );
  NAND2X0 U3471 ( .IN1(n3186), .IN2(g1580), .QN(n3235) );
  OR2X1 U3472 ( .IN1(n3186), .IN2(n2160), .Q(n3234) );
  NAND2X0 U3473 ( .IN1(n3236), .IN2(n3237), .QN(g6481) );
  OR2X1 U3474 ( .IN1(n3189), .IN2(n2144), .Q(n3237) );
  OR2X1 U3475 ( .IN1(n3186), .IN2(n2325), .Q(n3236) );
  NAND2X0 U3476 ( .IN1(n3238), .IN2(n3239), .QN(g6480) );
  OR2X1 U3477 ( .IN1(n3189), .IN2(n2147), .Q(n3239) );
  NAND2X0 U3478 ( .IN1(n3189), .IN2(g1419), .QN(n3238) );
  NAND2X0 U3479 ( .IN1(n3240), .IN2(n3241), .QN(g6479) );
  NAND2X0 U3480 ( .IN1(n3186), .IN2(g1595), .QN(n3241) );
  OR2X1 U3481 ( .IN1(n3186), .IN2(n2263), .Q(n3240) );
  NAND2X0 U3482 ( .IN1(n3242), .IN2(n3243), .QN(g6478) );
  NAND2X0 U3483 ( .IN1(n3186), .IN2(g1574), .QN(n3243) );
  OR2X1 U3484 ( .IN1(n3186), .IN2(n1627), .Q(n3242) );
  NOR2X0 U3485 ( .IN1(n3244), .IN2(n3167), .QN(g6471) );
  NOR2X0 U3486 ( .IN1(n3245), .IN2(n3169), .QN(n3244) );
  AND2X1 U3487 ( .IN1(n2338), .IN2(n3033), .Q(n3169) );
  NOR2X0 U3488 ( .IN1(n2338), .IN2(n3033), .QN(n3245) );
  NAND2X0 U3489 ( .IN1(n3246), .IN2(n3247), .QN(g6470) );
  NAND2X0 U3490 ( .IN1(n3186), .IN2(g1592), .QN(n3247) );
  OR2X1 U3491 ( .IN1(n3186), .IN2(n2264), .Q(n3246) );
  NAND2X0 U3492 ( .IN1(n3248), .IN2(n3249), .QN(g6469) );
  OR2X1 U3493 ( .IN1(n3189), .IN2(n2154), .Q(n3249) );
  OR2X1 U3494 ( .IN1(n3186), .IN2(n1710), .Q(n3248) );
  NAND2X0 U3495 ( .IN1(n3250), .IN2(n3251), .QN(g6468) );
  NAND2X0 U3496 ( .IN1(n3186), .IN2(g1567), .QN(n3251) );
  NAND2X0 U3497 ( .IN1(n3189), .IN2(g1415), .QN(n3250) );
  INVX0 U3498 ( .INP(n3186), .ZN(n3189) );
  NOR2X0 U3499 ( .IN1(n2363), .IN2(n1159), .QN(n3186) );
  NOR2X0 U3500 ( .IN1(n2364), .IN2(n3252), .QN(g6439) );
  XOR3X1 U3501 ( .IN1(n2278), .IN2(n2277), .IN3(n3253), .Q(n3252) );
  XNOR2X1 U3502 ( .IN1(n2279), .IN2(n2280), .Q(n3253) );
  NOR2X0 U3503 ( .IN1(n3254), .IN2(n3255), .QN(g6392) );
  NOR2X0 U3504 ( .IN1(n2362), .IN2(n2961), .QN(n3255) );
  INVX0 U3505 ( .INP(g881), .ZN(n2961) );
  NOR2X0 U3506 ( .IN1(n1678), .IN2(n2362), .QN(g6333) );
  NOR2X0 U3507 ( .IN1(n4122), .IN2(n2365), .QN(g6332) );
  NAND2X0 U3508 ( .IN1(n3256), .IN2(n3257), .QN(g6243) );
  INVX0 U3509 ( .INP(n2937), .ZN(n3257) );
  XNOR2X1 U3510 ( .IN1(n1717), .IN2(n2242), .Q(n3256) );
  NOR2X0 U3511 ( .IN1(n1710), .IN2(n2363), .QN(g6224) );
  NOR2X0 U3512 ( .IN1(n1627), .IN2(n2364), .QN(g6205) );
  NOR2X0 U3513 ( .IN1(n4129), .IN2(n2556), .QN(g6179) );
  NAND2X0 U3514 ( .IN1(n280), .IN2(n3258), .QN(n2556) );
  NOR2X0 U3515 ( .IN1(n2365), .IN2(n1619), .QN(n280) );
  NAND2X0 U3516 ( .IN1(n3259), .IN2(n3260), .QN(g6155) );
  NAND2X0 U3517 ( .IN1(g4076), .IN2(g1690), .QN(n3260) );
  NAND3X0 U3518 ( .IN1(g1700), .IN2(g1707), .IN3(n1653), .QN(n3259) );
  NOR2X0 U3519 ( .IN1(n2937), .IN2(n3261), .QN(g6126) );
  XOR2X1 U3520 ( .IN1(n2332), .IN2(n2567), .Q(n3261) );
  NOR2X0 U3521 ( .IN1(n2940), .IN2(n3262), .QN(g6123) );
  XOR2X1 U3522 ( .IN1(n2132), .IN2(n1193), .Q(n3262) );
  NAND2X0 U3523 ( .IN1(n3263), .IN2(n3264), .QN(g6099) );
  NAND2X0 U3524 ( .IN1(n3265), .IN2(g342), .QN(n3264) );
  NAND2X0 U3525 ( .IN1(n3266), .IN2(g1074), .QN(n3263) );
  NAND2X0 U3526 ( .IN1(n3267), .IN2(n3268), .QN(g6096) );
  NAND2X0 U3527 ( .IN1(n3265), .IN2(g366), .QN(n3268) );
  NAND2X0 U3528 ( .IN1(n3266), .IN2(g1098), .QN(n3267) );
  NAND2X0 U3529 ( .IN1(n3269), .IN2(n3270), .QN(g6093) );
  NAND2X0 U3530 ( .IN1(n3265), .IN2(g363), .QN(n3270) );
  NAND2X0 U3531 ( .IN1(n3266), .IN2(g1095), .QN(n3269) );
  NAND2X0 U3532 ( .IN1(n3271), .IN2(n3272), .QN(g6088) );
  NAND2X0 U3533 ( .IN1(n3265), .IN2(g360), .QN(n3272) );
  NAND2X0 U3534 ( .IN1(n3266), .IN2(g1092), .QN(n3271) );
  NAND2X0 U3535 ( .IN1(n3273), .IN2(n3274), .QN(g6080) );
  NAND2X0 U3536 ( .IN1(n3265), .IN2(g357), .QN(n3274) );
  NAND2X0 U3537 ( .IN1(n3266), .IN2(g1089), .QN(n3273) );
  NAND2X0 U3538 ( .IN1(n3275), .IN2(n3276), .QN(g6071) );
  NAND2X0 U3539 ( .IN1(n3265), .IN2(g354), .QN(n3276) );
  NAND2X0 U3540 ( .IN1(n3266), .IN2(g1086), .QN(n3275) );
  NAND2X0 U3541 ( .IN1(n3277), .IN2(n3278), .QN(g6068) );
  NAND2X0 U3542 ( .IN1(n3265), .IN2(g351), .QN(n3278) );
  NAND2X0 U3543 ( .IN1(n3266), .IN2(g1083), .QN(n3277) );
  NAND2X0 U3544 ( .IN1(n3279), .IN2(n3280), .QN(g6059) );
  NAND2X0 U3545 ( .IN1(n3265), .IN2(g348), .QN(n3280) );
  NAND2X0 U3546 ( .IN1(n3266), .IN2(g1080), .QN(n3279) );
  NAND2X0 U3547 ( .IN1(n3281), .IN2(n3282), .QN(g6054) );
  NAND2X0 U3548 ( .IN1(n3265), .IN2(g336), .QN(n3282) );
  NAND2X0 U3549 ( .IN1(test_so7), .IN2(n3266), .QN(n3281) );
  NAND2X0 U3550 ( .IN1(n3283), .IN2(n3284), .QN(g6049) );
  NAND2X0 U3551 ( .IN1(n2569), .IN2(g549), .QN(n3283) );
  NAND2X0 U3552 ( .IN1(n3285), .IN2(n3286), .QN(g6045) );
  NAND2X0 U3553 ( .IN1(n2569), .IN2(g575), .QN(n3285) );
  NAND2X0 U3554 ( .IN1(n3287), .IN2(n3288), .QN(g6042) );
  NAND2X0 U3555 ( .IN1(n2569), .IN2(g572), .QN(n3287) );
  NAND2X0 U3556 ( .IN1(n2844), .IN2(n3289), .QN(g6038) );
  NAND2X0 U3557 ( .IN1(n2569), .IN2(g569), .QN(n3289) );
  NAND2X0 U3558 ( .IN1(n2832), .IN2(n3290), .QN(g6035) );
  NAND2X0 U3559 ( .IN1(n2569), .IN2(g566), .QN(n3290) );
  NAND2X0 U3560 ( .IN1(n2815), .IN2(n3291), .QN(g6026) );
  NAND2X0 U3561 ( .IN1(n2569), .IN2(g563), .QN(n3291) );
  NAND2X0 U3562 ( .IN1(n2806), .IN2(n3292), .QN(g6015) );
  NAND2X0 U3563 ( .IN1(n2569), .IN2(g560), .QN(n3292) );
  NAND2X0 U3564 ( .IN1(n2849), .IN2(n3293), .QN(g6002) );
  NAND2X0 U3565 ( .IN1(n2569), .IN2(g557), .QN(n3293) );
  NAND2X0 U3566 ( .IN1(n2838), .IN2(n3294), .QN(g6000) );
  NAND2X0 U3567 ( .IN1(n2569), .IN2(g554), .QN(n3294) );
  NAND2X0 U3568 ( .IN1(n2826), .IN2(n3295), .QN(g5996) );
  NAND2X0 U3569 ( .IN1(n2569), .IN2(g546), .QN(n3295) );
  NAND2X0 U3570 ( .IN1(n3296), .IN2(n3297), .QN(g5918) );
  OR2X1 U3571 ( .IN1(n2365), .IN2(n1613), .Q(n3297) );
  NAND2X0 U3572 ( .IN1(n3298), .IN2(n3299), .QN(g5914) );
  NAND2X0 U3573 ( .IN1(n3265), .IN2(g345), .QN(n3299) );
  NAND2X0 U3574 ( .IN1(n3266), .IN2(g1077), .QN(n3298) );
  NAND2X0 U3575 ( .IN1(n3300), .IN2(n3301), .QN(g5910) );
  NAND2X0 U3576 ( .IN1(n3265), .IN2(g339), .QN(n3301) );
  NAND2X0 U3577 ( .IN1(n3266), .IN2(g1071), .QN(n3300) );
  NAND2X0 U3578 ( .IN1(n3302), .IN2(n3303), .QN(g5770) );
  OR3X1 U3579 ( .IN1(g1453), .IN2(n2363), .IN3(n3304), .Q(n3303) );
  NAND2X0 U3580 ( .IN1(g6180), .IN2(n3304), .QN(n3302) );
  XOR3X1 U3581 ( .IN1(n2293), .IN2(n2281), .IN3(n1707), .Q(n3304) );
  NOR2X0 U3582 ( .IN1(n2363), .IN2(n1628), .QN(g6180) );
  NOR2X0 U3583 ( .IN1(n3305), .IN2(n3306), .QN(g5763) );
  NOR2X0 U3584 ( .IN1(n4131), .IN2(n2362), .QN(n3306) );
  NAND2X0 U3585 ( .IN1(n3307), .IN2(n3308), .QN(g5755) );
  NAND3X0 U3586 ( .IN1(n1603), .IN2(g109), .IN3(n3309), .QN(n3308) );
  NAND2X0 U3587 ( .IN1(g6334), .IN2(n3310), .QN(n3307) );
  INVX0 U3588 ( .INP(n3309), .ZN(n3310) );
  XOR3X1 U3589 ( .IN1(n1678), .IN2(n1619), .IN3(n3311), .Q(n3309) );
  NAND2X0 U3590 ( .IN1(n2276), .IN2(n2558), .QN(n3311) );
  NAND2X0 U3591 ( .IN1(n1619), .IN2(n3258), .QN(n2558) );
  AND4X1 U3592 ( .IN1(n3312), .IN2(n3313), .IN3(n3314), .IN4(n3315), .Q(n3258)
         );
  AND4X1 U3593 ( .IN1(n3316), .IN2(n1711), .IN3(n1629), .IN4(n1678), .Q(n3315)
         );
  AND3X1 U3594 ( .IN1(n1598), .IN2(n4112), .IN3(n1603), .Q(n3316) );
  NOR4X0 U3595 ( .IN1(n3317), .IN2(g1386), .IN3(g219), .IN4(g192), .QN(n3314)
         );
  NAND3X0 U3596 ( .IN1(n2122), .IN2(n2121), .IN3(n2123), .QN(n3317) );
  NOR4X0 U3597 ( .IN1(n3318), .IN2(g1371), .IN3(g243), .IN4(g1383), .QN(n3313)
         );
  NAND3X0 U3598 ( .IN1(n2283), .IN2(n2282), .IN3(n2284), .QN(n3318) );
  AND4X1 U3599 ( .IN1(n4125), .IN2(n3319), .IN3(n4122), .IN4(n4118), .Q(n3312)
         );
  AND2X1 U3600 ( .IN1(n4126), .IN2(n4127), .Q(n3319) );
  NOR2X0 U3601 ( .IN1(n2364), .IN2(n1603), .QN(g6334) );
  AND3X1 U3602 ( .IN1(g743), .IN2(g109), .IN3(g744), .Q(g5659) );
  AND3X1 U3603 ( .IN1(g741), .IN2(g109), .IN3(g742), .Q(g5658) );
  NOR2X0 U3604 ( .IN1(n3320), .IN2(n3321), .QN(g5556) );
  OR4X1 U3605 ( .IN1(g1781), .IN2(n3113), .IN3(n3112), .IN4(n1626), .Q(n3321)
         );
  NAND3X0 U3606 ( .IN1(g1776), .IN2(g1766), .IN3(test_so5), .QN(n3113) );
  NAND4X0 U3607 ( .IN1(g1690), .IN2(g1801), .IN3(g1806), .IN4(g1707), .QN(
        n3320) );
  NOR2X0 U3608 ( .IN1(n2567), .IN2(n3322), .QN(g5543) );
  NOR2X0 U3609 ( .IN1(n3323), .IN2(n3324), .QN(n3322) );
  NOR2X0 U3610 ( .IN1(n1717), .IN2(g5849), .QN(n3324) );
  OR2X1 U3611 ( .IN1(n2937), .IN2(n2242), .Q(g5849) );
  NOR2X0 U3612 ( .IN1(n1622), .IN2(n2937), .QN(n3323) );
  NAND3X0 U3613 ( .IN1(g746), .IN2(g745), .IN3(g109), .QN(n2937) );
  NOR3X0 U3614 ( .IN1(n1717), .IN2(n2242), .IN3(n1622), .QN(n2567) );
  NOR3X0 U3615 ( .IN1(n2940), .IN2(n1213), .IN3(n1193), .QN(g5536) );
  NAND2X0 U3616 ( .IN1(n3325), .IN2(n3326), .QN(g5529) );
  NAND2X0 U3617 ( .IN1(g4940), .IN2(g4174), .QN(n3326) );
  NAND3X0 U3618 ( .IN1(n3327), .IN2(g4173), .IN3(n2130), .QN(n3325) );
  NAND2X0 U3619 ( .IN1(n3296), .IN2(n3328), .QN(g5445) );
  OR2X1 U3620 ( .IN1(n2362), .IN2(n2232), .Q(n3328) );
  NAND2X0 U3621 ( .IN1(n3296), .IN2(n3329), .QN(g5421) );
  OR2X1 U3622 ( .IN1(n2365), .IN2(n2233), .Q(n3329) );
  INVX0 U3623 ( .INP(n1195), .ZN(n3296) );
  NAND2X0 U3624 ( .IN1(n3330), .IN2(n3331), .QN(g5404) );
  NAND2X0 U3625 ( .IN1(n2795), .IN2(g1713), .QN(n3331) );
  NAND2X0 U3626 ( .IN1(n968), .IN2(g1718), .QN(n3330) );
  NAND2X0 U3627 ( .IN1(n3332), .IN2(n3333), .QN(g5396) );
  NAND2X0 U3628 ( .IN1(n2795), .IN2(g1710), .QN(n3333) );
  NAND2X0 U3629 ( .IN1(n968), .IN2(g1713), .QN(n3332) );
  NOR2X0 U3630 ( .IN1(n1654), .IN2(n3334), .QN(g5390) );
  NOR2X0 U3631 ( .IN1(n1677), .IN2(n3334), .QN(g5173) );
  NOR2X0 U3632 ( .IN1(n1614), .IN2(n3334), .QN(g5148) );
  NOR2X0 U3633 ( .IN1(n1658), .IN2(n3334), .QN(g5126) );
  NAND2X0 U3634 ( .IN1(g109), .IN2(DFF_126_n1), .QN(n3334) );
  NOR3X0 U3635 ( .IN1(n2795), .IN2(g4089), .IN3(n3335), .QN(g5083) );
  NOR2X0 U3636 ( .IN1(g4173), .IN2(n2940), .QN(g4940) );
  INVX0 U3637 ( .INP(n3327), .ZN(n2940) );
  NOR2X0 U3638 ( .IN1(n2362), .IN2(test_so1), .QN(n3327) );
  NOR2X0 U3639 ( .IN1(n2358), .IN2(DFF_489_n1), .QN(g4905) );
  NOR2X0 U3640 ( .IN1(n2358), .IN2(DFF_330_n1), .QN(g4903) );
  NOR2X0 U3641 ( .IN1(n2358), .IN2(DFF_385_n1), .QN(g4902) );
  NOR2X0 U3642 ( .IN1(n2356), .IN2(DFF_157_n1), .QN(g4893) );
  AND2X1 U3643 ( .IN1(n3177), .IN2(n3059), .Q(g4892) );
  INVX0 U3644 ( .INP(n2356), .ZN(n3177) );
  NOR2X0 U3645 ( .IN1(n2356), .IN2(DFF_136_n1), .QN(g4891) );
  NOR2X0 U3646 ( .IN1(n2356), .IN2(DFF_336_n1), .QN(g4890) );
  NAND2X0 U3647 ( .IN1(n2788), .IN2(n3336), .QN(n2356) );
  NAND2X0 U3648 ( .IN1(n1607), .IN2(g611), .QN(n3336) );
  NAND4X0 U3649 ( .IN1(n1609), .IN2(n1644), .IN3(n1593), .IN4(n1607), .QN(
        n2788) );
  NAND2X0 U3650 ( .IN1(n2348), .IN2(n2347), .QN(g4556) );
  NOR2X0 U3651 ( .IN1(n4124), .IN2(n2365), .QN(g4506) );
  NOR2X0 U3652 ( .IN1(n4130), .IN2(n2795), .QN(g4500) );
  NOR2X0 U3653 ( .IN1(n1617), .IN2(n2363), .QN(g4498) );
  NOR2X0 U3654 ( .IN1(n1660), .IN2(n2364), .QN(g4490) );
  NOR2X0 U3655 ( .IN1(n1597), .IN2(n2362), .QN(g4484) );
  NOR2X0 U3656 ( .IN1(n1706), .IN2(n2365), .QN(g4480) );
  NOR2X0 U3657 ( .IN1(n1705), .IN2(n2363), .QN(g4477) );
  NOR2X0 U3658 ( .IN1(n1708), .IN2(n2364), .QN(g4473) );
  NOR2X0 U3659 ( .IN1(n1618), .IN2(n2362), .QN(g4471) );
  NOR2X0 U3660 ( .IN1(n2365), .IN2(n2360), .QN(g4465) );
  NOR2X0 U3661 ( .IN1(n1685), .IN2(n2365), .QN(g4342) );
  NOR2X0 U3662 ( .IN1(n1686), .IN2(n2363), .QN(g4340) );
  NAND2X0 U3663 ( .IN1(n3337), .IN2(n3338), .QN(g4309) );
  NAND2X0 U3664 ( .IN1(n3339), .IN2(g1806), .QN(n3338) );
  NAND2X0 U3665 ( .IN1(n3340), .IN2(g1762), .QN(n3337) );
  NAND2X0 U3666 ( .IN1(n3341), .IN2(n3342), .QN(g4293) );
  NAND2X0 U3667 ( .IN1(n3339), .IN2(g1801), .QN(n3342) );
  NAND2X0 U3668 ( .IN1(n3340), .IN2(g1759), .QN(n3341) );
  NAND2X0 U3669 ( .IN1(n3343), .IN2(n3344), .QN(g4283) );
  NAND2X0 U3670 ( .IN1(n3339), .IN2(g1796), .QN(n3344) );
  NAND2X0 U3671 ( .IN1(n3340), .IN2(g1756), .QN(n3343) );
  NAND2X0 U3672 ( .IN1(n3345), .IN2(n3346), .QN(g4274) );
  NAND2X0 U3673 ( .IN1(n3339), .IN2(g1791), .QN(n3346) );
  NAND2X0 U3674 ( .IN1(n3340), .IN2(g1753), .QN(n3345) );
  NAND2X0 U3675 ( .IN1(n3347), .IN2(n3348), .QN(g4264) );
  NAND2X0 U3676 ( .IN1(n3339), .IN2(g1786), .QN(n3348) );
  NAND2X0 U3677 ( .IN1(n3340), .IN2(g1750), .QN(n3347) );
  NAND2X0 U3678 ( .IN1(n3349), .IN2(n3350), .QN(g4255) );
  NAND2X0 U3679 ( .IN1(n3339), .IN2(g1781), .QN(n3350) );
  NAND2X0 U3680 ( .IN1(n3340), .IN2(g1747), .QN(n3349) );
  NAND2X0 U3681 ( .IN1(n3351), .IN2(n3352), .QN(g4239) );
  NAND2X0 U3682 ( .IN1(n3339), .IN2(g1776), .QN(n3352) );
  NAND2X0 U3683 ( .IN1(n3340), .IN2(g1744), .QN(n3351) );
  NAND2X0 U3684 ( .IN1(n3353), .IN2(n3354), .QN(g4238) );
  NAND2X0 U3685 ( .IN1(n3339), .IN2(test_so5), .QN(n3354) );
  NAND2X0 U3686 ( .IN1(n3340), .IN2(g1741), .QN(n3353) );
  NAND2X0 U3687 ( .IN1(n3355), .IN2(n3356), .QN(g4231) );
  NAND2X0 U3688 ( .IN1(n3339), .IN2(g1766), .QN(n3356) );
  INVX0 U3689 ( .INP(n3340), .ZN(n3339) );
  NAND2X0 U3690 ( .IN1(n3340), .IN2(g1738), .QN(n3355) );
  NAND2X0 U3691 ( .IN1(g1700), .IN2(DFF_275_n1), .QN(g4089) );
  NOR2X0 U3692 ( .IN1(g1707), .IN2(n374), .QN(g4076) );
  INVX0 U3693 ( .INP(g1700), .ZN(n374) );
  NOR2X0 U3694 ( .IN1(n2337), .IN2(n3357), .QN(g3462) );
  NOR2X0 U3695 ( .IN1(n3358), .IN2(n3183), .QN(n3357) );
  NOR2X0 U3696 ( .IN1(n1647), .IN2(g750), .QN(n3358) );
  NOR4X0 U3697 ( .IN1(n1712), .IN2(n1630), .IN3(n1604), .IN4(n1591), .QN(g3381) );
  INVX0 U3698 ( .INP(g23), .ZN(g3327) );
  NOR2X0 U3699 ( .IN1(g1610), .IN2(g1737), .QN(g2478) );
  NAND2X0 U3700 ( .IN1(n3359), .IN2(n3360), .QN(g11647) );
  NAND2X0 U3701 ( .IN1(n3092), .IN2(g336), .QN(n3360) );
  NAND2X0 U3702 ( .IN1(n3183), .IN2(n3361), .QN(n3359) );
  NAND2X0 U3703 ( .IN1(n3362), .IN2(n3363), .QN(n3361) );
  NAND2X0 U3704 ( .IN1(n3364), .IN2(n3365), .QN(n3363) );
  NAND2X0 U3705 ( .IN1(n3366), .IN2(n3367), .QN(n3362) );
  NOR2X0 U3706 ( .IN1(n3368), .IN2(n3369), .QN(g11641) );
  NOR2X0 U3707 ( .IN1(n3370), .IN2(n3371), .QN(n3368) );
  NOR2X0 U3708 ( .IN1(n1721), .IN2(n1226), .QN(n3371) );
  AND2X1 U3709 ( .IN1(n2357), .IN2(n2), .Q(n1226) );
  NOR3X0 U3710 ( .IN1(n2566), .IN2(n2357), .IN3(n1227), .QN(n3370) );
  NOR2X0 U3711 ( .IN1(n2566), .IN2(n1721), .QN(n2357) );
  NAND3X0 U3712 ( .IN1(g1346), .IN2(g1336), .IN3(g1341), .QN(n2566) );
  NOR2X0 U3713 ( .IN1(n3372), .IN2(n3369), .QN(g11640) );
  AND2X1 U3714 ( .IN1(n3373), .IN2(n3374), .Q(n3372) );
  NAND2X0 U3715 ( .IN1(n3375), .IN2(g1346), .QN(n3374) );
  NAND3X0 U3716 ( .IN1(g1341), .IN2(g1336), .IN3(n2), .QN(n3375) );
  NAND2X0 U3717 ( .IN1(n1232), .IN2(n1231), .QN(n3373) );
  NOR2X0 U3718 ( .IN1(n3369), .IN2(n3376), .QN(g11639) );
  XOR2X1 U3719 ( .IN1(n2311), .IN2(n1231), .Q(n3376) );
  NOR2X0 U3720 ( .IN1(n3369), .IN2(n3377), .QN(g11636) );
  XOR2X1 U3721 ( .IN1(g1336), .IN2(n1227), .Q(n3377) );
  NAND2X0 U3722 ( .IN1(n3378), .IN2(g109), .QN(n3369) );
  OR3X1 U3723 ( .IN1(n3305), .IN2(n2347), .IN3(n3036), .Q(n3378) );
  NAND2X0 U3724 ( .IN1(n3379), .IN2(n3380), .QN(g11625) );
  NAND2X0 U3725 ( .IN1(n3092), .IN2(g345), .QN(n3380) );
  NAND2X0 U3726 ( .IN1(n3183), .IN2(n3381), .QN(n3379) );
  XOR2X1 U3727 ( .IN1(n3364), .IN2(n3367), .Q(n3381) );
  AND2X1 U3728 ( .IN1(n3382), .IN2(n3383), .Q(n3367) );
  OR2X1 U3729 ( .IN1(n14), .IN2(n1681), .Q(n3383) );
  NAND2X0 U3730 ( .IN1(n3384), .IN2(n14), .QN(n3382) );
  XNOR2X1 U3731 ( .IN1(n3385), .IN2(n3386), .Q(n3384) );
  OR2X1 U3732 ( .IN1(g466), .IN2(n3387), .Q(n3385) );
  XNOR3X1 U3733 ( .IN1(n3388), .IN2(n3389), .IN3(n3390), .Q(n3364) );
  XOR3X1 U3734 ( .IN1(n3391), .IN2(n3392), .IN3(n3393), .Q(n3390) );
  XNOR2X1 U3735 ( .IN1(n3394), .IN2(n3395), .Q(n3393) );
  XOR3X1 U3736 ( .IN1(n3396), .IN2(n3397), .IN3(n3398), .Q(n3388) );
  XOR2X1 U3737 ( .IN1(n3399), .IN2(n3400), .Q(n3398) );
  NAND2X0 U3738 ( .IN1(n3401), .IN2(n3402), .QN(g11610) );
  NAND2X0 U3739 ( .IN1(n3403), .IN2(g1806), .QN(n3402) );
  NAND2X0 U3740 ( .IN1(n3404), .IN2(g1333), .QN(n3401) );
  NAND2X0 U3741 ( .IN1(n3405), .IN2(n3406), .QN(g11609) );
  NAND2X0 U3742 ( .IN1(n3403), .IN2(g1801), .QN(n3406) );
  NAND2X0 U3743 ( .IN1(n3404), .IN2(g1330), .QN(n3405) );
  NAND2X0 U3744 ( .IN1(n3407), .IN2(n3408), .QN(g11608) );
  NAND2X0 U3745 ( .IN1(n3403), .IN2(g1796), .QN(n3408) );
  NAND2X0 U3746 ( .IN1(n3404), .IN2(g1327), .QN(n3407) );
  NAND2X0 U3747 ( .IN1(n3409), .IN2(n3410), .QN(g11607) );
  NAND2X0 U3748 ( .IN1(n3403), .IN2(g1791), .QN(n3410) );
  NAND2X0 U3749 ( .IN1(n3404), .IN2(g1324), .QN(n3409) );
  NAND2X0 U3750 ( .IN1(n3411), .IN2(n3412), .QN(g11606) );
  NAND2X0 U3751 ( .IN1(n3403), .IN2(g1786), .QN(n3412) );
  NAND2X0 U3752 ( .IN1(n3404), .IN2(g1321), .QN(n3411) );
  NAND2X0 U3753 ( .IN1(n3413), .IN2(n3414), .QN(g11605) );
  NAND2X0 U3754 ( .IN1(n3403), .IN2(g1781), .QN(n3414) );
  NAND2X0 U3755 ( .IN1(n3404), .IN2(g1318), .QN(n3413) );
  NAND2X0 U3756 ( .IN1(n3415), .IN2(n3416), .QN(g11604) );
  NAND2X0 U3757 ( .IN1(n3403), .IN2(g1776), .QN(n3416) );
  NAND2X0 U3758 ( .IN1(n3404), .IN2(g1314), .QN(n3415) );
  NAND2X0 U3759 ( .IN1(n3417), .IN2(n3418), .QN(g11603) );
  NAND2X0 U3760 ( .IN1(test_so9), .IN2(n3404), .QN(n3418) );
  NAND2X0 U3761 ( .IN1(n3403), .IN2(test_so5), .QN(n3417) );
  NAND2X0 U3762 ( .IN1(n3419), .IN2(n3420), .QN(g11602) );
  NAND2X0 U3763 ( .IN1(n3403), .IN2(g1766), .QN(n3420) );
  INVX0 U3764 ( .INP(n3404), .ZN(n3403) );
  NAND2X0 U3765 ( .IN1(n3404), .IN2(g1308), .QN(n3419) );
  NAND2X0 U3766 ( .IN1(n2), .IN2(g1317), .QN(n3404) );
  INVX0 U3767 ( .INP(n1227), .ZN(n2) );
  NAND3X0 U3768 ( .IN1(n3014), .IN2(n3421), .IN3(n3012), .QN(n1227) );
  NAND4X0 U3769 ( .IN1(n3422), .IN2(n3423), .IN3(n3424), .IN4(n3425), .QN(
        n3421) );
  NOR4X0 U3770 ( .IN1(n3426), .IN2(n3427), .IN3(n3428), .IN4(n3429), .QN(n3425) );
  XOR2X1 U3771 ( .IN1(n2243), .IN2(n2228), .Q(n3429) );
  XOR2X1 U3772 ( .IN1(n2268), .IN2(n2267), .Q(n3428) );
  XOR2X1 U3773 ( .IN1(n2240), .IN2(n2229), .Q(n3427) );
  NAND2X0 U3774 ( .IN1(n3430), .IN2(n3431), .QN(n3426) );
  XOR2X1 U3775 ( .IN1(n2304), .IN2(g1275), .Q(n3431) );
  XOR2X1 U3776 ( .IN1(n2306), .IN2(g1240), .Q(n3430) );
  NOR3X0 U3777 ( .IN1(n3432), .IN2(n3433), .IN3(n3434), .QN(n3424) );
  XNOR2X1 U3778 ( .IN1(n3435), .IN2(n3436), .Q(n3434) );
  XOR2X1 U3779 ( .IN1(test_so2), .IN2(g1255), .Q(n3433) );
  XNOR2X1 U3780 ( .IN1(n2203), .IN2(test_so6), .Q(n3432) );
  XOR2X1 U3781 ( .IN1(test_so8), .IN2(n2265), .Q(n3423) );
  XOR2X1 U3782 ( .IN1(n1871), .IN2(g1235), .Q(n3422) );
  NAND2X0 U3783 ( .IN1(n3437), .IN2(n3438), .QN(g11579) );
  NAND2X0 U3784 ( .IN1(n968), .IN2(g1618), .QN(n3438) );
  NAND2X0 U3785 ( .IN1(n3439), .IN2(n2795), .QN(n3437) );
  XOR2X1 U3786 ( .IN1(g1610), .IN2(n3440), .Q(n3439) );
  NAND2X0 U3787 ( .IN1(n3441), .IN2(n3442), .QN(n3440) );
  NAND2X0 U3788 ( .IN1(n3443), .IN2(n3444), .QN(n3442) );
  NAND2X0 U3789 ( .IN1(n1262), .IN2(n2557), .QN(n3444) );
  NAND3X0 U3790 ( .IN1(n3445), .IN2(n3446), .IN3(n3447), .QN(n2557) );
  NAND3X0 U3791 ( .IN1(n1658), .IN2(n2830), .IN3(n1677), .QN(n3447) );
  NAND2X0 U3792 ( .IN1(n1686), .IN2(g1149), .QN(n3446) );
  NAND2X0 U3793 ( .IN1(n1685), .IN2(n3448), .QN(n3445) );
  NAND4X0 U3794 ( .IN1(n3449), .IN2(n3450), .IN3(n1677), .IN4(n3451), .QN(
        n1262) );
  AND2X1 U3795 ( .IN1(n2830), .IN2(n1658), .Q(n3451) );
  NOR2X0 U3796 ( .IN1(g1107), .IN2(n1654), .QN(n2830) );
  OR2X1 U3797 ( .IN1(n1685), .IN2(n1686), .Q(n3450) );
  OR2X1 U3798 ( .IN1(g1149), .IN2(n3448), .Q(n3449) );
  NAND2X0 U3799 ( .IN1(n1686), .IN2(n3452), .QN(n3448) );
  NAND4X0 U3800 ( .IN1(n3453), .IN2(n1706), .IN3(n3454), .IN4(n3455), .QN(
        n3452) );
  NOR4X0 U3801 ( .IN1(n3456), .IN2(n3016), .IN3(g1163), .IN4(g1160), .QN(n3455) );
  NAND3X0 U3802 ( .IN1(n2275), .IN2(n1708), .IN3(n4132), .QN(n3456) );
  AND4X1 U3803 ( .IN1(n2360), .IN2(n1597), .IN3(n1617), .IN4(n1618), .Q(n3454)
         );
  AND2X1 U3804 ( .IN1(n1660), .IN2(n1705), .Q(n3453) );
  NAND2X0 U3805 ( .IN1(n1260), .IN2(n3457), .QN(n3441) );
  INVX0 U3806 ( .INP(n3443), .ZN(n3457) );
  NAND2X0 U3807 ( .IN1(n3458), .IN2(n3459), .QN(g11514) );
  OR3X1 U3808 ( .IN1(g1419), .IN2(n2364), .IN3(n3460), .Q(n3459) );
  NAND2X0 U3809 ( .IN1(g6193), .IN2(n3460), .QN(n3458) );
  XOR3X1 U3810 ( .IN1(n1627), .IN2(n3461), .IN3(n3443), .Q(n3460) );
  NAND2X0 U3811 ( .IN1(n3462), .IN2(n3463), .QN(n3443) );
  OR2X1 U3812 ( .IN1(n2569), .IN2(n1619), .Q(n3463) );
  NAND2X0 U3813 ( .IN1(n3464), .IN2(n2569), .QN(n3462) );
  NAND2X0 U3814 ( .IN1(n3465), .IN2(n3466), .QN(n3464) );
  OR2X1 U3815 ( .IN1(n3467), .IN2(g1811), .Q(n3466) );
  NAND2X0 U3816 ( .IN1(n3467), .IN2(n3468), .QN(n3465) );
  NAND2X0 U3817 ( .IN1(n3469), .IN2(n3470), .QN(n3468) );
  NAND4X0 U3818 ( .IN1(n4117), .IN2(n4119), .IN3(n4120), .IN4(n4123), .QN(
        n3467) );
  XOR2X1 U3819 ( .IN1(n2262), .IN2(n2137), .Q(n3461) );
  NOR2X0 U3820 ( .IN1(n2363), .IN2(n1602), .QN(g6193) );
  NAND2X0 U3821 ( .IN1(n3471), .IN2(n3472), .QN(g11488) );
  NAND2X0 U3822 ( .IN1(n3092), .IN2(g342), .QN(n3472) );
  NAND2X0 U3823 ( .IN1(n3183), .IN2(n3397), .QN(n3471) );
  NAND2X0 U3824 ( .IN1(n3473), .IN2(n3474), .QN(n3397) );
  OR2X1 U3825 ( .IN1(n14), .IN2(n2072), .Q(n3474) );
  NAND2X0 U3826 ( .IN1(n3475), .IN2(n14), .QN(n3473) );
  XOR2X1 U3827 ( .IN1(n3476), .IN2(n1620), .Q(n3475) );
  NAND4X0 U3828 ( .IN1(n1646), .IN2(n1594), .IN3(g471), .IN4(g456), .QN(n3476)
         );
  NAND2X0 U3829 ( .IN1(n3477), .IN2(n3478), .QN(g11487) );
  NAND2X0 U3830 ( .IN1(n3092), .IN2(g366), .QN(n3478) );
  NAND2X0 U3831 ( .IN1(n3183), .IN2(n3396), .QN(n3477) );
  NAND2X0 U3832 ( .IN1(n3479), .IN2(n3480), .QN(n3396) );
  OR2X1 U3833 ( .IN1(n14), .IN2(n2291), .Q(n3480) );
  NAND2X0 U3834 ( .IN1(n3481), .IN2(n14), .QN(n3479) );
  XOR2X1 U3835 ( .IN1(g511), .IN2(n3482), .Q(n3481) );
  NOR2X0 U3836 ( .IN1(g461), .IN2(n3483), .QN(n3482) );
  NAND2X0 U3837 ( .IN1(n3484), .IN2(n3485), .QN(g11486) );
  NAND2X0 U3838 ( .IN1(n3092), .IN2(g363), .QN(n3485) );
  NAND2X0 U3839 ( .IN1(n3183), .IN2(n3400), .QN(n3484) );
  NAND2X0 U3840 ( .IN1(n3486), .IN2(n3487), .QN(n3400) );
  OR2X1 U3841 ( .IN1(n14), .IN2(n2071), .Q(n3487) );
  NAND2X0 U3842 ( .IN1(n3488), .IN2(n14), .QN(n3486) );
  XOR2X1 U3843 ( .IN1(n3489), .IN2(n1600), .Q(n3488) );
  NAND2X0 U3844 ( .IN1(n3490), .IN2(n1606), .QN(n3489) );
  NAND2X0 U3845 ( .IN1(n3491), .IN2(n3492), .QN(g11485) );
  NAND2X0 U3846 ( .IN1(n3092), .IN2(g360), .QN(n3492) );
  NAND2X0 U3847 ( .IN1(n3183), .IN2(n3392), .QN(n3491) );
  NAND2X0 U3848 ( .IN1(n3493), .IN2(n3494), .QN(n3392) );
  OR2X1 U3849 ( .IN1(n14), .IN2(n2273), .Q(n3494) );
  NAND2X0 U3850 ( .IN1(n3495), .IN2(n14), .QN(n3493) );
  XOR2X1 U3851 ( .IN1(g501), .IN2(n3496), .Q(n3495) );
  NOR2X0 U3852 ( .IN1(n1594), .IN2(n3497), .QN(n3496) );
  NAND2X0 U3853 ( .IN1(n3498), .IN2(n3499), .QN(g11484) );
  NAND2X0 U3854 ( .IN1(n3092), .IN2(g357), .QN(n3499) );
  NAND2X0 U3855 ( .IN1(n3183), .IN2(n3391), .QN(n3498) );
  NAND2X0 U3856 ( .IN1(n3500), .IN2(n3501), .QN(n3391) );
  OR2X1 U3857 ( .IN1(n14), .IN2(n2269), .Q(n3501) );
  NAND2X0 U3858 ( .IN1(n3502), .IN2(n14), .QN(n3500) );
  XOR2X1 U3859 ( .IN1(g496), .IN2(n3503), .Q(n3502) );
  NOR2X0 U3860 ( .IN1(n1646), .IN2(n3387), .QN(n3503) );
  NAND3X0 U3861 ( .IN1(n1594), .IN2(g456), .IN3(n1606), .QN(n3387) );
  NAND2X0 U3862 ( .IN1(n3504), .IN2(n3505), .QN(g11483) );
  NAND2X0 U3863 ( .IN1(n3092), .IN2(g354), .QN(n3505) );
  NAND2X0 U3864 ( .IN1(n3183), .IN2(n3394), .QN(n3504) );
  NAND2X0 U3865 ( .IN1(n3506), .IN2(n3507), .QN(n3394) );
  OR2X1 U3866 ( .IN1(n14), .IN2(n2310), .Q(n3507) );
  NAND2X0 U3867 ( .IN1(n3508), .IN2(n14), .QN(n3506) );
  XOR2X1 U3868 ( .IN1(g491), .IN2(n3509), .Q(n3508) );
  NOR2X0 U3869 ( .IN1(g461), .IN2(n3497), .QN(n3509) );
  NAND3X0 U3870 ( .IN1(n1606), .IN2(g466), .IN3(n1641), .QN(n3497) );
  NAND2X0 U3871 ( .IN1(n3510), .IN2(n3511), .QN(g11482) );
  NAND2X0 U3872 ( .IN1(n3092), .IN2(g351), .QN(n3511) );
  NAND2X0 U3873 ( .IN1(n3183), .IN2(n3389), .QN(n3510) );
  NAND2X0 U3874 ( .IN1(n3512), .IN2(n3513), .QN(n3389) );
  OR2X1 U3875 ( .IN1(n14), .IN2(n2271), .Q(n3513) );
  NAND2X0 U3876 ( .IN1(n3514), .IN2(n14), .QN(n3512) );
  XOR2X1 U3877 ( .IN1(g486), .IN2(n3515), .Q(n3514) );
  NOR2X0 U3878 ( .IN1(n1641), .IN2(n3516), .QN(n3515) );
  NAND2X0 U3879 ( .IN1(n3517), .IN2(n3518), .QN(g11481) );
  NAND2X0 U3880 ( .IN1(n3092), .IN2(g348), .QN(n3518) );
  NAND2X0 U3881 ( .IN1(n3183), .IN2(n3395), .QN(n3517) );
  NAND2X0 U3882 ( .IN1(n3519), .IN2(n3520), .QN(n3395) );
  OR2X1 U3883 ( .IN1(n14), .IN2(n2308), .Q(n3520) );
  NAND2X0 U3884 ( .IN1(n3521), .IN2(n14), .QN(n3519) );
  XOR2X1 U3885 ( .IN1(g481), .IN2(n3522), .Q(n3521) );
  NOR2X0 U3886 ( .IN1(n3516), .IN2(g456), .QN(n3522) );
  NAND3X0 U3887 ( .IN1(n1606), .IN2(g461), .IN3(n1646), .QN(n3516) );
  NAND2X0 U3888 ( .IN1(n3523), .IN2(n3524), .QN(g11478) );
  NAND2X0 U3889 ( .IN1(n3092), .IN2(g339), .QN(n3524) );
  NAND2X0 U3890 ( .IN1(n3183), .IN2(n3399), .QN(n3523) );
  NAND2X0 U3891 ( .IN1(n3525), .IN2(n3526), .QN(n3399) );
  OR2X1 U3892 ( .IN1(n14), .IN2(n2289), .Q(n3526) );
  NAND2X0 U3893 ( .IN1(n3527), .IN2(n14), .QN(n3525) );
  XOR2X1 U3894 ( .IN1(g476), .IN2(n3528), .Q(n3527) );
  NOR2X0 U3895 ( .IN1(n1594), .IN2(n3483), .QN(n3528) );
  NAND3X0 U3896 ( .IN1(n1646), .IN2(g471), .IN3(n1641), .QN(n3483) );
  INVX0 U3897 ( .INP(n3092), .ZN(n3183) );
  NAND2X0 U3898 ( .IN1(n1647), .IN2(g750), .QN(n3092) );
  NAND2X0 U3899 ( .IN1(n3529), .IN2(n3530), .QN(g11443) );
  NAND2X0 U3900 ( .IN1(n3043), .IN2(g1275), .QN(n3530) );
  NOR2X0 U3901 ( .IN1(n3012), .IN2(n2364), .QN(n3043) );
  NAND2X0 U3902 ( .IN1(n3012), .IN2(n3435), .QN(n3529) );
  NAND2X0 U3903 ( .IN1(n3531), .IN2(n3532), .QN(n3435) );
  OR2X1 U3904 ( .IN1(n3436), .IN2(n3014), .Q(n3532) );
  XOR2X1 U3905 ( .IN1(n2350), .IN2(n3533), .Q(n3436) );
  NOR2X0 U3906 ( .IN1(n3366), .IN2(n2201), .QN(n3533) );
  INVX0 U3907 ( .INP(n3365), .ZN(n3366) );
  NAND2X0 U3908 ( .IN1(n3534), .IN2(n3014), .QN(n3531) );
  NOR2X0 U3909 ( .IN1(n3010), .IN2(n2117), .QN(n3014) );
  OR3X1 U3910 ( .IN1(n2119), .IN2(n2120), .IN3(n2118), .Q(n3010) );
  NAND2X0 U3911 ( .IN1(n3535), .IN2(n3536), .QN(n3534) );
  NAND2X0 U3912 ( .IN1(n1864), .IN2(g1280), .QN(n3536) );
  NAND2X0 U3913 ( .IN1(n1862), .IN2(n3537), .QN(n3535) );
  NAND2X0 U3914 ( .IN1(n1864), .IN2(n3538), .QN(n3537) );
  NAND4X0 U3915 ( .IN1(n3539), .IN2(n2246), .IN3(n3540), .IN4(n3541), .QN(
        n3538) );
  NOR4X0 U3916 ( .IN1(n3542), .IN2(g1240), .IN3(g1250), .IN4(g1275), .QN(n3541) );
  NAND3X0 U3917 ( .IN1(n2265), .IN2(n2247), .IN3(n2266), .QN(n3542) );
  NOR4X0 U3918 ( .IN1(test_so6), .IN2(g1255), .IN3(g1260), .IN4(g1265), .QN(
        n3540) );
  NOR2X0 U3919 ( .IN1(g1292), .IN2(g1296), .QN(n3539) );
  NOR3X0 U3920 ( .IN1(n968), .IN2(n2348), .IN3(g1713), .QN(n3012) );
  NOR2X0 U3921 ( .IN1(n3543), .IN2(n3544), .QN(g11393) );
  NOR2X0 U3922 ( .IN1(n3545), .IN2(n3546), .QN(n3543) );
  NOR2X0 U3923 ( .IN1(n1722), .IN2(n3547), .QN(n3546) );
  AND2X1 U3924 ( .IN1(n11), .IN2(n33), .Q(n3547) );
  INVX0 U3925 ( .INP(n3548), .ZN(n11) );
  NOR3X0 U3926 ( .IN1(n3549), .IN2(n1720), .IN3(n33), .QN(n3545) );
  NOR4X0 U3927 ( .IN1(n1720), .IN2(n1722), .IN3(n2314), .IN4(n2315), .QN(n33)
         );
  NOR2X0 U3928 ( .IN1(n3544), .IN2(n3550), .QN(g11392) );
  XNOR2X1 U3929 ( .IN1(n1720), .IN2(n3549), .Q(n3550) );
  NAND2X0 U3930 ( .IN1(n3551), .IN2(g976), .QN(n3549) );
  NOR2X0 U3931 ( .IN1(n3544), .IN2(n3552), .QN(g11391) );
  XOR2X1 U3932 ( .IN1(n2314), .IN2(n3551), .Q(n3552) );
  NOR2X0 U3933 ( .IN1(n3553), .IN2(n3554), .QN(g11380) );
  NOR2X0 U3934 ( .IN1(n3555), .IN2(g471), .QN(n3553) );
  NOR2X0 U3935 ( .IN1(n3556), .IN2(n3554), .QN(g11376) );
  NOR2X0 U3936 ( .IN1(n3557), .IN2(n3558), .QN(n3556) );
  NOR2X0 U3937 ( .IN1(n1646), .IN2(n3555), .QN(n3558) );
  NOR2X0 U3938 ( .IN1(n3559), .IN2(n3560), .QN(n3555) );
  AND3X1 U3939 ( .IN1(n3560), .IN2(g461), .IN3(n3561), .Q(n3557) );
  NOR2X0 U3940 ( .IN1(n3554), .IN2(n3562), .QN(g11372) );
  XOR2X1 U3941 ( .IN1(n1594), .IN2(n3561), .Q(n3562) );
  NOR2X0 U3942 ( .IN1(n3559), .IN2(n1641), .QN(n3561) );
  NOR3X0 U3943 ( .IN1(n3544), .IN2(n3551), .IN3(n3563), .QN(g11349) );
  AND2X1 U3944 ( .IN1(n3548), .IN2(n2315), .Q(n3563) );
  NOR2X0 U3945 ( .IN1(n3548), .IN2(n2315), .QN(n3551) );
  NAND3X0 U3946 ( .IN1(n3564), .IN2(n14), .IN3(n1420), .QN(n3548) );
  NAND4X0 U3947 ( .IN1(n3565), .IN2(n3566), .IN3(n3567), .IN4(n3568), .QN(
        n3564) );
  NOR4X0 U3948 ( .IN1(n3569), .IN2(n3570), .IN3(n3571), .IN4(n3572), .QN(n3568) );
  XOR2X1 U3949 ( .IN1(n2274), .IN2(n2273), .Q(n3572) );
  XOR2X1 U3950 ( .IN1(n2292), .IN2(n2291), .Q(n3571) );
  XOR2X1 U3951 ( .IN1(n2290), .IN2(n2289), .Q(n3570) );
  NAND2X0 U3952 ( .IN1(n3573), .IN2(n3574), .QN(n3569) );
  XOR2X1 U3953 ( .IN1(n2308), .IN2(g426), .Q(n3574) );
  XOR2X1 U3954 ( .IN1(n2310), .IN2(g391), .Q(n3573) );
  NOR3X0 U3955 ( .IN1(n3575), .IN2(n3576), .IN3(n3577), .QN(n3567) );
  XNOR2X1 U3956 ( .IN1(n1681), .IN2(n3578), .Q(n3577) );
  XOR2X1 U3957 ( .IN1(n2248), .IN2(n2072), .Q(n3576) );
  XOR2X1 U3958 ( .IN1(n2241), .IN2(n2071), .Q(n3575) );
  XOR2X1 U3959 ( .IN1(n2269), .IN2(g396), .Q(n3566) );
  XOR2X1 U3960 ( .IN1(n2271), .IN2(g386), .Q(n3565) );
  NAND2X0 U3961 ( .IN1(n3579), .IN2(g109), .QN(n3544) );
  OR3X1 U3962 ( .IN1(n2555), .IN2(n2116), .IN3(n3064), .Q(n3579) );
  NOR2X0 U3963 ( .IN1(n3554), .IN2(n3580), .QN(g11340) );
  XOR2X1 U3964 ( .IN1(g456), .IN2(n3559), .Q(n3580) );
  NAND2X0 U3965 ( .IN1(n14), .IN2(n3581), .QN(n3559) );
  NAND2X0 U3966 ( .IN1(n3490), .IN2(g471), .QN(n3581) );
  INVX0 U3967 ( .INP(n3560), .ZN(n3490) );
  NAND3X0 U3968 ( .IN1(g456), .IN2(g466), .IN3(g461), .QN(n3560) );
  NAND2X0 U3969 ( .IN1(g109), .IN2(DFF_441_n1), .QN(n3554) );
  NAND2X0 U3970 ( .IN1(n3582), .IN2(n3583), .QN(g11338) );
  NAND2X0 U3971 ( .IN1(n2351), .IN2(g476), .QN(n3583) );
  NAND2X0 U3972 ( .IN1(n14), .IN2(g516), .QN(n3582) );
  NAND2X0 U3973 ( .IN1(n3584), .IN2(n3585), .QN(g11337) );
  NAND2X0 U3974 ( .IN1(n2351), .IN2(g516), .QN(n3585) );
  NAND2X0 U3975 ( .IN1(n14), .IN2(g511), .QN(n3584) );
  NAND2X0 U3976 ( .IN1(n3586), .IN2(n3587), .QN(g11336) );
  NAND2X0 U3977 ( .IN1(n2351), .IN2(g511), .QN(n3587) );
  NAND2X0 U3978 ( .IN1(n14), .IN2(g506), .QN(n3586) );
  NAND2X0 U3979 ( .IN1(n3588), .IN2(n3589), .QN(g11335) );
  NAND2X0 U3980 ( .IN1(n2351), .IN2(g506), .QN(n3589) );
  NAND2X0 U3981 ( .IN1(n14), .IN2(g501), .QN(n3588) );
  NAND2X0 U3982 ( .IN1(n3590), .IN2(n3591), .QN(g11334) );
  NAND2X0 U3983 ( .IN1(n2351), .IN2(g501), .QN(n3591) );
  NAND2X0 U3984 ( .IN1(n14), .IN2(g496), .QN(n3590) );
  NAND2X0 U3985 ( .IN1(n3592), .IN2(n3593), .QN(g11333) );
  NAND2X0 U3986 ( .IN1(n2351), .IN2(g496), .QN(n3593) );
  NAND2X0 U3987 ( .IN1(n14), .IN2(g491), .QN(n3592) );
  NAND2X0 U3988 ( .IN1(n3594), .IN2(n3595), .QN(g11332) );
  NAND2X0 U3989 ( .IN1(n2351), .IN2(g491), .QN(n3595) );
  NAND2X0 U3990 ( .IN1(n14), .IN2(g486), .QN(n3594) );
  NAND2X0 U3991 ( .IN1(n3596), .IN2(n3597), .QN(g11331) );
  NAND2X0 U3992 ( .IN1(n2351), .IN2(g486), .QN(n3597) );
  NAND2X0 U3993 ( .IN1(n14), .IN2(g481), .QN(n3596) );
  NAND2X0 U3994 ( .IN1(n3598), .IN2(n3599), .QN(g11330) );
  NAND2X0 U3995 ( .IN1(n2351), .IN2(g521), .QN(n3599) );
  NAND2X0 U3996 ( .IN1(n14), .IN2(g525), .QN(n3598) );
  NAND2X0 U3997 ( .IN1(n3600), .IN2(n3601), .QN(g11329) );
  NAND2X0 U3998 ( .IN1(n2351), .IN2(g525), .QN(n3601) );
  NAND2X0 U3999 ( .IN1(n14), .IN2(g530), .QN(n3600) );
  NAND2X0 U4000 ( .IN1(n3602), .IN2(n3603), .QN(g11328) );
  NAND2X0 U4001 ( .IN1(n2351), .IN2(g530), .QN(n3603) );
  NAND2X0 U4002 ( .IN1(n14), .IN2(g534), .QN(n3602) );
  NAND2X0 U4003 ( .IN1(n3604), .IN2(n3605), .QN(g11327) );
  NAND2X0 U4004 ( .IN1(n2351), .IN2(g534), .QN(n3605) );
  NAND2X0 U4005 ( .IN1(n14), .IN2(g538), .QN(n3604) );
  NAND2X0 U4006 ( .IN1(n3606), .IN2(n3607), .QN(g11326) );
  NAND2X0 U4007 ( .IN1(n2351), .IN2(g538), .QN(n3607) );
  NAND2X0 U4008 ( .IN1(n14), .IN2(g542), .QN(n3606) );
  NAND2X0 U4009 ( .IN1(n3608), .IN2(n3609), .QN(g11325) );
  NAND2X0 U4010 ( .IN1(n2351), .IN2(g542), .QN(n3609) );
  NAND2X0 U4011 ( .IN1(n14), .IN2(g476), .QN(n3608) );
  NAND2X0 U4012 ( .IN1(n3610), .IN2(n3611), .QN(g11324) );
  NAND2X0 U4013 ( .IN1(n2351), .IN2(g481), .QN(n3611) );
  NAND2X0 U4014 ( .IN1(n3386), .IN2(n14), .QN(n3610) );
  NAND2X0 U4015 ( .IN1(n3612), .IN2(n3613), .QN(n3386) );
  NAND2X0 U4016 ( .IN1(n1695), .IN2(g521), .QN(n3613) );
  NAND2X0 U4017 ( .IN1(n1698), .IN2(n3614), .QN(n3612) );
  NAND2X0 U4018 ( .IN1(n1695), .IN2(n3615), .QN(n3614) );
  NAND2X0 U4019 ( .IN1(n3616), .IN2(n3617), .QN(n3615) );
  NOR4X0 U4020 ( .IN1(n3618), .IN2(g496), .IN3(g511), .IN4(g481), .QN(n3617)
         );
  NAND4X0 U4021 ( .IN1(n1621), .IN2(n1620), .IN3(n1600), .IN4(n1599), .QN(
        n3618) );
  NOR4X0 U4022 ( .IN1(n3619), .IN2(g542), .IN3(g534), .IN4(g538), .QN(n3616)
         );
  NAND3X0 U4023 ( .IN1(n1691), .IN2(n1690), .IN3(n2296), .QN(n3619) );
  AND3X1 U4024 ( .IN1(n3620), .IN2(n3621), .IN3(n3622), .Q(g11320) );
  INVX0 U4025 ( .INP(n3623), .ZN(n3622) );
  NAND2X0 U4026 ( .IN1(n2226), .IN2(n3624), .QN(n3620) );
  NAND2X0 U4027 ( .IN1(n14), .IN2(n3625), .QN(n3624) );
  NAND2X0 U4028 ( .IN1(n3626), .IN2(n3627), .QN(g11314) );
  NAND2X0 U4029 ( .IN1(n1855), .IN2(g861), .QN(n3627) );
  NAND2X0 U4030 ( .IN1(n3628), .IN2(g968), .QN(n3626) );
  NAND2X0 U4031 ( .IN1(n3629), .IN2(n3630), .QN(g11312) );
  NAND2X0 U4032 ( .IN1(n1855), .IN2(g857), .QN(n3630) );
  NAND2X0 U4033 ( .IN1(g965), .IN2(n3628), .QN(n3629) );
  NAND2X0 U4034 ( .IN1(n3631), .IN2(n3632), .QN(g11310) );
  OR2X1 U4035 ( .IN1(n3628), .IN2(n2079), .Q(n3632) );
  NAND2X0 U4036 ( .IN1(g962), .IN2(n3628), .QN(n3631) );
  NAND2X0 U4037 ( .IN1(n3633), .IN2(n3634), .QN(g11308) );
  OR2X1 U4038 ( .IN1(n3628), .IN2(n2102), .Q(n3634) );
  NAND2X0 U4039 ( .IN1(n3628), .IN2(g959), .QN(n3633) );
  NAND2X0 U4040 ( .IN1(n3635), .IN2(n3636), .QN(g11306) );
  OR2X1 U4041 ( .IN1(n3628), .IN2(n2103), .Q(n3636) );
  OR2X1 U4042 ( .IN1(n1855), .IN2(n2085), .Q(n3635) );
  NAND2X0 U4043 ( .IN1(n3637), .IN2(n3638), .QN(g11305) );
  NAND2X0 U4044 ( .IN1(n1855), .IN2(g841), .QN(n3638) );
  NAND2X0 U4045 ( .IN1(n3628), .IN2(g953), .QN(n3637) );
  NAND2X0 U4046 ( .IN1(n3639), .IN2(n3640), .QN(g11303) );
  NAND2X0 U4047 ( .IN1(n1855), .IN2(g837), .QN(n3640) );
  NAND2X0 U4048 ( .IN1(n3628), .IN2(g950), .QN(n3639) );
  NAND2X0 U4049 ( .IN1(n3641), .IN2(n3642), .QN(g11300) );
  OR2X1 U4050 ( .IN1(n3628), .IN2(n2074), .Q(n3642) );
  OR2X1 U4051 ( .IN1(n1855), .IN2(n2073), .Q(n3641) );
  NAND2X0 U4052 ( .IN1(n3643), .IN2(n3644), .QN(g11298) );
  NAND2X0 U4053 ( .IN1(n3628), .IN2(g944), .QN(n3644) );
  OR2X1 U4054 ( .IN1(n3628), .IN2(n1651), .Q(n3643) );
  INVX0 U4055 ( .INP(n1855), .ZN(n3628) );
  NAND3X0 U4056 ( .IN1(n3645), .IN2(n3646), .IN3(n3647), .QN(g11294) );
  NAND3X0 U4057 ( .IN1(n3648), .IN2(n3649), .IN3(n2741), .QN(n3647) );
  NAND3X0 U4058 ( .IN1(n3650), .IN2(n3651), .IN3(g1690), .QN(n3649) );
  NAND2X0 U4059 ( .IN1(n3652), .IN2(n3653), .QN(n3651) );
  NAND2X0 U4060 ( .IN1(n25), .IN2(n38), .QN(n3653) );
  NAND2X0 U4061 ( .IN1(n32), .IN2(n16), .QN(n3652) );
  NAND2X0 U4062 ( .IN1(n3654), .IN2(n3655), .QN(n3650) );
  NAND2X0 U4063 ( .IN1(n114), .IN2(n44), .QN(n3655) );
  NAND2X0 U4064 ( .IN1(g10726), .IN2(n42), .QN(n3654) );
  NAND3X0 U4065 ( .IN1(n3656), .IN2(n3657), .IN3(n1653), .QN(n3648) );
  NAND2X0 U4066 ( .IN1(n3112), .IN2(n3658), .QN(n3657) );
  NAND2X0 U4067 ( .IN1(g1796), .IN2(g1801), .QN(n3658) );
  NAND2X0 U4068 ( .IN1(g1791), .IN2(g1786), .QN(n3112) );
  NAND2X0 U4069 ( .IN1(n3659), .IN2(n3660), .QN(n3656) );
  NAND2X0 U4070 ( .IN1(g1781), .IN2(g1776), .QN(n3660) );
  NAND2X0 U4071 ( .IN1(test_so5), .IN2(g1766), .QN(n3659) );
  NAND2X0 U4072 ( .IN1(n3142), .IN2(g1857), .QN(n3646) );
  INVX0 U4073 ( .INP(n3167), .ZN(n3142) );
  NAND2X0 U4074 ( .IN1(n2587), .IN2(n367), .QN(n3167) );
  INVX0 U4075 ( .INP(n926), .ZN(n367) );
  NAND3X0 U4076 ( .IN1(n926), .IN2(n3661), .IN3(n1682), .QN(n3645) );
  NAND4X0 U4077 ( .IN1(n817), .IN2(n822), .IN3(n2602), .IN4(n2591), .QN(n3661)
         );
  NAND2X0 U4078 ( .IN1(g1814), .IN2(g1828), .QN(n817) );
  NAND2X0 U4079 ( .IN1(n3662), .IN2(n3663), .QN(g11293) );
  NAND2X0 U4080 ( .IN1(n3664), .IN2(n2587), .QN(n3663) );
  NAND2X0 U4081 ( .IN1(n2591), .IN2(n3665), .QN(n3664) );
  NAND2X0 U4082 ( .IN1(n3666), .IN2(g1854), .QN(n3665) );
  NAND4X0 U4083 ( .IN1(g4904), .IN2(n3667), .IN3(n3668), .IN4(n3669), .QN(
        n3666) );
  NAND2X0 U4084 ( .IN1(n3670), .IN2(g1857), .QN(n3669) );
  XOR2X1 U4085 ( .IN1(n2602), .IN2(n3671), .Q(n3670) );
  NAND2X0 U4086 ( .IN1(n1682), .IN2(n3672), .QN(n3668) );
  XOR2X1 U4087 ( .IN1(n1380), .IN2(n3671), .Q(n3672) );
  NAND4X0 U4088 ( .IN1(n1380), .IN2(n822), .IN3(n2602), .IN4(n2917), .QN(n3667) );
  NAND4X0 U4089 ( .IN1(n2301), .IN2(n1655), .IN3(n1605), .IN4(g1814), .QN(
        n2917) );
  NAND2X0 U4090 ( .IN1(n1608), .IN2(g1822), .QN(n2602) );
  NAND2X0 U4091 ( .IN1(n1605), .IN2(g1822), .QN(n822) );
  AND2X1 U4092 ( .IN1(n3170), .IN2(n3044), .Q(g4904) );
  INVX0 U4093 ( .INP(n2358), .ZN(n3170) );
  NAND2X0 U4094 ( .IN1(n2587), .IN2(n3673), .QN(n2358) );
  NAND2X0 U4095 ( .IN1(n1608), .IN2(g1834), .QN(n3673) );
  NAND3X0 U4096 ( .IN1(n1643), .IN2(g1828), .IN3(n1608), .QN(n2591) );
  NAND2X0 U4097 ( .IN1(n3674), .IN2(n2741), .QN(n3662) );
  INVX0 U4098 ( .INP(n2587), .ZN(n2741) );
  NAND4X0 U4099 ( .IN1(n1608), .IN2(n1643), .IN3(n1655), .IN4(n1605), .QN(
        n2587) );
  NAND2X0 U4100 ( .IN1(n3675), .IN2(n3676), .QN(n3674) );
  NAND2X0 U4101 ( .IN1(n3677), .IN2(g1690), .QN(n3676) );
  NAND2X0 U4102 ( .IN1(n1653), .IN2(n2340), .QN(n3675) );
  NOR2X0 U4103 ( .IN1(n3678), .IN2(n3623), .QN(g11292) );
  NOR2X0 U4104 ( .IN1(n3679), .IN2(g382), .QN(n3678) );
  NOR2X0 U4105 ( .IN1(n3680), .IN2(n3623), .QN(g11291) );
  NOR2X0 U4106 ( .IN1(n3681), .IN2(n3682), .QN(n3680) );
  NOR2X0 U4107 ( .IN1(n2225), .IN2(n3679), .QN(n3682) );
  NOR3X0 U4108 ( .IN1(n40), .IN2(n1420), .IN3(n2351), .QN(n3679) );
  INVX0 U4109 ( .INP(n3683), .ZN(n40) );
  NOR3X0 U4110 ( .IN1(n3621), .IN2(n2227), .IN3(n3683), .QN(n3681) );
  NOR3X0 U4111 ( .IN1(n2226), .IN2(n2227), .IN3(n2225), .QN(n3683) );
  NOR2X0 U4112 ( .IN1(n3623), .IN2(n3684), .QN(g11290) );
  XNOR2X1 U4113 ( .IN1(n2227), .IN2(n3621), .Q(n3684) );
  OR3X1 U4114 ( .IN1(n1420), .IN2(n2226), .IN3(n2351), .Q(n3621) );
  NAND2X0 U4115 ( .IN1(n2116), .IN2(g109), .QN(n3623) );
  NAND2X0 U4116 ( .IN1(n3685), .IN2(n3686), .QN(g11270) );
  NAND2X0 U4117 ( .IN1(n2351), .IN2(g421), .QN(n3686) );
  NAND2X0 U4118 ( .IN1(n14), .IN2(g416), .QN(n3685) );
  NAND2X0 U4119 ( .IN1(n3687), .IN2(n3688), .QN(g11269) );
  NAND2X0 U4120 ( .IN1(n2351), .IN2(g416), .QN(n3688) );
  NAND2X0 U4121 ( .IN1(n14), .IN2(g411), .QN(n3687) );
  NAND2X0 U4122 ( .IN1(n3689), .IN2(n3690), .QN(g11268) );
  NAND2X0 U4123 ( .IN1(n2351), .IN2(g411), .QN(n3690) );
  NAND2X0 U4124 ( .IN1(n14), .IN2(g406), .QN(n3689) );
  NAND2X0 U4125 ( .IN1(n3691), .IN2(n3692), .QN(g11267) );
  NAND2X0 U4126 ( .IN1(n2351), .IN2(g406), .QN(n3692) );
  NAND2X0 U4127 ( .IN1(n14), .IN2(g401), .QN(n3691) );
  NAND2X0 U4128 ( .IN1(n3693), .IN2(n3694), .QN(g11266) );
  NAND2X0 U4129 ( .IN1(n2351), .IN2(g401), .QN(n3694) );
  NAND2X0 U4130 ( .IN1(n14), .IN2(g396), .QN(n3693) );
  NAND2X0 U4131 ( .IN1(n3695), .IN2(n3696), .QN(g11265) );
  NAND2X0 U4132 ( .IN1(n2351), .IN2(g396), .QN(n3696) );
  NAND2X0 U4133 ( .IN1(n14), .IN2(g391), .QN(n3695) );
  NAND2X0 U4134 ( .IN1(n3697), .IN2(n3698), .QN(g11264) );
  NAND2X0 U4135 ( .IN1(n2351), .IN2(g391), .QN(n3698) );
  NAND2X0 U4136 ( .IN1(n14), .IN2(g386), .QN(n3697) );
  NAND2X0 U4137 ( .IN1(n3699), .IN2(n3700), .QN(g11263) );
  NAND2X0 U4138 ( .IN1(n2351), .IN2(g386), .QN(n3700) );
  NAND2X0 U4139 ( .IN1(n14), .IN2(g426), .QN(n3699) );
  NAND2X0 U4140 ( .IN1(n3701), .IN2(n3702), .QN(g11262) );
  NAND2X0 U4141 ( .IN1(n2351), .IN2(g431), .QN(n3702) );
  NAND2X0 U4142 ( .IN1(n14), .IN2(g435), .QN(n3701) );
  NAND2X0 U4143 ( .IN1(n3703), .IN2(n3704), .QN(g11261) );
  NAND2X0 U4144 ( .IN1(n2351), .IN2(g435), .QN(n3704) );
  NAND2X0 U4145 ( .IN1(n14), .IN2(g440), .QN(n3703) );
  NAND2X0 U4146 ( .IN1(n3705), .IN2(n3706), .QN(g11260) );
  NAND2X0 U4147 ( .IN1(n2351), .IN2(g440), .QN(n3706) );
  NAND2X0 U4148 ( .IN1(n14), .IN2(g444), .QN(n3705) );
  NAND2X0 U4149 ( .IN1(n3707), .IN2(n3708), .QN(g11259) );
  NAND2X0 U4150 ( .IN1(n2351), .IN2(g444), .QN(n3708) );
  NAND2X0 U4151 ( .IN1(n14), .IN2(g448), .QN(n3707) );
  NAND2X0 U4152 ( .IN1(n3709), .IN2(n3710), .QN(g11258) );
  NAND2X0 U4153 ( .IN1(n2351), .IN2(g448), .QN(n3710) );
  NAND2X0 U4154 ( .IN1(n14), .IN2(g452), .QN(n3709) );
  NAND2X0 U4155 ( .IN1(n3711), .IN2(n3712), .QN(g11257) );
  NAND2X0 U4156 ( .IN1(n2351), .IN2(g452), .QN(n3712) );
  NAND2X0 U4157 ( .IN1(n14), .IN2(g421), .QN(n3711) );
  NAND2X0 U4158 ( .IN1(n3713), .IN2(n3714), .QN(g11256) );
  NAND2X0 U4159 ( .IN1(n2351), .IN2(g426), .QN(n3714) );
  NAND2X0 U4160 ( .IN1(n3578), .IN2(n14), .QN(n3713) );
  NOR4X0 U4161 ( .IN1(g837), .IN2(g861), .IN3(n3715), .IN4(n3716), .QN(n2351)
         );
  NAND4X0 U4162 ( .IN1(n2103), .IN2(n2102), .IN3(n3717), .IN4(n2079), .QN(
        n3716) );
  NOR2X0 U4163 ( .IN1(g841), .IN2(g857), .QN(n3717) );
  NAND3X0 U4164 ( .IN1(n1651), .IN2(n3718), .IN3(n2074), .QN(n3715) );
  NAND3X0 U4165 ( .IN1(n3719), .IN2(n3720), .IN3(n3721), .QN(n3718) );
  NAND2X0 U4166 ( .IN1(n3722), .IN2(g109), .QN(n3721) );
  NAND2X0 U4167 ( .IN1(n3723), .IN2(n3724), .QN(n3722) );
  AND2X1 U4168 ( .IN1(n3725), .IN2(n3726), .Q(n3578) );
  NAND2X0 U4169 ( .IN1(n1681), .IN2(n3625), .QN(n3726) );
  INVX0 U4170 ( .INP(n1420), .ZN(n3625) );
  NAND2X0 U4171 ( .IN1(n3727), .IN2(n1420), .QN(n3725) );
  NAND2X0 U4172 ( .IN1(n3728), .IN2(n3729), .QN(n3727) );
  NAND2X0 U4173 ( .IN1(g431), .IN2(g435), .QN(n3729) );
  NAND3X0 U4174 ( .IN1(n1876), .IN2(n3730), .IN3(n1878), .QN(n3728) );
  NAND4X0 U4175 ( .IN1(n3731), .IN2(n2309), .IN3(n3732), .IN4(n3733), .QN(
        n3730) );
  NOR4X0 U4176 ( .IN1(n3734), .IN2(g396), .IN3(g448), .IN4(g452), .QN(n3733)
         );
  NAND4X0 U4177 ( .IN1(n2250), .IN2(n2249), .IN3(n2241), .IN4(n2248), .QN(
        n3734) );
  AND3X1 U4178 ( .IN1(n2274), .IN2(n2272), .IN3(n2290), .Q(n3732) );
  NOR2X0 U4179 ( .IN1(g411), .IN2(g426), .QN(n3731) );
  NOR2X0 U4180 ( .IN1(n3735), .IN2(n3736), .QN(g11206) );
  XOR2X1 U4181 ( .IN1(n3737), .IN2(n3735), .Q(g11163) );
  NAND3X0 U4182 ( .IN1(n3738), .IN2(n3739), .IN3(n3740), .QN(n3735) );
  NAND2X0 U4183 ( .IN1(g5392), .IN2(n44), .QN(n3740) );
  NOR2X0 U4184 ( .IN1(n3340), .IN2(n2362), .QN(g5392) );
  NAND2X0 U4185 ( .IN1(g1765), .IN2(g1610), .QN(n3340) );
  NAND2X0 U4186 ( .IN1(n3741), .IN2(g109), .QN(n3739) );
  NAND3X0 U4187 ( .IN1(n3742), .IN2(n3743), .IN3(n3744), .QN(n3741) );
  NAND2X0 U4188 ( .IN1(n2095), .IN2(g10726), .QN(n3744) );
  NAND2X0 U4189 ( .IN1(n114), .IN2(g2648), .QN(n3743) );
  NAND2X0 U4190 ( .IN1(n3745), .IN2(n3036), .QN(n3742) );
  NAND2X0 U4191 ( .IN1(n3305), .IN2(n42), .QN(n3738) );
  AND3X1 U4192 ( .IN1(DFF_194_n1), .IN2(g3069), .IN3(g109), .Q(n3305) );
  NAND2X0 U4193 ( .IN1(n3746), .IN2(n3747), .QN(g10936) );
  NAND2X0 U4194 ( .IN1(n1054), .IN2(g1811), .QN(n3747) );
  NAND2X0 U4195 ( .IN1(n1391), .IN2(n263), .QN(n3746) );
  NAND4X0 U4196 ( .IN1(n3745), .IN2(n3724), .IN3(n3469), .IN4(n3748), .QN(
        n1391) );
  INVX0 U4197 ( .INP(n3749), .ZN(n3724) );
  NAND2X0 U4198 ( .IN1(n3750), .IN2(n3751), .QN(g10898) );
  OR2X1 U4199 ( .IN1(n2795), .IN2(n2095), .Q(n3751) );
  NAND2X0 U4200 ( .IN1(n3752), .IN2(n2795), .QN(n3750) );
  NAND2X0 U4201 ( .IN1(n3753), .IN2(n3365), .QN(n3752) );
  NAND2X0 U4202 ( .IN1(n3469), .IN2(n3754), .QN(n3365) );
  NAND2X0 U4203 ( .IN1(n2563), .IN2(n2565), .QN(n3469) );
  AND3X1 U4204 ( .IN1(g42), .IN2(n2562), .IN3(n2560), .Q(n2563) );
  AND4X1 U4205 ( .IN1(n2583), .IN2(n3755), .IN3(n3756), .IN4(n3757), .Q(n2560)
         );
  NOR2X0 U4206 ( .IN1(g48), .IN2(g45), .QN(n3756) );
  XOR3X1 U4207 ( .IN1(test_so8), .IN2(n2229), .IN3(n3758), .Q(n3753) );
  XOR2X1 U4208 ( .IN1(n3759), .IN2(n3760), .Q(n3758) );
  XOR3X1 U4209 ( .IN1(n2306), .IN2(n2304), .IN3(n3761), .Q(n3760) );
  XOR2X1 U4210 ( .IN1(test_so2), .IN2(n2350), .Q(n3761) );
  XOR3X1 U4211 ( .IN1(n2203), .IN2(n1871), .IN3(n3762), .Q(n3759) );
  XNOR2X1 U4212 ( .IN1(n2228), .IN2(n2267), .Q(n3762) );
  NAND2X0 U4213 ( .IN1(n3763), .IN2(n3764), .QN(g10866) );
  NAND2X0 U4214 ( .IN1(n968), .IN2(g1684), .QN(n3764) );
  NAND2X0 U4215 ( .IN1(n3765), .IN2(n3766), .QN(g10865) );
  NAND2X0 U4216 ( .IN1(n3266), .IN2(g1669), .QN(n3766) );
  NAND3X0 U4217 ( .IN1(n1404), .IN2(n3767), .IN3(n3265), .QN(n3765) );
  NAND2X0 U4218 ( .IN1(n3768), .IN2(g109), .QN(n3767) );
  NAND2X0 U4219 ( .IN1(n3769), .IN2(n3770), .QN(g10864) );
  NAND2X0 U4220 ( .IN1(n968), .IN2(g1681), .QN(n3770) );
  NAND2X0 U4221 ( .IN1(n3771), .IN2(n3772), .QN(g10863) );
  NAND2X0 U4222 ( .IN1(n3266), .IN2(g1666), .QN(n3772) );
  NAND3X0 U4223 ( .IN1(n3773), .IN2(n3774), .IN3(n3265), .QN(n3771) );
  NAND2X0 U4224 ( .IN1(n1611), .IN2(n3720), .QN(n3773) );
  NAND2X0 U4225 ( .IN1(n3775), .IN2(n3776), .QN(g10862) );
  NAND2X0 U4226 ( .IN1(n968), .IN2(g1678), .QN(n3776) );
  NAND2X0 U4227 ( .IN1(n3777), .IN2(n3778), .QN(g10861) );
  NAND2X0 U4228 ( .IN1(n3266), .IN2(g1663), .QN(n3778) );
  NAND2X0 U4229 ( .IN1(n3265), .IN2(n3779), .QN(n3777) );
  NAND2X0 U4230 ( .IN1(n3780), .IN2(n3781), .QN(g10860) );
  NAND2X0 U4231 ( .IN1(n968), .IN2(g1675), .QN(n3781) );
  NAND2X0 U4232 ( .IN1(n3782), .IN2(n3783), .QN(g10859) );
  NAND2X0 U4233 ( .IN1(n3266), .IN2(g1660), .QN(n3783) );
  NAND2X0 U4234 ( .IN1(n3265), .IN2(n3784), .QN(n3782) );
  NAND2X0 U4235 ( .IN1(n3785), .IN2(n3786), .QN(g10858) );
  NAND2X0 U4236 ( .IN1(n968), .IN2(g1672), .QN(n3786) );
  NAND2X0 U4237 ( .IN1(n3787), .IN2(n3788), .QN(g10855) );
  NAND2X0 U4238 ( .IN1(n968), .IN2(g549), .QN(n3788) );
  NAND2X0 U4239 ( .IN1(n3779), .IN2(n2795), .QN(n3787) );
  NAND3X0 U4240 ( .IN1(n3789), .IN2(n3790), .IN3(n1611), .QN(n3779) );
  NAND3X0 U4241 ( .IN1(g109), .IN2(n32), .IN3(n3774), .QN(n3790) );
  NAND2X0 U4242 ( .IN1(n2985), .IN2(n3791), .QN(n3789) );
  NAND2X0 U4243 ( .IN1(n3792), .IN2(n3284), .QN(n2985) );
  NAND2X0 U4244 ( .IN1(g18), .IN2(g192), .QN(n3284) );
  NAND2X0 U4245 ( .IN1(n2569), .IN2(g1512), .QN(n3792) );
  NAND2X0 U4246 ( .IN1(n2359), .IN2(n3737), .QN(g10801) );
  INVX0 U4247 ( .INP(n17), .ZN(n3737) );
  XNOR3X1 U4248 ( .IN1(n1858), .IN2(n3793), .IN3(n3794), .Q(n17) );
  NAND3X0 U4249 ( .IN1(n3795), .IN2(n3796), .IN3(n3749), .QN(n3794) );
  NAND3X0 U4250 ( .IN1(n3797), .IN2(n3798), .IN3(n3677), .QN(n3749) );
  NAND2X0 U4251 ( .IN1(n3799), .IN2(n16), .QN(n3796) );
  XOR2X1 U4252 ( .IN1(n32), .IN2(n42), .Q(n3799) );
  NAND3X0 U4253 ( .IN1(n42), .IN2(n32), .IN3(n3677), .QN(n3795) );
  XOR2X1 U4254 ( .IN1(n3800), .IN2(n3801), .Q(n3793) );
  NAND3X0 U4255 ( .IN1(n3802), .IN2(n3803), .IN3(n3804), .QN(n3801) );
  INVX0 U4256 ( .INP(n3723), .ZN(n3804) );
  NOR3X0 U4257 ( .IN1(n114), .IN2(n44), .IN3(g10726), .QN(n3723) );
  NAND2X0 U4258 ( .IN1(n3805), .IN2(g10726), .QN(n3803) );
  XOR2X1 U4259 ( .IN1(n44), .IN2(n114), .Q(n3805) );
  NAND3X0 U4260 ( .IN1(n114), .IN2(n44), .IN3(n3470), .QN(n3802) );
  NAND2X0 U4261 ( .IN1(n4113), .IN2(n3806), .QN(n3800) );
  XOR2X1 U4262 ( .IN1(n3768), .IN2(n38), .Q(n1858) );
  NAND2X0 U4263 ( .IN1(n3807), .IN2(n3808), .QN(g10800) );
  NAND2X0 U4264 ( .IN1(n968), .IN2(g575), .QN(n3808) );
  NAND2X0 U4265 ( .IN1(n3784), .IN2(n2795), .QN(n3807) );
  NAND3X0 U4266 ( .IN1(n3809), .IN2(n3810), .IN3(n1611), .QN(n3784) );
  NAND2X0 U4267 ( .IN1(n3811), .IN2(n3774), .QN(n3810) );
  NAND2X0 U4268 ( .IN1(n3677), .IN2(g109), .QN(n3811) );
  NAND2X0 U4269 ( .IN1(n2980), .IN2(n3791), .QN(n3809) );
  NAND2X0 U4270 ( .IN1(n3812), .IN2(n3286), .QN(n2980) );
  NAND2X0 U4271 ( .IN1(g18), .IN2(g248), .QN(n3286) );
  NAND2X0 U4272 ( .IN1(n2569), .IN2(g1636), .QN(n3812) );
  NAND2X0 U4273 ( .IN1(n3813), .IN2(n3814), .QN(g10799) );
  NAND2X0 U4274 ( .IN1(n968), .IN2(g566), .QN(n3814) );
  NAND2X0 U4275 ( .IN1(n3763), .IN2(n3815), .QN(g10798) );
  NAND2X0 U4276 ( .IN1(n968), .IN2(g563), .QN(n3815) );
  NAND2X0 U4277 ( .IN1(n3816), .IN2(n2795), .QN(n3763) );
  NAND2X0 U4278 ( .IN1(n3817), .IN2(n3818), .QN(n3816) );
  NAND2X0 U4279 ( .IN1(n3791), .IN2(n2983), .QN(n3818) );
  NAND2X0 U4280 ( .IN1(n2815), .IN2(n3819), .QN(n2983) );
  NAND2X0 U4281 ( .IN1(n2569), .IN2(g1624), .QN(n3819) );
  OR2X1 U4282 ( .IN1(n2569), .IN2(n2282), .Q(n2815) );
  NAND2X0 U4283 ( .IN1(n1404), .IN2(n3671), .QN(n3817) );
  NAND2X0 U4284 ( .IN1(n3769), .IN2(n3820), .QN(g10797) );
  NAND2X0 U4285 ( .IN1(n968), .IN2(g560), .QN(n3820) );
  NAND2X0 U4286 ( .IN1(n3821), .IN2(n2795), .QN(n3769) );
  NAND2X0 U4287 ( .IN1(n3822), .IN2(n3823), .QN(n3821) );
  NAND2X0 U4288 ( .IN1(n3791), .IN2(n2978), .QN(n3823) );
  NAND2X0 U4289 ( .IN1(n2806), .IN2(n3824), .QN(n2978) );
  NAND2X0 U4290 ( .IN1(n2569), .IN2(g1621), .QN(n3824) );
  NAND2X0 U4291 ( .IN1(g18), .IN2(g219), .QN(n2806) );
  NAND2X0 U4292 ( .IN1(n1404), .IN2(n3745), .QN(n3822) );
  NAND2X0 U4293 ( .IN1(n3775), .IN2(n3825), .QN(g10795) );
  NAND2X0 U4294 ( .IN1(n968), .IN2(g557), .QN(n3825) );
  NAND2X0 U4295 ( .IN1(n3826), .IN2(n2795), .QN(n3775) );
  NAND2X0 U4296 ( .IN1(n3827), .IN2(n3828), .QN(n3826) );
  NAND2X0 U4297 ( .IN1(n3791), .IN2(n2970), .QN(n3828) );
  NAND2X0 U4298 ( .IN1(n2849), .IN2(n3829), .QN(n2970) );
  NAND2X0 U4299 ( .IN1(n2569), .IN2(g1615), .QN(n3829) );
  OR2X1 U4300 ( .IN1(n2569), .IN2(n2123), .Q(n2849) );
  NAND2X0 U4301 ( .IN1(n1404), .IN2(n3830), .QN(n3827) );
  NAND2X0 U4302 ( .IN1(n3780), .IN2(n3831), .QN(g10793) );
  NAND2X0 U4303 ( .IN1(n968), .IN2(g554), .QN(n3831) );
  NAND3X0 U4304 ( .IN1(n3832), .IN2(n2795), .IN3(n3833), .QN(n3780) );
  NAND2X0 U4305 ( .IN1(n3791), .IN2(n2966), .QN(n3833) );
  AND2X1 U4306 ( .IN1(n2838), .IN2(n3834), .Q(n2966) );
  NAND2X0 U4307 ( .IN1(n2569), .IN2(g1639), .QN(n3834) );
  OR2X1 U4308 ( .IN1(n2569), .IN2(n2122), .Q(n2838) );
  NAND3X0 U4309 ( .IN1(n3797), .IN2(g109), .IN3(n1404), .QN(n3832) );
  NAND2X0 U4310 ( .IN1(n3785), .IN2(n3835), .QN(g10791) );
  NAND2X0 U4311 ( .IN1(n968), .IN2(g546), .QN(n3835) );
  NAND2X0 U4312 ( .IN1(n3836), .IN2(n2795), .QN(n3785) );
  NAND2X0 U4313 ( .IN1(n3837), .IN2(n3838), .QN(n3836) );
  NAND3X0 U4314 ( .IN1(n16), .IN2(g109), .IN3(n1404), .QN(n3838) );
  NAND2X0 U4315 ( .IN1(n3791), .IN2(n2987), .QN(n3837) );
  NAND2X0 U4316 ( .IN1(n2826), .IN2(n3839), .QN(n2987) );
  NAND2X0 U4317 ( .IN1(n2569), .IN2(g1618), .QN(n3839) );
  OR2X1 U4318 ( .IN1(n2569), .IN2(n2121), .Q(n2826) );
  NOR2X0 U4319 ( .IN1(n4120), .IN2(n263), .QN(g10785) );
  NOR2X0 U4320 ( .IN1(n4119), .IN2(n263), .QN(g10784) );
  NOR2X0 U4321 ( .IN1(n4117), .IN2(n263), .QN(g10782) );
  NOR2X0 U4322 ( .IN1(n4123), .IN2(n263), .QN(g10780) );
  INVX0 U4323 ( .INP(n1054), .ZN(n263) );
  NAND2X0 U4324 ( .IN1(g1696), .IN2(n2349), .QN(n1054) );
  NAND2X0 U4325 ( .IN1(n3813), .IN2(n3840), .QN(g10776) );
  NAND2X0 U4326 ( .IN1(n968), .IN2(g1687), .QN(n3840) );
  NAND2X0 U4327 ( .IN1(n3841), .IN2(n2795), .QN(n3813) );
  NAND3X0 U4328 ( .IN1(n3842), .IN2(n3843), .IN3(n3844), .QN(n3841) );
  NAND2X0 U4329 ( .IN1(n1404), .IN2(g10726), .QN(n3844) );
  NAND2X0 U4330 ( .IN1(n3791), .IN2(n2989), .QN(n3842) );
  NAND2X0 U4331 ( .IN1(n2832), .IN2(n3845), .QN(n2989) );
  NAND2X0 U4332 ( .IN1(n2569), .IN2(g1627), .QN(n3845) );
  OR2X1 U4333 ( .IN1(n2569), .IN2(n2283), .Q(n2832) );
  NAND2X0 U4334 ( .IN1(n3846), .IN2(n3847), .QN(g10773) );
  NAND2X0 U4335 ( .IN1(n3848), .IN2(g1727), .QN(n3847) );
  NAND2X0 U4336 ( .IN1(n3335), .IN2(n3830), .QN(n3846) );
  NAND2X0 U4337 ( .IN1(n3849), .IN2(n3850), .QN(g10771) );
  NAND2X0 U4338 ( .IN1(n3848), .IN2(g1724), .QN(n3850) );
  NAND3X0 U4339 ( .IN1(g109), .IN2(n32), .IN3(n3335), .QN(n3849) );
  NAND2X0 U4340 ( .IN1(n3851), .IN2(n3852), .QN(g10770) );
  NAND2X0 U4341 ( .IN1(n3848), .IN2(g1721), .QN(n3852) );
  NAND3X0 U4342 ( .IN1(g109), .IN2(n16), .IN3(n3335), .QN(n3851) );
  NAND2X0 U4343 ( .IN1(n3853), .IN2(n3854), .QN(g10767) );
  NAND2X0 U4344 ( .IN1(n3266), .IN2(g1657), .QN(n3854) );
  NAND2X0 U4345 ( .IN1(n3265), .IN2(n3855), .QN(n3853) );
  NAND2X0 U4346 ( .IN1(n3856), .IN2(n3857), .QN(g10765) );
  NAND2X0 U4347 ( .IN1(n3266), .IN2(g1654), .QN(n3857) );
  INVX0 U4348 ( .INP(n3265), .ZN(n3266) );
  NAND2X0 U4349 ( .IN1(n3265), .IN2(n3858), .QN(n3856) );
  NOR2X0 U4350 ( .IN1(g1696), .IN2(n2349), .QN(n3265) );
  INVX0 U4351 ( .INP(n3470), .ZN(g10726) );
  NAND2X0 U4352 ( .IN1(n3859), .IN2(n3860), .QN(g10718) );
  NAND2X0 U4353 ( .IN1(n968), .IN2(g572), .QN(n3860) );
  NAND2X0 U4354 ( .IN1(n3855), .IN2(n2795), .QN(n3859) );
  NAND3X0 U4355 ( .IN1(n3861), .IN2(n3862), .IN3(n1611), .QN(n3855) );
  NAND3X0 U4356 ( .IN1(g109), .IN2(n114), .IN3(n3774), .QN(n3862) );
  NAND4X0 U4357 ( .IN1(n3863), .IN2(n3864), .IN3(n3865), .IN4(n3866), .QN(n114) );
  NOR4X0 U4358 ( .IN1(n3867), .IN2(n3868), .IN3(n3869), .IN4(n3870), .QN(n3866) );
  NOR2X0 U4359 ( .IN1(n2073), .IN2(n3871), .QN(n3870) );
  NOR2X0 U4360 ( .IN1(n4115), .IN2(n3872), .QN(n3869) );
  NAND2X0 U4361 ( .IN1(n3873), .IN2(n3874), .QN(n3868) );
  NAND2X0 U4362 ( .IN1(n1486), .IN2(g1546), .QN(n3874) );
  NAND2X0 U4363 ( .IN1(g1191), .IN2(n3875), .QN(n3873) );
  NOR2X0 U4364 ( .IN1(n2175), .IN2(n3876), .QN(n3867) );
  AND3X1 U4365 ( .IN1(n3877), .IN2(n3878), .IN3(n3879), .Q(n3865) );
  NAND2X0 U4366 ( .IN1(test_so9), .IN2(n3880), .QN(n3879) );
  NAND4X0 U4367 ( .IN1(n3881), .IN2(n3882), .IN3(n1478), .IN4(n3883), .QN(
        n3878) );
  NAND2X0 U4368 ( .IN1(n3884), .IN2(g1741), .QN(n3877) );
  NAND2X0 U4369 ( .IN1(g919), .IN2(n3885), .QN(n3864) );
  NAND2X0 U4370 ( .IN1(n1485), .IN2(g1589), .QN(n3863) );
  NAND2X0 U4371 ( .IN1(n2972), .IN2(n3791), .QN(n3861) );
  NAND2X0 U4372 ( .IN1(n3886), .IN2(n3288), .QN(n2972) );
  NAND2X0 U4373 ( .IN1(g18), .IN2(g243), .QN(n3288) );
  NAND2X0 U4374 ( .IN1(n2569), .IN2(g1633), .QN(n3886) );
  NAND2X0 U4375 ( .IN1(n3887), .IN2(n3888), .QN(g10717) );
  NAND2X0 U4376 ( .IN1(n968), .IN2(g569), .QN(n3888) );
  NAND2X0 U4377 ( .IN1(n3858), .IN2(n2795), .QN(n3887) );
  INVX0 U4378 ( .INP(n968), .ZN(n2795) );
  NAND2X0 U4379 ( .IN1(n2349), .IN2(n3889), .QN(n968) );
  NAND3X0 U4380 ( .IN1(n3890), .IN2(n3843), .IN3(n3891), .QN(n3858) );
  NAND2X0 U4381 ( .IN1(n1404), .IN2(n44), .QN(n3891) );
  INVX0 U4382 ( .INP(n3754), .ZN(n44) );
  NOR2X0 U4383 ( .IN1(g1718), .IN2(n3791), .QN(n1404) );
  INVX0 U4384 ( .INP(n1450), .ZN(n3843) );
  NAND2X0 U4385 ( .IN1(n3791), .IN2(n2991), .QN(n3890) );
  NAND2X0 U4386 ( .IN1(n2844), .IN2(n3892), .QN(n2991) );
  NAND2X0 U4387 ( .IN1(n2569), .IN2(g1630), .QN(n3892) );
  OR2X1 U4388 ( .IN1(n2569), .IN2(n2284), .Q(n2844) );
  INVX0 U4389 ( .INP(g18), .ZN(n2569) );
  INVX0 U4390 ( .INP(n3774), .ZN(n3791) );
  NAND2X0 U4391 ( .IN1(n4130), .IN2(n1611), .QN(n3774) );
  NAND2X0 U4392 ( .IN1(n3893), .IN2(n3894), .QN(g10711) );
  NAND2X0 U4393 ( .IN1(n3848), .IN2(g1733), .QN(n3894) );
  NAND2X0 U4394 ( .IN1(n3335), .IN2(n3671), .QN(n3893) );
  NAND2X0 U4395 ( .IN1(g109), .IN2(n3798), .QN(n3671) );
  NAND2X0 U4396 ( .IN1(n3895), .IN2(n3896), .QN(g10707) );
  NAND2X0 U4397 ( .IN1(n3848), .IN2(g1730), .QN(n3896) );
  INVX0 U4398 ( .INP(n3335), .ZN(n3848) );
  NAND2X0 U4399 ( .IN1(n3335), .IN2(n3745), .QN(n3895) );
  NOR2X0 U4400 ( .IN1(n3889), .IN2(n2349), .QN(n3335) );
  INVX0 U4401 ( .INP(g1696), .ZN(n3889) );
  INVX0 U4402 ( .INP(n3736), .ZN(g10628) );
  NAND2X0 U4403 ( .IN1(n3897), .IN2(n3898), .QN(n3736) );
  NAND2X0 U4404 ( .IN1(n3899), .IN2(g109), .QN(n3898) );
  NAND4X0 U4405 ( .IN1(n3900), .IN2(n3901), .IN3(n3902), .IN4(n3903), .QN(
        n3899) );
  NAND2X0 U4406 ( .IN1(n2555), .IN2(n42), .QN(n3903) );
  INVX0 U4407 ( .INP(n3798), .ZN(n42) );
  AND2X1 U4408 ( .IN1(n2094), .IN2(g3007), .Q(n2555) );
  NAND2X0 U4409 ( .IN1(n3745), .IN2(n3064), .QN(n3902) );
  INVX0 U4410 ( .INP(n3719), .ZN(n3745) );
  NAND2X0 U4411 ( .IN1(n25), .IN2(g109), .QN(n3719) );
  INVX0 U4412 ( .INP(n3768), .ZN(n25) );
  NOR4X0 U4413 ( .IN1(n3904), .IN2(n3905), .IN3(n3906), .IN4(n3907), .QN(n3768) );
  NAND4X0 U4414 ( .IN1(n3908), .IN2(n3909), .IN3(n3910), .IN4(n3911), .QN(
        n3907) );
  NOR4X0 U4415 ( .IN1(n3912), .IN2(n3913), .IN3(n3914), .IN4(n3915), .QN(n3911) );
  NOR2X0 U4416 ( .IN1(n1722), .IN2(n3871), .QN(n3915) );
  NOR2X0 U4417 ( .IN1(n4114), .IN2(n3916), .QN(n3914) );
  NAND2X0 U4418 ( .IN1(n3917), .IN2(n3918), .QN(n3913) );
  NAND2X0 U4419 ( .IN1(n3919), .IN2(g8), .QN(n3918) );
  NAND2X0 U4420 ( .IN1(g895), .IN2(n3920), .QN(n3917) );
  NOR2X0 U4421 ( .IN1(n1712), .IN2(n3921), .QN(n3912) );
  AND3X1 U4422 ( .IN1(n3922), .IN2(n3923), .IN3(n3924), .Q(n3910) );
  NAND2X0 U4423 ( .IN1(n3884), .IN2(g1730), .QN(n3924) );
  NAND2X0 U4424 ( .IN1(n3925), .IN2(g1324), .QN(n3923) );
  NAND2X0 U4425 ( .IN1(g907), .IN2(n3885), .QN(n3922) );
  OR2X1 U4426 ( .IN1(n3882), .IN2(n1721), .Q(n3909) );
  NAND2X0 U4427 ( .IN1(g1179), .IN2(n3875), .QN(n3908) );
  NAND4X0 U4428 ( .IN1(n3926), .IN2(n3927), .IN3(n3928), .IN4(n3929), .QN(
        n3906) );
  NOR2X0 U4429 ( .IN1(n3930), .IN2(n3931), .QN(n3929) );
  AND2X1 U4430 ( .IN1(g1534), .IN2(n1486), .Q(n3931) );
  NOR2X0 U4431 ( .IN1(n2147), .IN2(n3932), .QN(n3930) );
  NAND2X0 U4432 ( .IN1(n1479), .IN2(g1558), .QN(n3928) );
  NAND2X0 U4433 ( .IN1(n382), .IN2(g1601), .QN(n3927) );
  NAND2X0 U4434 ( .IN1(g1203), .IN2(n1512), .QN(n3926) );
  NAND3X0 U4435 ( .IN1(n3933), .IN2(n3934), .IN3(n3935), .QN(n3905) );
  NAND2X0 U4436 ( .IN1(n3936), .IN2(g959), .QN(n3935) );
  NAND2X0 U4437 ( .IN1(n3937), .IN2(g1753), .QN(n3934) );
  NAND2X0 U4438 ( .IN1(n3048), .IN2(n3806), .QN(n3933) );
  NAND3X0 U4439 ( .IN1(n3938), .IN2(n3939), .IN3(n3940), .QN(n3904) );
  NAND2X0 U4440 ( .IN1(n3941), .IN2(g296), .QN(n3940) );
  NAND2X0 U4441 ( .IN1(n3942), .IN2(g272), .QN(n3938) );
  NAND2X0 U4442 ( .IN1(g881), .IN2(n32), .QN(n3901) );
  INVX0 U4443 ( .INP(n3797), .ZN(n32) );
  NAND2X0 U4444 ( .IN1(g877), .IN2(n16), .QN(n3900) );
  INVX0 U4445 ( .INP(n3677), .ZN(n16) );
  NAND2X0 U4446 ( .IN1(n3830), .IN2(n3254), .QN(n3897) );
  INVX0 U4447 ( .INP(n2962), .ZN(n3254) );
  NAND3X0 U4448 ( .IN1(DFF_121_n1), .IN2(g2986), .IN3(g109), .QN(n2962) );
  INVX0 U4449 ( .INP(n3720), .ZN(n3830) );
  NAND2X0 U4450 ( .IN1(n38), .IN2(g109), .QN(n3720) );
  INVX0 U4451 ( .INP(n3748), .ZN(n38) );
  NAND2X0 U4452 ( .IN1(n2359), .IN2(n3470), .QN(g10465) );
  NOR4X0 U4453 ( .IN1(n3943), .IN2(n3944), .IN3(n3945), .IN4(n3946), .QN(n3470) );
  NAND3X0 U4454 ( .IN1(n3947), .IN2(n3948), .IN3(n3949), .QN(n3946) );
  NAND2X0 U4455 ( .IN1(n3941), .IN2(g302), .QN(n3949) );
  NAND2X0 U4456 ( .IN1(g1185), .IN2(n3875), .QN(n3948) );
  NAND2X0 U4457 ( .IN1(n3942), .IN2(g278), .QN(n3947) );
  NAND4X0 U4458 ( .IN1(n3950), .IN2(n3951), .IN3(n3952), .IN4(n3953), .QN(
        n3945) );
  NAND2X0 U4459 ( .IN1(n1478), .IN2(n3954), .QN(n3953) );
  NAND2X0 U4460 ( .IN1(n382), .IN2(g1607), .QN(n3952) );
  NAND2X0 U4461 ( .IN1(n3925), .IN2(g1330), .QN(n3951) );
  NAND2X0 U4462 ( .IN1(g913), .IN2(n3885), .QN(n3950) );
  NAND3X0 U4463 ( .IN1(n3955), .IN2(n3956), .IN3(n3957), .QN(n3944) );
  NAND2X0 U4464 ( .IN1(n1486), .IN2(g1540), .QN(n3957) );
  NAND2X0 U4465 ( .IN1(n1479), .IN2(g1564), .QN(n3956) );
  NAND2X0 U4466 ( .IN1(n1485), .IN2(g1583), .QN(n3955) );
  NAND3X0 U4467 ( .IN1(n3958), .IN2(n3959), .IN3(n3960), .QN(n3943) );
  NAND2X0 U4468 ( .IN1(n3936), .IN2(g965), .QN(n3960) );
  NAND2X0 U4469 ( .IN1(n3937), .IN2(g1759), .QN(n3959) );
  NAND2X0 U4470 ( .IN1(n3806), .IN2(n1650), .QN(n3958) );
  NAND2X0 U4471 ( .IN1(n2359), .IN2(n3798), .QN(g10463) );
  NOR4X0 U4472 ( .IN1(n3961), .IN2(n3962), .IN3(n3963), .IN4(n3964), .QN(n3798) );
  NAND4X0 U4473 ( .IN1(n3965), .IN2(n3966), .IN3(n3967), .IN4(n3968), .QN(
        n3964) );
  NAND2X0 U4474 ( .IN1(n382), .IN2(g1604), .QN(n3968) );
  NAND2X0 U4475 ( .IN1(n1479), .IN2(g1561), .QN(n3967) );
  NAND2X0 U4476 ( .IN1(n1485), .IN2(g1580), .QN(n3966) );
  NAND2X0 U4477 ( .IN1(n1486), .IN2(g1537), .QN(n3965) );
  NAND4X0 U4478 ( .IN1(n3969), .IN2(n3970), .IN3(n3971), .IN4(n3972), .QN(
        n3963) );
  NAND2X0 U4479 ( .IN1(n3941), .IN2(g299), .QN(n3972) );
  NAND2X0 U4480 ( .IN1(n3937), .IN2(g1756), .QN(n3971) );
  NAND2X0 U4481 ( .IN1(n3806), .IN2(n3034), .QN(n3970) );
  NAND2X0 U4482 ( .IN1(n3936), .IN2(g962), .QN(n3969) );
  NAND4X0 U4483 ( .IN1(n3973), .IN2(n3974), .IN3(n3975), .IN4(n3976), .QN(
        n3962) );
  NAND2X0 U4484 ( .IN1(n3919), .IN2(n3025), .QN(n3976) );
  NAND2X0 U4485 ( .IN1(n3977), .IN2(n3978), .QN(n3975) );
  NAND2X0 U4486 ( .IN1(g1182), .IN2(n3875), .QN(n3974) );
  NAND2X0 U4487 ( .IN1(n3942), .IN2(g275), .QN(n3973) );
  NAND4X0 U4488 ( .IN1(n3979), .IN2(n3980), .IN3(n3981), .IN4(n3982), .QN(
        n3961) );
  NAND2X0 U4489 ( .IN1(n3983), .IN2(n3057), .QN(n3982) );
  INVX0 U4490 ( .INP(n3916), .ZN(n3983) );
  NAND2X0 U4491 ( .IN1(g910), .IN2(n3885), .QN(n3981) );
  NAND2X0 U4492 ( .IN1(n3925), .IN2(g1327), .QN(n3980) );
  NAND2X0 U4493 ( .IN1(n3884), .IN2(g1733), .QN(n3979) );
  NAND2X0 U4494 ( .IN1(n2359), .IN2(n3748), .QN(g10459) );
  NOR4X0 U4495 ( .IN1(n3984), .IN2(n3985), .IN3(n3986), .IN4(n3987), .QN(n3748) );
  NAND4X0 U4496 ( .IN1(n3939), .IN2(n3988), .IN3(n3989), .IN4(n3990), .QN(
        n3987) );
  NOR4X0 U4497 ( .IN1(n3991), .IN2(n3992), .IN3(n3993), .IN4(n3994), .QN(n3990) );
  NOR2X0 U4498 ( .IN1(n2085), .IN2(n1472), .QN(n3994) );
  NOR2X0 U4499 ( .IN1(n3872), .IN2(DFF_242_n1), .QN(n3993) );
  NOR2X0 U4500 ( .IN1(n2144), .IN2(n3995), .QN(n3992) );
  NAND3X0 U4501 ( .IN1(n3996), .IN2(n3997), .IN3(n3998), .QN(n3991) );
  NAND2X0 U4502 ( .IN1(n3937), .IN2(g1750), .QN(n3998) );
  NAND2X0 U4503 ( .IN1(n3942), .IN2(g269), .QN(n3997) );
  NAND2X0 U4504 ( .IN1(n3941), .IN2(g293), .QN(n3996) );
  AND3X1 U4505 ( .IN1(n3999), .IN2(n4000), .IN3(n4001), .Q(n3989) );
  NAND2X0 U4506 ( .IN1(n1485), .IN2(g1574), .QN(n4001) );
  NAND2X0 U4507 ( .IN1(n1512), .IN2(g1200), .QN(n4000) );
  NAND2X0 U4508 ( .IN1(n1479), .IN2(g1555), .QN(n3999) );
  NAND2X0 U4509 ( .IN1(n1486), .IN2(g1531), .QN(n3988) );
  NAND4X0 U4510 ( .IN1(n4002), .IN2(n4003), .IN3(n4004), .IN4(n4005), .QN(
        n3986) );
  NOR2X0 U4511 ( .IN1(n4006), .IN2(n4007), .QN(n4005) );
  NOR2X0 U4512 ( .IN1(n1720), .IN2(n3871), .QN(n4007) );
  NOR2X0 U4513 ( .IN1(n2233), .IN2(n3916), .QN(n4006) );
  OR2X1 U4514 ( .IN1(n3921), .IN2(n1630), .Q(n4004) );
  NAND2X0 U4515 ( .IN1(n3919), .IN2(g1), .QN(n4003) );
  NAND2X0 U4516 ( .IN1(g892), .IN2(n3920), .QN(n4002) );
  NAND2X0 U4517 ( .IN1(n4008), .IN2(n4009), .QN(n3985) );
  NAND2X0 U4518 ( .IN1(n3880), .IN2(g1346), .QN(n4009) );
  NAND2X0 U4519 ( .IN1(g1176), .IN2(n3875), .QN(n4008) );
  NAND3X0 U4520 ( .IN1(n4010), .IN2(n4011), .IN3(n4012), .QN(n3984) );
  NAND2X0 U4521 ( .IN1(n3884), .IN2(g1727), .QN(n4012) );
  NAND2X0 U4522 ( .IN1(n3925), .IN2(g1321), .QN(n4011) );
  NAND2X0 U4523 ( .IN1(g904), .IN2(n3885), .QN(n4010) );
  NAND2X0 U4524 ( .IN1(n2359), .IN2(n3797), .QN(g10457) );
  NOR4X0 U4525 ( .IN1(n4013), .IN2(n4014), .IN3(n4015), .IN4(n4016), .QN(n3797) );
  NAND4X0 U4526 ( .IN1(n4017), .IN2(n4018), .IN3(n4019), .IN4(n4020), .QN(
        n4016) );
  NOR4X0 U4527 ( .IN1(n4021), .IN2(n4022), .IN3(n4023), .IN4(n4024), .QN(n4020) );
  NOR2X0 U4528 ( .IN1(n2232), .IN2(n3916), .QN(n4024) );
  NOR2X0 U4529 ( .IN1(n1591), .IN2(n3921), .QN(n4023) );
  NOR2X0 U4530 ( .IN1(n2314), .IN2(n3871), .QN(n4022) );
  NAND3X0 U4531 ( .IN1(n4025), .IN2(n4026), .IN3(n4027), .QN(n4021) );
  NAND2X0 U4532 ( .IN1(g889), .IN2(n3920), .QN(n4027) );
  NAND2X0 U4533 ( .IN1(n1486), .IN2(g1528), .QN(n4026) );
  NAND2X0 U4534 ( .IN1(n3919), .IN2(g4), .QN(n4025) );
  AND3X1 U4535 ( .IN1(n4028), .IN2(n4029), .IN3(n4030), .Q(n4019) );
  NAND2X0 U4536 ( .IN1(n3884), .IN2(g1724), .QN(n4030) );
  NAND2X0 U4537 ( .IN1(n3925), .IN2(g1318), .QN(n4029) );
  NAND2X0 U4538 ( .IN1(g901), .IN2(n3885), .QN(n4028) );
  NAND2X0 U4539 ( .IN1(n3880), .IN2(g1341), .QN(n4018) );
  NAND2X0 U4540 ( .IN1(g1173), .IN2(n3875), .QN(n4017) );
  NAND4X0 U4541 ( .IN1(n4031), .IN2(n4032), .IN3(n4033), .IN4(n4034), .QN(
        n4015) );
  NOR2X0 U4542 ( .IN1(n4035), .IN2(n4036), .QN(n4034) );
  NOR2X0 U4543 ( .IN1(n2154), .IN2(n3932), .QN(n4036) );
  NOR2X0 U4544 ( .IN1(n2143), .IN2(n4037), .QN(n4035) );
  NAND2X0 U4545 ( .IN1(n1530), .IN2(g925), .QN(n4033) );
  NAND2X0 U4546 ( .IN1(n3936), .IN2(g953), .QN(n4032) );
  NAND2X0 U4547 ( .IN1(g1197), .IN2(n1512), .QN(n4031) );
  NAND3X0 U4548 ( .IN1(n4038), .IN2(n4039), .IN3(n4040), .QN(n4014) );
  NAND2X0 U4549 ( .IN1(n3806), .IN2(n3031), .QN(n4040) );
  NAND2X0 U4550 ( .IN1(n3937), .IN2(g1747), .QN(n4039) );
  NAND2X0 U4551 ( .IN1(n382), .IN2(g1595), .QN(n4038) );
  NAND3X0 U4552 ( .IN1(n4041), .IN2(n3939), .IN3(n4042), .QN(n4013) );
  NAND2X0 U4553 ( .IN1(n3941), .IN2(g290), .QN(n4042) );
  NAND2X0 U4554 ( .IN1(n3942), .IN2(g266), .QN(n4041) );
  NAND2X0 U4555 ( .IN1(n2359), .IN2(n3677), .QN(g10455) );
  NOR4X0 U4556 ( .IN1(n4043), .IN2(n4044), .IN3(n4045), .IN4(n4046), .QN(n3677) );
  NAND4X0 U4557 ( .IN1(n4047), .IN2(n4048), .IN3(n4049), .IN4(n4050), .QN(
        n4046) );
  NOR4X0 U4558 ( .IN1(n4051), .IN2(n4052), .IN3(n4053), .IN4(n4054), .QN(n4050) );
  NOR2X0 U4559 ( .IN1(n1613), .IN2(n3916), .QN(n4054) );
  NOR2X0 U4560 ( .IN1(n1604), .IN2(n3921), .QN(n4053) );
  NOR2X0 U4561 ( .IN1(n2315), .IN2(n3871), .QN(n4052) );
  NAND3X0 U4562 ( .IN1(n4055), .IN2(n4056), .IN3(n4057), .QN(n4051) );
  NAND2X0 U4563 ( .IN1(g886), .IN2(n3920), .QN(n4057) );
  INVX0 U4564 ( .INP(n4058), .ZN(n3920) );
  NAND2X0 U4565 ( .IN1(n1486), .IN2(g1524), .QN(n4056) );
  NAND2X0 U4566 ( .IN1(n3919), .IN2(g123), .QN(n4055) );
  INVX0 U4567 ( .INP(n3978), .ZN(n3919) );
  AND3X1 U4568 ( .IN1(n4059), .IN2(n4060), .IN3(n4061), .Q(n4049) );
  NAND2X0 U4569 ( .IN1(n3884), .IN2(g1721), .QN(n4061) );
  NAND2X0 U4570 ( .IN1(n3925), .IN2(g1314), .QN(n4060) );
  NAND2X0 U4571 ( .IN1(g898), .IN2(n3885), .QN(n4059) );
  NAND2X0 U4572 ( .IN1(n3880), .IN2(g1336), .QN(n4048) );
  NAND2X0 U4573 ( .IN1(g1170), .IN2(n3875), .QN(n4047) );
  NAND4X0 U4574 ( .IN1(n4062), .IN2(n4063), .IN3(n4064), .IN4(n4065), .QN(
        n4045) );
  AND3X1 U4575 ( .IN1(n4066), .IN2(n4067), .IN3(n4068), .Q(n4065) );
  NAND2X0 U4576 ( .IN1(n1485), .IN2(g1567), .QN(n4068) );
  NAND2X0 U4577 ( .IN1(g922), .IN2(n1530), .QN(n4067) );
  NAND2X0 U4578 ( .IN1(n1479), .IN2(g1549), .QN(n4066) );
  NAND2X0 U4579 ( .IN1(g1194), .IN2(n1512), .QN(n4064) );
  NAND2X0 U4580 ( .IN1(n3806), .IN2(n3051), .QN(n4063) );
  NAND2X0 U4581 ( .IN1(n3936), .IN2(g950), .QN(n4062) );
  NAND3X0 U4582 ( .IN1(n4069), .IN2(n4070), .IN3(n4071), .QN(n4044) );
  NAND2X0 U4583 ( .IN1(n3937), .IN2(g1744), .QN(n4071) );
  NAND2X0 U4584 ( .IN1(n3942), .IN2(g263), .QN(n4070) );
  NAND2X0 U4585 ( .IN1(n3941), .IN2(g287), .QN(n4069) );
  INVX0 U4586 ( .INP(n4072), .ZN(n3941) );
  NAND3X0 U4587 ( .IN1(n3939), .IN2(n2553), .IN3(n4073), .QN(n4043) );
  NAND2X0 U4588 ( .IN1(n382), .IN2(g1592), .QN(n4073) );
  INVX0 U4589 ( .INP(n3995), .ZN(n382) );
  NAND4X0 U4590 ( .IN1(n3977), .IN2(n3978), .IN3(n3882), .IN4(n4074), .QN(
        n3939) );
  INVX0 U4591 ( .INP(n1512), .ZN(n4074) );
  NAND2X0 U4592 ( .IN1(n4075), .IN2(g42), .QN(n3978) );
  AND4X1 U4593 ( .IN1(n1546), .IN2(n3954), .IN3(n3916), .IN4(n2553), .Q(n3977)
         );
  NAND2X0 U4594 ( .IN1(n4075), .IN2(n2561), .QN(n3916) );
  AND4X1 U4595 ( .IN1(n1548), .IN2(g43), .IN3(n3757), .IN4(n4076), .Q(n4075)
         );
  AND4X1 U4596 ( .IN1(n4058), .IN2(n3921), .IN3(n4077), .IN4(n4078), .Q(n1546)
         );
  NOR4X0 U4597 ( .IN1(n4079), .IN2(n4080), .IN3(n3936), .IN4(n3806), .QN(n4078) );
  INVX0 U4598 ( .INP(n1472), .ZN(n3936) );
  NAND2X0 U4599 ( .IN1(n4081), .IN2(n1574), .QN(n1472) );
  NOR2X0 U4600 ( .IN1(n1530), .IN2(n3885), .QN(n4077) );
  NAND4X0 U4601 ( .IN1(n1574), .IN2(g45), .IN3(n4082), .IN4(g44), .QN(n3921)
         );
  NOR2X0 U4602 ( .IN1(g43), .IN2(n2561), .QN(n4082) );
  NAND4X0 U4603 ( .IN1(n1574), .IN2(n4083), .IN3(g43), .IN4(g42), .QN(n4058)
         );
  NAND2X0 U4604 ( .IN1(n2359), .IN2(n3754), .QN(g10377) );
  NOR3X0 U4605 ( .IN1(n4084), .IN2(n4085), .IN3(n4086), .QN(n3754) );
  NAND4X0 U4606 ( .IN1(n4087), .IN2(n4088), .IN3(n2553), .IN4(n4089), .QN(
        n4086) );
  NOR4X0 U4607 ( .IN1(n1564), .IN2(n4090), .IN3(n4091), .IN4(n4092), .QN(n4089) );
  AND2X1 U4608 ( .IN1(g1188), .IN2(n3875), .Q(n4092) );
  NOR2X0 U4609 ( .IN1(n2141), .IN2(n3932), .QN(n4091) );
  INVX0 U4610 ( .INP(n1485), .ZN(n3932) );
  NOR2X0 U4611 ( .IN1(n4116), .IN2(n3872), .QN(n4090) );
  INVX0 U4612 ( .INP(n3806), .ZN(n3872) );
  NAND4X0 U4613 ( .IN1(g46), .IN2(g47), .IN3(n4093), .IN4(n4094), .QN(n2553)
         );
  INVX0 U4614 ( .INP(n1545), .ZN(n4094) );
  NAND4X0 U4615 ( .IN1(g44), .IN2(g43), .IN3(n2561), .IN4(n4076), .QN(n1545)
         );
  NAND2X0 U4616 ( .IN1(n3942), .IN2(g281), .QN(n4088) );
  INVX0 U4617 ( .INP(n3876), .ZN(n3942) );
  NAND2X0 U4618 ( .IN1(n4079), .IN2(n4072), .QN(n3876) );
  NAND2X0 U4619 ( .IN1(n4079), .IN2(n2561), .QN(n4072) );
  AND4X1 U4620 ( .IN1(n1548), .IN2(g44), .IN3(n3755), .IN4(n4076), .Q(n4079)
         );
  NAND2X0 U4621 ( .IN1(n3937), .IN2(g1762), .QN(n4087) );
  INVX0 U4622 ( .INP(n4095), .ZN(n3937) );
  NAND4X0 U4623 ( .IN1(n4096), .IN2(n4097), .IN3(n4098), .IN4(n4099), .QN(
        n4085) );
  NAND2X0 U4624 ( .IN1(n3880), .IN2(g1308), .QN(n4099) );
  INVX0 U4625 ( .INP(n3882), .ZN(n3880) );
  NAND3X0 U4626 ( .IN1(n1478), .IN2(n3954), .IN3(n3882), .QN(n4098) );
  NAND2X0 U4627 ( .IN1(n4100), .IN2(n1544), .QN(n3882) );
  AND4X1 U4628 ( .IN1(n3881), .IN2(n4101), .IN3(n3883), .IN4(n4095), .Q(n3954)
         );
  NAND2X0 U4629 ( .IN1(n4102), .IN2(n2561), .QN(n4095) );
  NOR3X0 U4630 ( .IN1(n1566), .IN2(n1567), .IN3(n3875), .QN(n3881) );
  AND2X1 U4631 ( .IN1(n1544), .IN2(n4103), .Q(n3875) );
  NAND2X0 U4632 ( .IN1(n3995), .IN2(n4104), .QN(n1567) );
  NAND2X0 U4633 ( .IN1(n4100), .IN2(n1548), .QN(n4104) );
  NAND2X0 U4634 ( .IN1(n4081), .IN2(n1548), .QN(n3995) );
  NAND2X0 U4635 ( .IN1(n4037), .IN2(n4105), .QN(n1566) );
  NAND2X0 U4636 ( .IN1(n1548), .IN2(n4103), .QN(n4105) );
  AND3X1 U4637 ( .IN1(n2565), .IN2(n2562), .IN3(n4093), .Q(n1548) );
  INVX0 U4638 ( .INP(n1479), .ZN(n4037) );
  NAND2X0 U4639 ( .IN1(n3884), .IN2(g1738), .QN(n4097) );
  INVX0 U4640 ( .INP(n3883), .ZN(n3884) );
  NAND2X0 U4641 ( .IN1(n4102), .IN2(g42), .QN(n3883) );
  AND4X1 U4642 ( .IN1(g45), .IN2(n1544), .IN3(g44), .IN4(g43), .Q(n4102) );
  NAND2X0 U4643 ( .IN1(n1486), .IN2(g1543), .QN(n4096) );
  NAND3X0 U4644 ( .IN1(n4106), .IN2(n4107), .IN3(n4108), .QN(n4084) );
  NAND2X0 U4645 ( .IN1(g916), .IN2(n3885), .QN(n4108) );
  AND2X1 U4646 ( .IN1(n1574), .IN2(n4103), .Q(n3885) );
  NOR4X0 U4647 ( .IN1(n3757), .IN2(n3755), .IN3(n2561), .IN4(g45), .QN(n4103)
         );
  INVX0 U4648 ( .INP(g44), .ZN(n3757) );
  NAND2X0 U4649 ( .IN1(n4080), .IN2(g944), .QN(n4107) );
  INVX0 U4650 ( .INP(n3871), .ZN(n4080) );
  NAND2X0 U4651 ( .IN1(n1574), .IN2(n4100), .QN(n3871) );
  AND3X1 U4652 ( .IN1(g42), .IN2(n3755), .IN3(n4083), .Q(n4100) );
  AND3X1 U4653 ( .IN1(n4093), .IN2(n2562), .IN3(g46), .Q(n1574) );
  INVX0 U4654 ( .INP(g47), .ZN(n2562) );
  NAND2X0 U4655 ( .IN1(n3925), .IN2(g1333), .QN(n4106) );
  INVX0 U4656 ( .INP(n4101), .ZN(n3925) );
  NAND2X0 U4657 ( .IN1(n4081), .IN2(n1544), .QN(n4101) );
  AND3X1 U4658 ( .IN1(n4093), .IN2(n2565), .IN3(g47), .Q(n1544) );
  INVX0 U4659 ( .INP(g46), .ZN(n2565) );
  AND2X1 U4660 ( .IN1(n2583), .IN2(g48), .Q(n4093) );
  NOR3X0 U4661 ( .IN1(n4109), .IN2(n4110), .IN3(g41), .QN(n2583) );
  AND2X1 U4662 ( .IN1(n3806), .IN2(g48), .Q(n4110) );
  NOR2X0 U4663 ( .IN1(g48), .IN2(n2581), .QN(n4109) );
  INVX0 U4664 ( .INP(g30), .ZN(n2581) );
  AND3X1 U4665 ( .IN1(n2561), .IN2(n3755), .IN3(n4083), .Q(n4081) );
  NOR2X0 U4666 ( .IN1(n4076), .IN2(g44), .QN(n4083) );
  INVX0 U4667 ( .INP(g45), .ZN(n4076) );
  INVX0 U4668 ( .INP(g43), .ZN(n3755) );
  INVX0 U4669 ( .INP(g42), .ZN(n2561) );
  NOR2X0 U4670 ( .IN1(n3806), .IN2(g30), .QN(n2359) );
  NAND2X0 U4671 ( .IN1(g48), .IN2(n2582), .QN(n3806) );
  INVX0 U4672 ( .INP(g31), .ZN(n2582) );
  XOR2X1 U4673 ( .IN1(test_so1), .IN2(n2941), .Q(N599) );
  NOR3X0 U4674 ( .IN1(n2129), .IN2(n2134), .IN3(n2944), .QN(n2941) );
  INVX0 U4675 ( .INP(n1093), .ZN(n2944) );
  OR2X1 U1550_U1 ( .IN1(n25), .IN2(n2359), .Q(g10461) );
  OR2X1 U1551_U1 ( .IN1(n114), .IN2(n2359), .Q(g10379) );
  INVX0 U1586_U2 ( .INP(n11), .ZN(U1586_n1) );
  NOR2X0 U1586_U1 ( .IN1(n2353), .IN2(U1586_n1), .QN(n1855) );
  INVX0 U1754_U2 ( .INP(n1548), .ZN(U1754_n1) );
  NOR2X0 U1754_U1 ( .IN1(n1545), .IN2(U1754_n1), .QN(n1479) );
  INVX0 U1798_U2 ( .INP(n1567), .ZN(U1798_n1) );
  NOR2X0 U1798_U1 ( .IN1(n382), .IN2(U1798_n1), .QN(n1485) );
  INVX0 U1839_U2 ( .INP(n1566), .ZN(U1839_n1) );
  NOR2X0 U1839_U1 ( .IN1(n1479), .IN2(U1839_n1), .QN(n1486) );
  INVX0 U1843_U2 ( .INP(n1546), .ZN(U1843_n1) );
  NOR2X0 U1843_U1 ( .IN1(n387), .IN2(U1843_n1), .QN(n1478) );
  INVX0 U1877_U2 ( .INP(n1137), .ZN(U1877_n1) );
  NOR2X0 U1877_U1 ( .IN1(n2365), .IN2(U1877_n1), .QN(n1195) );
  INVX0 U1908_U2 ( .INP(n1544), .ZN(U1908_n1) );
  NOR2X0 U1908_U1 ( .IN1(n1545), .IN2(U1908_n1), .QN(n1512) );
  INVX0 U1909_U2 ( .INP(n1574), .ZN(U1909_n1) );
  NOR2X0 U1909_U1 ( .IN1(n1545), .IN2(U1909_n1), .QN(n1530) );
  INVX0 U1987_U2 ( .INP(n822), .ZN(U1987_n1) );
  NOR2X0 U1987_U1 ( .IN1(n177), .IN2(U1987_n1), .QN(n916) );
  INVX0 U2031_U2 ( .INP(n1057), .ZN(U2031_n1) );
  NOR2X0 U2031_U1 ( .IN1(n1054), .IN2(U2031_n1), .QN(n1056) );
  INVX0 U2035_U2 ( .INP(n1404), .ZN(U2035_n1) );
  NOR2X0 U2035_U1 ( .IN1(g109), .IN2(U2035_n1), .QN(n1450) );
  INVX0 U2418_U2 ( .INP(g968), .ZN(U2418_n1) );
  NOR2X0 U2418_U1 ( .IN1(n1472), .IN2(U2418_n1), .QN(n1564) );
  INVX0 U2468_U2 ( .INP(g1336), .ZN(U2468_n1) );
  NOR2X0 U2468_U1 ( .IN1(n1227), .IN2(U2468_n1), .QN(n1231) );
  INVX0 U2478_U2 ( .INP(g1341), .ZN(U2478_n1) );
  NOR2X0 U2478_U1 ( .IN1(n1229), .IN2(U2478_n1), .QN(n1232) );
  INVX0 U2488_U2 ( .INP(n1262), .ZN(U2488_n1) );
  NOR2X0 U2488_U1 ( .IN1(n22), .IN2(U2488_n1), .QN(n1260) );
  INVX0 U2533_U2 ( .INP(g178), .ZN(U2533_n1) );
  NOR2X0 U2533_U1 ( .IN1(n2363), .IN2(U2533_n1), .QN(g6786) );
  INVX0 U2534_U2 ( .INP(g1424), .ZN(U2534_n1) );
  NOR2X0 U2534_U1 ( .IN1(n2364), .IN2(U2534_n1), .QN(g6234) );
  INVX0 U2639_U2 ( .INP(n962), .ZN(U2639_n1) );
  NOR2X0 U2639_U1 ( .IN1(n958), .IN2(U2639_n1), .QN(n804) );
  INVX0 U2641_U2 ( .INP(n39), .ZN(U2641_n1) );
  NOR2X0 U2641_U1 ( .IN1(g1868), .IN2(U2641_n1), .QN(n926) );
  INVX0 U2654_U2 ( .INP(g746), .ZN(U2654_n1) );
  NOR2X0 U2654_U1 ( .IN1(g750), .IN2(U2654_n1), .QN(g4171) );
  INVX0 U2658_U2 ( .INP(n917), .ZN(U2658_n1) );
  NOR2X0 U2658_U1 ( .IN1(n918), .IN2(U2658_n1), .QN(n812) );
  INVX0 U2683_U2 ( .INP(g382), .ZN(U2683_n1) );
  NOR2X0 U2683_U1 ( .IN1(n40), .IN2(U2683_n1), .QN(n1420) );
  INVX0 U2699_U2 ( .INP(n808), .ZN(U2699_n1) );
  NOR2X0 U2699_U1 ( .IN1(n367), .IN2(U2699_n1), .QN(n806) );
  INVX0 U2846_U2 ( .INP(g4175), .ZN(U2846_n1) );
  NOR2X0 U2846_U1 ( .IN1(n1214), .IN2(U2846_n1), .QN(n1193) );
  INVX0 U2847_U2 ( .INP(g4177), .ZN(U2847_n1) );
  NOR2X0 U2847_U1 ( .IN1(n1153), .IN2(U2847_n1), .QN(n1125) );
  INVX0 U2848_U2 ( .INP(g4179), .ZN(U2848_n1) );
  NOR2X0 U2848_U1 ( .IN1(n1099), .IN2(U2848_n1), .QN(n1093) );
  INVX0 U2859_U2 ( .INP(n1137), .ZN(U2859_n1) );
  NOR2X0 U2859_U1 ( .IN1(g12), .IN2(U2859_n1), .QN(n1159) );
  INVX0 U2860_U2 ( .INP(g810), .ZN(U2860_n1) );
  NOR2X0 U2860_U1 ( .IN1(n1151), .IN2(U2860_n1), .QN(n1123) );
  INVX0 U2861_U2 ( .INP(g818), .ZN(U2861_n1) );
  NOR2X0 U2861_U1 ( .IN1(n1097), .IN2(U2861_n1), .QN(n1090) );
  INVX0 U2867_U2 ( .INP(n817), .ZN(U2867_n1) );
  NOR2X0 U2867_U1 ( .IN1(g1834), .IN2(U2867_n1), .QN(n1380) );
  INVX0 U2879_U2 ( .INP(g713), .ZN(U2879_n1) );
  NOR2X0 U2879_U1 ( .IN1(n1656), .IN2(U2879_n1), .QN(n967) );
  INVX0 U2881_U2 ( .INP(g1927), .ZN(U2881_n1) );
  NOR2X0 U2881_U1 ( .IN1(n1657), .IN2(U2881_n1), .QN(n921) );
  INVX0 U2882_U2 ( .INP(g1160), .ZN(U2882_n1) );
  NOR2X0 U2882_U1 ( .IN1(n2362), .IN2(U2882_n1), .QN(g4334) );
  INVX0 U2883_U2 ( .INP(g1166), .ZN(U2883_n1) );
  NOR2X0 U2883_U1 ( .IN1(n2365), .IN2(U2883_n1), .QN(g4325) );
  INVX0 U2884_U2 ( .INP(g148), .ZN(U2884_n1) );
  NOR2X0 U2884_U1 ( .IN1(n2363), .IN2(U2884_n1), .QN(g6759) );
  INVX0 U2885_U2 ( .INP(g1157), .ZN(U2885_n1) );
  NOR2X0 U2885_U1 ( .IN1(n2364), .IN2(U2885_n1), .QN(g4338) );
  INVX0 U2886_U2 ( .INP(g1163), .ZN(U2886_n1) );
  NOR2X0 U2886_U1 ( .IN1(n2362), .IN2(U2886_n1), .QN(g4330) );
  INVX0 U2887_U2 ( .INP(g237), .ZN(U2887_n1) );
  NOR2X0 U2887_U1 ( .IN1(n2365), .IN2(U2887_n1), .QN(g6821) );
  INVX0 U2888_U2 ( .INP(g1499), .ZN(U2888_n1) );
  NOR2X0 U2888_U1 ( .IN1(n2363), .IN2(U2888_n1), .QN(g6198) );
  INVX0 U2889_U2 ( .INP(g1411), .ZN(U2889_n1) );
  NOR2X0 U2889_U1 ( .IN1(n2364), .IN2(U2889_n1), .QN(g6244) );
  INVX0 U2890_U2 ( .INP(g225), .ZN(U2890_n1) );
  NOR2X0 U2890_U1 ( .IN1(n2362), .IN2(U2890_n1), .QN(g6826) );
  INVX0 U2891_U2 ( .INP(g1407), .ZN(U2891_n1) );
  NOR2X0 U2891_U1 ( .IN1(n2365), .IN2(U2891_n1), .QN(g6216) );
  INVX0 U2892_U2 ( .INP(g213), .ZN(U2892_n1) );
  NOR2X0 U2892_U1 ( .IN1(n2363), .IN2(U2892_n1), .QN(g6829) );
  INVX0 U2893_U2 ( .INP(g186), .ZN(U2893_n1) );
  NOR2X0 U2893_U1 ( .IN1(n2364), .IN2(U2893_n1), .QN(g6833) );
  INVX0 U2894_U2 ( .INP(g219), .ZN(U2894_n1) );
  NOR2X0 U2894_U1 ( .IN1(n2362), .IN2(U2894_n1), .QN(g6827) );
  INVX0 U2895_U2 ( .INP(g143), .ZN(U2895_n1) );
  NOR2X0 U2895_U1 ( .IN1(n2365), .IN2(U2895_n1), .QN(g6757) );
  INVX0 U2896_U2 ( .INP(g207), .ZN(U2896_n1) );
  NOR2X0 U2896_U1 ( .IN1(n2363), .IN2(U2896_n1), .QN(g6831) );
  INVX0 U2897_U2 ( .INP(g231), .ZN(U2897_n1) );
  NOR2X0 U2897_U1 ( .IN1(n2364), .IN2(U2897_n1), .QN(g6822) );
  INVX0 U2898_U2 ( .INP(g192), .ZN(U2898_n1) );
  NOR2X0 U2898_U1 ( .IN1(n2362), .IN2(U2898_n1), .QN(g6838) );
  INVX0 U2899_U2 ( .INP(test_so3), .ZN(U2899_n1) );
  NOR2X0 U2899_U1 ( .IN1(n2365), .IN2(U2899_n1), .QN(g6823) );
  INVX0 U2900_U2 ( .INP(g1371), .ZN(U2900_n1) );
  NOR2X0 U2900_U1 ( .IN1(n2363), .IN2(U2900_n1), .QN(g6824) );
  INVX0 U2901_U2 ( .INP(g1383), .ZN(U2901_n1) );
  NOR2X0 U2901_U1 ( .IN1(n2364), .IN2(U2901_n1), .QN(g6832) );
  INVX0 U2902_U2 ( .INP(g243), .ZN(U2902_n1) );
  NOR2X0 U2902_U1 ( .IN1(n2362), .IN2(U2902_n1), .QN(g6819) );
  INVX0 U3090_U2 ( .INP(n1151), .ZN(U3090_n1) );
  NOR2X0 U3090_U1 ( .IN1(g810), .IN2(U3090_n1), .QN(n1150) );
  INVX0 U3092_U2 ( .INP(n1097), .ZN(U3092_n1) );
  NOR2X0 U3092_U1 ( .IN1(g818), .IN2(U3092_n1), .QN(n1096) );
  INVX0 U3094_U2 ( .INP(n1099), .ZN(U3094_n1) );
  NOR2X0 U3094_U1 ( .IN1(g4179), .IN2(U3094_n1), .QN(n1098) );
  INVX0 U3096_U2 ( .INP(n1214), .ZN(U3096_n1) );
  NOR2X0 U3096_U1 ( .IN1(g4175), .IN2(U3096_n1), .QN(n1213) );
  INVX0 U3098_U2 ( .INP(n1153), .ZN(U3098_n1) );
  NOR2X0 U3098_U1 ( .IN1(g4177), .IN2(U3098_n1), .QN(n1152) );
  INVX0 U3124_U2 ( .INP(n837), .ZN(U3124_n1) );
  NOR2X0 U3124_U1 ( .IN1(n838), .IN2(U3124_n1), .QN(n836) );
  INVX0 U3171_U2 ( .INP(g1610), .ZN(U3171_n1) );
  NOR2X0 U3171_U1 ( .IN1(n263), .IN2(U3171_n1), .QN(g5194) );
endmodule

