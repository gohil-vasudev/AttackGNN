module add_mul_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, 
        b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation, Result_0_, 
        Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, 
        Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, 
        Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951;

  OR2_X1 U482 ( .A1(n466), .A2(n467), .ZN(Result_9_) );
  AND2_X1 U483 ( .A1(n468), .A2(operation), .ZN(n467) );
  XNOR2_X1 U484 ( .A(n469), .B(n470), .ZN(n468) );
  XOR2_X1 U485 ( .A(n471), .B(n472), .Z(n470) );
  AND2_X1 U486 ( .A1(n473), .A2(n474), .ZN(n466) );
  OR2_X1 U487 ( .A1(n475), .A2(n476), .ZN(n473) );
  OR2_X1 U488 ( .A1(n477), .A2(n478), .ZN(n476) );
  AND2_X1 U489 ( .A1(n479), .A2(n480), .ZN(n478) );
  XNOR2_X1 U490 ( .A(n481), .B(n482), .ZN(n479) );
  AND2_X1 U491 ( .A1(n483), .A2(b_1_), .ZN(n477) );
  AND2_X1 U492 ( .A1(n484), .A2(n481), .ZN(n483) );
  AND2_X1 U493 ( .A1(n485), .A2(n482), .ZN(n475) );
  OR2_X1 U494 ( .A1(n486), .A2(n487), .ZN(Result_8_) );
  AND2_X1 U495 ( .A1(n488), .A2(operation), .ZN(n487) );
  XNOR2_X1 U496 ( .A(n489), .B(n490), .ZN(n488) );
  XOR2_X1 U497 ( .A(n491), .B(n492), .Z(n490) );
  AND2_X1 U498 ( .A1(n493), .A2(n474), .ZN(n486) );
  XOR2_X1 U499 ( .A(n494), .B(n495), .Z(n493) );
  XNOR2_X1 U500 ( .A(n496), .B(a_0_), .ZN(n495) );
  AND2_X1 U501 ( .A1(n497), .A2(n498), .ZN(n494) );
  OR2_X1 U502 ( .A1(n485), .A2(n482), .ZN(n498) );
  INV_X1 U503 ( .A(n484), .ZN(n482) );
  OR2_X1 U504 ( .A1(n499), .A2(n500), .ZN(n484) );
  INV_X1 U505 ( .A(n501), .ZN(n500) );
  AND2_X1 U506 ( .A1(n502), .A2(n503), .ZN(n499) );
  OR2_X1 U507 ( .A1(b_1_), .A2(a_1_), .ZN(n497) );
  AND2_X1 U508 ( .A1(operation), .A2(n504), .ZN(Result_7_) );
  XOR2_X1 U509 ( .A(n505), .B(n506), .Z(n504) );
  AND2_X1 U510 ( .A1(n507), .A2(operation), .ZN(Result_6_) );
  AND2_X1 U511 ( .A1(n508), .A2(n509), .ZN(n507) );
  OR2_X1 U512 ( .A1(n510), .A2(n511), .ZN(n508) );
  XOR2_X1 U513 ( .A(n512), .B(n513), .Z(n511) );
  INV_X1 U514 ( .A(n514), .ZN(n510) );
  AND2_X1 U515 ( .A1(operation), .A2(n515), .ZN(Result_5_) );
  XOR2_X1 U516 ( .A(n516), .B(n517), .Z(n515) );
  OR2_X1 U517 ( .A1(n518), .A2(n519), .ZN(n516) );
  AND2_X1 U518 ( .A1(n520), .A2(operation), .ZN(Result_4_) );
  XOR2_X1 U519 ( .A(n521), .B(n522), .Z(n520) );
  AND2_X1 U520 ( .A1(operation), .A2(n523), .ZN(Result_3_) );
  XOR2_X1 U521 ( .A(n524), .B(n525), .Z(n523) );
  AND2_X1 U522 ( .A1(n526), .A2(n527), .ZN(n525) );
  OR2_X1 U523 ( .A1(n528), .A2(n529), .ZN(n527) );
  INV_X1 U524 ( .A(n530), .ZN(n526) );
  AND2_X1 U525 ( .A1(n531), .A2(operation), .ZN(Result_2_) );
  XOR2_X1 U526 ( .A(n532), .B(n533), .Z(n531) );
  AND2_X1 U527 ( .A1(operation), .A2(n534), .ZN(Result_1_) );
  XOR2_X1 U528 ( .A(n535), .B(n536), .Z(n534) );
  AND2_X1 U529 ( .A1(n537), .A2(n538), .ZN(n536) );
  OR2_X1 U530 ( .A1(n539), .A2(n540), .ZN(n538) );
  AND2_X1 U531 ( .A1(n541), .A2(n542), .ZN(n539) );
  INV_X1 U532 ( .A(n543), .ZN(n537) );
  OR2_X1 U533 ( .A1(n544), .A2(n545), .ZN(Result_15_) );
  AND2_X1 U534 ( .A1(n546), .A2(operation), .ZN(n545) );
  AND2_X1 U535 ( .A1(n547), .A2(n474), .ZN(n544) );
  XNOR2_X1 U536 ( .A(n548), .B(a_7_), .ZN(n547) );
  OR2_X1 U537 ( .A1(n549), .A2(n550), .ZN(Result_14_) );
  AND2_X1 U538 ( .A1(n551), .A2(operation), .ZN(n550) );
  XNOR2_X1 U539 ( .A(n552), .B(n553), .ZN(n551) );
  AND2_X1 U540 ( .A1(b_7_), .A2(a_6_), .ZN(n553) );
  AND2_X1 U541 ( .A1(n554), .A2(n474), .ZN(n549) );
  XOR2_X1 U542 ( .A(n546), .B(n555), .Z(n554) );
  XNOR2_X1 U543 ( .A(n556), .B(a_6_), .ZN(n555) );
  OR2_X1 U544 ( .A1(n557), .A2(n558), .ZN(Result_13_) );
  AND2_X1 U545 ( .A1(n559), .A2(operation), .ZN(n558) );
  XOR2_X1 U546 ( .A(n560), .B(n561), .Z(n559) );
  XNOR2_X1 U547 ( .A(n562), .B(n563), .ZN(n561) );
  AND2_X1 U548 ( .A1(n564), .A2(n474), .ZN(n557) );
  OR2_X1 U549 ( .A1(n565), .A2(n566), .ZN(n564) );
  AND2_X1 U550 ( .A1(n567), .A2(n568), .ZN(n566) );
  XNOR2_X1 U551 ( .A(n569), .B(a_5_), .ZN(n567) );
  AND2_X1 U552 ( .A1(n570), .A2(n571), .ZN(n565) );
  INV_X1 U553 ( .A(n568), .ZN(n571) );
  OR2_X1 U554 ( .A1(n572), .A2(n573), .ZN(n570) );
  OR2_X1 U555 ( .A1(n574), .A2(n575), .ZN(Result_12_) );
  AND2_X1 U556 ( .A1(n576), .A2(operation), .ZN(n575) );
  XNOR2_X1 U557 ( .A(n577), .B(n578), .ZN(n576) );
  XOR2_X1 U558 ( .A(n579), .B(n580), .Z(n578) );
  AND2_X1 U559 ( .A1(n581), .A2(n474), .ZN(n574) );
  XNOR2_X1 U560 ( .A(n582), .B(n583), .ZN(n581) );
  AND2_X1 U561 ( .A1(n584), .A2(n585), .ZN(n583) );
  OR2_X1 U562 ( .A1(n586), .A2(n587), .ZN(Result_11_) );
  AND2_X1 U563 ( .A1(n588), .A2(operation), .ZN(n587) );
  XNOR2_X1 U564 ( .A(n589), .B(n590), .ZN(n588) );
  XOR2_X1 U565 ( .A(n591), .B(n592), .Z(n590) );
  AND2_X1 U566 ( .A1(n593), .A2(n474), .ZN(n586) );
  OR2_X1 U567 ( .A1(n594), .A2(n595), .ZN(n593) );
  OR2_X1 U568 ( .A1(n596), .A2(n597), .ZN(n595) );
  AND2_X1 U569 ( .A1(n598), .A2(n599), .ZN(n597) );
  XNOR2_X1 U570 ( .A(n600), .B(n601), .ZN(n598) );
  AND2_X1 U571 ( .A1(n602), .A2(b_3_), .ZN(n596) );
  AND2_X1 U572 ( .A1(n603), .A2(n600), .ZN(n602) );
  AND2_X1 U573 ( .A1(n601), .A2(n604), .ZN(n594) );
  OR2_X1 U574 ( .A1(n605), .A2(n606), .ZN(Result_10_) );
  AND2_X1 U575 ( .A1(n607), .A2(operation), .ZN(n606) );
  XNOR2_X1 U576 ( .A(n608), .B(n609), .ZN(n607) );
  XOR2_X1 U577 ( .A(n610), .B(n611), .Z(n609) );
  AND2_X1 U578 ( .A1(n612), .A2(n474), .ZN(n605) );
  INV_X1 U579 ( .A(operation), .ZN(n474) );
  XNOR2_X1 U580 ( .A(n502), .B(n613), .ZN(n612) );
  AND2_X1 U581 ( .A1(n503), .A2(n501), .ZN(n613) );
  OR2_X1 U582 ( .A1(a_2_), .A2(b_2_), .ZN(n501) );
  OR2_X1 U583 ( .A1(n614), .A2(n615), .ZN(n502) );
  AND2_X1 U584 ( .A1(n600), .A2(n599), .ZN(n615) );
  AND2_X1 U585 ( .A1(n603), .A2(n616), .ZN(n614) );
  INV_X1 U586 ( .A(n601), .ZN(n603) );
  AND2_X1 U587 ( .A1(n617), .A2(n585), .ZN(n601) );
  OR2_X1 U588 ( .A1(a_4_), .A2(b_4_), .ZN(n585) );
  INV_X1 U589 ( .A(n618), .ZN(n617) );
  AND2_X1 U590 ( .A1(n584), .A2(n582), .ZN(n618) );
  OR2_X1 U591 ( .A1(n572), .A2(n619), .ZN(n582) );
  AND2_X1 U592 ( .A1(n568), .A2(n620), .ZN(n619) );
  AND2_X1 U593 ( .A1(n621), .A2(n622), .ZN(n568) );
  OR2_X1 U594 ( .A1(n548), .A2(n552), .ZN(n622) );
  INV_X1 U595 ( .A(n623), .ZN(n621) );
  AND2_X1 U596 ( .A1(a_6_), .A2(n624), .ZN(n623) );
  OR2_X1 U597 ( .A1(n546), .A2(b_6_), .ZN(n624) );
  AND2_X1 U598 ( .A1(a_7_), .A2(b_7_), .ZN(n546) );
  AND2_X1 U599 ( .A1(n625), .A2(n569), .ZN(n572) );
  AND2_X1 U600 ( .A1(operation), .A2(n626), .ZN(Result_0_) );
  OR2_X1 U601 ( .A1(n627), .A2(n628), .ZN(n626) );
  OR2_X1 U602 ( .A1(n543), .A2(n629), .ZN(n628) );
  AND2_X1 U603 ( .A1(n535), .A2(n540), .ZN(n629) );
  AND2_X1 U604 ( .A1(n532), .A2(n533), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n542), .B(n630), .ZN(n533) );
  OR2_X1 U606 ( .A1(n631), .A2(n632), .ZN(n532) );
  OR2_X1 U607 ( .A1(n633), .A2(n530), .ZN(n631) );
  AND2_X1 U608 ( .A1(n528), .A2(n529), .ZN(n530) );
  AND2_X1 U609 ( .A1(n634), .A2(n635), .ZN(n529) );
  INV_X1 U610 ( .A(n636), .ZN(n634) );
  AND2_X1 U611 ( .A1(n524), .A2(n528), .ZN(n633) );
  INV_X1 U612 ( .A(n637), .ZN(n528) );
  OR2_X1 U613 ( .A1(n638), .A2(n632), .ZN(n637) );
  INV_X1 U614 ( .A(n639), .ZN(n632) );
  OR2_X1 U615 ( .A1(n640), .A2(n641), .ZN(n639) );
  AND2_X1 U616 ( .A1(n640), .A2(n641), .ZN(n638) );
  OR2_X1 U617 ( .A1(n642), .A2(n643), .ZN(n641) );
  AND2_X1 U618 ( .A1(n644), .A2(n645), .ZN(n643) );
  AND2_X1 U619 ( .A1(n646), .A2(n647), .ZN(n642) );
  OR2_X1 U620 ( .A1(n645), .A2(n644), .ZN(n647) );
  XOR2_X1 U621 ( .A(n648), .B(n649), .Z(n640) );
  XOR2_X1 U622 ( .A(n650), .B(n651), .Z(n649) );
  AND2_X1 U623 ( .A1(n521), .A2(n522), .ZN(n524) );
  XNOR2_X1 U624 ( .A(n635), .B(n636), .ZN(n522) );
  OR2_X1 U625 ( .A1(n652), .A2(n653), .ZN(n636) );
  AND2_X1 U626 ( .A1(n654), .A2(n655), .ZN(n653) );
  AND2_X1 U627 ( .A1(n656), .A2(n657), .ZN(n652) );
  OR2_X1 U628 ( .A1(n655), .A2(n654), .ZN(n657) );
  XOR2_X1 U629 ( .A(n658), .B(n646), .Z(n635) );
  XOR2_X1 U630 ( .A(n659), .B(n660), .Z(n646) );
  XOR2_X1 U631 ( .A(n661), .B(n662), .Z(n660) );
  XNOR2_X1 U632 ( .A(n645), .B(n644), .ZN(n658) );
  OR2_X1 U633 ( .A1(n663), .A2(n664), .ZN(n644) );
  AND2_X1 U634 ( .A1(n665), .A2(n666), .ZN(n664) );
  AND2_X1 U635 ( .A1(n667), .A2(n668), .ZN(n663) );
  OR2_X1 U636 ( .A1(n666), .A2(n665), .ZN(n668) );
  OR2_X1 U637 ( .A1(n599), .A2(n669), .ZN(n645) );
  OR2_X1 U638 ( .A1(n670), .A2(n671), .ZN(n521) );
  INV_X1 U639 ( .A(n672), .ZN(n671) );
  OR2_X1 U640 ( .A1(n673), .A2(n674), .ZN(n670) );
  AND2_X1 U641 ( .A1(n518), .A2(n517), .ZN(n674) );
  AND2_X1 U642 ( .A1(n519), .A2(n517), .ZN(n673) );
  AND2_X1 U643 ( .A1(n675), .A2(n672), .ZN(n517) );
  OR2_X1 U644 ( .A1(n676), .A2(n677), .ZN(n672) );
  INV_X1 U645 ( .A(n678), .ZN(n675) );
  AND2_X1 U646 ( .A1(n676), .A2(n677), .ZN(n678) );
  OR2_X1 U647 ( .A1(n679), .A2(n680), .ZN(n677) );
  AND2_X1 U648 ( .A1(n681), .A2(n682), .ZN(n680) );
  AND2_X1 U649 ( .A1(n683), .A2(n684), .ZN(n679) );
  OR2_X1 U650 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U651 ( .A(n656), .B(n685), .Z(n676) );
  XOR2_X1 U652 ( .A(n655), .B(n654), .Z(n685) );
  OR2_X1 U653 ( .A1(n686), .A2(n669), .ZN(n654) );
  OR2_X1 U654 ( .A1(n687), .A2(n688), .ZN(n655) );
  AND2_X1 U655 ( .A1(n689), .A2(n690), .ZN(n688) );
  AND2_X1 U656 ( .A1(n691), .A2(n692), .ZN(n687) );
  OR2_X1 U657 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U658 ( .A(n693), .B(n667), .ZN(n656) );
  XNOR2_X1 U659 ( .A(n694), .B(n695), .ZN(n667) );
  XNOR2_X1 U660 ( .A(n503), .B(n696), .ZN(n694) );
  XNOR2_X1 U661 ( .A(n666), .B(n665), .ZN(n693) );
  OR2_X1 U662 ( .A1(n697), .A2(n698), .ZN(n665) );
  AND2_X1 U663 ( .A1(n699), .A2(n700), .ZN(n698) );
  AND2_X1 U664 ( .A1(n701), .A2(n702), .ZN(n697) );
  OR2_X1 U665 ( .A1(n700), .A2(n699), .ZN(n702) );
  OR2_X1 U666 ( .A1(n599), .A2(n481), .ZN(n666) );
  INV_X1 U667 ( .A(n509), .ZN(n519) );
  OR2_X1 U668 ( .A1(n703), .A2(n514), .ZN(n509) );
  OR2_X1 U669 ( .A1(n506), .A2(n505), .ZN(n514) );
  OR2_X1 U670 ( .A1(n704), .A2(n705), .ZN(n505) );
  AND2_X1 U671 ( .A1(n492), .A2(n491), .ZN(n705) );
  AND2_X1 U672 ( .A1(n489), .A2(n706), .ZN(n704) );
  OR2_X1 U673 ( .A1(n491), .A2(n492), .ZN(n706) );
  OR2_X1 U674 ( .A1(n548), .A2(n669), .ZN(n492) );
  OR2_X1 U675 ( .A1(n707), .A2(n708), .ZN(n491) );
  AND2_X1 U676 ( .A1(n472), .A2(n471), .ZN(n708) );
  AND2_X1 U677 ( .A1(n469), .A2(n709), .ZN(n707) );
  OR2_X1 U678 ( .A1(n471), .A2(n472), .ZN(n709) );
  OR2_X1 U679 ( .A1(n548), .A2(n481), .ZN(n472) );
  OR2_X1 U680 ( .A1(n710), .A2(n711), .ZN(n471) );
  AND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n711) );
  AND2_X1 U682 ( .A1(n608), .A2(n712), .ZN(n710) );
  OR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n712) );
  OR2_X1 U684 ( .A1(n713), .A2(n714), .ZN(n610) );
  AND2_X1 U685 ( .A1(n592), .A2(n591), .ZN(n714) );
  AND2_X1 U686 ( .A1(n589), .A2(n715), .ZN(n713) );
  OR2_X1 U687 ( .A1(n592), .A2(n591), .ZN(n715) );
  OR2_X1 U688 ( .A1(n716), .A2(n717), .ZN(n591) );
  AND2_X1 U689 ( .A1(n580), .A2(n579), .ZN(n717) );
  AND2_X1 U690 ( .A1(n577), .A2(n718), .ZN(n716) );
  OR2_X1 U691 ( .A1(n580), .A2(n579), .ZN(n718) );
  OR2_X1 U692 ( .A1(n719), .A2(n720), .ZN(n579) );
  AND2_X1 U693 ( .A1(n562), .A2(n563), .ZN(n720) );
  AND2_X1 U694 ( .A1(n560), .A2(n721), .ZN(n719) );
  OR2_X1 U695 ( .A1(n562), .A2(n563), .ZN(n721) );
  OR2_X1 U696 ( .A1(n548), .A2(n722), .ZN(n563) );
  OR2_X1 U697 ( .A1(n723), .A2(n552), .ZN(n722) );
  OR2_X1 U698 ( .A1(n625), .A2(n548), .ZN(n562) );
  XNOR2_X1 U699 ( .A(n724), .B(n725), .ZN(n560) );
  OR2_X1 U700 ( .A1(n723), .A2(n556), .ZN(n724) );
  OR2_X1 U701 ( .A1(n726), .A2(n548), .ZN(n580) );
  XNOR2_X1 U702 ( .A(n727), .B(n728), .ZN(n577) );
  XNOR2_X1 U703 ( .A(n729), .B(n730), .ZN(n727) );
  OR2_X1 U704 ( .A1(n600), .A2(n548), .ZN(n592) );
  XOR2_X1 U705 ( .A(n731), .B(n732), .Z(n589) );
  XOR2_X1 U706 ( .A(n733), .B(n734), .Z(n732) );
  OR2_X1 U707 ( .A1(n735), .A2(n548), .ZN(n611) );
  INV_X1 U708 ( .A(b_7_), .ZN(n548) );
  XOR2_X1 U709 ( .A(n736), .B(n737), .Z(n608) );
  XOR2_X1 U710 ( .A(n738), .B(n739), .Z(n737) );
  XOR2_X1 U711 ( .A(n740), .B(n741), .Z(n469) );
  XOR2_X1 U712 ( .A(n742), .B(n743), .Z(n741) );
  XOR2_X1 U713 ( .A(n744), .B(n745), .Z(n489) );
  XOR2_X1 U714 ( .A(n746), .B(n747), .Z(n745) );
  XOR2_X1 U715 ( .A(n748), .B(n749), .Z(n506) );
  XOR2_X1 U716 ( .A(n750), .B(n751), .Z(n749) );
  OR2_X1 U717 ( .A1(n518), .A2(n752), .ZN(n703) );
  AND2_X1 U718 ( .A1(n512), .A2(n513), .ZN(n752) );
  INV_X1 U719 ( .A(n753), .ZN(n518) );
  OR2_X1 U720 ( .A1(n512), .A2(n513), .ZN(n753) );
  OR2_X1 U721 ( .A1(n754), .A2(n755), .ZN(n513) );
  AND2_X1 U722 ( .A1(n751), .A2(n750), .ZN(n755) );
  AND2_X1 U723 ( .A1(n748), .A2(n756), .ZN(n754) );
  OR2_X1 U724 ( .A1(n750), .A2(n751), .ZN(n756) );
  OR2_X1 U725 ( .A1(n556), .A2(n669), .ZN(n751) );
  OR2_X1 U726 ( .A1(n757), .A2(n758), .ZN(n750) );
  AND2_X1 U727 ( .A1(n747), .A2(n746), .ZN(n758) );
  AND2_X1 U728 ( .A1(n744), .A2(n759), .ZN(n757) );
  OR2_X1 U729 ( .A1(n746), .A2(n747), .ZN(n759) );
  OR2_X1 U730 ( .A1(n556), .A2(n481), .ZN(n747) );
  OR2_X1 U731 ( .A1(n760), .A2(n761), .ZN(n746) );
  AND2_X1 U732 ( .A1(n743), .A2(n742), .ZN(n761) );
  AND2_X1 U733 ( .A1(n740), .A2(n762), .ZN(n760) );
  OR2_X1 U734 ( .A1(n742), .A2(n743), .ZN(n762) );
  OR2_X1 U735 ( .A1(n556), .A2(n735), .ZN(n743) );
  OR2_X1 U736 ( .A1(n763), .A2(n764), .ZN(n742) );
  AND2_X1 U737 ( .A1(n739), .A2(n738), .ZN(n764) );
  AND2_X1 U738 ( .A1(n736), .A2(n765), .ZN(n763) );
  OR2_X1 U739 ( .A1(n739), .A2(n738), .ZN(n765) );
  OR2_X1 U740 ( .A1(n766), .A2(n767), .ZN(n738) );
  AND2_X1 U741 ( .A1(n734), .A2(n733), .ZN(n767) );
  AND2_X1 U742 ( .A1(n731), .A2(n768), .ZN(n766) );
  OR2_X1 U743 ( .A1(n734), .A2(n733), .ZN(n768) );
  OR2_X1 U744 ( .A1(n769), .A2(n770), .ZN(n733) );
  AND2_X1 U745 ( .A1(n729), .A2(n730), .ZN(n770) );
  AND2_X1 U746 ( .A1(n728), .A2(n771), .ZN(n769) );
  OR2_X1 U747 ( .A1(n729), .A2(n730), .ZN(n771) );
  OR2_X1 U748 ( .A1(n552), .A2(n772), .ZN(n730) );
  OR2_X1 U749 ( .A1(n773), .A2(n556), .ZN(n552) );
  OR2_X1 U750 ( .A1(n625), .A2(n556), .ZN(n729) );
  XNOR2_X1 U751 ( .A(n774), .B(n772), .ZN(n728) );
  OR2_X1 U752 ( .A1(n723), .A2(n569), .ZN(n772) );
  OR2_X1 U753 ( .A1(n773), .A2(n686), .ZN(n774) );
  OR2_X1 U754 ( .A1(n726), .A2(n556), .ZN(n734) );
  XOR2_X1 U755 ( .A(n775), .B(n776), .Z(n731) );
  XNOR2_X1 U756 ( .A(n777), .B(n573), .ZN(n776) );
  OR2_X1 U757 ( .A1(n600), .A2(n556), .ZN(n739) );
  INV_X1 U758 ( .A(b_6_), .ZN(n556) );
  XOR2_X1 U759 ( .A(n778), .B(n779), .Z(n736) );
  XOR2_X1 U760 ( .A(n780), .B(n781), .Z(n779) );
  XOR2_X1 U761 ( .A(n782), .B(n783), .Z(n740) );
  XOR2_X1 U762 ( .A(n784), .B(n785), .Z(n783) );
  XOR2_X1 U763 ( .A(n786), .B(n787), .Z(n744) );
  XOR2_X1 U764 ( .A(n788), .B(n789), .Z(n787) );
  XOR2_X1 U765 ( .A(n790), .B(n791), .Z(n748) );
  XOR2_X1 U766 ( .A(n792), .B(n793), .Z(n791) );
  XOR2_X1 U767 ( .A(n681), .B(n794), .Z(n512) );
  XOR2_X1 U768 ( .A(n684), .B(n682), .Z(n794) );
  OR2_X1 U769 ( .A1(n569), .A2(n669), .ZN(n682) );
  OR2_X1 U770 ( .A1(n795), .A2(n796), .ZN(n684) );
  AND2_X1 U771 ( .A1(n793), .A2(n792), .ZN(n796) );
  AND2_X1 U772 ( .A1(n790), .A2(n797), .ZN(n795) );
  OR2_X1 U773 ( .A1(n792), .A2(n793), .ZN(n797) );
  OR2_X1 U774 ( .A1(n569), .A2(n481), .ZN(n793) );
  OR2_X1 U775 ( .A1(n798), .A2(n799), .ZN(n792) );
  AND2_X1 U776 ( .A1(n789), .A2(n788), .ZN(n799) );
  AND2_X1 U777 ( .A1(n786), .A2(n800), .ZN(n798) );
  OR2_X1 U778 ( .A1(n788), .A2(n789), .ZN(n800) );
  OR2_X1 U779 ( .A1(n569), .A2(n735), .ZN(n789) );
  OR2_X1 U780 ( .A1(n801), .A2(n802), .ZN(n788) );
  AND2_X1 U781 ( .A1(n785), .A2(n784), .ZN(n802) );
  AND2_X1 U782 ( .A1(n782), .A2(n803), .ZN(n801) );
  OR2_X1 U783 ( .A1(n784), .A2(n785), .ZN(n803) );
  OR2_X1 U784 ( .A1(n569), .A2(n600), .ZN(n785) );
  OR2_X1 U785 ( .A1(n804), .A2(n805), .ZN(n784) );
  AND2_X1 U786 ( .A1(n781), .A2(n780), .ZN(n805) );
  AND2_X1 U787 ( .A1(n778), .A2(n806), .ZN(n804) );
  OR2_X1 U788 ( .A1(n781), .A2(n780), .ZN(n806) );
  OR2_X1 U789 ( .A1(n807), .A2(n808), .ZN(n780) );
  AND2_X1 U790 ( .A1(n620), .A2(n777), .ZN(n808) );
  AND2_X1 U791 ( .A1(n809), .A2(n775), .ZN(n807) );
  OR2_X1 U792 ( .A1(n810), .A2(n811), .ZN(n775) );
  INV_X1 U793 ( .A(n812), .ZN(n811) );
  AND2_X1 U794 ( .A1(n813), .A2(n814), .ZN(n810) );
  OR2_X1 U795 ( .A1(n620), .A2(n777), .ZN(n809) );
  OR2_X1 U796 ( .A1(n814), .A2(n725), .ZN(n777) );
  OR2_X1 U797 ( .A1(n773), .A2(n569), .ZN(n725) );
  INV_X1 U798 ( .A(n573), .ZN(n620) );
  AND2_X1 U799 ( .A1(a_5_), .A2(b_5_), .ZN(n573) );
  OR2_X1 U800 ( .A1(n726), .A2(n569), .ZN(n781) );
  INV_X1 U801 ( .A(b_5_), .ZN(n569) );
  XNOR2_X1 U802 ( .A(n815), .B(n816), .ZN(n778) );
  XNOR2_X1 U803 ( .A(n817), .B(n812), .ZN(n815) );
  XNOR2_X1 U804 ( .A(n818), .B(n819), .ZN(n782) );
  XNOR2_X1 U805 ( .A(n584), .B(n820), .ZN(n818) );
  XOR2_X1 U806 ( .A(n821), .B(n822), .Z(n786) );
  XOR2_X1 U807 ( .A(n823), .B(n824), .Z(n822) );
  XOR2_X1 U808 ( .A(n825), .B(n826), .Z(n790) );
  XOR2_X1 U809 ( .A(n827), .B(n828), .Z(n826) );
  XOR2_X1 U810 ( .A(n689), .B(n829), .Z(n681) );
  XOR2_X1 U811 ( .A(n692), .B(n690), .Z(n829) );
  OR2_X1 U812 ( .A1(n686), .A2(n481), .ZN(n690) );
  OR2_X1 U813 ( .A1(n830), .A2(n831), .ZN(n692) );
  AND2_X1 U814 ( .A1(n828), .A2(n827), .ZN(n831) );
  AND2_X1 U815 ( .A1(n825), .A2(n832), .ZN(n830) );
  OR2_X1 U816 ( .A1(n827), .A2(n828), .ZN(n832) );
  OR2_X1 U817 ( .A1(n686), .A2(n735), .ZN(n828) );
  OR2_X1 U818 ( .A1(n833), .A2(n834), .ZN(n827) );
  AND2_X1 U819 ( .A1(n824), .A2(n823), .ZN(n834) );
  AND2_X1 U820 ( .A1(n821), .A2(n835), .ZN(n833) );
  OR2_X1 U821 ( .A1(n823), .A2(n824), .ZN(n835) );
  OR2_X1 U822 ( .A1(n686), .A2(n600), .ZN(n824) );
  OR2_X1 U823 ( .A1(n836), .A2(n837), .ZN(n823) );
  AND2_X1 U824 ( .A1(n820), .A2(n584), .ZN(n837) );
  AND2_X1 U825 ( .A1(n819), .A2(n838), .ZN(n836) );
  OR2_X1 U826 ( .A1(n584), .A2(n820), .ZN(n838) );
  OR2_X1 U827 ( .A1(n839), .A2(n840), .ZN(n820) );
  AND2_X1 U828 ( .A1(n816), .A2(n812), .ZN(n840) );
  AND2_X1 U829 ( .A1(n841), .A2(n817), .ZN(n839) );
  OR2_X1 U830 ( .A1(n842), .A2(n843), .ZN(n817) );
  AND2_X1 U831 ( .A1(n844), .A2(n845), .ZN(n842) );
  OR2_X1 U832 ( .A1(n816), .A2(n812), .ZN(n841) );
  OR2_X1 U833 ( .A1(n813), .A2(n814), .ZN(n812) );
  OR2_X1 U834 ( .A1(n723), .A2(n686), .ZN(n814) );
  OR2_X1 U835 ( .A1(n773), .A2(n599), .ZN(n813) );
  OR2_X1 U836 ( .A1(n625), .A2(n686), .ZN(n816) );
  OR2_X1 U837 ( .A1(n726), .A2(n686), .ZN(n584) );
  INV_X1 U838 ( .A(b_4_), .ZN(n686) );
  XOR2_X1 U839 ( .A(n846), .B(n843), .Z(n819) );
  INV_X1 U840 ( .A(n847), .ZN(n843) );
  XNOR2_X1 U841 ( .A(n848), .B(n849), .ZN(n846) );
  XNOR2_X1 U842 ( .A(n850), .B(n851), .ZN(n821) );
  XNOR2_X1 U843 ( .A(n852), .B(n853), .ZN(n850) );
  XNOR2_X1 U844 ( .A(n854), .B(n855), .ZN(n825) );
  XNOR2_X1 U845 ( .A(n616), .B(n856), .ZN(n854) );
  XNOR2_X1 U846 ( .A(n857), .B(n701), .ZN(n689) );
  XNOR2_X1 U847 ( .A(n858), .B(n859), .ZN(n701) );
  XNOR2_X1 U848 ( .A(n860), .B(n861), .ZN(n858) );
  XNOR2_X1 U849 ( .A(n700), .B(n699), .ZN(n857) );
  OR2_X1 U850 ( .A1(n862), .A2(n863), .ZN(n699) );
  AND2_X1 U851 ( .A1(n856), .A2(n616), .ZN(n863) );
  AND2_X1 U852 ( .A1(n855), .A2(n864), .ZN(n862) );
  OR2_X1 U853 ( .A1(n616), .A2(n856), .ZN(n864) );
  OR2_X1 U854 ( .A1(n865), .A2(n866), .ZN(n856) );
  AND2_X1 U855 ( .A1(n853), .A2(n852), .ZN(n866) );
  AND2_X1 U856 ( .A1(n851), .A2(n867), .ZN(n865) );
  OR2_X1 U857 ( .A1(n852), .A2(n853), .ZN(n867) );
  OR2_X1 U858 ( .A1(n868), .A2(n869), .ZN(n853) );
  AND2_X1 U859 ( .A1(n847), .A2(n849), .ZN(n869) );
  AND2_X1 U860 ( .A1(n870), .A2(n848), .ZN(n868) );
  OR2_X1 U861 ( .A1(n871), .A2(n872), .ZN(n848) );
  INV_X1 U862 ( .A(n873), .ZN(n872) );
  AND2_X1 U863 ( .A1(n874), .A2(n875), .ZN(n871) );
  OR2_X1 U864 ( .A1(n849), .A2(n847), .ZN(n870) );
  OR2_X1 U865 ( .A1(n844), .A2(n845), .ZN(n847) );
  OR2_X1 U866 ( .A1(n773), .A2(n876), .ZN(n845) );
  OR2_X1 U867 ( .A1(n723), .A2(n599), .ZN(n844) );
  OR2_X1 U868 ( .A1(n599), .A2(n625), .ZN(n849) );
  OR2_X1 U869 ( .A1(n599), .A2(n726), .ZN(n852) );
  XNOR2_X1 U870 ( .A(n877), .B(n878), .ZN(n851) );
  XNOR2_X1 U871 ( .A(n879), .B(n873), .ZN(n877) );
  INV_X1 U872 ( .A(n604), .ZN(n616) );
  AND2_X1 U873 ( .A1(b_3_), .A2(a_3_), .ZN(n604) );
  XOR2_X1 U874 ( .A(n880), .B(n881), .Z(n855) );
  XOR2_X1 U875 ( .A(n882), .B(n883), .Z(n881) );
  OR2_X1 U876 ( .A1(n599), .A2(n735), .ZN(n700) );
  INV_X1 U877 ( .A(b_3_), .ZN(n599) );
  AND2_X1 U878 ( .A1(n541), .A2(n884), .ZN(n543) );
  AND2_X1 U879 ( .A1(n542), .A2(n540), .ZN(n884) );
  XOR2_X1 U880 ( .A(n885), .B(n886), .Z(n540) );
  OR2_X1 U881 ( .A1(n496), .A2(n669), .ZN(n885) );
  XNOR2_X1 U882 ( .A(n887), .B(n888), .ZN(n542) );
  XOR2_X1 U883 ( .A(n889), .B(n890), .Z(n888) );
  INV_X1 U884 ( .A(n630), .ZN(n541) );
  OR2_X1 U885 ( .A1(n891), .A2(n892), .ZN(n630) );
  AND2_X1 U886 ( .A1(n651), .A2(n650), .ZN(n892) );
  AND2_X1 U887 ( .A1(n648), .A2(n893), .ZN(n891) );
  OR2_X1 U888 ( .A1(n650), .A2(n651), .ZN(n893) );
  OR2_X1 U889 ( .A1(n876), .A2(n669), .ZN(n651) );
  OR2_X1 U890 ( .A1(n894), .A2(n895), .ZN(n650) );
  AND2_X1 U891 ( .A1(n662), .A2(n661), .ZN(n895) );
  AND2_X1 U892 ( .A1(n659), .A2(n896), .ZN(n894) );
  OR2_X1 U893 ( .A1(n661), .A2(n662), .ZN(n896) );
  OR2_X1 U894 ( .A1(n876), .A2(n481), .ZN(n662) );
  OR2_X1 U895 ( .A1(n897), .A2(n898), .ZN(n661) );
  AND2_X1 U896 ( .A1(n696), .A2(n503), .ZN(n898) );
  AND2_X1 U897 ( .A1(n695), .A2(n899), .ZN(n897) );
  OR2_X1 U898 ( .A1(n503), .A2(n696), .ZN(n899) );
  OR2_X1 U899 ( .A1(n900), .A2(n901), .ZN(n696) );
  AND2_X1 U900 ( .A1(n861), .A2(n860), .ZN(n901) );
  AND2_X1 U901 ( .A1(n859), .A2(n902), .ZN(n900) );
  OR2_X1 U902 ( .A1(n860), .A2(n861), .ZN(n902) );
  OR2_X1 U903 ( .A1(n903), .A2(n904), .ZN(n861) );
  AND2_X1 U904 ( .A1(n883), .A2(n882), .ZN(n904) );
  AND2_X1 U905 ( .A1(n880), .A2(n905), .ZN(n903) );
  OR2_X1 U906 ( .A1(n882), .A2(n883), .ZN(n905) );
  OR2_X1 U907 ( .A1(n876), .A2(n726), .ZN(n883) );
  OR2_X1 U908 ( .A1(n906), .A2(n907), .ZN(n882) );
  AND2_X1 U909 ( .A1(n878), .A2(n873), .ZN(n907) );
  AND2_X1 U910 ( .A1(n908), .A2(n879), .ZN(n906) );
  OR2_X1 U911 ( .A1(n909), .A2(n910), .ZN(n879) );
  INV_X1 U912 ( .A(n911), .ZN(n910) );
  AND2_X1 U913 ( .A1(n912), .A2(n913), .ZN(n909) );
  OR2_X1 U914 ( .A1(n873), .A2(n878), .ZN(n908) );
  OR2_X1 U915 ( .A1(n876), .A2(n625), .ZN(n878) );
  OR2_X1 U916 ( .A1(n874), .A2(n875), .ZN(n873) );
  OR2_X1 U917 ( .A1(n876), .A2(n723), .ZN(n875) );
  OR2_X1 U918 ( .A1(n773), .A2(n480), .ZN(n874) );
  XNOR2_X1 U919 ( .A(n914), .B(n911), .ZN(n880) );
  OR2_X1 U920 ( .A1(n915), .A2(n916), .ZN(n914) );
  INV_X1 U921 ( .A(n917), .ZN(n916) );
  AND2_X1 U922 ( .A1(n918), .A2(n919), .ZN(n915) );
  OR2_X1 U923 ( .A1(n876), .A2(n600), .ZN(n860) );
  XOR2_X1 U924 ( .A(n920), .B(n921), .Z(n859) );
  XOR2_X1 U925 ( .A(n922), .B(n923), .Z(n920) );
  OR2_X1 U926 ( .A1(n876), .A2(n735), .ZN(n503) );
  INV_X1 U927 ( .A(b_2_), .ZN(n876) );
  XOR2_X1 U928 ( .A(n924), .B(n925), .Z(n695) );
  XOR2_X1 U929 ( .A(n926), .B(n927), .Z(n925) );
  XOR2_X1 U930 ( .A(n928), .B(n929), .Z(n659) );
  XOR2_X1 U931 ( .A(n930), .B(n931), .Z(n929) );
  XNOR2_X1 U932 ( .A(n932), .B(n933), .ZN(n648) );
  XNOR2_X1 U933 ( .A(n934), .B(n935), .ZN(n932) );
  AND2_X1 U934 ( .A1(n936), .A2(a_0_), .ZN(n627) );
  INV_X1 U935 ( .A(n886), .ZN(n936) );
  OR2_X1 U936 ( .A1(n937), .A2(n938), .ZN(n886) );
  AND2_X1 U937 ( .A1(n887), .A2(n889), .ZN(n938) );
  AND2_X1 U938 ( .A1(n939), .A2(n890), .ZN(n937) );
  OR2_X1 U939 ( .A1(n480), .A2(n669), .ZN(n890) );
  INV_X1 U940 ( .A(a_0_), .ZN(n669) );
  OR2_X1 U941 ( .A1(n889), .A2(n887), .ZN(n939) );
  OR2_X1 U942 ( .A1(n481), .A2(n496), .ZN(n887) );
  INV_X1 U943 ( .A(a_1_), .ZN(n481) );
  OR2_X1 U944 ( .A1(n940), .A2(n941), .ZN(n889) );
  AND2_X1 U945 ( .A1(n933), .A2(n935), .ZN(n941) );
  AND2_X1 U946 ( .A1(n942), .A2(n934), .ZN(n940) );
  INV_X1 U947 ( .A(n485), .ZN(n934) );
  AND2_X1 U948 ( .A1(b_1_), .A2(a_1_), .ZN(n485) );
  OR2_X1 U949 ( .A1(n935), .A2(n933), .ZN(n942) );
  OR2_X1 U950 ( .A1(n735), .A2(n496), .ZN(n933) );
  OR2_X1 U951 ( .A1(n943), .A2(n944), .ZN(n935) );
  AND2_X1 U952 ( .A1(n928), .A2(n930), .ZN(n944) );
  AND2_X1 U953 ( .A1(n945), .A2(n931), .ZN(n943) );
  OR2_X1 U954 ( .A1(n600), .A2(n496), .ZN(n931) );
  OR2_X1 U955 ( .A1(n930), .A2(n928), .ZN(n945) );
  OR2_X1 U956 ( .A1(n480), .A2(n735), .ZN(n928) );
  INV_X1 U957 ( .A(a_2_), .ZN(n735) );
  OR2_X1 U958 ( .A1(n946), .A2(n947), .ZN(n930) );
  AND2_X1 U959 ( .A1(n924), .A2(n926), .ZN(n947) );
  AND2_X1 U960 ( .A1(n948), .A2(n927), .ZN(n946) );
  OR2_X1 U961 ( .A1(n480), .A2(n600), .ZN(n927) );
  INV_X1 U962 ( .A(a_3_), .ZN(n600) );
  OR2_X1 U963 ( .A1(n926), .A2(n924), .ZN(n948) );
  OR2_X1 U964 ( .A1(n726), .A2(n496), .ZN(n924) );
  OR2_X1 U965 ( .A1(n949), .A2(n950), .ZN(n926) );
  AND2_X1 U966 ( .A1(n921), .A2(n923), .ZN(n950) );
  AND2_X1 U967 ( .A1(n922), .A2(n951), .ZN(n949) );
  OR2_X1 U968 ( .A1(n923), .A2(n921), .ZN(n951) );
  OR2_X1 U969 ( .A1(n625), .A2(n496), .ZN(n921) );
  OR2_X1 U970 ( .A1(n480), .A2(n726), .ZN(n923) );
  INV_X1 U971 ( .A(a_4_), .ZN(n726) );
  AND2_X1 U972 ( .A1(n917), .A2(n911), .ZN(n922) );
  OR2_X1 U973 ( .A1(n913), .A2(n912), .ZN(n911) );
  OR2_X1 U974 ( .A1(n773), .A2(n496), .ZN(n912) );
  INV_X1 U975 ( .A(a_7_), .ZN(n773) );
  OR2_X1 U976 ( .A1(n723), .A2(n480), .ZN(n913) );
  OR2_X1 U977 ( .A1(n919), .A2(n918), .ZN(n917) );
  OR2_X1 U978 ( .A1(n723), .A2(n496), .ZN(n918) );
  INV_X1 U979 ( .A(b_0_), .ZN(n496) );
  INV_X1 U980 ( .A(a_6_), .ZN(n723) );
  OR2_X1 U981 ( .A1(n480), .A2(n625), .ZN(n919) );
  INV_X1 U982 ( .A(a_5_), .ZN(n625) );
  INV_X1 U983 ( .A(b_1_), .ZN(n480) );
endmodule

