module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n1009_, new_n238_, new_n479_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n1017_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n1033_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n172_, keyIn_0_45 );
not g001 ( new_n173_, keyIn_0_28 );
not g002 ( new_n174_, N108 );
not g003 ( new_n175_, N102 );
and g004 ( new_n176_, new_n175_, keyIn_0_16 );
not g005 ( new_n177_, keyIn_0_16 );
and g006 ( new_n178_, new_n177_, N102 );
or g007 ( new_n179_, new_n176_, new_n178_, new_n174_ );
and g008 ( new_n180_, new_n179_, new_n173_ );
not g009 ( new_n181_, new_n176_ );
not g010 ( new_n182_, new_n178_ );
and g011 ( new_n183_, new_n181_, new_n182_, keyIn_0_28, N108 );
or g012 ( new_n184_, new_n180_, new_n183_ );
not g013 ( new_n185_, keyIn_0_27 );
not g014 ( new_n186_, N95 );
or g015 ( new_n187_, keyIn_0_14, N89 );
not g016 ( new_n188_, new_n187_ );
and g017 ( new_n189_, keyIn_0_14, N89 );
or g018 ( new_n190_, new_n188_, new_n186_, new_n189_ );
and g019 ( new_n191_, new_n190_, new_n185_ );
not g020 ( new_n192_, new_n189_ );
and g021 ( new_n193_, new_n192_, keyIn_0_27, N95, new_n187_ );
or g022 ( new_n194_, new_n191_, new_n193_ );
not g023 ( new_n195_, N76 );
and g024 ( new_n196_, new_n195_, keyIn_0_12 );
not g025 ( new_n197_, new_n196_ );
or g026 ( new_n198_, new_n195_, keyIn_0_12 );
and g027 ( new_n199_, new_n197_, new_n198_, N82 );
or g028 ( new_n200_, new_n199_, keyIn_0_26 );
not g029 ( new_n201_, keyIn_0_26 );
not g030 ( new_n202_, N82 );
not g031 ( new_n203_, new_n198_ );
or g032 ( new_n204_, new_n203_, new_n201_, new_n202_, new_n196_ );
and g033 ( new_n205_, new_n200_, new_n204_ );
and g034 ( new_n206_, new_n194_, new_n205_, new_n184_ );
not g035 ( new_n207_, N4 );
not g036 ( new_n208_, N1 );
and g037 ( new_n209_, new_n208_, keyIn_0_0 );
not g038 ( new_n210_, keyIn_0_0 );
and g039 ( new_n211_, new_n210_, N1 );
or g040 ( new_n212_, new_n209_, new_n211_, new_n207_ );
and g041 ( new_n213_, new_n212_, keyIn_0_18 );
not g042 ( new_n214_, keyIn_0_18 );
not g043 ( new_n215_, new_n209_ );
not g044 ( new_n216_, new_n211_ );
and g045 ( new_n217_, new_n215_, new_n216_, new_n214_, N4 );
or g046 ( new_n218_, new_n213_, new_n217_ );
not g047 ( new_n219_, keyIn_0_21 );
not g048 ( new_n220_, N17 );
not g049 ( new_n221_, N11 );
and g050 ( new_n222_, new_n221_, keyIn_0_2 );
not g051 ( new_n223_, keyIn_0_2 );
and g052 ( new_n224_, new_n223_, N11 );
or g053 ( new_n225_, new_n222_, new_n224_, new_n220_ );
and g054 ( new_n226_, new_n225_, new_n219_ );
not g055 ( new_n227_, new_n222_ );
not g056 ( new_n228_, new_n224_ );
and g057 ( new_n229_, new_n227_, new_n228_, keyIn_0_21, N17 );
or g058 ( new_n230_, new_n226_, new_n229_ );
and g059 ( new_n231_, new_n218_, new_n230_ );
not g060 ( new_n232_, keyIn_0_22 );
not g061 ( new_n233_, N30 );
not g062 ( new_n234_, N24 );
and g063 ( new_n235_, new_n234_, keyIn_0_4 );
not g064 ( new_n236_, keyIn_0_4 );
and g065 ( new_n237_, new_n236_, N24 );
or g066 ( new_n238_, new_n235_, new_n237_, new_n233_ );
and g067 ( new_n239_, new_n238_, new_n232_ );
not g068 ( new_n240_, new_n235_ );
not g069 ( new_n241_, new_n237_ );
and g070 ( new_n242_, new_n240_, new_n241_, keyIn_0_22, N30 );
or g071 ( new_n243_, new_n239_, new_n242_ );
not g072 ( new_n244_, keyIn_0_23 );
and g073 ( new_n245_, keyIn_0_6, N37 );
not g074 ( new_n246_, new_n245_ );
or g075 ( new_n247_, keyIn_0_6, N37 );
and g076 ( new_n248_, new_n246_, new_n247_ );
not g077 ( new_n249_, new_n248_ );
and g078 ( new_n250_, new_n249_, new_n244_, N43 );
not g079 ( new_n251_, N43 );
or g080 ( new_n252_, new_n248_, new_n251_ );
and g081 ( new_n253_, new_n252_, keyIn_0_23 );
or g082 ( new_n254_, new_n253_, new_n250_ );
and g083 ( new_n255_, new_n254_, new_n243_ );
not g084 ( new_n256_, keyIn_0_10 );
or g085 ( new_n257_, new_n256_, N63 );
not g086 ( new_n258_, N63 );
or g087 ( new_n259_, new_n258_, keyIn_0_10 );
and g088 ( new_n260_, new_n257_, new_n259_, N69 );
or g089 ( new_n261_, new_n260_, keyIn_0_25 );
not g090 ( new_n262_, keyIn_0_25 );
not g091 ( new_n263_, N69 );
not g092 ( new_n264_, new_n257_ );
not g093 ( new_n265_, new_n259_ );
or g094 ( new_n266_, new_n264_, new_n265_, new_n262_, new_n263_ );
and g095 ( new_n267_, new_n266_, new_n261_ );
not g096 ( new_n268_, keyIn_0_8 );
or g097 ( new_n269_, new_n268_, N50 );
not g098 ( new_n270_, N50 );
or g099 ( new_n271_, new_n270_, keyIn_0_8 );
and g100 ( new_n272_, new_n269_, new_n271_, N56 );
or g101 ( new_n273_, new_n272_, keyIn_0_24 );
not g102 ( new_n274_, keyIn_0_24 );
not g103 ( new_n275_, N56 );
not g104 ( new_n276_, new_n269_ );
not g105 ( new_n277_, new_n271_ );
or g106 ( new_n278_, new_n276_, new_n277_, new_n274_, new_n275_ );
and g107 ( new_n279_, new_n278_, new_n273_ );
and g108 ( new_n280_, new_n267_, new_n279_ );
and g109 ( new_n281_, new_n255_, new_n206_, new_n231_, new_n280_ );
or g110 ( new_n282_, new_n281_, new_n172_ );
and g111 ( new_n283_, new_n280_, new_n243_, new_n254_ );
and g112 ( new_n284_, new_n283_, new_n172_, new_n206_, new_n231_ );
not g113 ( new_n285_, new_n284_ );
and g114 ( N223, new_n282_, new_n285_ );
not g115 ( new_n287_, keyIn_0_63 );
not g116 ( new_n288_, keyIn_0_52 );
not g117 ( new_n289_, new_n279_ );
and g118 ( new_n290_, new_n282_, new_n285_, keyIn_0_46 );
not g119 ( new_n291_, new_n290_ );
or g120 ( new_n292_, N223, keyIn_0_46 );
and g121 ( new_n293_, new_n292_, new_n291_ );
or g122 ( new_n294_, new_n293_, new_n289_ );
and g123 ( new_n295_, new_n293_, new_n289_ );
not g124 ( new_n296_, new_n295_ );
and g125 ( new_n297_, new_n296_, new_n288_, new_n294_ );
not g126 ( new_n298_, new_n297_ );
and g127 ( new_n299_, new_n296_, new_n294_ );
or g128 ( new_n300_, new_n299_, new_n288_ );
not g129 ( new_n301_, N60 );
and g130 ( new_n302_, new_n275_, keyIn_0_9 );
not g131 ( new_n303_, new_n302_ );
or g132 ( new_n304_, new_n275_, keyIn_0_9 );
and g133 ( new_n305_, new_n303_, new_n304_ );
not g134 ( new_n306_, new_n305_ );
and g135 ( new_n307_, new_n306_, new_n301_ );
or g136 ( new_n308_, new_n307_, keyIn_0_35 );
not g137 ( new_n309_, keyIn_0_35 );
or g138 ( new_n310_, new_n305_, new_n309_, N60 );
and g139 ( new_n311_, new_n308_, new_n310_ );
and g140 ( new_n312_, new_n300_, new_n298_, new_n311_ );
not g141 ( new_n313_, new_n312_ );
and g142 ( new_n314_, new_n313_, new_n287_ );
and g143 ( new_n315_, new_n312_, keyIn_0_63 );
or g144 ( new_n316_, new_n314_, new_n315_ );
not g145 ( new_n317_, keyIn_0_67 );
not g146 ( new_n318_, keyIn_0_56 );
or g147 ( new_n319_, new_n293_, new_n184_ );
and g148 ( new_n320_, new_n292_, new_n184_, new_n291_ );
not g149 ( new_n321_, new_n320_ );
and g150 ( new_n322_, new_n319_, new_n318_, new_n321_ );
not g151 ( new_n323_, new_n322_ );
and g152 ( new_n324_, new_n319_, new_n321_ );
or g153 ( new_n325_, new_n324_, new_n318_ );
and g154 ( new_n326_, new_n325_, new_n323_ );
not g155 ( new_n327_, keyIn_0_43 );
not g156 ( new_n328_, N112 );
or g157 ( new_n329_, keyIn_0_17, N108 );
and g158 ( new_n330_, keyIn_0_17, N108 );
not g159 ( new_n331_, new_n330_ );
and g160 ( new_n332_, new_n331_, new_n329_ );
not g161 ( new_n333_, new_n332_ );
and g162 ( new_n334_, new_n333_, new_n328_ );
and g163 ( new_n335_, new_n334_, new_n327_ );
not g164 ( new_n336_, new_n335_ );
or g165 ( new_n337_, new_n334_, new_n327_ );
and g166 ( new_n338_, new_n336_, new_n337_ );
or g167 ( new_n339_, new_n326_, new_n338_ );
and g168 ( new_n340_, new_n339_, new_n317_ );
not g169 ( new_n341_, new_n326_ );
not g170 ( new_n342_, new_n338_ );
and g171 ( new_n343_, new_n341_, keyIn_0_67, new_n342_ );
or g172 ( new_n344_, new_n340_, new_n343_ );
not g173 ( new_n345_, keyIn_0_64 );
not g174 ( new_n346_, keyIn_0_53 );
not g175 ( new_n347_, new_n267_ );
or g176 ( new_n348_, new_n293_, new_n347_ );
and g177 ( new_n349_, new_n293_, new_n347_ );
not g178 ( new_n350_, new_n349_ );
and g179 ( new_n351_, new_n350_, new_n348_ );
and g180 ( new_n352_, new_n351_, new_n346_ );
not g181 ( new_n353_, new_n352_ );
or g182 ( new_n354_, new_n351_, new_n346_ );
not g183 ( new_n355_, N73 );
and g184 ( new_n356_, new_n263_, keyIn_0_11 );
not g185 ( new_n357_, new_n356_ );
or g186 ( new_n358_, new_n263_, keyIn_0_11 );
and g187 ( new_n359_, new_n357_, new_n358_ );
not g188 ( new_n360_, new_n359_ );
and g189 ( new_n361_, new_n360_, new_n355_ );
or g190 ( new_n362_, new_n361_, keyIn_0_37 );
not g191 ( new_n363_, keyIn_0_37 );
or g192 ( new_n364_, new_n359_, new_n363_, N73 );
and g193 ( new_n365_, new_n362_, new_n364_ );
and g194 ( new_n366_, new_n353_, new_n354_, new_n365_ );
or g195 ( new_n367_, new_n366_, new_n345_ );
and g196 ( new_n368_, new_n353_, new_n345_, new_n354_, new_n365_ );
not g197 ( new_n369_, new_n368_ );
and g198 ( new_n370_, new_n367_, new_n369_ );
and g199 ( new_n371_, new_n344_, new_n316_, new_n370_ );
not g200 ( new_n372_, keyIn_0_65 );
not g201 ( new_n373_, keyIn_0_54 );
not g202 ( new_n374_, new_n293_ );
and g203 ( new_n375_, new_n374_, new_n205_ );
not g204 ( new_n376_, new_n375_ );
not g205 ( new_n377_, new_n205_ );
and g206 ( new_n378_, new_n293_, new_n377_ );
not g207 ( new_n379_, new_n378_ );
and g208 ( new_n380_, new_n376_, new_n379_ );
and g209 ( new_n381_, new_n380_, new_n373_ );
or g210 ( new_n382_, new_n375_, new_n378_ );
and g211 ( new_n383_, new_n382_, keyIn_0_54 );
or g212 ( new_n384_, new_n381_, new_n383_ );
not g213 ( new_n385_, keyIn_0_39 );
not g214 ( new_n386_, N86 );
and g215 ( new_n387_, new_n202_, keyIn_0_13 );
not g216 ( new_n388_, new_n387_ );
or g217 ( new_n389_, new_n202_, keyIn_0_13 );
and g218 ( new_n390_, new_n388_, new_n389_ );
not g219 ( new_n391_, new_n390_ );
and g220 ( new_n392_, new_n391_, new_n386_ );
not g221 ( new_n393_, new_n392_ );
and g222 ( new_n394_, new_n393_, new_n385_ );
and g223 ( new_n395_, new_n392_, keyIn_0_39 );
or g224 ( new_n396_, new_n394_, new_n395_ );
not g225 ( new_n397_, new_n396_ );
and g226 ( new_n398_, new_n384_, new_n397_ );
or g227 ( new_n399_, new_n398_, new_n372_ );
not g228 ( new_n400_, new_n384_ );
or g229 ( new_n401_, new_n400_, keyIn_0_65, new_n396_ );
or g230 ( new_n402_, new_n293_, new_n194_ );
and g231 ( new_n403_, new_n293_, new_n194_ );
not g232 ( new_n404_, new_n403_ );
and g233 ( new_n405_, new_n404_, new_n402_ );
or g234 ( new_n406_, new_n405_, keyIn_0_55 );
and g235 ( new_n407_, new_n405_, keyIn_0_55 );
not g236 ( new_n408_, new_n407_ );
not g237 ( new_n409_, keyIn_0_41 );
not g238 ( new_n410_, N99 );
or g239 ( new_n411_, keyIn_0_15, N95 );
and g240 ( new_n412_, keyIn_0_15, N95 );
not g241 ( new_n413_, new_n412_ );
and g242 ( new_n414_, new_n413_, new_n411_ );
not g243 ( new_n415_, new_n414_ );
and g244 ( new_n416_, new_n415_, new_n410_ );
and g245 ( new_n417_, new_n416_, new_n409_ );
not g246 ( new_n418_, new_n416_ );
and g247 ( new_n419_, new_n418_, keyIn_0_41 );
or g248 ( new_n420_, new_n419_, new_n417_ );
and g249 ( new_n421_, new_n408_, new_n406_, new_n420_ );
or g250 ( new_n422_, new_n421_, keyIn_0_66 );
and g251 ( new_n423_, new_n408_, keyIn_0_66, new_n406_, new_n420_ );
not g252 ( new_n424_, new_n423_ );
and g253 ( new_n425_, new_n422_, new_n424_ );
and g254 ( new_n426_, new_n425_, new_n399_, new_n401_ );
not g255 ( new_n427_, new_n243_ );
or g256 ( new_n428_, new_n293_, new_n427_ );
and g257 ( new_n429_, new_n292_, new_n427_, new_n291_ );
not g258 ( new_n430_, new_n429_ );
and g259 ( new_n431_, new_n428_, keyIn_0_50, new_n430_ );
not g260 ( new_n432_, new_n431_ );
and g261 ( new_n433_, new_n428_, new_n430_ );
or g262 ( new_n434_, new_n433_, keyIn_0_50 );
and g263 ( new_n435_, new_n434_, new_n432_ );
not g264 ( new_n436_, new_n435_ );
not g265 ( new_n437_, keyIn_0_31 );
not g266 ( new_n438_, N34 );
and g267 ( new_n439_, keyIn_0_5, N30 );
not g268 ( new_n440_, new_n439_ );
or g269 ( new_n441_, keyIn_0_5, N30 );
and g270 ( new_n442_, new_n440_, new_n438_, new_n441_ );
not g271 ( new_n443_, new_n442_ );
and g272 ( new_n444_, new_n443_, new_n437_ );
and g273 ( new_n445_, new_n442_, keyIn_0_31 );
or g274 ( new_n446_, new_n444_, new_n445_ );
and g275 ( new_n447_, new_n436_, keyIn_0_61, new_n446_ );
not g276 ( new_n448_, keyIn_0_61 );
not g277 ( new_n449_, new_n446_ );
or g278 ( new_n450_, new_n435_, new_n449_ );
and g279 ( new_n451_, new_n450_, new_n448_ );
or g280 ( new_n452_, new_n451_, new_n447_ );
not g281 ( new_n453_, new_n254_ );
or g282 ( new_n454_, new_n293_, new_n453_ );
and g283 ( new_n455_, new_n293_, new_n453_ );
not g284 ( new_n456_, new_n455_ );
and g285 ( new_n457_, new_n456_, new_n454_ );
and g286 ( new_n458_, new_n457_, keyIn_0_51 );
not g287 ( new_n459_, new_n458_ );
or g288 ( new_n460_, new_n457_, keyIn_0_51 );
not g289 ( new_n461_, keyIn_0_33 );
not g290 ( new_n462_, N47 );
or g291 ( new_n463_, keyIn_0_7, N43 );
and g292 ( new_n464_, keyIn_0_7, N43 );
not g293 ( new_n465_, new_n464_ );
and g294 ( new_n466_, new_n465_, new_n463_ );
not g295 ( new_n467_, new_n466_ );
and g296 ( new_n468_, new_n467_, new_n462_ );
and g297 ( new_n469_, new_n468_, new_n461_ );
not g298 ( new_n470_, new_n468_ );
and g299 ( new_n471_, new_n470_, keyIn_0_33 );
or g300 ( new_n472_, new_n471_, new_n469_ );
and g301 ( new_n473_, new_n459_, new_n460_, new_n472_ );
or g302 ( new_n474_, new_n473_, keyIn_0_62 );
and g303 ( new_n475_, new_n459_, keyIn_0_62, new_n460_, new_n472_ );
not g304 ( new_n476_, new_n475_ );
and g305 ( new_n477_, new_n474_, new_n476_ );
not g306 ( new_n478_, keyIn_0_60 );
not g307 ( new_n479_, keyIn_0_49 );
or g308 ( new_n480_, new_n293_, new_n230_ );
and g309 ( new_n481_, new_n293_, new_n230_ );
not g310 ( new_n482_, new_n481_ );
and g311 ( new_n483_, new_n482_, new_n479_, new_n480_ );
not g312 ( new_n484_, new_n483_ );
and g313 ( new_n485_, new_n482_, new_n480_ );
or g314 ( new_n486_, new_n485_, new_n479_ );
not g315 ( new_n487_, N21 );
or g316 ( new_n488_, keyIn_0_3, N17 );
and g317 ( new_n489_, keyIn_0_3, N17 );
not g318 ( new_n490_, new_n489_ );
and g319 ( new_n491_, new_n490_, new_n488_ );
not g320 ( new_n492_, new_n491_ );
and g321 ( new_n493_, new_n492_, new_n487_ );
or g322 ( new_n494_, new_n493_, keyIn_0_29 );
not g323 ( new_n495_, keyIn_0_29 );
or g324 ( new_n496_, new_n491_, new_n495_, N21 );
and g325 ( new_n497_, new_n494_, new_n496_ );
and g326 ( new_n498_, new_n486_, new_n484_, new_n497_ );
or g327 ( new_n499_, new_n498_, new_n478_ );
and g328 ( new_n500_, new_n498_, new_n478_ );
not g329 ( new_n501_, new_n500_ );
and g330 ( new_n502_, new_n501_, new_n499_ );
not g331 ( new_n503_, keyIn_0_48 );
not g332 ( new_n504_, new_n218_ );
and g333 ( new_n505_, new_n292_, new_n504_, new_n291_ );
not g334 ( new_n506_, new_n505_ );
or g335 ( new_n507_, new_n293_, new_n504_ );
and g336 ( new_n508_, new_n507_, new_n503_, new_n506_ );
not g337 ( new_n509_, new_n508_ );
and g338 ( new_n510_, new_n507_, new_n506_ );
or g339 ( new_n511_, new_n510_, new_n503_ );
not g340 ( new_n512_, N8 );
and g341 ( new_n513_, new_n207_, keyIn_0_1 );
not g342 ( new_n514_, new_n513_ );
or g343 ( new_n515_, new_n207_, keyIn_0_1 );
and g344 ( new_n516_, new_n514_, new_n515_ );
not g345 ( new_n517_, new_n516_ );
and g346 ( new_n518_, new_n517_, new_n512_ );
or g347 ( new_n519_, new_n518_, keyIn_0_19 );
not g348 ( new_n520_, keyIn_0_19 );
or g349 ( new_n521_, new_n516_, new_n520_, N8 );
and g350 ( new_n522_, new_n519_, new_n521_ );
and g351 ( new_n523_, new_n511_, new_n509_, new_n522_ );
not g352 ( new_n524_, new_n523_ );
and g353 ( new_n525_, new_n524_, keyIn_0_58 );
not g354 ( new_n526_, keyIn_0_58 );
and g355 ( new_n527_, new_n523_, new_n526_ );
or g356 ( new_n528_, new_n525_, new_n527_ );
and g357 ( new_n529_, new_n452_, new_n477_, new_n502_, new_n528_ );
and g358 ( new_n530_, new_n529_, new_n371_, keyIn_0_76, new_n426_ );
not g359 ( new_n531_, new_n530_ );
and g360 ( new_n532_, new_n529_, new_n371_, new_n426_ );
or g361 ( new_n533_, new_n532_, keyIn_0_76 );
and g362 ( new_n534_, new_n533_, new_n531_ );
not g363 ( N329, new_n534_ );
not g364 ( new_n536_, keyIn_0_107 );
not g365 ( new_n537_, keyIn_0_90 );
not g366 ( new_n538_, keyIn_0_86 );
and g367 ( new_n539_, new_n533_, new_n538_, new_n531_ );
not g368 ( new_n540_, new_n539_ );
or g369 ( new_n541_, new_n534_, new_n538_ );
and g370 ( new_n542_, new_n541_, new_n540_ );
or g371 ( new_n543_, new_n542_, new_n452_ );
and g372 ( new_n544_, new_n541_, new_n452_, new_n540_ );
not g373 ( new_n545_, new_n544_ );
and g374 ( new_n546_, new_n543_, new_n537_, new_n545_ );
not g375 ( new_n547_, new_n546_ );
and g376 ( new_n548_, new_n543_, new_n545_ );
or g377 ( new_n549_, new_n548_, new_n537_ );
not g378 ( new_n550_, keyIn_0_79 );
not g379 ( new_n551_, keyIn_0_69 );
not g380 ( new_n552_, keyIn_0_32 );
not g381 ( new_n553_, N40 );
and g382 ( new_n554_, new_n440_, new_n553_, new_n441_ );
not g383 ( new_n555_, new_n554_ );
and g384 ( new_n556_, new_n555_, new_n552_ );
and g385 ( new_n557_, new_n554_, keyIn_0_32 );
or g386 ( new_n558_, new_n556_, new_n557_ );
and g387 ( new_n559_, new_n436_, new_n558_ );
and g388 ( new_n560_, new_n559_, new_n551_ );
not g389 ( new_n561_, new_n560_ );
or g390 ( new_n562_, new_n559_, new_n551_ );
and g391 ( new_n563_, new_n561_, new_n562_ );
and g392 ( new_n564_, new_n563_, new_n550_ );
not g393 ( new_n565_, new_n563_ );
and g394 ( new_n566_, new_n565_, keyIn_0_79 );
or g395 ( new_n567_, new_n566_, new_n564_ );
and g396 ( new_n568_, new_n549_, new_n547_, new_n567_ );
not g397 ( new_n569_, new_n568_ );
and g398 ( new_n570_, new_n569_, keyIn_0_100 );
not g399 ( new_n571_, keyIn_0_100 );
and g400 ( new_n572_, new_n568_, new_n571_ );
or g401 ( new_n573_, new_n570_, new_n572_ );
or g402 ( new_n574_, new_n542_, new_n528_ );
and g403 ( new_n575_, new_n541_, new_n528_, new_n540_ );
not g404 ( new_n576_, new_n575_ );
and g405 ( new_n577_, new_n574_, keyIn_0_88, new_n576_ );
not g406 ( new_n578_, new_n577_ );
and g407 ( new_n579_, new_n574_, new_n576_ );
or g408 ( new_n580_, new_n579_, keyIn_0_88 );
not g409 ( new_n581_, keyIn_0_77 );
or g410 ( new_n582_, new_n516_, N14 );
or g411 ( new_n583_, new_n582_, keyIn_0_20 );
not g412 ( new_n584_, keyIn_0_20 );
not g413 ( new_n585_, new_n582_ );
or g414 ( new_n586_, new_n585_, new_n584_ );
and g415 ( new_n587_, new_n511_, new_n509_, new_n583_, new_n586_ );
or g416 ( new_n588_, new_n587_, keyIn_0_59 );
and g417 ( new_n589_, new_n587_, keyIn_0_59 );
not g418 ( new_n590_, new_n589_ );
and g419 ( new_n591_, new_n590_, new_n588_ );
not g420 ( new_n592_, new_n591_ );
and g421 ( new_n593_, new_n592_, new_n581_ );
and g422 ( new_n594_, new_n591_, keyIn_0_77 );
or g423 ( new_n595_, new_n593_, new_n594_ );
and g424 ( new_n596_, new_n580_, new_n578_, new_n595_ );
not g425 ( new_n597_, new_n596_ );
and g426 ( new_n598_, new_n597_, keyIn_0_98 );
not g427 ( new_n599_, keyIn_0_98 );
and g428 ( new_n600_, new_n596_, new_n599_ );
or g429 ( new_n601_, new_n598_, new_n600_ );
not g430 ( new_n602_, keyIn_0_102 );
or g431 ( new_n603_, new_n542_, new_n316_ );
and g432 ( new_n604_, new_n542_, new_n316_ );
not g433 ( new_n605_, new_n604_ );
and g434 ( new_n606_, new_n605_, keyIn_0_92, new_n603_ );
not g435 ( new_n607_, new_n606_ );
and g436 ( new_n608_, new_n605_, new_n603_ );
or g437 ( new_n609_, new_n608_, keyIn_0_92 );
not g438 ( new_n610_, keyIn_0_81 );
not g439 ( new_n611_, keyIn_0_71 );
or g440 ( new_n612_, new_n305_, N66 );
not g441 ( new_n613_, new_n612_ );
or g442 ( new_n614_, new_n613_, keyIn_0_36 );
not g443 ( new_n615_, keyIn_0_36 );
or g444 ( new_n616_, new_n612_, new_n615_ );
and g445 ( new_n617_, new_n300_, new_n298_, new_n614_, new_n616_ );
and g446 ( new_n618_, new_n617_, new_n611_ );
not g447 ( new_n619_, new_n618_ );
or g448 ( new_n620_, new_n617_, new_n611_ );
and g449 ( new_n621_, new_n619_, new_n620_ );
and g450 ( new_n622_, new_n621_, new_n610_ );
not g451 ( new_n623_, new_n621_ );
and g452 ( new_n624_, new_n623_, keyIn_0_81 );
or g453 ( new_n625_, new_n624_, new_n622_ );
and g454 ( new_n626_, new_n609_, new_n602_, new_n607_, new_n625_ );
not g455 ( new_n627_, new_n626_ );
and g456 ( new_n628_, new_n609_, new_n607_, new_n625_ );
or g457 ( new_n629_, new_n628_, new_n602_ );
and g458 ( new_n630_, new_n629_, new_n627_ );
and g459 ( new_n631_, new_n573_, new_n601_, new_n630_ );
not g460 ( new_n632_, keyIn_0_89 );
not g461 ( new_n633_, new_n502_ );
or g462 ( new_n634_, new_n542_, new_n633_ );
and g463 ( new_n635_, new_n542_, new_n633_ );
not g464 ( new_n636_, new_n635_ );
and g465 ( new_n637_, new_n636_, new_n634_ );
and g466 ( new_n638_, new_n637_, new_n632_ );
not g467 ( new_n639_, new_n634_ );
or g468 ( new_n640_, new_n639_, new_n635_ );
and g469 ( new_n641_, new_n640_, keyIn_0_89 );
or g470 ( new_n642_, new_n641_, new_n638_ );
not g471 ( new_n643_, new_n642_ );
or g472 ( new_n644_, new_n491_, N27 );
or g473 ( new_n645_, new_n644_, keyIn_0_30 );
not g474 ( new_n646_, keyIn_0_30 );
not g475 ( new_n647_, new_n644_ );
or g476 ( new_n648_, new_n647_, new_n646_ );
and g477 ( new_n649_, new_n486_, new_n484_, new_n645_, new_n648_ );
or g478 ( new_n650_, new_n649_, keyIn_0_68 );
and g479 ( new_n651_, new_n649_, keyIn_0_68 );
not g480 ( new_n652_, new_n651_ );
and g481 ( new_n653_, new_n652_, new_n650_ );
or g482 ( new_n654_, new_n653_, keyIn_0_78 );
and g483 ( new_n655_, new_n653_, keyIn_0_78 );
not g484 ( new_n656_, new_n655_ );
and g485 ( new_n657_, new_n656_, new_n654_ );
or g486 ( new_n658_, new_n643_, keyIn_0_99, new_n657_ );
not g487 ( new_n659_, keyIn_0_91 );
not g488 ( new_n660_, new_n477_ );
or g489 ( new_n661_, new_n542_, new_n660_ );
and g490 ( new_n662_, new_n542_, new_n660_ );
not g491 ( new_n663_, new_n662_ );
and g492 ( new_n664_, new_n663_, new_n661_ );
and g493 ( new_n665_, new_n664_, new_n659_ );
not g494 ( new_n666_, new_n542_ );
and g495 ( new_n667_, new_n666_, new_n477_ );
or g496 ( new_n668_, new_n667_, new_n662_ );
and g497 ( new_n669_, new_n668_, keyIn_0_91 );
or g498 ( new_n670_, new_n669_, new_n665_ );
not g499 ( new_n671_, new_n670_ );
not g500 ( new_n672_, keyIn_0_70 );
not g501 ( new_n673_, keyIn_0_34 );
or g502 ( new_n674_, new_n466_, N53 );
not g503 ( new_n675_, new_n674_ );
and g504 ( new_n676_, new_n675_, new_n673_ );
and g505 ( new_n677_, new_n674_, keyIn_0_34 );
or g506 ( new_n678_, new_n676_, new_n677_ );
and g507 ( new_n679_, new_n459_, new_n460_, new_n678_ );
and g508 ( new_n680_, new_n679_, new_n672_ );
not g509 ( new_n681_, new_n680_ );
or g510 ( new_n682_, new_n679_, new_n672_ );
and g511 ( new_n683_, new_n681_, new_n682_ );
or g512 ( new_n684_, new_n683_, keyIn_0_80 );
and g513 ( new_n685_, new_n683_, keyIn_0_80 );
not g514 ( new_n686_, new_n685_ );
and g515 ( new_n687_, new_n686_, new_n684_ );
or g516 ( new_n688_, new_n671_, keyIn_0_101, new_n687_ );
not g517 ( new_n689_, keyIn_0_99 );
not g518 ( new_n690_, new_n657_ );
and g519 ( new_n691_, new_n642_, new_n690_ );
or g520 ( new_n692_, new_n691_, new_n689_ );
not g521 ( new_n693_, keyIn_0_101 );
not g522 ( new_n694_, new_n687_ );
and g523 ( new_n695_, new_n670_, new_n694_ );
or g524 ( new_n696_, new_n695_, new_n693_ );
and g525 ( new_n697_, new_n692_, new_n696_, new_n658_, new_n688_ );
not g526 ( new_n698_, keyIn_0_105 );
or g527 ( new_n699_, new_n542_, new_n425_ );
and g528 ( new_n700_, new_n541_, new_n425_, new_n540_ );
not g529 ( new_n701_, new_n700_ );
and g530 ( new_n702_, new_n699_, new_n701_ );
or g531 ( new_n703_, new_n702_, keyIn_0_96 );
not g532 ( new_n704_, keyIn_0_84 );
not g533 ( new_n705_, keyIn_0_74 );
not g534 ( new_n706_, keyIn_0_42 );
or g535 ( new_n707_, new_n414_, N105 );
and g536 ( new_n708_, new_n707_, new_n706_ );
not g537 ( new_n709_, new_n707_ );
and g538 ( new_n710_, new_n709_, keyIn_0_42 );
or g539 ( new_n711_, new_n710_, new_n708_ );
and g540 ( new_n712_, new_n408_, new_n406_, new_n711_ );
and g541 ( new_n713_, new_n712_, new_n705_ );
not g542 ( new_n714_, new_n713_ );
or g543 ( new_n715_, new_n712_, new_n705_ );
and g544 ( new_n716_, new_n714_, new_n715_ );
and g545 ( new_n717_, new_n716_, new_n704_ );
not g546 ( new_n718_, new_n717_ );
or g547 ( new_n719_, new_n716_, new_n704_ );
and g548 ( new_n720_, new_n718_, new_n719_ );
not g549 ( new_n721_, new_n720_ );
and g550 ( new_n722_, new_n699_, keyIn_0_96, new_n701_ );
not g551 ( new_n723_, new_n722_ );
and g552 ( new_n724_, new_n703_, new_n721_, new_n723_ );
or g553 ( new_n725_, new_n724_, new_n698_ );
not g554 ( new_n726_, keyIn_0_103 );
and g555 ( new_n727_, new_n541_, new_n370_, new_n540_ );
not g556 ( new_n728_, new_n727_ );
or g557 ( new_n729_, new_n542_, new_n370_ );
and g558 ( new_n730_, new_n729_, keyIn_0_93, new_n728_ );
not g559 ( new_n731_, new_n730_ );
and g560 ( new_n732_, new_n729_, new_n728_ );
or g561 ( new_n733_, new_n732_, keyIn_0_93 );
and g562 ( new_n734_, new_n733_, new_n731_ );
not g563 ( new_n735_, keyIn_0_82 );
not g564 ( new_n736_, keyIn_0_72 );
or g565 ( new_n737_, new_n359_, N79 );
not g566 ( new_n738_, new_n737_ );
or g567 ( new_n739_, new_n738_, keyIn_0_38 );
not g568 ( new_n740_, keyIn_0_38 );
or g569 ( new_n741_, new_n737_, new_n740_ );
and g570 ( new_n742_, new_n353_, new_n354_, new_n739_, new_n741_ );
and g571 ( new_n743_, new_n742_, new_n736_ );
not g572 ( new_n744_, new_n743_ );
or g573 ( new_n745_, new_n742_, new_n736_ );
and g574 ( new_n746_, new_n744_, new_n745_ );
and g575 ( new_n747_, new_n746_, new_n735_ );
not g576 ( new_n748_, new_n747_ );
or g577 ( new_n749_, new_n746_, new_n735_ );
and g578 ( new_n750_, new_n748_, new_n749_ );
or g579 ( new_n751_, new_n734_, new_n726_, new_n750_ );
not g580 ( new_n752_, keyIn_0_104 );
and g581 ( new_n753_, new_n399_, new_n401_ );
or g582 ( new_n754_, new_n542_, new_n753_ );
not g583 ( new_n755_, new_n754_ );
and g584 ( new_n756_, new_n542_, new_n753_ );
or g585 ( new_n757_, new_n755_, new_n756_ );
and g586 ( new_n758_, new_n757_, keyIn_0_94 );
not g587 ( new_n759_, keyIn_0_94 );
not g588 ( new_n760_, new_n756_ );
and g589 ( new_n761_, new_n760_, new_n759_, new_n754_ );
not g590 ( new_n762_, keyIn_0_83 );
not g591 ( new_n763_, keyIn_0_73 );
not g592 ( new_n764_, keyIn_0_40 );
or g593 ( new_n765_, new_n390_, N92 );
not g594 ( new_n766_, new_n765_ );
and g595 ( new_n767_, new_n766_, new_n764_ );
and g596 ( new_n768_, new_n765_, keyIn_0_40 );
or g597 ( new_n769_, new_n767_, new_n768_ );
and g598 ( new_n770_, new_n384_, new_n769_ );
and g599 ( new_n771_, new_n770_, new_n763_ );
not g600 ( new_n772_, new_n771_ );
or g601 ( new_n773_, new_n770_, new_n763_ );
and g602 ( new_n774_, new_n772_, new_n773_ );
and g603 ( new_n775_, new_n774_, new_n762_ );
not g604 ( new_n776_, new_n775_ );
or g605 ( new_n777_, new_n774_, new_n762_ );
and g606 ( new_n778_, new_n776_, new_n777_ );
or g607 ( new_n779_, new_n758_, new_n752_, new_n761_, new_n778_ );
not g608 ( new_n780_, new_n703_ );
or g609 ( new_n781_, new_n780_, keyIn_0_105, new_n720_, new_n722_ );
and g610 ( new_n782_, new_n751_, new_n725_, new_n779_, new_n781_ );
not g611 ( new_n783_, new_n734_ );
not g612 ( new_n784_, new_n750_ );
and g613 ( new_n785_, new_n783_, new_n784_ );
or g614 ( new_n786_, new_n785_, keyIn_0_103 );
not g615 ( new_n787_, new_n758_ );
not g616 ( new_n788_, new_n761_ );
not g617 ( new_n789_, new_n778_ );
and g618 ( new_n790_, new_n787_, new_n788_, new_n789_ );
or g619 ( new_n791_, new_n790_, keyIn_0_104 );
not g620 ( new_n792_, keyIn_0_106 );
and g621 ( new_n793_, new_n541_, new_n344_, new_n540_ );
not g622 ( new_n794_, new_n793_ );
or g623 ( new_n795_, new_n542_, new_n344_ );
and g624 ( new_n796_, new_n795_, keyIn_0_97, new_n794_ );
not g625 ( new_n797_, new_n796_ );
and g626 ( new_n798_, new_n795_, new_n794_ );
or g627 ( new_n799_, new_n798_, keyIn_0_97 );
not g628 ( new_n800_, keyIn_0_85 );
not g629 ( new_n801_, keyIn_0_75 );
not g630 ( new_n802_, keyIn_0_44 );
or g631 ( new_n803_, new_n332_, N115 );
not g632 ( new_n804_, new_n803_ );
and g633 ( new_n805_, new_n804_, new_n802_ );
and g634 ( new_n806_, new_n803_, keyIn_0_44 );
or g635 ( new_n807_, new_n805_, new_n806_ );
and g636 ( new_n808_, new_n341_, new_n807_ );
and g637 ( new_n809_, new_n808_, new_n801_ );
not g638 ( new_n810_, new_n809_ );
or g639 ( new_n811_, new_n808_, new_n801_ );
and g640 ( new_n812_, new_n810_, new_n811_ );
and g641 ( new_n813_, new_n812_, new_n800_ );
not g642 ( new_n814_, new_n812_ );
and g643 ( new_n815_, new_n814_, keyIn_0_85 );
or g644 ( new_n816_, new_n815_, new_n813_ );
and g645 ( new_n817_, new_n799_, new_n797_, new_n816_ );
not g646 ( new_n818_, new_n817_ );
and g647 ( new_n819_, new_n818_, new_n792_ );
and g648 ( new_n820_, new_n817_, keyIn_0_106 );
or g649 ( new_n821_, new_n819_, new_n820_ );
and g650 ( new_n822_, new_n821_, new_n782_, new_n786_, new_n791_ );
and g651 ( new_n823_, new_n822_, new_n697_, new_n631_, new_n536_ );
not g652 ( new_n824_, new_n823_ );
or g653 ( new_n825_, new_n758_, new_n752_, new_n761_, new_n778_ );
or g654 ( new_n826_, new_n780_, keyIn_0_105, new_n720_, new_n722_ );
and g655 ( new_n827_, new_n751_, new_n725_, new_n825_, new_n826_ );
and g656 ( new_n828_, new_n821_, new_n827_, new_n786_, new_n791_ );
and g657 ( new_n829_, new_n828_, new_n631_, new_n697_ );
or g658 ( new_n830_, new_n829_, new_n536_ );
and g659 ( N370, new_n830_, new_n824_ );
not g660 ( new_n832_, keyIn_0_120 );
not g661 ( new_n833_, keyIn_0_109 );
and g662 ( new_n834_, new_n830_, keyIn_0_108, new_n824_ );
not g663 ( new_n835_, new_n834_ );
or g664 ( new_n836_, N370, keyIn_0_108 );
and g665 ( new_n837_, new_n836_, N53, new_n835_ );
not g666 ( new_n838_, new_n837_ );
and g667 ( new_n839_, new_n838_, new_n833_ );
not g668 ( new_n840_, keyIn_0_87 );
and g669 ( new_n841_, new_n534_, new_n840_ );
and g670 ( new_n842_, N329, keyIn_0_87 );
or g671 ( new_n843_, new_n842_, new_n841_ );
and g672 ( new_n844_, new_n843_, N47 );
not g673 ( new_n845_, new_n844_ );
and g674 ( new_n846_, new_n845_, keyIn_0_95 );
or g675 ( new_n847_, new_n845_, keyIn_0_95 );
not g676 ( new_n848_, new_n847_ );
not g677 ( new_n849_, keyIn_0_57 );
or g678 ( new_n850_, N223, keyIn_0_47 );
and g679 ( new_n851_, N223, keyIn_0_47 );
not g680 ( new_n852_, new_n851_ );
and g681 ( new_n853_, new_n852_, new_n850_ );
and g682 ( new_n854_, new_n853_, N37 );
and g683 ( new_n855_, new_n854_, new_n849_ );
not g684 ( new_n856_, new_n855_ );
or g685 ( new_n857_, new_n854_, new_n849_ );
and g686 ( new_n858_, new_n856_, new_n857_ );
or g687 ( new_n859_, new_n848_, new_n251_, new_n846_, new_n858_ );
not g688 ( new_n860_, keyIn_0_108 );
and g689 ( new_n861_, new_n822_, new_n631_, new_n697_ );
not g690 ( new_n862_, new_n861_ );
and g691 ( new_n863_, new_n862_, keyIn_0_107 );
or g692 ( new_n864_, new_n863_, new_n860_, new_n823_ );
and g693 ( new_n865_, new_n836_, keyIn_0_109, N53, new_n864_ );
or g694 ( new_n866_, new_n865_, new_n859_ );
or g695 ( new_n867_, new_n839_, new_n866_, keyIn_0_113 );
not g696 ( new_n868_, keyIn_0_113 );
or g697 ( new_n869_, new_n837_, keyIn_0_109 );
not g698 ( new_n870_, new_n859_ );
not g699 ( new_n871_, new_n865_ );
and g700 ( new_n872_, new_n869_, new_n870_, new_n871_ );
or g701 ( new_n873_, new_n872_, new_n868_ );
and g702 ( new_n874_, new_n873_, new_n867_ );
not g703 ( new_n875_, keyIn_0_114 );
and g704 ( new_n876_, new_n836_, N66, new_n864_ );
not g705 ( new_n877_, new_n876_ );
and g706 ( new_n878_, new_n843_, N60 );
and g707 ( new_n879_, new_n853_, N50 );
or g708 ( new_n880_, new_n878_, new_n275_, new_n879_ );
not g709 ( new_n881_, new_n880_ );
and g710 ( new_n882_, new_n877_, new_n875_, new_n881_ );
or g711 ( new_n883_, new_n876_, new_n880_ );
and g712 ( new_n884_, new_n883_, keyIn_0_114 );
or g713 ( new_n885_, new_n884_, new_n882_ );
and g714 ( new_n886_, new_n874_, new_n885_ );
not g715 ( new_n887_, keyIn_0_112 );
and g716 ( new_n888_, new_n836_, N40, new_n864_ );
and g717 ( new_n889_, new_n843_, N34 );
and g718 ( new_n890_, new_n853_, N24 );
or g719 ( new_n891_, new_n889_, new_n233_, new_n890_ );
or g720 ( new_n892_, new_n888_, new_n891_ );
and g721 ( new_n893_, new_n892_, new_n887_ );
not g722 ( new_n894_, new_n888_ );
not g723 ( new_n895_, new_n891_ );
and g724 ( new_n896_, new_n894_, keyIn_0_112, new_n895_ );
or g725 ( new_n897_, new_n893_, new_n896_ );
not g726 ( new_n898_, keyIn_0_111 );
and g727 ( new_n899_, new_n836_, new_n864_ );
and g728 ( new_n900_, new_n899_, N27 );
and g729 ( new_n901_, new_n843_, N21 );
and g730 ( new_n902_, new_n853_, N11 );
or g731 ( new_n903_, new_n901_, new_n220_, new_n902_ );
or g732 ( new_n904_, new_n900_, new_n903_ );
not g733 ( new_n905_, new_n904_ );
and g734 ( new_n906_, new_n905_, new_n898_ );
and g735 ( new_n907_, new_n904_, keyIn_0_111 );
or g736 ( new_n908_, new_n906_, new_n907_ );
and g737 ( new_n909_, new_n908_, new_n897_ );
not g738 ( new_n910_, keyIn_0_117 );
and g739 ( new_n911_, new_n836_, N105, new_n864_ );
not g740 ( new_n912_, new_n911_ );
and g741 ( new_n913_, new_n843_, N99 );
and g742 ( new_n914_, new_n853_, N89 );
or g743 ( new_n915_, new_n913_, new_n186_, new_n914_ );
not g744 ( new_n916_, new_n915_ );
and g745 ( new_n917_, new_n912_, new_n910_, new_n916_ );
not g746 ( new_n918_, new_n917_ );
or g747 ( new_n919_, new_n911_, new_n915_ );
and g748 ( new_n920_, new_n919_, keyIn_0_117 );
not g749 ( new_n921_, new_n920_ );
and g750 ( new_n922_, new_n899_, N115 );
and g751 ( new_n923_, new_n843_, N112 );
and g752 ( new_n924_, new_n853_, N102 );
or g753 ( new_n925_, new_n923_, new_n174_, new_n924_ );
or g754 ( new_n926_, new_n922_, keyIn_0_118, new_n925_ );
not g755 ( new_n927_, keyIn_0_118 );
not g756 ( new_n928_, new_n922_ );
not g757 ( new_n929_, new_n923_ );
not g758 ( new_n930_, new_n924_ );
and g759 ( new_n931_, new_n928_, N108, new_n929_, new_n930_ );
or g760 ( new_n932_, new_n931_, new_n927_ );
and g761 ( new_n933_, new_n932_, new_n918_, new_n921_, new_n926_ );
not g762 ( new_n934_, keyIn_0_115 );
and g763 ( new_n935_, new_n836_, N79, new_n864_ );
not g764 ( new_n936_, new_n935_ );
and g765 ( new_n937_, new_n843_, N73 );
and g766 ( new_n938_, new_n853_, N63 );
or g767 ( new_n939_, new_n937_, new_n263_, new_n938_ );
not g768 ( new_n940_, new_n939_ );
and g769 ( new_n941_, new_n936_, new_n934_, new_n940_ );
not g770 ( new_n942_, new_n941_ );
or g771 ( new_n943_, new_n935_, new_n939_ );
and g772 ( new_n944_, new_n943_, keyIn_0_115 );
not g773 ( new_n945_, new_n944_ );
not g774 ( new_n946_, keyIn_0_116 );
and g775 ( new_n947_, new_n836_, N92, new_n864_ );
and g776 ( new_n948_, new_n843_, N86 );
and g777 ( new_n949_, new_n853_, N76 );
or g778 ( new_n950_, new_n948_, new_n202_, new_n949_ );
or g779 ( new_n951_, new_n947_, new_n950_ );
not g780 ( new_n952_, new_n951_ );
and g781 ( new_n953_, new_n952_, new_n946_ );
not g782 ( new_n954_, new_n953_ );
and g783 ( new_n955_, new_n951_, keyIn_0_116 );
not g784 ( new_n956_, new_n955_ );
and g785 ( new_n957_, new_n954_, new_n942_, new_n945_, new_n956_ );
and g786 ( new_n958_, new_n933_, new_n957_ );
and g787 ( new_n959_, new_n958_, keyIn_0_119, new_n886_, new_n909_ );
not g788 ( new_n960_, new_n959_ );
and g789 ( new_n961_, new_n909_, new_n886_, new_n933_, new_n957_ );
or g790 ( new_n962_, new_n961_, keyIn_0_119 );
not g791 ( new_n963_, keyIn_0_110 );
and g792 ( new_n964_, new_n899_, N14 );
and g793 ( new_n965_, new_n843_, N8 );
and g794 ( new_n966_, new_n853_, N1 );
or g795 ( new_n967_, new_n964_, new_n207_, new_n965_, new_n966_ );
and g796 ( new_n968_, new_n967_, new_n963_ );
not g797 ( new_n969_, new_n967_ );
and g798 ( new_n970_, new_n969_, keyIn_0_110 );
or g799 ( new_n971_, new_n970_, new_n968_ );
and g800 ( new_n972_, new_n962_, new_n960_, new_n971_ );
not g801 ( new_n973_, new_n972_ );
and g802 ( new_n974_, new_n973_, new_n832_ );
and g803 ( new_n975_, new_n972_, keyIn_0_120 );
or g804 ( N421, new_n974_, new_n975_ );
not g805 ( new_n977_, keyIn_0_125 );
not g806 ( new_n978_, keyIn_0_121 );
not g807 ( new_n979_, new_n897_ );
and g808 ( new_n980_, new_n899_, N53 );
or g809 ( new_n981_, new_n980_, keyIn_0_109 );
and g810 ( new_n982_, new_n981_, new_n870_, new_n871_ );
or g811 ( new_n983_, new_n982_, new_n868_ );
and g812 ( new_n984_, new_n983_, new_n867_ );
or g813 ( new_n985_, new_n984_, new_n978_, new_n979_ );
not g814 ( new_n986_, new_n867_ );
or g815 ( new_n987_, new_n839_, new_n866_ );
and g816 ( new_n988_, new_n987_, keyIn_0_113 );
or g817 ( new_n989_, new_n988_, new_n986_ );
and g818 ( new_n990_, new_n989_, new_n897_ );
or g819 ( new_n991_, new_n990_, keyIn_0_121 );
and g820 ( new_n992_, new_n991_, new_n985_ );
and g821 ( new_n993_, new_n909_, new_n885_ );
not g822 ( new_n994_, new_n993_ );
or g823 ( new_n995_, new_n992_, new_n994_ );
and g824 ( new_n996_, new_n995_, new_n977_ );
not g825 ( new_n997_, new_n992_ );
and g826 ( new_n998_, new_n997_, keyIn_0_125, new_n993_ );
or g827 ( N430, new_n996_, new_n998_ );
not g828 ( new_n1000_, keyIn_0_126 );
not g829 ( new_n1001_, new_n908_ );
and g830 ( new_n1002_, new_n873_, new_n867_, new_n897_ );
or g831 ( new_n1003_, new_n944_, new_n941_ );
and g832 ( new_n1004_, new_n885_, new_n1003_ );
and g833 ( new_n1005_, new_n1002_, new_n1004_ );
not g834 ( new_n1006_, new_n1005_ );
and g835 ( new_n1007_, new_n1006_, keyIn_0_122 );
not g836 ( new_n1008_, keyIn_0_122 );
and g837 ( new_n1009_, new_n897_, new_n1008_ );
and g838 ( new_n1010_, new_n984_, new_n1004_, new_n1009_ );
or g839 ( new_n1011_, new_n1007_, new_n1010_ );
not g840 ( new_n1012_, keyIn_0_123 );
or g841 ( new_n1013_, new_n953_, new_n955_ );
and g842 ( new_n1014_, new_n874_, new_n885_, new_n1013_ );
or g843 ( new_n1015_, new_n1014_, new_n1012_ );
and g844 ( new_n1016_, new_n1013_, new_n1012_, new_n885_ );
and g845 ( new_n1017_, new_n984_, new_n1016_ );
not g846 ( new_n1018_, new_n1017_ );
and g847 ( new_n1019_, new_n1018_, new_n1015_ );
or g848 ( new_n1020_, new_n1011_, new_n1019_, new_n979_, new_n1001_ );
and g849 ( new_n1021_, new_n1020_, new_n1000_ );
not g850 ( new_n1022_, new_n1011_ );
not g851 ( new_n1023_, new_n1019_ );
and g852 ( new_n1024_, new_n1022_, keyIn_0_126, new_n909_, new_n1023_ );
or g853 ( N431, new_n1021_, new_n1024_ );
not g854 ( new_n1026_, keyIn_0_127 );
not g855 ( new_n1027_, keyIn_0_124 );
or g856 ( new_n1028_, new_n920_, new_n917_ );
and g857 ( new_n1029_, new_n1028_, new_n954_, new_n956_ );
and g858 ( new_n1030_, new_n1002_, new_n1027_, new_n1029_ );
not g859 ( new_n1031_, new_n1030_ );
and g860 ( new_n1032_, new_n1002_, new_n1029_ );
or g861 ( new_n1033_, new_n1032_, new_n1027_ );
and g862 ( new_n1034_, new_n1033_, new_n1031_ );
not g863 ( new_n1035_, new_n1034_ );
and g864 ( new_n1036_, new_n997_, new_n908_ );
and g865 ( new_n1037_, new_n1036_, new_n1026_, new_n1022_, new_n1035_ );
or g866 ( new_n1038_, new_n1011_, new_n992_, new_n1034_, new_n1001_ );
and g867 ( new_n1039_, new_n1038_, keyIn_0_127 );
or g868 ( N432, new_n1039_, new_n1037_ );
endmodule