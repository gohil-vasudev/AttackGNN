module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n246_, new_n170_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n562_, new_n578_, new_n177_, new_n493_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n148_, new_n662_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n405_;

not g000 ( new_n138_, keyIn_0_38 );
not g001 ( new_n139_, keyIn_0_30 );
not g002 ( new_n140_, keyIn_0_26 );
xnor g003 ( new_n141_, N65, N69 );
nand g004 ( new_n142_, new_n141_, keyIn_0_5 );
not g005 ( new_n143_, keyIn_0_5 );
or g006 ( new_n144_, N65, N69 );
nand g007 ( new_n145_, N65, N69 );
nand g008 ( new_n146_, new_n144_, new_n143_, new_n145_ );
nand g009 ( new_n147_, new_n142_, new_n146_ );
xnor g010 ( new_n148_, N73, N77 );
xnor g011 ( new_n149_, new_n147_, new_n148_ );
xnor g012 ( new_n150_, new_n149_, keyIn_0_10 );
xor g013 ( new_n151_, N81, N85 );
xnor g014 ( new_n152_, N89, N93 );
xnor g015 ( new_n153_, new_n151_, new_n152_ );
xnor g016 ( new_n154_, new_n153_, keyIn_0_11 );
nand g017 ( new_n155_, new_n150_, new_n154_ );
not g018 ( new_n156_, keyIn_0_10 );
xnor g019 ( new_n157_, new_n149_, new_n156_ );
not g020 ( new_n158_, keyIn_0_11 );
xnor g021 ( new_n159_, new_n153_, new_n158_ );
nand g022 ( new_n160_, new_n157_, new_n159_ );
nand g023 ( new_n161_, new_n155_, new_n160_ );
nand g024 ( new_n162_, new_n161_, new_n140_ );
nand g025 ( new_n163_, new_n155_, new_n160_, keyIn_0_26 );
nand g026 ( new_n164_, new_n162_, new_n163_ );
nand g027 ( new_n165_, N129, N137 );
nand g028 ( new_n166_, new_n164_, new_n165_ );
nand g029 ( new_n167_, new_n162_, N129, N137, new_n163_ );
nand g030 ( new_n168_, new_n166_, new_n167_ );
nand g031 ( new_n169_, new_n168_, new_n139_ );
nand g032 ( new_n170_, new_n166_, keyIn_0_30, new_n167_ );
nand g033 ( new_n171_, new_n169_, new_n170_ );
xor g034 ( new_n172_, N1, N17 );
xnor g035 ( new_n173_, N33, N49 );
xnor g036 ( new_n174_, new_n172_, new_n173_ );
xor g037 ( new_n175_, new_n174_, keyIn_0_14 );
not g038 ( new_n176_, new_n175_ );
nand g039 ( new_n177_, new_n171_, new_n176_ );
nand g040 ( new_n178_, new_n169_, new_n170_, new_n175_ );
nand g041 ( new_n179_, new_n177_, new_n178_ );
nand g042 ( new_n180_, new_n179_, new_n138_ );
nand g043 ( new_n181_, new_n177_, keyIn_0_38, new_n178_ );
nand g044 ( new_n182_, new_n180_, new_n181_ );
not g045 ( new_n183_, new_n182_ );
not g046 ( new_n184_, keyIn_0_56 );
not g047 ( new_n185_, keyIn_0_54 );
not g048 ( new_n186_, keyIn_0_32 );
not g049 ( new_n187_, keyIn_0_12 );
xnor g050 ( new_n188_, N105, N109 );
xor g051 ( new_n189_, N97, N101 );
xnor g052 ( new_n190_, new_n189_, new_n188_ );
xnor g053 ( new_n191_, new_n190_, new_n187_ );
nand g054 ( new_n192_, new_n150_, new_n191_ );
xnor g055 ( new_n193_, new_n190_, keyIn_0_12 );
nand g056 ( new_n194_, new_n157_, new_n193_ );
nand g057 ( new_n195_, new_n192_, new_n194_ );
nand g058 ( new_n196_, new_n195_, keyIn_0_28 );
not g059 ( new_n197_, keyIn_0_28 );
nand g060 ( new_n198_, new_n192_, new_n194_, new_n197_ );
nand g061 ( new_n199_, new_n196_, new_n198_ );
nand g062 ( new_n200_, N131, N137 );
nand g063 ( new_n201_, new_n199_, new_n200_ );
nand g064 ( new_n202_, new_n196_, N131, N137, new_n198_ );
nand g065 ( new_n203_, new_n201_, new_n202_ );
nand g066 ( new_n204_, new_n203_, new_n186_ );
nand g067 ( new_n205_, new_n201_, keyIn_0_32, new_n202_ );
nand g068 ( new_n206_, new_n204_, new_n205_ );
xor g069 ( new_n207_, N9, N25 );
xnor g070 ( new_n208_, N41, N57 );
xnor g071 ( new_n209_, new_n207_, new_n208_ );
xnor g072 ( new_n210_, new_n209_, keyIn_0_16 );
not g073 ( new_n211_, new_n210_ );
nand g074 ( new_n212_, new_n206_, new_n211_ );
nand g075 ( new_n213_, new_n204_, new_n205_, new_n210_ );
nand g076 ( new_n214_, new_n212_, new_n213_ );
nand g077 ( new_n215_, new_n214_, keyIn_0_40 );
not g078 ( new_n216_, keyIn_0_40 );
nand g079 ( new_n217_, new_n212_, new_n216_, new_n213_ );
nand g080 ( new_n218_, new_n215_, new_n217_ );
not g081 ( new_n219_, keyIn_0_41 );
not g082 ( new_n220_, keyIn_0_33 );
xor g083 ( new_n221_, N113, N117 );
xnor g084 ( new_n222_, N121, N125 );
xnor g085 ( new_n223_, new_n221_, new_n222_ );
xnor g086 ( new_n224_, new_n223_, keyIn_0_13 );
nand g087 ( new_n225_, new_n154_, new_n224_ );
not g088 ( new_n226_, keyIn_0_13 );
xnor g089 ( new_n227_, new_n223_, new_n226_ );
nand g090 ( new_n228_, new_n159_, new_n227_ );
nand g091 ( new_n229_, new_n225_, new_n228_ );
nand g092 ( new_n230_, new_n229_, keyIn_0_29 );
not g093 ( new_n231_, keyIn_0_29 );
nand g094 ( new_n232_, new_n225_, new_n228_, new_n231_ );
nand g095 ( new_n233_, new_n230_, new_n232_ );
nand g096 ( new_n234_, N132, N137 );
nand g097 ( new_n235_, new_n233_, new_n234_ );
nand g098 ( new_n236_, new_n230_, N132, N137, new_n232_ );
nand g099 ( new_n237_, new_n235_, new_n236_ );
nand g100 ( new_n238_, new_n237_, new_n220_ );
nand g101 ( new_n239_, new_n235_, keyIn_0_33, new_n236_ );
nand g102 ( new_n240_, new_n238_, new_n239_ );
xor g103 ( new_n241_, N13, N29 );
xnor g104 ( new_n242_, N45, N61 );
xnor g105 ( new_n243_, new_n241_, new_n242_ );
xor g106 ( new_n244_, new_n243_, keyIn_0_17 );
not g107 ( new_n245_, new_n244_ );
nand g108 ( new_n246_, new_n240_, new_n245_ );
nand g109 ( new_n247_, new_n238_, new_n239_, new_n244_ );
nand g110 ( new_n248_, new_n246_, new_n247_ );
xnor g111 ( new_n249_, new_n248_, new_n219_ );
not g112 ( new_n250_, keyIn_0_39 );
not g113 ( new_n251_, keyIn_0_31 );
not g114 ( new_n252_, keyIn_0_27 );
nand g115 ( new_n253_, new_n193_, new_n227_ );
nand g116 ( new_n254_, new_n191_, new_n224_ );
nand g117 ( new_n255_, new_n253_, new_n254_ );
nand g118 ( new_n256_, new_n255_, new_n252_ );
nand g119 ( new_n257_, new_n253_, new_n254_, keyIn_0_27 );
nand g120 ( new_n258_, new_n256_, new_n257_ );
nand g121 ( new_n259_, N130, N137 );
nand g122 ( new_n260_, new_n258_, new_n259_ );
nand g123 ( new_n261_, new_n256_, N130, N137, new_n257_ );
nand g124 ( new_n262_, new_n260_, new_n261_ );
nand g125 ( new_n263_, new_n262_, new_n251_ );
nand g126 ( new_n264_, new_n260_, keyIn_0_31, new_n261_ );
nand g127 ( new_n265_, new_n263_, new_n264_ );
xor g128 ( new_n266_, N5, N21 );
xnor g129 ( new_n267_, N37, N53 );
xnor g130 ( new_n268_, new_n266_, new_n267_ );
xnor g131 ( new_n269_, new_n268_, keyIn_0_15 );
not g132 ( new_n270_, new_n269_ );
nand g133 ( new_n271_, new_n265_, new_n270_ );
nand g134 ( new_n272_, new_n263_, new_n264_, new_n269_ );
nand g135 ( new_n273_, new_n271_, new_n272_ );
xnor g136 ( new_n274_, new_n273_, new_n250_ );
not g137 ( new_n275_, new_n274_ );
nand g138 ( new_n276_, new_n182_, new_n218_, new_n275_, new_n249_ );
xnor g139 ( new_n277_, new_n276_, keyIn_0_48 );
xnor g140 ( new_n278_, new_n248_, keyIn_0_41 );
nand g141 ( new_n279_, new_n182_, new_n218_, new_n278_, new_n274_ );
xnor g142 ( new_n280_, new_n279_, keyIn_0_46 );
not g143 ( new_n281_, keyIn_0_47 );
and g144 ( new_n282_, new_n215_, new_n217_ );
nand g145 ( new_n283_, new_n282_, new_n182_, new_n249_, new_n274_ );
nand g146 ( new_n284_, new_n283_, new_n281_ );
nor g147 ( new_n285_, new_n218_, new_n278_ );
nand g148 ( new_n286_, new_n285_, keyIn_0_47, new_n182_, new_n274_ );
nand g149 ( new_n287_, new_n284_, new_n286_ );
and g150 ( new_n288_, new_n280_, new_n287_ );
nand g151 ( new_n289_, new_n274_, new_n249_, new_n180_, new_n181_ );
nor g152 ( new_n290_, new_n289_, new_n282_ );
xnor g153 ( new_n291_, new_n290_, keyIn_0_49 );
nand g154 ( new_n292_, new_n288_, new_n185_, new_n277_, new_n291_ );
nand g155 ( new_n293_, new_n291_, new_n277_, new_n280_, new_n287_ );
nand g156 ( new_n294_, new_n293_, keyIn_0_54 );
not g157 ( new_n295_, keyIn_0_45 );
not g158 ( new_n296_, keyIn_0_37 );
not g159 ( new_n297_, keyIn_0_25 );
not g160 ( new_n298_, N29 );
nand g161 ( new_n299_, new_n298_, N25 );
not g162 ( new_n300_, N25 );
nand g163 ( new_n301_, new_n300_, N29 );
nand g164 ( new_n302_, new_n299_, new_n301_ );
nand g165 ( new_n303_, new_n302_, keyIn_0_0 );
not g166 ( new_n304_, keyIn_0_0 );
nand g167 ( new_n305_, new_n299_, new_n301_, new_n304_ );
nand g168 ( new_n306_, new_n303_, new_n305_ );
xor g169 ( new_n307_, N17, N21 );
nand g170 ( new_n308_, new_n306_, new_n307_ );
not g171 ( new_n309_, new_n307_ );
nand g172 ( new_n310_, new_n309_, new_n303_, new_n305_ );
nand g173 ( new_n311_, new_n308_, new_n310_ );
nand g174 ( new_n312_, new_n311_, keyIn_0_7 );
not g175 ( new_n313_, keyIn_0_7 );
nand g176 ( new_n314_, new_n308_, new_n313_, new_n310_ );
nand g177 ( new_n315_, new_n312_, new_n314_ );
not g178 ( new_n316_, new_n315_ );
xor g179 ( new_n317_, N57, N61 );
nand g180 ( new_n318_, new_n317_, keyIn_0_4 );
not g181 ( new_n319_, keyIn_0_4 );
xnor g182 ( new_n320_, N57, N61 );
nand g183 ( new_n321_, new_n320_, new_n319_ );
nand g184 ( new_n322_, new_n318_, new_n321_ );
xnor g185 ( new_n323_, N49, N53 );
xnor g186 ( new_n324_, new_n323_, keyIn_0_3 );
nand g187 ( new_n325_, new_n324_, new_n322_ );
not g188 ( new_n326_, N53 );
nand g189 ( new_n327_, new_n326_, N49 );
not g190 ( new_n328_, N49 );
nand g191 ( new_n329_, new_n328_, N53 );
nand g192 ( new_n330_, new_n327_, new_n329_ );
nand g193 ( new_n331_, new_n330_, keyIn_0_3 );
not g194 ( new_n332_, keyIn_0_3 );
nand g195 ( new_n333_, new_n323_, new_n332_ );
nand g196 ( new_n334_, new_n331_, new_n333_ );
nand g197 ( new_n335_, new_n334_, new_n318_, new_n321_ );
nand g198 ( new_n336_, new_n325_, new_n335_ );
nand g199 ( new_n337_, new_n336_, keyIn_0_9 );
not g200 ( new_n338_, keyIn_0_9 );
nand g201 ( new_n339_, new_n325_, new_n335_, new_n338_ );
nand g202 ( new_n340_, new_n337_, new_n339_ );
nand g203 ( new_n341_, new_n316_, new_n340_ );
nand g204 ( new_n342_, new_n315_, new_n337_, new_n339_ );
nand g205 ( new_n343_, new_n341_, new_n342_ );
nand g206 ( new_n344_, new_n343_, new_n297_ );
nand g207 ( new_n345_, new_n341_, keyIn_0_25, new_n342_ );
nand g208 ( new_n346_, new_n344_, new_n345_ );
nand g209 ( new_n347_, N136, N137 );
not g210 ( new_n348_, new_n347_ );
nand g211 ( new_n349_, new_n346_, new_n348_ );
nand g212 ( new_n350_, new_n344_, new_n345_, new_n347_ );
nand g213 ( new_n351_, new_n349_, new_n350_ );
nand g214 ( new_n352_, new_n351_, new_n296_ );
nand g215 ( new_n353_, new_n349_, keyIn_0_37, new_n350_ );
nand g216 ( new_n354_, new_n352_, new_n353_ );
xor g217 ( new_n355_, N77, N93 );
xnor g218 ( new_n356_, N109, N125 );
xnor g219 ( new_n357_, new_n355_, new_n356_ );
xnor g220 ( new_n358_, new_n357_, keyIn_0_21 );
nand g221 ( new_n359_, new_n354_, new_n358_ );
not g222 ( new_n360_, new_n358_ );
nand g223 ( new_n361_, new_n352_, new_n353_, new_n360_ );
nand g224 ( new_n362_, new_n359_, new_n361_ );
nand g225 ( new_n363_, new_n362_, new_n295_ );
nand g226 ( new_n364_, new_n359_, keyIn_0_45, new_n361_ );
nand g227 ( new_n365_, new_n363_, new_n364_ );
not g228 ( new_n366_, keyIn_0_44 );
not g229 ( new_n367_, keyIn_0_24 );
xnor g230 ( new_n368_, N1, N5 );
xnor g231 ( new_n369_, N9, N13 );
xnor g232 ( new_n370_, new_n368_, new_n369_ );
xnor g233 ( new_n371_, new_n370_, keyIn_0_6 );
not g234 ( new_n372_, keyIn_0_8 );
not g235 ( new_n373_, N37 );
nand g236 ( new_n374_, new_n373_, N33 );
not g237 ( new_n375_, N33 );
nand g238 ( new_n376_, new_n375_, N37 );
nand g239 ( new_n377_, new_n374_, new_n376_ );
nand g240 ( new_n378_, new_n377_, keyIn_0_1 );
not g241 ( new_n379_, keyIn_0_1 );
nand g242 ( new_n380_, new_n374_, new_n376_, new_n379_ );
nand g243 ( new_n381_, new_n378_, new_n380_ );
not g244 ( new_n382_, keyIn_0_2 );
not g245 ( new_n383_, N45 );
nand g246 ( new_n384_, new_n383_, N41 );
not g247 ( new_n385_, N41 );
nand g248 ( new_n386_, new_n385_, N45 );
nand g249 ( new_n387_, new_n384_, new_n386_ );
nand g250 ( new_n388_, new_n387_, new_n382_ );
nand g251 ( new_n389_, new_n384_, new_n386_, keyIn_0_2 );
nand g252 ( new_n390_, new_n388_, new_n389_ );
nand g253 ( new_n391_, new_n381_, new_n390_ );
nand g254 ( new_n392_, new_n378_, new_n388_, new_n380_, new_n389_ );
nand g255 ( new_n393_, new_n391_, new_n392_ );
nand g256 ( new_n394_, new_n393_, new_n372_ );
nand g257 ( new_n395_, new_n391_, keyIn_0_8, new_n392_ );
nand g258 ( new_n396_, new_n394_, new_n395_ );
nand g259 ( new_n397_, new_n396_, new_n371_ );
not g260 ( new_n398_, keyIn_0_6 );
xnor g261 ( new_n399_, new_n370_, new_n398_ );
nand g262 ( new_n400_, new_n399_, new_n394_, new_n395_ );
nand g263 ( new_n401_, new_n397_, new_n400_ );
nand g264 ( new_n402_, new_n401_, new_n367_ );
nand g265 ( new_n403_, new_n397_, keyIn_0_24, new_n400_ );
nand g266 ( new_n404_, new_n402_, new_n403_ );
nand g267 ( new_n405_, N135, N137 );
not g268 ( new_n406_, new_n405_ );
nand g269 ( new_n407_, new_n404_, new_n406_ );
nand g270 ( new_n408_, new_n402_, new_n403_, new_n405_ );
nand g271 ( new_n409_, new_n407_, new_n408_ );
nand g272 ( new_n410_, new_n409_, keyIn_0_36 );
not g273 ( new_n411_, keyIn_0_36 );
nand g274 ( new_n412_, new_n407_, new_n411_, new_n408_ );
nand g275 ( new_n413_, new_n410_, new_n412_ );
xor g276 ( new_n414_, N73, N89 );
xnor g277 ( new_n415_, N105, N121 );
xnor g278 ( new_n416_, new_n414_, new_n415_ );
xor g279 ( new_n417_, new_n416_, keyIn_0_20 );
not g280 ( new_n418_, new_n417_ );
nand g281 ( new_n419_, new_n413_, new_n418_ );
nand g282 ( new_n420_, new_n410_, new_n412_, new_n417_ );
nand g283 ( new_n421_, new_n419_, new_n420_ );
nand g284 ( new_n422_, new_n421_, new_n366_ );
nand g285 ( new_n423_, new_n419_, keyIn_0_44, new_n420_ );
nand g286 ( new_n424_, new_n422_, new_n423_ );
nor g287 ( new_n425_, new_n365_, new_n424_ );
not g288 ( new_n426_, new_n425_ );
not g289 ( new_n427_, keyIn_0_42 );
nand g290 ( new_n428_, new_n315_, new_n399_ );
nand g291 ( new_n429_, new_n371_, new_n312_, new_n314_ );
nand g292 ( new_n430_, new_n428_, new_n429_ );
nand g293 ( new_n431_, new_n430_, keyIn_0_22 );
not g294 ( new_n432_, keyIn_0_22 );
nand g295 ( new_n433_, new_n428_, new_n432_, new_n429_ );
nand g296 ( new_n434_, new_n431_, new_n433_ );
nand g297 ( new_n435_, N133, N137 );
not g298 ( new_n436_, new_n435_ );
nand g299 ( new_n437_, new_n434_, new_n436_ );
nand g300 ( new_n438_, new_n431_, new_n433_, new_n435_ );
nand g301 ( new_n439_, new_n437_, new_n438_ );
nand g302 ( new_n440_, new_n439_, keyIn_0_34 );
not g303 ( new_n441_, keyIn_0_34 );
nand g304 ( new_n442_, new_n437_, new_n441_, new_n438_ );
nand g305 ( new_n443_, new_n440_, new_n442_ );
xor g306 ( new_n444_, N65, N81 );
xnor g307 ( new_n445_, N97, N113 );
xnor g308 ( new_n446_, new_n444_, new_n445_ );
xor g309 ( new_n447_, new_n446_, keyIn_0_18 );
nand g310 ( new_n448_, new_n443_, new_n447_ );
not g311 ( new_n449_, new_n447_ );
nand g312 ( new_n450_, new_n440_, new_n442_, new_n449_ );
nand g313 ( new_n451_, new_n448_, new_n450_ );
nand g314 ( new_n452_, new_n451_, new_n427_ );
nand g315 ( new_n453_, new_n448_, keyIn_0_42, new_n450_ );
nand g316 ( new_n454_, new_n452_, new_n453_ );
not g317 ( new_n455_, keyIn_0_43 );
not g318 ( new_n456_, keyIn_0_35 );
nand g319 ( new_n457_, new_n340_, new_n396_ );
nand g320 ( new_n458_, new_n337_, new_n339_, new_n394_, new_n395_ );
nand g321 ( new_n459_, new_n457_, new_n458_ );
nand g322 ( new_n460_, new_n459_, keyIn_0_23 );
not g323 ( new_n461_, keyIn_0_23 );
nand g324 ( new_n462_, new_n457_, new_n461_, new_n458_ );
nand g325 ( new_n463_, new_n460_, new_n462_ );
nand g326 ( new_n464_, N134, N137 );
nand g327 ( new_n465_, new_n463_, new_n464_ );
nand g328 ( new_n466_, new_n460_, N134, N137, new_n462_ );
nand g329 ( new_n467_, new_n465_, new_n466_ );
nand g330 ( new_n468_, new_n467_, new_n456_ );
nand g331 ( new_n469_, new_n465_, keyIn_0_35, new_n466_ );
nand g332 ( new_n470_, new_n468_, new_n469_ );
xor g333 ( new_n471_, N69, N85 );
xnor g334 ( new_n472_, N101, N117 );
xnor g335 ( new_n473_, new_n471_, new_n472_ );
xnor g336 ( new_n474_, new_n473_, keyIn_0_19 );
not g337 ( new_n475_, new_n474_ );
nand g338 ( new_n476_, new_n470_, new_n475_ );
nand g339 ( new_n477_, new_n468_, new_n469_, new_n474_ );
nand g340 ( new_n478_, new_n476_, new_n477_ );
nand g341 ( new_n479_, new_n478_, new_n455_ );
nand g342 ( new_n480_, new_n476_, keyIn_0_43, new_n477_ );
and g343 ( new_n481_, new_n479_, new_n480_ );
nor g344 ( new_n482_, new_n426_, new_n454_, new_n481_ );
nand g345 ( new_n483_, new_n292_, new_n294_, new_n482_ );
nand g346 ( new_n484_, new_n483_, new_n184_ );
nand g347 ( new_n485_, new_n292_, new_n294_, keyIn_0_56, new_n482_ );
nand g348 ( new_n486_, new_n484_, new_n485_ );
nand g349 ( new_n487_, new_n486_, new_n183_ );
nand g350 ( new_n488_, new_n487_, N1 );
not g351 ( new_n489_, N1 );
nand g352 ( new_n490_, new_n486_, new_n489_, new_n183_ );
nand g353 ( N724, new_n488_, new_n490_ );
nand g354 ( new_n492_, new_n486_, new_n275_ );
nand g355 ( new_n493_, new_n492_, N5 );
not g356 ( new_n494_, N5 );
nand g357 ( new_n495_, new_n486_, new_n494_, new_n275_ );
nand g358 ( N725, new_n493_, new_n495_ );
nand g359 ( new_n497_, new_n486_, new_n282_ );
nand g360 ( new_n498_, new_n497_, N9 );
not g361 ( new_n499_, N9 );
nand g362 ( new_n500_, new_n486_, new_n499_, new_n282_ );
nand g363 ( N726, new_n498_, new_n500_ );
nand g364 ( new_n502_, new_n486_, new_n278_ );
nand g365 ( new_n503_, new_n502_, N13 );
not g366 ( new_n504_, N13 );
nand g367 ( new_n505_, new_n486_, new_n504_, new_n278_ );
nand g368 ( N727, new_n503_, new_n505_ );
not g369 ( new_n507_, keyIn_0_57 );
and g370 ( new_n508_, new_n363_, new_n364_ );
nand g371 ( new_n509_, new_n479_, new_n480_ );
nand g372 ( new_n510_, new_n509_, new_n424_ );
nor g373 ( new_n511_, new_n510_, new_n508_, new_n454_ );
nand g374 ( new_n512_, new_n292_, new_n294_, new_n511_ );
nand g375 ( new_n513_, new_n512_, new_n507_ );
nand g376 ( new_n514_, new_n292_, new_n294_, keyIn_0_57, new_n511_ );
nand g377 ( new_n515_, new_n513_, new_n514_ );
nand g378 ( new_n516_, new_n515_, new_n183_ );
nand g379 ( new_n517_, new_n516_, N17 );
not g380 ( new_n518_, N17 );
nand g381 ( new_n519_, new_n515_, new_n518_, new_n183_ );
nand g382 ( N728, new_n517_, new_n519_ );
nand g383 ( new_n521_, new_n515_, new_n275_ );
nand g384 ( new_n522_, new_n521_, N21 );
not g385 ( new_n523_, N21 );
nand g386 ( new_n524_, new_n515_, new_n523_, new_n275_ );
nand g387 ( N729, new_n522_, new_n524_ );
nand g388 ( new_n526_, new_n515_, new_n282_ );
nand g389 ( new_n527_, new_n526_, N25 );
nand g390 ( new_n528_, new_n515_, new_n300_, new_n282_ );
nand g391 ( N730, new_n527_, new_n528_ );
nand g392 ( new_n530_, new_n515_, new_n278_ );
nand g393 ( new_n531_, new_n530_, N29 );
nand g394 ( new_n532_, new_n515_, new_n298_, new_n278_ );
nand g395 ( N731, new_n531_, new_n532_ );
not g396 ( new_n534_, keyIn_0_58 );
not g397 ( new_n535_, new_n454_ );
nor g398 ( new_n536_, new_n426_, new_n535_, new_n509_ );
nand g399 ( new_n537_, new_n292_, new_n294_, new_n534_, new_n536_ );
nand g400 ( new_n538_, new_n292_, new_n294_, new_n536_ );
nand g401 ( new_n539_, new_n538_, keyIn_0_58 );
nand g402 ( new_n540_, new_n539_, new_n183_, new_n537_ );
xnor g403 ( N732, new_n540_, N33 );
nand g404 ( new_n542_, new_n539_, new_n275_, new_n537_ );
xnor g405 ( N733, new_n542_, N37 );
nand g406 ( new_n544_, new_n539_, new_n282_, new_n537_ );
xnor g407 ( N734, new_n544_, N41 );
nand g408 ( new_n546_, new_n539_, new_n278_, new_n537_ );
xnor g409 ( N735, new_n546_, N45 );
not g410 ( new_n548_, keyIn_0_59 );
not g411 ( new_n549_, new_n424_ );
nand g412 ( new_n550_, new_n454_, new_n479_, new_n480_ );
nor g413 ( new_n551_, new_n508_, new_n550_, new_n549_ );
nand g414 ( new_n552_, new_n292_, new_n294_, new_n551_ );
nand g415 ( new_n553_, new_n552_, new_n548_ );
nand g416 ( new_n554_, new_n292_, new_n294_, keyIn_0_59, new_n551_ );
nand g417 ( new_n555_, new_n553_, new_n554_ );
nand g418 ( new_n556_, new_n555_, new_n183_ );
nand g419 ( new_n557_, new_n556_, N49 );
nand g420 ( new_n558_, new_n555_, new_n328_, new_n183_ );
nand g421 ( N736, new_n557_, new_n558_ );
nand g422 ( new_n560_, new_n555_, new_n275_ );
nand g423 ( new_n561_, new_n560_, N53 );
nand g424 ( new_n562_, new_n555_, new_n326_, new_n275_ );
nand g425 ( N737, new_n561_, new_n562_ );
nand g426 ( new_n564_, new_n555_, new_n282_ );
nand g427 ( new_n565_, new_n564_, N57 );
not g428 ( new_n566_, N57 );
nand g429 ( new_n567_, new_n555_, new_n566_, new_n282_ );
nand g430 ( N738, new_n565_, new_n567_ );
nand g431 ( new_n569_, new_n555_, new_n278_ );
nand g432 ( new_n570_, new_n569_, N61 );
not g433 ( new_n571_, N61 );
nand g434 ( new_n572_, new_n555_, new_n571_, new_n278_ );
nand g435 ( N739, new_n570_, new_n572_ );
not g436 ( new_n574_, keyIn_0_55 );
not g437 ( new_n575_, keyIn_0_50 );
nand g438 ( new_n576_, new_n365_, new_n509_, new_n424_, new_n454_ );
xnor g439 ( new_n577_, new_n576_, new_n575_ );
nand g440 ( new_n578_, new_n508_, new_n549_, new_n454_, new_n509_ );
nand g441 ( new_n579_, new_n578_, keyIn_0_51 );
not g442 ( new_n580_, keyIn_0_51 );
nand g443 ( new_n581_, new_n425_, new_n580_, new_n454_, new_n509_ );
nand g444 ( new_n582_, new_n579_, new_n581_ );
nand g445 ( new_n583_, new_n424_, new_n363_, new_n364_ );
nor g446 ( new_n584_, new_n583_, new_n550_ );
nand g447 ( new_n585_, new_n584_, keyIn_0_52 );
not g448 ( new_n586_, keyIn_0_52 );
nand g449 ( new_n587_, new_n508_, new_n481_, new_n424_, new_n454_ );
nand g450 ( new_n588_, new_n587_, new_n586_ );
nand g451 ( new_n589_, new_n588_, new_n585_ );
nand g452 ( new_n590_, new_n363_, new_n364_, new_n452_, new_n453_ );
nor g453 ( new_n591_, new_n510_, new_n590_ );
nor g454 ( new_n592_, new_n591_, keyIn_0_53 );
not g455 ( new_n593_, keyIn_0_53 );
nor g456 ( new_n594_, new_n510_, new_n590_, new_n593_ );
nor g457 ( new_n595_, new_n592_, new_n594_ );
nand g458 ( new_n596_, new_n595_, new_n577_, new_n582_, new_n589_ );
nand g459 ( new_n597_, new_n596_, new_n574_ );
nor g460 ( new_n598_, new_n583_, new_n550_, new_n586_ );
nor g461 ( new_n599_, new_n584_, keyIn_0_52 );
nor g462 ( new_n600_, new_n599_, new_n598_ );
nand g463 ( new_n601_, new_n508_, new_n424_, new_n535_, new_n509_ );
nand g464 ( new_n602_, new_n601_, new_n593_ );
nand g465 ( new_n603_, new_n591_, keyIn_0_53 );
nand g466 ( new_n604_, new_n602_, new_n603_ );
nor g467 ( new_n605_, new_n600_, new_n604_ );
nand g468 ( new_n606_, new_n605_, keyIn_0_55, new_n577_, new_n582_ );
nand g469 ( new_n607_, new_n606_, new_n597_ );
nor g470 ( new_n608_, new_n289_, new_n218_ );
nand g471 ( new_n609_, new_n607_, keyIn_0_60, new_n608_ );
not g472 ( new_n610_, keyIn_0_60 );
nand g473 ( new_n611_, new_n607_, new_n608_ );
nand g474 ( new_n612_, new_n611_, new_n610_ );
nand g475 ( new_n613_, new_n612_, new_n535_, new_n609_ );
xnor g476 ( N740, new_n613_, N65 );
nand g477 ( new_n615_, new_n612_, new_n481_, new_n609_ );
xnor g478 ( N741, new_n615_, N69 );
nand g479 ( new_n617_, new_n612_, new_n549_, new_n609_ );
xnor g480 ( N742, new_n617_, N73 );
nand g481 ( new_n619_, new_n612_, new_n365_, new_n609_ );
xnor g482 ( N743, new_n619_, N77 );
nand g483 ( new_n621_, new_n218_, new_n278_ );
nor g484 ( new_n622_, new_n621_, new_n182_, new_n275_ );
nand g485 ( new_n623_, new_n607_, new_n622_ );
nand g486 ( new_n624_, new_n623_, keyIn_0_61 );
not g487 ( new_n625_, keyIn_0_61 );
nand g488 ( new_n626_, new_n607_, new_n625_, new_n622_ );
nand g489 ( new_n627_, new_n624_, new_n626_ );
nand g490 ( new_n628_, new_n627_, new_n535_ );
nand g491 ( new_n629_, new_n628_, N81 );
not g492 ( new_n630_, N81 );
nand g493 ( new_n631_, new_n627_, new_n630_, new_n535_ );
nand g494 ( N744, new_n629_, new_n631_ );
nand g495 ( new_n633_, new_n627_, new_n481_ );
nand g496 ( new_n634_, new_n633_, N85 );
not g497 ( new_n635_, N85 );
nand g498 ( new_n636_, new_n627_, new_n635_, new_n481_ );
nand g499 ( N745, new_n634_, new_n636_ );
nand g500 ( new_n638_, new_n627_, new_n549_ );
nand g501 ( new_n639_, new_n638_, N89 );
not g502 ( new_n640_, N89 );
nand g503 ( new_n641_, new_n627_, new_n640_, new_n549_ );
nand g504 ( N746, new_n639_, new_n641_ );
nand g505 ( new_n643_, new_n627_, new_n365_ );
nand g506 ( new_n644_, new_n643_, N93 );
not g507 ( new_n645_, N93 );
nand g508 ( new_n646_, new_n627_, new_n645_, new_n365_ );
nand g509 ( N747, new_n644_, new_n646_ );
nand g510 ( new_n648_, new_n182_, new_n275_ );
nor g511 ( new_n649_, new_n648_, new_n218_, new_n278_ );
nand g512 ( new_n650_, new_n607_, keyIn_0_62, new_n649_ );
not g513 ( new_n651_, keyIn_0_62 );
nand g514 ( new_n652_, new_n607_, new_n649_ );
nand g515 ( new_n653_, new_n652_, new_n651_ );
nand g516 ( new_n654_, new_n653_, new_n535_, new_n650_ );
xnor g517 ( N748, new_n654_, N97 );
nand g518 ( new_n656_, new_n653_, new_n481_, new_n650_ );
xnor g519 ( N749, new_n656_, N101 );
nand g520 ( new_n658_, new_n653_, new_n549_, new_n650_ );
xnor g521 ( N750, new_n658_, N105 );
nand g522 ( new_n660_, new_n653_, new_n365_, new_n650_ );
xnor g523 ( N751, new_n660_, N109 );
nor g524 ( new_n662_, new_n648_, new_n621_ );
nand g525 ( new_n663_, new_n607_, new_n662_ );
nand g526 ( new_n664_, new_n663_, keyIn_0_63 );
not g527 ( new_n665_, keyIn_0_63 );
nand g528 ( new_n666_, new_n607_, new_n665_, new_n662_ );
nand g529 ( new_n667_, new_n664_, new_n666_ );
nand g530 ( new_n668_, new_n667_, new_n535_ );
nand g531 ( new_n669_, new_n668_, N113 );
not g532 ( new_n670_, N113 );
nand g533 ( new_n671_, new_n667_, new_n670_, new_n535_ );
nand g534 ( N752, new_n669_, new_n671_ );
nand g535 ( new_n673_, new_n667_, new_n481_ );
nand g536 ( new_n674_, new_n673_, N117 );
not g537 ( new_n675_, N117 );
nand g538 ( new_n676_, new_n667_, new_n675_, new_n481_ );
nand g539 ( N753, new_n674_, new_n676_ );
nand g540 ( new_n678_, new_n667_, new_n549_ );
nand g541 ( new_n679_, new_n678_, N121 );
not g542 ( new_n680_, N121 );
nand g543 ( new_n681_, new_n667_, new_n680_, new_n549_ );
nand g544 ( N754, new_n679_, new_n681_ );
nand g545 ( new_n683_, new_n667_, new_n365_ );
nand g546 ( new_n684_, new_n683_, N125 );
not g547 ( new_n685_, N125 );
nand g548 ( new_n686_, new_n667_, new_n685_, new_n365_ );
nand g549 ( N755, new_n684_, new_n686_ );
endmodule