module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n374_, new_n375_, new_n376_, new_n377_, new_n379_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n403_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n415_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n458_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_;
  INV_X1 g000 ( .A(KEYINPUT0), .ZN(new_n123_) );
  INV_X1 g001 ( .A(G953), .ZN(new_n124_) );
  NAND2_X1 g002 ( .A1(G234), .A2(G237), .ZN(new_n125_) );
  XNOR2_X1 g003 ( .A(new_n125_), .B(KEYINPUT14), .ZN(new_n126_) );
  AND2_X1 g004 ( .A1(new_n126_), .A2(G952), .ZN(new_n127_) );
  NAND2_X1 g005 ( .A1(new_n127_), .A2(new_n124_), .ZN(new_n128_) );
  INV_X1 g006 ( .A(G898), .ZN(new_n129_) );
  NAND4_X1 g007 ( .A1(new_n126_), .A2(new_n129_), .A3(G902), .A4(G953), .ZN(new_n130_) );
  NAND2_X1 g008 ( .A1(new_n128_), .A2(new_n130_), .ZN(new_n131_) );
  INV_X1 g009 ( .A(KEYINPUT19), .ZN(new_n132_) );
  NOR2_X1 g010 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n133_) );
  AND2_X1 g011 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n134_) );
  OR2_X1 g012 ( .A1(new_n134_), .A2(new_n133_), .ZN(new_n135_) );
  INV_X1 g013 ( .A(G116), .ZN(new_n136_) );
  NAND2_X1 g014 ( .A1(new_n136_), .A2(G113), .ZN(new_n137_) );
  INV_X1 g015 ( .A(G113), .ZN(new_n138_) );
  NAND2_X1 g016 ( .A1(new_n138_), .A2(G116), .ZN(new_n139_) );
  NAND2_X1 g017 ( .A1(new_n137_), .A2(new_n139_), .ZN(new_n140_) );
  XNOR2_X1 g018 ( .A(G119), .B(KEYINPUT3), .ZN(new_n141_) );
  NAND2_X1 g019 ( .A1(new_n140_), .A2(new_n141_), .ZN(new_n142_) );
  OR2_X1 g020 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n143_) );
  NAND2_X1 g021 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n144_) );
  NAND4_X1 g022 ( .A1(new_n143_), .A2(new_n137_), .A3(new_n139_), .A4(new_n144_), .ZN(new_n145_) );
  NAND2_X1 g023 ( .A1(new_n142_), .A2(new_n145_), .ZN(new_n146_) );
  XOR2_X1 g024 ( .A(G122), .B(KEYINPUT16), .Z(new_n147_) );
  INV_X1 g025 ( .A(new_n147_), .ZN(new_n148_) );
  NAND2_X1 g026 ( .A1(new_n146_), .A2(new_n148_), .ZN(new_n149_) );
  NAND3_X1 g027 ( .A1(new_n142_), .A2(new_n145_), .A3(new_n147_), .ZN(new_n150_) );
  NAND2_X1 g028 ( .A1(new_n149_), .A2(new_n150_), .ZN(new_n151_) );
  INV_X1 g029 ( .A(KEYINPUT18), .ZN(new_n152_) );
  NAND2_X1 g030 ( .A1(new_n152_), .A2(KEYINPUT17), .ZN(new_n153_) );
  INV_X1 g031 ( .A(KEYINPUT17), .ZN(new_n154_) );
  NAND2_X1 g032 ( .A1(new_n154_), .A2(KEYINPUT18), .ZN(new_n155_) );
  NAND2_X1 g033 ( .A1(new_n153_), .A2(new_n155_), .ZN(new_n156_) );
  NAND2_X1 g034 ( .A1(new_n124_), .A2(G224), .ZN(new_n157_) );
  NAND2_X1 g035 ( .A1(new_n156_), .A2(new_n157_), .ZN(new_n158_) );
  NAND4_X1 g036 ( .A1(new_n153_), .A2(new_n155_), .A3(G224), .A4(new_n124_), .ZN(new_n159_) );
  NAND2_X1 g037 ( .A1(new_n158_), .A2(new_n159_), .ZN(new_n160_) );
  XNOR2_X1 g038 ( .A(G125), .B(G146), .ZN(new_n161_) );
  INV_X1 g039 ( .A(new_n161_), .ZN(new_n162_) );
  NAND2_X1 g040 ( .A1(new_n160_), .A2(new_n162_), .ZN(new_n163_) );
  NAND3_X1 g041 ( .A1(new_n158_), .A2(new_n159_), .A3(new_n161_), .ZN(new_n164_) );
  NAND2_X1 g042 ( .A1(new_n163_), .A2(new_n164_), .ZN(new_n165_) );
  NAND2_X1 g043 ( .A1(new_n151_), .A2(new_n165_), .ZN(new_n166_) );
  NAND4_X1 g044 ( .A1(new_n149_), .A2(new_n163_), .A3(new_n150_), .A4(new_n164_), .ZN(new_n167_) );
  NAND2_X1 g045 ( .A1(new_n166_), .A2(new_n167_), .ZN(new_n168_) );
  INV_X1 g046 ( .A(G101), .ZN(new_n169_) );
  INV_X1 g047 ( .A(KEYINPUT4), .ZN(new_n170_) );
  INV_X1 g048 ( .A(G128), .ZN(new_n171_) );
  NAND2_X1 g049 ( .A1(new_n171_), .A2(G143), .ZN(new_n172_) );
  INV_X1 g050 ( .A(G143), .ZN(new_n173_) );
  NAND2_X1 g051 ( .A1(new_n173_), .A2(G128), .ZN(new_n174_) );
  NAND2_X1 g052 ( .A1(new_n172_), .A2(new_n174_), .ZN(new_n175_) );
  NAND2_X1 g053 ( .A1(new_n175_), .A2(new_n170_), .ZN(new_n176_) );
  NAND3_X1 g054 ( .A1(new_n172_), .A2(new_n174_), .A3(KEYINPUT4), .ZN(new_n177_) );
  NAND2_X1 g055 ( .A1(new_n176_), .A2(new_n177_), .ZN(new_n178_) );
  NAND2_X1 g056 ( .A1(new_n178_), .A2(new_n169_), .ZN(new_n179_) );
  NAND3_X1 g057 ( .A1(new_n176_), .A2(G101), .A3(new_n177_), .ZN(new_n180_) );
  NAND2_X1 g058 ( .A1(new_n179_), .A2(new_n180_), .ZN(new_n181_) );
  XNOR2_X1 g059 ( .A(G104), .B(G110), .ZN(new_n182_) );
  XNOR2_X1 g060 ( .A(new_n182_), .B(G107), .ZN(new_n183_) );
  INV_X1 g061 ( .A(new_n183_), .ZN(new_n184_) );
  NAND2_X1 g062 ( .A1(new_n181_), .A2(new_n184_), .ZN(new_n185_) );
  NAND3_X1 g063 ( .A1(new_n179_), .A2(new_n180_), .A3(new_n183_), .ZN(new_n186_) );
  NAND2_X1 g064 ( .A1(new_n185_), .A2(new_n186_), .ZN(new_n187_) );
  NAND2_X1 g065 ( .A1(new_n168_), .A2(new_n187_), .ZN(new_n188_) );
  NAND4_X1 g066 ( .A1(new_n166_), .A2(new_n185_), .A3(new_n167_), .A4(new_n186_), .ZN(new_n189_) );
  NAND2_X1 g067 ( .A1(new_n188_), .A2(new_n189_), .ZN(new_n190_) );
  NAND2_X1 g068 ( .A1(new_n190_), .A2(new_n135_), .ZN(new_n191_) );
  INV_X1 g069 ( .A(G210), .ZN(new_n192_) );
  NOR2_X1 g070 ( .A1(G237), .A2(G902), .ZN(new_n193_) );
  NOR2_X1 g071 ( .A1(new_n193_), .A2(new_n192_), .ZN(new_n194_) );
  NAND2_X1 g072 ( .A1(new_n191_), .A2(new_n194_), .ZN(new_n195_) );
  INV_X1 g073 ( .A(new_n194_), .ZN(new_n196_) );
  NAND3_X1 g074 ( .A1(new_n190_), .A2(new_n135_), .A3(new_n196_), .ZN(new_n197_) );
  NAND2_X1 g075 ( .A1(new_n195_), .A2(new_n197_), .ZN(new_n198_) );
  INV_X1 g076 ( .A(G214), .ZN(new_n199_) );
  OR2_X1 g077 ( .A1(new_n193_), .A2(new_n199_), .ZN(new_n200_) );
  NAND2_X1 g078 ( .A1(new_n198_), .A2(new_n200_), .ZN(new_n201_) );
  NAND2_X1 g079 ( .A1(new_n201_), .A2(new_n132_), .ZN(new_n202_) );
  NAND3_X1 g080 ( .A1(new_n198_), .A2(KEYINPUT19), .A3(new_n200_), .ZN(new_n203_) );
  NAND3_X1 g081 ( .A1(new_n202_), .A2(new_n131_), .A3(new_n203_), .ZN(new_n204_) );
  NAND2_X1 g082 ( .A1(new_n204_), .A2(new_n123_), .ZN(new_n205_) );
  NAND4_X1 g083 ( .A1(new_n202_), .A2(KEYINPUT0), .A3(new_n131_), .A4(new_n203_), .ZN(new_n206_) );
  NAND2_X1 g084 ( .A1(new_n205_), .A2(new_n206_), .ZN(new_n207_) );
  NAND2_X1 g085 ( .A1(new_n135_), .A2(G234), .ZN(new_n208_) );
  XNOR2_X1 g086 ( .A(new_n208_), .B(KEYINPUT20), .ZN(new_n209_) );
  NAND2_X1 g087 ( .A1(new_n209_), .A2(G221), .ZN(new_n210_) );
  XNOR2_X1 g088 ( .A(new_n210_), .B(KEYINPUT21), .ZN(new_n211_) );
  XOR2_X1 g089 ( .A(G475), .B(KEYINPUT13), .Z(new_n212_) );
  INV_X1 g090 ( .A(G902), .ZN(new_n213_) );
  XNOR2_X1 g091 ( .A(G125), .B(KEYINPUT10), .ZN(new_n214_) );
  INV_X1 g092 ( .A(new_n214_), .ZN(new_n215_) );
  XNOR2_X1 g093 ( .A(G140), .B(KEYINPUT11), .ZN(new_n216_) );
  XNOR2_X1 g094 ( .A(G113), .B(G122), .ZN(new_n217_) );
  XNOR2_X1 g095 ( .A(new_n216_), .B(new_n217_), .ZN(new_n218_) );
  OR2_X1 g096 ( .A1(new_n218_), .A2(new_n215_), .ZN(new_n219_) );
  NAND2_X1 g097 ( .A1(new_n218_), .A2(new_n215_), .ZN(new_n220_) );
  NAND2_X1 g098 ( .A1(new_n219_), .A2(new_n220_), .ZN(new_n221_) );
  XOR2_X1 g099 ( .A(G104), .B(G143), .Z(new_n222_) );
  INV_X1 g100 ( .A(new_n222_), .ZN(new_n223_) );
  NAND2_X1 g101 ( .A1(new_n221_), .A2(new_n223_), .ZN(new_n224_) );
  NAND3_X1 g102 ( .A1(new_n219_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n225_) );
  NAND2_X1 g103 ( .A1(new_n224_), .A2(new_n225_), .ZN(new_n226_) );
  XNOR2_X1 g104 ( .A(G131), .B(G146), .ZN(new_n227_) );
  XNOR2_X1 g105 ( .A(new_n227_), .B(KEYINPUT12), .ZN(new_n228_) );
  NOR3_X1 g106 ( .A1(new_n199_), .A2(G237), .A3(G953), .ZN(new_n229_) );
  XNOR2_X1 g107 ( .A(new_n228_), .B(new_n229_), .ZN(new_n230_) );
  INV_X1 g108 ( .A(new_n230_), .ZN(new_n231_) );
  NAND2_X1 g109 ( .A1(new_n226_), .A2(new_n231_), .ZN(new_n232_) );
  NAND3_X1 g110 ( .A1(new_n224_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n233_) );
  NAND3_X1 g111 ( .A1(new_n232_), .A2(new_n213_), .A3(new_n233_), .ZN(new_n234_) );
  XNOR2_X1 g112 ( .A(new_n234_), .B(new_n212_), .ZN(new_n235_) );
  INV_X1 g113 ( .A(KEYINPUT8), .ZN(new_n236_) );
  NAND2_X1 g114 ( .A1(new_n124_), .A2(G234), .ZN(new_n237_) );
  XNOR2_X1 g115 ( .A(new_n237_), .B(new_n236_), .ZN(new_n238_) );
  NAND2_X1 g116 ( .A1(new_n238_), .A2(G217), .ZN(new_n239_) );
  XNOR2_X1 g117 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(new_n240_) );
  INV_X1 g118 ( .A(new_n240_), .ZN(new_n241_) );
  NAND2_X1 g119 ( .A1(new_n239_), .A2(new_n241_), .ZN(new_n242_) );
  NAND3_X1 g120 ( .A1(new_n238_), .A2(G217), .A3(new_n240_), .ZN(new_n243_) );
  NAND2_X1 g121 ( .A1(new_n242_), .A2(new_n243_), .ZN(new_n244_) );
  NAND2_X1 g122 ( .A1(new_n244_), .A2(new_n136_), .ZN(new_n245_) );
  NAND3_X1 g123 ( .A1(new_n242_), .A2(G116), .A3(new_n243_), .ZN(new_n246_) );
  NAND2_X1 g124 ( .A1(new_n245_), .A2(new_n246_), .ZN(new_n247_) );
  XOR2_X1 g125 ( .A(new_n175_), .B(G107), .Z(new_n248_) );
  INV_X1 g126 ( .A(new_n248_), .ZN(new_n249_) );
  NAND2_X1 g127 ( .A1(new_n247_), .A2(new_n249_), .ZN(new_n250_) );
  NAND3_X1 g128 ( .A1(new_n245_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n251_) );
  NAND2_X1 g129 ( .A1(new_n250_), .A2(new_n251_), .ZN(new_n252_) );
  XNOR2_X1 g130 ( .A(G122), .B(G134), .ZN(new_n253_) );
  INV_X1 g131 ( .A(new_n253_), .ZN(new_n254_) );
  NAND2_X1 g132 ( .A1(new_n252_), .A2(new_n254_), .ZN(new_n255_) );
  NAND3_X1 g133 ( .A1(new_n250_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n256_) );
  NAND3_X1 g134 ( .A1(new_n255_), .A2(new_n213_), .A3(new_n256_), .ZN(new_n257_) );
  NAND2_X1 g135 ( .A1(new_n257_), .A2(G478), .ZN(new_n258_) );
  INV_X1 g136 ( .A(G478), .ZN(new_n259_) );
  NAND4_X1 g137 ( .A1(new_n255_), .A2(new_n259_), .A3(new_n213_), .A4(new_n256_), .ZN(new_n260_) );
  NAND2_X1 g138 ( .A1(new_n258_), .A2(new_n260_), .ZN(new_n261_) );
  NOR2_X1 g139 ( .A1(new_n261_), .A2(new_n235_), .ZN(new_n262_) );
  INV_X1 g140 ( .A(new_n262_), .ZN(new_n263_) );
  NOR2_X1 g141 ( .A1(new_n263_), .A2(new_n211_), .ZN(new_n264_) );
  NAND2_X1 g142 ( .A1(new_n207_), .A2(new_n264_), .ZN(new_n265_) );
  NAND2_X1 g143 ( .A1(new_n265_), .A2(KEYINPUT22), .ZN(new_n266_) );
  INV_X1 g144 ( .A(KEYINPUT22), .ZN(new_n267_) );
  NAND3_X1 g145 ( .A1(new_n207_), .A2(new_n267_), .A3(new_n264_), .ZN(new_n268_) );
  AND2_X1 g146 ( .A1(new_n266_), .A2(new_n268_), .ZN(new_n269_) );
  INV_X1 g147 ( .A(G131), .ZN(new_n270_) );
  NAND2_X1 g148 ( .A1(new_n270_), .A2(G146), .ZN(new_n271_) );
  INV_X1 g149 ( .A(G146), .ZN(new_n272_) );
  NAND2_X1 g150 ( .A1(new_n272_), .A2(G131), .ZN(new_n273_) );
  NAND2_X1 g151 ( .A1(new_n271_), .A2(new_n273_), .ZN(new_n274_) );
  NAND2_X1 g152 ( .A1(new_n274_), .A2(G134), .ZN(new_n275_) );
  INV_X1 g153 ( .A(G134), .ZN(new_n276_) );
  NAND2_X1 g154 ( .A1(new_n227_), .A2(new_n276_), .ZN(new_n277_) );
  NAND2_X1 g155 ( .A1(new_n275_), .A2(new_n277_), .ZN(new_n278_) );
  XNOR2_X1 g156 ( .A(G137), .B(G140), .ZN(new_n279_) );
  INV_X1 g157 ( .A(new_n279_), .ZN(new_n280_) );
  NAND2_X1 g158 ( .A1(new_n278_), .A2(new_n280_), .ZN(new_n281_) );
  NAND3_X1 g159 ( .A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n282_) );
  NAND2_X1 g160 ( .A1(new_n281_), .A2(new_n282_), .ZN(new_n283_) );
  NAND2_X1 g161 ( .A1(new_n124_), .A2(G227), .ZN(new_n284_) );
  INV_X1 g162 ( .A(new_n284_), .ZN(new_n285_) );
  NAND2_X1 g163 ( .A1(new_n283_), .A2(new_n285_), .ZN(new_n286_) );
  NAND3_X1 g164 ( .A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n287_) );
  NAND2_X1 g165 ( .A1(new_n286_), .A2(new_n287_), .ZN(new_n288_) );
  NAND2_X1 g166 ( .A1(new_n288_), .A2(new_n187_), .ZN(new_n289_) );
  NAND4_X1 g167 ( .A1(new_n286_), .A2(new_n185_), .A3(new_n186_), .A4(new_n287_), .ZN(new_n290_) );
  NAND3_X1 g168 ( .A1(new_n289_), .A2(new_n213_), .A3(new_n290_), .ZN(new_n291_) );
  NAND2_X1 g169 ( .A1(new_n291_), .A2(G469), .ZN(new_n292_) );
  INV_X1 g170 ( .A(G469), .ZN(new_n293_) );
  NAND4_X1 g171 ( .A1(new_n289_), .A2(new_n293_), .A3(new_n213_), .A4(new_n290_), .ZN(new_n294_) );
  NAND2_X1 g172 ( .A1(new_n292_), .A2(new_n294_), .ZN(new_n295_) );
  NAND2_X1 g173 ( .A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n296_) );
  INV_X1 g174 ( .A(KEYINPUT1), .ZN(new_n297_) );
  NAND3_X1 g175 ( .A1(new_n292_), .A2(new_n297_), .A3(new_n294_), .ZN(new_n298_) );
  NAND2_X1 g176 ( .A1(new_n296_), .A2(new_n298_), .ZN(new_n299_) );
  INV_X1 g177 ( .A(new_n299_), .ZN(new_n300_) );
  INV_X1 g178 ( .A(G472), .ZN(new_n301_) );
  INV_X1 g179 ( .A(KEYINPUT5), .ZN(new_n302_) );
  NAND2_X1 g180 ( .A1(new_n302_), .A2(G137), .ZN(new_n303_) );
  INV_X1 g181 ( .A(G137), .ZN(new_n304_) );
  NAND2_X1 g182 ( .A1(new_n304_), .A2(KEYINPUT5), .ZN(new_n305_) );
  NAND2_X1 g183 ( .A1(new_n303_), .A2(new_n305_), .ZN(new_n306_) );
  INV_X1 g184 ( .A(G237), .ZN(new_n307_) );
  NAND3_X1 g185 ( .A1(new_n307_), .A2(new_n124_), .A3(G210), .ZN(new_n308_) );
  NAND2_X1 g186 ( .A1(new_n306_), .A2(new_n308_), .ZN(new_n309_) );
  NOR3_X1 g187 ( .A1(new_n192_), .A2(G237), .A3(G953), .ZN(new_n310_) );
  NAND3_X1 g188 ( .A1(new_n310_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n311_) );
  NAND2_X1 g189 ( .A1(new_n309_), .A2(new_n311_), .ZN(new_n312_) );
  NAND2_X1 g190 ( .A1(new_n146_), .A2(new_n312_), .ZN(new_n313_) );
  NAND4_X1 g191 ( .A1(new_n142_), .A2(new_n309_), .A3(new_n145_), .A4(new_n311_), .ZN(new_n314_) );
  NAND2_X1 g192 ( .A1(new_n313_), .A2(new_n314_), .ZN(new_n315_) );
  NAND2_X1 g193 ( .A1(new_n315_), .A2(new_n278_), .ZN(new_n316_) );
  NAND4_X1 g194 ( .A1(new_n313_), .A2(new_n275_), .A3(new_n277_), .A4(new_n314_), .ZN(new_n317_) );
  NAND2_X1 g195 ( .A1(new_n316_), .A2(new_n317_), .ZN(new_n318_) );
  NAND2_X1 g196 ( .A1(new_n318_), .A2(new_n181_), .ZN(new_n319_) );
  NAND4_X1 g197 ( .A1(new_n316_), .A2(new_n179_), .A3(new_n180_), .A4(new_n317_), .ZN(new_n320_) );
  NAND3_X1 g198 ( .A1(new_n319_), .A2(new_n213_), .A3(new_n320_), .ZN(new_n321_) );
  NAND2_X1 g199 ( .A1(new_n321_), .A2(new_n301_), .ZN(new_n322_) );
  NAND4_X1 g200 ( .A1(new_n319_), .A2(G472), .A3(new_n213_), .A4(new_n320_), .ZN(new_n323_) );
  NAND2_X1 g201 ( .A1(new_n322_), .A2(new_n323_), .ZN(new_n324_) );
  NAND2_X1 g202 ( .A1(new_n324_), .A2(KEYINPUT6), .ZN(new_n325_) );
  INV_X1 g203 ( .A(KEYINPUT6), .ZN(new_n326_) );
  NAND3_X1 g204 ( .A1(new_n322_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n327_) );
  NAND2_X1 g205 ( .A1(new_n325_), .A2(new_n327_), .ZN(new_n328_) );
  INV_X1 g206 ( .A(new_n328_), .ZN(new_n329_) );
  INV_X1 g207 ( .A(KEYINPUT25), .ZN(new_n330_) );
  NAND2_X1 g208 ( .A1(new_n209_), .A2(G217), .ZN(new_n331_) );
  NAND2_X1 g209 ( .A1(new_n214_), .A2(new_n279_), .ZN(new_n332_) );
  NAND2_X1 g210 ( .A1(new_n215_), .A2(new_n280_), .ZN(new_n333_) );
  NAND2_X1 g211 ( .A1(new_n333_), .A2(new_n332_), .ZN(new_n334_) );
  XOR2_X1 g212 ( .A(G119), .B(G146), .Z(new_n335_) );
  XNOR2_X1 g213 ( .A(G110), .B(G128), .ZN(new_n336_) );
  NAND2_X1 g214 ( .A1(new_n335_), .A2(new_n336_), .ZN(new_n337_) );
  OR2_X1 g215 ( .A1(new_n335_), .A2(new_n336_), .ZN(new_n338_) );
  NAND2_X1 g216 ( .A1(new_n338_), .A2(new_n337_), .ZN(new_n339_) );
  NAND2_X1 g217 ( .A1(new_n339_), .A2(new_n334_), .ZN(new_n340_) );
  NAND4_X1 g218 ( .A1(new_n338_), .A2(new_n332_), .A3(new_n333_), .A4(new_n337_), .ZN(new_n341_) );
  NAND2_X1 g219 ( .A1(new_n340_), .A2(new_n341_), .ZN(new_n342_) );
  NAND2_X1 g220 ( .A1(new_n238_), .A2(G221), .ZN(new_n343_) );
  XOR2_X1 g221 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n344_) );
  NAND2_X1 g222 ( .A1(new_n343_), .A2(new_n344_), .ZN(new_n345_) );
  OR2_X1 g223 ( .A1(new_n343_), .A2(new_n344_), .ZN(new_n346_) );
  NAND2_X1 g224 ( .A1(new_n346_), .A2(new_n345_), .ZN(new_n347_) );
  NAND2_X1 g225 ( .A1(new_n347_), .A2(new_n342_), .ZN(new_n348_) );
  NAND4_X1 g226 ( .A1(new_n346_), .A2(new_n340_), .A3(new_n341_), .A4(new_n345_), .ZN(new_n349_) );
  NAND4_X1 g227 ( .A1(new_n348_), .A2(new_n213_), .A3(new_n331_), .A4(new_n349_), .ZN(new_n350_) );
  INV_X1 g228 ( .A(new_n331_), .ZN(new_n351_) );
  NAND3_X1 g229 ( .A1(new_n348_), .A2(new_n213_), .A3(new_n349_), .ZN(new_n352_) );
  NAND2_X1 g230 ( .A1(new_n352_), .A2(new_n351_), .ZN(new_n353_) );
  NAND2_X1 g231 ( .A1(new_n353_), .A2(new_n350_), .ZN(new_n354_) );
  NAND2_X1 g232 ( .A1(new_n354_), .A2(new_n330_), .ZN(new_n355_) );
  NAND3_X1 g233 ( .A1(new_n353_), .A2(KEYINPUT25), .A3(new_n350_), .ZN(new_n356_) );
  NAND2_X1 g234 ( .A1(new_n355_), .A2(new_n356_), .ZN(new_n357_) );
  INV_X1 g235 ( .A(new_n357_), .ZN(new_n358_) );
  NAND4_X1 g236 ( .A1(new_n269_), .A2(new_n300_), .A3(new_n329_), .A4(new_n358_), .ZN(new_n359_) );
  XNOR2_X1 g237 ( .A(new_n359_), .B(G101), .ZN(G3) );
  AND2_X1 g238 ( .A1(new_n292_), .A2(new_n294_), .ZN(new_n361_) );
  INV_X1 g239 ( .A(new_n324_), .ZN(new_n362_) );
  INV_X1 g240 ( .A(new_n211_), .ZN(new_n363_) );
  AND3_X1 g241 ( .A1(new_n355_), .A2(new_n363_), .A3(new_n356_), .ZN(new_n364_) );
  INV_X1 g242 ( .A(new_n364_), .ZN(new_n365_) );
  NOR3_X1 g243 ( .A1(new_n365_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n366_) );
  NAND2_X1 g244 ( .A1(new_n207_), .A2(new_n366_), .ZN(new_n367_) );
  INV_X1 g245 ( .A(new_n212_), .ZN(new_n368_) );
  XNOR2_X1 g246 ( .A(new_n234_), .B(new_n368_), .ZN(new_n369_) );
  NOR2_X1 g247 ( .A1(new_n261_), .A2(new_n369_), .ZN(new_n370_) );
  INV_X1 g248 ( .A(new_n370_), .ZN(new_n371_) );
  NOR2_X1 g249 ( .A1(new_n367_), .A2(new_n371_), .ZN(new_n372_) );
  XOR2_X1 g250 ( .A(new_n372_), .B(G104), .Z(G6) );
  NAND2_X1 g251 ( .A1(new_n261_), .A2(new_n369_), .ZN(new_n374_) );
  NOR2_X1 g252 ( .A1(new_n367_), .A2(new_n374_), .ZN(new_n375_) );
  XNOR2_X1 g253 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(new_n376_) );
  XNOR2_X1 g254 ( .A(new_n375_), .B(new_n376_), .ZN(new_n377_) );
  XNOR2_X1 g255 ( .A(new_n377_), .B(G107), .ZN(G9) );
  NAND4_X1 g256 ( .A1(new_n269_), .A2(new_n300_), .A3(new_n324_), .A4(new_n357_), .ZN(new_n379_) );
  XNOR2_X1 g257 ( .A(new_n379_), .B(G110), .ZN(G12) );
  INV_X1 g258 ( .A(new_n374_), .ZN(new_n381_) );
  AND2_X1 g259 ( .A1(new_n202_), .A2(new_n203_), .ZN(new_n382_) );
  INV_X1 g260 ( .A(KEYINPUT28), .ZN(new_n383_) );
  NOR2_X1 g261 ( .A1(new_n124_), .A2(G900), .ZN(new_n384_) );
  NAND3_X1 g262 ( .A1(new_n126_), .A2(G902), .A3(new_n384_), .ZN(new_n385_) );
  NAND2_X1 g263 ( .A1(new_n128_), .A2(new_n385_), .ZN(new_n386_) );
  INV_X1 g264 ( .A(new_n386_), .ZN(new_n387_) );
  NOR2_X1 g265 ( .A1(new_n211_), .A2(new_n387_), .ZN(new_n388_) );
  NAND4_X1 g266 ( .A1(new_n357_), .A2(new_n383_), .A3(new_n362_), .A4(new_n388_), .ZN(new_n389_) );
  NAND3_X1 g267 ( .A1(new_n357_), .A2(new_n362_), .A3(new_n388_), .ZN(new_n390_) );
  NAND2_X1 g268 ( .A1(new_n390_), .A2(KEYINPUT28), .ZN(new_n391_) );
  AND3_X1 g269 ( .A1(new_n391_), .A2(new_n295_), .A3(new_n389_), .ZN(new_n392_) );
  AND2_X1 g270 ( .A1(new_n392_), .A2(new_n382_), .ZN(new_n393_) );
  NAND2_X1 g271 ( .A1(new_n393_), .A2(new_n381_), .ZN(new_n394_) );
  XOR2_X1 g272 ( .A(G128), .B(KEYINPUT29), .Z(new_n395_) );
  XNOR2_X1 g273 ( .A(new_n394_), .B(new_n395_), .ZN(G30) );
  NAND3_X1 g274 ( .A1(new_n322_), .A2(new_n200_), .A3(new_n323_), .ZN(new_n397_) );
  XOR2_X1 g275 ( .A(new_n397_), .B(KEYINPUT30), .Z(new_n398_) );
  NOR4_X1 g276 ( .A1(new_n357_), .A2(new_n361_), .A3(new_n211_), .A4(new_n387_), .ZN(new_n399_) );
  AND2_X1 g277 ( .A1(new_n261_), .A2(new_n235_), .ZN(new_n400_) );
  NAND4_X1 g278 ( .A1(new_n400_), .A2(new_n198_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n401_) );
  XNOR2_X1 g279 ( .A(new_n401_), .B(G143), .ZN(G45) );
  NAND2_X1 g280 ( .A1(new_n393_), .A2(new_n370_), .ZN(new_n403_) );
  XNOR2_X1 g281 ( .A(new_n403_), .B(G146), .ZN(G48) );
  INV_X1 g282 ( .A(KEYINPUT31), .ZN(new_n405_) );
  NOR2_X1 g283 ( .A1(new_n300_), .A2(new_n365_), .ZN(new_n406_) );
  INV_X1 g284 ( .A(new_n406_), .ZN(new_n407_) );
  NOR2_X1 g285 ( .A1(new_n407_), .A2(new_n324_), .ZN(new_n408_) );
  NAND2_X1 g286 ( .A1(new_n408_), .A2(new_n207_), .ZN(new_n409_) );
  NAND2_X1 g287 ( .A1(new_n409_), .A2(new_n405_), .ZN(new_n410_) );
  NAND3_X1 g288 ( .A1(new_n408_), .A2(new_n207_), .A3(KEYINPUT31), .ZN(new_n411_) );
  NAND2_X1 g289 ( .A1(new_n410_), .A2(new_n411_), .ZN(new_n412_) );
  NOR2_X1 g290 ( .A1(new_n412_), .A2(new_n371_), .ZN(new_n413_) );
  XNOR2_X1 g291 ( .A(new_n413_), .B(new_n138_), .ZN(G15) );
  NOR2_X1 g292 ( .A1(new_n412_), .A2(new_n374_), .ZN(new_n415_) );
  XNOR2_X1 g293 ( .A(new_n415_), .B(new_n136_), .ZN(G18) );
  NOR3_X1 g294 ( .A1(new_n300_), .A2(new_n328_), .A3(new_n358_), .ZN(new_n417_) );
  NAND3_X1 g295 ( .A1(new_n266_), .A2(new_n268_), .A3(new_n417_), .ZN(new_n418_) );
  NAND2_X1 g296 ( .A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n419_) );
  INV_X1 g297 ( .A(KEYINPUT32), .ZN(new_n420_) );
  NAND4_X1 g298 ( .A1(new_n266_), .A2(new_n420_), .A3(new_n268_), .A4(new_n417_), .ZN(new_n421_) );
  NAND2_X1 g299 ( .A1(new_n419_), .A2(new_n421_), .ZN(new_n422_) );
  XNOR2_X1 g300 ( .A(new_n422_), .B(G119), .ZN(G21) );
  INV_X1 g301 ( .A(KEYINPUT34), .ZN(new_n424_) );
  NAND3_X1 g302 ( .A1(new_n299_), .A2(new_n328_), .A3(new_n364_), .ZN(new_n425_) );
  XNOR2_X1 g303 ( .A(new_n425_), .B(KEYINPUT33), .ZN(new_n426_) );
  NAND2_X1 g304 ( .A1(new_n426_), .A2(new_n207_), .ZN(new_n427_) );
  NAND2_X1 g305 ( .A1(new_n427_), .A2(new_n424_), .ZN(new_n428_) );
  NAND3_X1 g306 ( .A1(new_n426_), .A2(new_n207_), .A3(KEYINPUT34), .ZN(new_n429_) );
  NAND2_X1 g307 ( .A1(new_n428_), .A2(new_n429_), .ZN(new_n430_) );
  NAND2_X1 g308 ( .A1(new_n430_), .A2(new_n400_), .ZN(new_n431_) );
  NAND2_X1 g309 ( .A1(new_n431_), .A2(KEYINPUT35), .ZN(new_n432_) );
  INV_X1 g310 ( .A(KEYINPUT35), .ZN(new_n433_) );
  NAND3_X1 g311 ( .A1(new_n430_), .A2(new_n433_), .A3(new_n400_), .ZN(new_n434_) );
  NAND2_X1 g312 ( .A1(new_n432_), .A2(new_n434_), .ZN(new_n435_) );
  XOR2_X1 g313 ( .A(new_n435_), .B(G122), .Z(G24) );
  NAND3_X1 g314 ( .A1(new_n328_), .A2(new_n357_), .A3(new_n388_), .ZN(new_n437_) );
  NOR2_X1 g315 ( .A1(new_n371_), .A2(new_n437_), .ZN(new_n438_) );
  NAND3_X1 g316 ( .A1(new_n438_), .A2(new_n198_), .A3(new_n200_), .ZN(new_n439_) );
  OR2_X1 g317 ( .A1(new_n439_), .A2(KEYINPUT36), .ZN(new_n440_) );
  NAND2_X1 g318 ( .A1(new_n439_), .A2(KEYINPUT36), .ZN(new_n441_) );
  NAND3_X1 g319 ( .A1(new_n440_), .A2(new_n299_), .A3(new_n441_), .ZN(new_n442_) );
  XOR2_X1 g320 ( .A(new_n442_), .B(G125), .Z(new_n443_) );
  XNOR2_X1 g321 ( .A(new_n443_), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 g322 ( .A(KEYINPUT40), .ZN(new_n445_) );
  INV_X1 g323 ( .A(KEYINPUT38), .ZN(new_n446_) );
  XNOR2_X1 g324 ( .A(new_n198_), .B(new_n446_), .ZN(new_n447_) );
  NAND3_X1 g325 ( .A1(new_n398_), .A2(new_n447_), .A3(new_n399_), .ZN(new_n448_) );
  NAND2_X1 g326 ( .A1(new_n448_), .A2(KEYINPUT39), .ZN(new_n449_) );
  INV_X1 g327 ( .A(KEYINPUT39), .ZN(new_n450_) );
  NAND4_X1 g328 ( .A1(new_n398_), .A2(new_n447_), .A3(new_n399_), .A4(new_n450_), .ZN(new_n451_) );
  NAND2_X1 g329 ( .A1(new_n449_), .A2(new_n451_), .ZN(new_n452_) );
  NAND2_X1 g330 ( .A1(new_n452_), .A2(new_n370_), .ZN(new_n453_) );
  NAND2_X1 g331 ( .A1(new_n453_), .A2(new_n445_), .ZN(new_n454_) );
  NAND3_X1 g332 ( .A1(new_n452_), .A2(KEYINPUT40), .A3(new_n370_), .ZN(new_n455_) );
  NAND2_X1 g333 ( .A1(new_n454_), .A2(new_n455_), .ZN(new_n456_) );
  XNOR2_X1 g334 ( .A(new_n456_), .B(new_n270_), .ZN(G33) );
  NAND2_X1 g335 ( .A1(new_n452_), .A2(new_n381_), .ZN(new_n458_) );
  XNOR2_X1 g336 ( .A(new_n458_), .B(G134), .ZN(G36) );
  INV_X1 g337 ( .A(KEYINPUT42), .ZN(new_n460_) );
  INV_X1 g338 ( .A(KEYINPUT41), .ZN(new_n461_) );
  AND4_X1 g339 ( .A1(new_n200_), .A2(new_n369_), .A3(new_n258_), .A4(new_n260_), .ZN(new_n462_) );
  NAND2_X1 g340 ( .A1(new_n462_), .A2(new_n447_), .ZN(new_n463_) );
  NAND2_X1 g341 ( .A1(new_n463_), .A2(new_n461_), .ZN(new_n464_) );
  NAND3_X1 g342 ( .A1(new_n462_), .A2(KEYINPUT41), .A3(new_n447_), .ZN(new_n465_) );
  NAND3_X1 g343 ( .A1(new_n464_), .A2(new_n392_), .A3(new_n465_), .ZN(new_n466_) );
  NAND2_X1 g344 ( .A1(new_n466_), .A2(new_n460_), .ZN(new_n467_) );
  NAND4_X1 g345 ( .A1(new_n464_), .A2(KEYINPUT42), .A3(new_n392_), .A4(new_n465_), .ZN(new_n468_) );
  AND2_X1 g346 ( .A1(new_n467_), .A2(new_n468_), .ZN(new_n469_) );
  XNOR2_X1 g347 ( .A(new_n469_), .B(G137), .ZN(G39) );
  INV_X1 g348 ( .A(KEYINPUT43), .ZN(new_n471_) );
  NAND3_X1 g349 ( .A1(new_n438_), .A2(new_n200_), .A3(new_n300_), .ZN(new_n472_) );
  OR2_X1 g350 ( .A1(new_n472_), .A2(new_n471_), .ZN(new_n473_) );
  NAND2_X1 g351 ( .A1(new_n472_), .A2(new_n471_), .ZN(new_n474_) );
  NAND4_X1 g352 ( .A1(new_n473_), .A2(new_n195_), .A3(new_n197_), .A4(new_n474_), .ZN(new_n475_) );
  XNOR2_X1 g353 ( .A(new_n475_), .B(G140), .ZN(G42) );
  INV_X1 g354 ( .A(KEYINPUT2), .ZN(new_n477_) );
  INV_X1 g355 ( .A(KEYINPUT48), .ZN(new_n478_) );
  INV_X1 g356 ( .A(KEYINPUT46), .ZN(new_n479_) );
  NAND4_X1 g357 ( .A1(new_n454_), .A2(new_n455_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n480_) );
  NAND2_X1 g358 ( .A1(new_n480_), .A2(new_n479_), .ZN(new_n481_) );
  NAND4_X1 g359 ( .A1(new_n469_), .A2(KEYINPUT46), .A3(new_n454_), .A4(new_n455_), .ZN(new_n482_) );
  NAND2_X1 g360 ( .A1(new_n482_), .A2(new_n481_), .ZN(new_n483_) );
  NAND2_X1 g361 ( .A1(new_n442_), .A2(new_n401_), .ZN(new_n484_) );
  NAND2_X1 g362 ( .A1(new_n371_), .A2(new_n374_), .ZN(new_n485_) );
  NAND2_X1 g363 ( .A1(new_n393_), .A2(new_n485_), .ZN(new_n486_) );
  XNOR2_X1 g364 ( .A(new_n486_), .B(KEYINPUT47), .ZN(new_n487_) );
  NOR2_X1 g365 ( .A1(new_n484_), .A2(new_n487_), .ZN(new_n488_) );
  NAND3_X1 g366 ( .A1(new_n483_), .A2(new_n488_), .A3(new_n478_), .ZN(new_n489_) );
  NAND2_X1 g367 ( .A1(new_n483_), .A2(new_n488_), .ZN(new_n490_) );
  NAND2_X1 g368 ( .A1(new_n490_), .A2(KEYINPUT48), .ZN(new_n491_) );
  AND2_X1 g369 ( .A1(new_n475_), .A2(new_n458_), .ZN(new_n492_) );
  AND3_X1 g370 ( .A1(new_n491_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_) );
  INV_X1 g371 ( .A(KEYINPUT45), .ZN(new_n494_) );
  NAND2_X1 g372 ( .A1(new_n422_), .A2(new_n379_), .ZN(new_n495_) );
  NAND2_X1 g373 ( .A1(new_n495_), .A2(KEYINPUT44), .ZN(new_n496_) );
  AND2_X1 g374 ( .A1(new_n422_), .A2(new_n379_), .ZN(new_n497_) );
  INV_X1 g375 ( .A(KEYINPUT44), .ZN(new_n498_) );
  AND3_X1 g376 ( .A1(new_n432_), .A2(new_n498_), .A3(new_n434_), .ZN(new_n499_) );
  NAND2_X1 g377 ( .A1(new_n499_), .A2(new_n497_), .ZN(new_n500_) );
  NAND2_X1 g378 ( .A1(new_n435_), .A2(KEYINPUT44), .ZN(new_n501_) );
  NAND2_X1 g379 ( .A1(new_n412_), .A2(new_n367_), .ZN(new_n502_) );
  NAND2_X1 g380 ( .A1(new_n502_), .A2(new_n485_), .ZN(new_n503_) );
  AND2_X1 g381 ( .A1(new_n503_), .A2(new_n359_), .ZN(new_n504_) );
  NAND4_X1 g382 ( .A1(new_n500_), .A2(new_n496_), .A3(new_n501_), .A4(new_n504_), .ZN(new_n505_) );
  NAND2_X1 g383 ( .A1(new_n505_), .A2(new_n494_), .ZN(new_n506_) );
  AND2_X1 g384 ( .A1(new_n501_), .A2(new_n504_), .ZN(new_n507_) );
  NAND4_X1 g385 ( .A1(new_n507_), .A2(KEYINPUT45), .A3(new_n496_), .A4(new_n500_), .ZN(new_n508_) );
  NAND3_X1 g386 ( .A1(new_n506_), .A2(new_n493_), .A3(new_n508_), .ZN(new_n509_) );
  NAND2_X1 g387 ( .A1(new_n509_), .A2(new_n477_), .ZN(new_n510_) );
  NAND4_X1 g388 ( .A1(new_n506_), .A2(new_n493_), .A3(new_n508_), .A4(KEYINPUT2), .ZN(new_n511_) );
  NAND2_X1 g389 ( .A1(new_n510_), .A2(new_n511_), .ZN(new_n512_) );
  INV_X1 g390 ( .A(new_n408_), .ZN(new_n513_) );
  NOR2_X1 g391 ( .A1(new_n299_), .A2(new_n364_), .ZN(new_n514_) );
  NAND2_X1 g392 ( .A1(new_n514_), .A2(KEYINPUT50), .ZN(new_n515_) );
  OR2_X1 g393 ( .A1(new_n514_), .A2(KEYINPUT50), .ZN(new_n516_) );
  NAND2_X1 g394 ( .A1(new_n357_), .A2(new_n211_), .ZN(new_n517_) );
  XOR2_X1 g395 ( .A(new_n517_), .B(KEYINPUT49), .Z(new_n518_) );
  NAND4_X1 g396 ( .A1(new_n518_), .A2(new_n516_), .A3(new_n324_), .A4(new_n515_), .ZN(new_n519_) );
  NAND2_X1 g397 ( .A1(new_n513_), .A2(new_n519_), .ZN(new_n520_) );
  OR2_X1 g398 ( .A1(new_n520_), .A2(KEYINPUT51), .ZN(new_n521_) );
  NAND2_X1 g399 ( .A1(new_n520_), .A2(KEYINPUT51), .ZN(new_n522_) );
  NAND4_X1 g400 ( .A1(new_n521_), .A2(new_n464_), .A3(new_n465_), .A4(new_n522_), .ZN(new_n523_) );
  NAND2_X1 g401 ( .A1(new_n485_), .A2(new_n200_), .ZN(new_n524_) );
  NAND2_X1 g402 ( .A1(new_n524_), .A2(new_n263_), .ZN(new_n525_) );
  OR2_X1 g403 ( .A1(new_n462_), .A2(new_n447_), .ZN(new_n526_) );
  NAND3_X1 g404 ( .A1(new_n525_), .A2(new_n426_), .A3(new_n526_), .ZN(new_n527_) );
  AND2_X1 g405 ( .A1(new_n523_), .A2(new_n527_), .ZN(new_n528_) );
  NAND2_X1 g406 ( .A1(new_n528_), .A2(KEYINPUT52), .ZN(new_n529_) );
  OR2_X1 g407 ( .A1(new_n528_), .A2(KEYINPUT52), .ZN(new_n530_) );
  NAND3_X1 g408 ( .A1(new_n530_), .A2(new_n127_), .A3(new_n529_), .ZN(new_n531_) );
  NAND3_X1 g409 ( .A1(new_n464_), .A2(new_n426_), .A3(new_n465_), .ZN(new_n532_) );
  NAND4_X1 g410 ( .A1(new_n512_), .A2(new_n124_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_) );
  XOR2_X1 g411 ( .A(new_n533_), .B(KEYINPUT53), .Z(G75) );
  INV_X1 g412 ( .A(KEYINPUT56), .ZN(new_n535_) );
  NOR2_X1 g413 ( .A1(new_n135_), .A2(new_n192_), .ZN(new_n536_) );
  XOR2_X1 g414 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(new_n537_) );
  XNOR2_X1 g415 ( .A(new_n190_), .B(new_n537_), .ZN(new_n538_) );
  NAND4_X1 g416 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n539_) );
  OR2_X1 g417 ( .A1(new_n124_), .A2(G952), .ZN(new_n540_) );
  NAND3_X1 g418 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n536_), .ZN(new_n541_) );
  INV_X1 g419 ( .A(new_n538_), .ZN(new_n542_) );
  NAND2_X1 g420 ( .A1(new_n541_), .A2(new_n542_), .ZN(new_n543_) );
  NAND3_X1 g421 ( .A1(new_n543_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n544_) );
  NAND2_X1 g422 ( .A1(new_n544_), .A2(new_n535_), .ZN(new_n545_) );
  NAND4_X1 g423 ( .A1(new_n543_), .A2(KEYINPUT56), .A3(new_n539_), .A4(new_n540_), .ZN(new_n546_) );
  NAND2_X1 g424 ( .A1(new_n545_), .A2(new_n546_), .ZN(G51) );
  NOR2_X1 g425 ( .A1(new_n135_), .A2(new_n293_), .ZN(new_n548_) );
  NAND3_X1 g426 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n548_), .ZN(new_n549_) );
  XNOR2_X1 g427 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(new_n550_) );
  INV_X1 g428 ( .A(new_n550_), .ZN(new_n551_) );
  NAND2_X1 g429 ( .A1(new_n549_), .A2(new_n551_), .ZN(new_n552_) );
  NAND4_X1 g430 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n548_), .A4(new_n550_), .ZN(new_n553_) );
  NAND4_X1 g431 ( .A1(new_n552_), .A2(new_n289_), .A3(new_n290_), .A4(new_n553_), .ZN(new_n554_) );
  NAND2_X1 g432 ( .A1(new_n289_), .A2(new_n290_), .ZN(new_n555_) );
  NAND2_X1 g433 ( .A1(new_n552_), .A2(new_n553_), .ZN(new_n556_) );
  NAND2_X1 g434 ( .A1(new_n556_), .A2(new_n555_), .ZN(new_n557_) );
  AND3_X1 g435 ( .A1(new_n557_), .A2(new_n540_), .A3(new_n554_), .ZN(G54) );
  INV_X1 g436 ( .A(KEYINPUT60), .ZN(new_n559_) );
  INV_X1 g437 ( .A(new_n135_), .ZN(new_n560_) );
  AND2_X1 g438 ( .A1(new_n560_), .A2(G475), .ZN(new_n561_) );
  NAND3_X1 g439 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n561_), .ZN(new_n562_) );
  NAND2_X1 g440 ( .A1(new_n232_), .A2(new_n233_), .ZN(new_n563_) );
  XNOR2_X1 g441 ( .A(new_n563_), .B(KEYINPUT59), .ZN(new_n564_) );
  INV_X1 g442 ( .A(new_n564_), .ZN(new_n565_) );
  NAND2_X1 g443 ( .A1(new_n562_), .A2(new_n565_), .ZN(new_n566_) );
  NAND4_X1 g444 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n561_), .A4(new_n564_), .ZN(new_n567_) );
  NAND3_X1 g445 ( .A1(new_n566_), .A2(new_n540_), .A3(new_n567_), .ZN(new_n568_) );
  NAND2_X1 g446 ( .A1(new_n568_), .A2(new_n559_), .ZN(new_n569_) );
  NAND4_X1 g447 ( .A1(new_n566_), .A2(KEYINPUT60), .A3(new_n540_), .A4(new_n567_), .ZN(new_n570_) );
  NAND2_X1 g448 ( .A1(new_n569_), .A2(new_n570_), .ZN(G60) );
  NAND2_X1 g449 ( .A1(new_n255_), .A2(new_n256_), .ZN(new_n572_) );
  INV_X1 g450 ( .A(new_n512_), .ZN(new_n573_) );
  NAND3_X1 g451 ( .A1(new_n573_), .A2(G478), .A3(new_n560_), .ZN(new_n574_) );
  NAND2_X1 g452 ( .A1(new_n574_), .A2(new_n572_), .ZN(new_n575_) );
  INV_X1 g453 ( .A(new_n572_), .ZN(new_n576_) );
  NAND4_X1 g454 ( .A1(new_n573_), .A2(G478), .A3(new_n560_), .A4(new_n576_), .ZN(new_n577_) );
  AND3_X1 g455 ( .A1(new_n575_), .A2(new_n540_), .A3(new_n577_), .ZN(G63) );
  NAND2_X1 g456 ( .A1(new_n348_), .A2(new_n349_), .ZN(new_n579_) );
  NAND3_X1 g457 ( .A1(new_n573_), .A2(G217), .A3(new_n560_), .ZN(new_n580_) );
  NAND2_X1 g458 ( .A1(new_n580_), .A2(new_n579_), .ZN(new_n581_) );
  INV_X1 g459 ( .A(new_n579_), .ZN(new_n582_) );
  NAND4_X1 g460 ( .A1(new_n573_), .A2(G217), .A3(new_n560_), .A4(new_n582_), .ZN(new_n583_) );
  AND3_X1 g461 ( .A1(new_n581_), .A2(new_n540_), .A3(new_n583_), .ZN(G66) );
  AND2_X1 g462 ( .A1(G224), .A2(G953), .ZN(new_n585_) );
  OR2_X1 g463 ( .A1(new_n585_), .A2(KEYINPUT61), .ZN(new_n586_) );
  NAND2_X1 g464 ( .A1(new_n585_), .A2(KEYINPUT61), .ZN(new_n587_) );
  NAND3_X1 g465 ( .A1(new_n586_), .A2(G898), .A3(new_n587_), .ZN(new_n588_) );
  NAND3_X1 g466 ( .A1(new_n506_), .A2(new_n124_), .A3(new_n508_), .ZN(new_n589_) );
  NAND2_X1 g467 ( .A1(new_n589_), .A2(new_n588_), .ZN(new_n590_) );
  NAND2_X1 g468 ( .A1(new_n129_), .A2(G953), .ZN(new_n591_) );
  XNOR2_X1 g469 ( .A(new_n183_), .B(G101), .ZN(new_n592_) );
  XNOR2_X1 g470 ( .A(new_n592_), .B(new_n151_), .ZN(new_n593_) );
  NAND2_X1 g471 ( .A1(new_n593_), .A2(new_n591_), .ZN(new_n594_) );
  XOR2_X1 g472 ( .A(new_n590_), .B(new_n594_), .Z(G69) );
  XNOR2_X1 g473 ( .A(new_n178_), .B(new_n215_), .ZN(new_n596_) );
  XNOR2_X1 g474 ( .A(new_n596_), .B(new_n283_), .ZN(new_n597_) );
  XOR2_X1 g475 ( .A(new_n493_), .B(new_n597_), .Z(new_n598_) );
  NAND2_X1 g476 ( .A1(new_n598_), .A2(new_n124_), .ZN(new_n599_) );
  XNOR2_X1 g477 ( .A(new_n597_), .B(G227), .ZN(new_n600_) );
  NAND2_X1 g478 ( .A1(new_n600_), .A2(G900), .ZN(new_n601_) );
  NAND2_X1 g479 ( .A1(new_n601_), .A2(G953), .ZN(new_n602_) );
  NAND2_X1 g480 ( .A1(new_n599_), .A2(new_n602_), .ZN(G72) );
  NOR2_X1 g481 ( .A1(new_n135_), .A2(new_n301_), .ZN(new_n604_) );
  NAND3_X1 g482 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n604_), .ZN(new_n605_) );
  NAND2_X1 g483 ( .A1(new_n319_), .A2(new_n320_), .ZN(new_n606_) );
  XOR2_X1 g484 ( .A(new_n606_), .B(KEYINPUT62), .Z(new_n607_) );
  INV_X1 g485 ( .A(new_n607_), .ZN(new_n608_) );
  NAND2_X1 g486 ( .A1(new_n605_), .A2(new_n608_), .ZN(new_n609_) );
  NAND4_X1 g487 ( .A1(new_n510_), .A2(new_n511_), .A3(new_n604_), .A4(new_n607_), .ZN(new_n610_) );
  NAND3_X1 g488 ( .A1(new_n609_), .A2(new_n540_), .A3(new_n610_), .ZN(new_n611_) );
  NAND2_X1 g489 ( .A1(new_n611_), .A2(KEYINPUT63), .ZN(new_n612_) );
  INV_X1 g490 ( .A(KEYINPUT63), .ZN(new_n613_) );
  NAND4_X1 g491 ( .A1(new_n609_), .A2(new_n613_), .A3(new_n540_), .A4(new_n610_), .ZN(new_n614_) );
  NAND2_X1 g492 ( .A1(new_n612_), .A2(new_n614_), .ZN(G57) );
endmodule


