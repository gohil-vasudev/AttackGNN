module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743;

  OR2_X1 U8014 ( .A1(n16335), .A2(n8935), .ZN(n7950) );
  OR2_X1 U8015 ( .A1(operation_1_), .A2(operation_0_), .ZN(n7951) );
  OR2_X1 U8016 ( .A1(n16560), .A2(operation_0_), .ZN(n7952) );
  INV_X2 U8017 ( .A(b_15_), .ZN(n8951) );
  INV_X2 U8018 ( .A(b_7_), .ZN(n8667) );
  INV_X2 U8019 ( .A(b_23_), .ZN(n8940) );
  INV_X2 U8020 ( .A(b_6_), .ZN(n8963) );
  INV_X2 U8021 ( .A(b_8_), .ZN(n8961) );
  AND2_X2 U8022 ( .A1(n16557), .A2(n16558), .ZN(n7956) );
  INV_X1 U8023 ( .A(n7950), .ZN(n7953) );
  INV_X2 U8024 ( .A(n7951), .ZN(n7954) );
  INV_X4 U8025 ( .A(a_20_), .ZN(n8944) );
  INV_X4 U8026 ( .A(a_24_), .ZN(n8939) );
  NAND2_X4 U8027 ( .A1(operation_0_), .A2(n16560), .ZN(n8013) );
  INV_X4 U8028 ( .A(n7952), .ZN(n7955) );
  AND2_X4 U8029 ( .A1(operation_0_), .A2(operation_1_), .ZN(n7959) );
  INV_X2 U8030 ( .A(b_5_), .ZN(n8964) );
  INV_X2 U8031 ( .A(b_27_), .ZN(n8102) );
  INV_X2 U8032 ( .A(b_25_), .ZN(n8938) );
  INV_X2 U8033 ( .A(b_29_), .ZN(n8936) );
  INV_X2 U8034 ( .A(b_0_), .ZN(n8975) );
  INV_X2 U8035 ( .A(b_13_), .ZN(n8954) );
  INV_X2 U8036 ( .A(b_17_), .ZN(n8948) );
  INV_X2 U8037 ( .A(b_24_), .ZN(n8185) );
  INV_X2 U8038 ( .A(b_22_), .ZN(n8240) );
  INV_X2 U8039 ( .A(b_19_), .ZN(n8945) );
  INV_X2 U8040 ( .A(b_4_), .ZN(n8965) );
  NAND2_X2 U8041 ( .A1(a_30_), .A2(n16335), .ZN(n9341) );
  INV_X2 U8042 ( .A(b_26_), .ZN(n8130) );
  NAND2_X2 U8043 ( .A1(a_31_), .A2(n8935), .ZN(n8003) );
  INV_X2 U8044 ( .A(b_28_), .ZN(n8069) );
  INV_X2 U8045 ( .A(b_21_), .ZN(n8942) );
  INV_X2 U8046 ( .A(a_25_), .ZN(n8158) );
  INV_X2 U8047 ( .A(a_28_), .ZN(n8055) );
  INV_X2 U8048 ( .A(a_2_), .ZN(n8792) );
  INV_X2 U8049 ( .A(b_31_), .ZN(n7999) );
  INV_X2 U8050 ( .A(a_23_), .ZN(n8213) );
  INV_X2 U8051 ( .A(a_6_), .ZN(n8681) );
  INV_X2 U8052 ( .A(a_7_), .ZN(n8962) );
  INV_X2 U8053 ( .A(a_29_), .ZN(n8041) );
  INV_X2 U8054 ( .A(a_17_), .ZN(n8385) );
  INV_X2 U8055 ( .A(a_15_), .ZN(n8440) );
  INV_X2 U8056 ( .A(a_13_), .ZN(n8495) );
  INV_X2 U8057 ( .A(a_14_), .ZN(n8953) );
  INV_X2 U8058 ( .A(a_21_), .ZN(n8268) );
  INV_X2 U8059 ( .A(a_19_), .ZN(n8324) );
  INV_X2 U8060 ( .A(a_12_), .ZN(n8956) );
  INV_X2 U8061 ( .A(a_9_), .ZN(n8605) );
  INV_X2 U8062 ( .A(a_3_), .ZN(n8778) );
  INV_X2 U8063 ( .A(a_0_), .ZN(n8974) );
  INV_X2 U8064 ( .A(b_30_), .ZN(n8002) );
  INV_X2 U8065 ( .A(a_4_), .ZN(n8966) );
  INV_X2 U8066 ( .A(a_11_), .ZN(n8550) );
  INV_X2 U8067 ( .A(a_10_), .ZN(n8959) );
  INV_X2 U8068 ( .A(a_18_), .ZN(n8947) );
  INV_X2 U8069 ( .A(a_16_), .ZN(n8950) );
  INV_X2 U8070 ( .A(a_8_), .ZN(n8619) );
  INV_X2 U8071 ( .A(a_5_), .ZN(n8723) );
  INV_X2 U8072 ( .A(a_22_), .ZN(n8941) );
  INV_X2 U8073 ( .A(a_1_), .ZN(n8969) );
  NAND2_X1 U8074 ( .A1(n7956), .A2(n7957), .ZN(Result_9_) );
  NAND2_X1 U8075 ( .A1(n7958), .A2(n7959), .ZN(n7957) );
  XOR2_X1 U8076 ( .A(n7960), .B(n7961), .Z(n7958) );
  AND2_X1 U8077 ( .A1(n7962), .A2(n7963), .ZN(n7961) );
  NAND2_X1 U8078 ( .A1(n7956), .A2(n7964), .ZN(Result_8_) );
  NAND2_X1 U8079 ( .A1(n7965), .A2(n7959), .ZN(n7964) );
  XOR2_X1 U8080 ( .A(n7966), .B(n7967), .Z(n7965) );
  AND2_X1 U8081 ( .A1(n7968), .A2(n7969), .ZN(n7967) );
  NAND2_X1 U8082 ( .A1(n7956), .A2(n7970), .ZN(Result_7_) );
  NAND2_X1 U8083 ( .A1(n7971), .A2(n7959), .ZN(n7970) );
  XOR2_X1 U8084 ( .A(n7972), .B(n7973), .Z(n7971) );
  AND2_X1 U8085 ( .A1(n7974), .A2(n7975), .ZN(n7973) );
  NAND2_X1 U8086 ( .A1(n7956), .A2(n7976), .ZN(Result_6_) );
  NAND2_X1 U8087 ( .A1(n7977), .A2(n7959), .ZN(n7976) );
  XOR2_X1 U8088 ( .A(n7978), .B(n7979), .Z(n7977) );
  AND2_X1 U8089 ( .A1(n7980), .A2(n7981), .ZN(n7979) );
  NAND2_X1 U8090 ( .A1(n7982), .A2(n7983), .ZN(Result_63_) );
  NAND2_X1 U8091 ( .A1(n7984), .A2(n7959), .ZN(n7983) );
  NAND2_X1 U8092 ( .A1(n7985), .A2(n7986), .ZN(n7982) );
  NAND2_X1 U8093 ( .A1(n7987), .A2(n7951), .ZN(n7986) );
  NOR2_X1 U8094 ( .A1(n7955), .A2(n7988), .ZN(n7987) );
  NAND2_X1 U8095 ( .A1(n7989), .A2(n7990), .ZN(n7985) );
  NAND2_X1 U8096 ( .A1(n7991), .A2(n7992), .ZN(Result_62_) );
  NAND2_X1 U8097 ( .A1(n7959), .A2(n7993), .ZN(n7992) );
  NAND2_X1 U8098 ( .A1(n7994), .A2(n7995), .ZN(n7993) );
  NAND2_X1 U8099 ( .A1(n7996), .A2(a_30_), .ZN(n7995) );
  NOR2_X1 U8100 ( .A1(n7997), .A2(n7998), .ZN(n7994) );
  NOR2_X1 U8101 ( .A1(n7999), .A2(n8000), .ZN(n7998) );
  NOR2_X1 U8102 ( .A1(n8001), .A2(n8002), .ZN(n7997) );
  AND2_X1 U8103 ( .A1(n8003), .A2(n7989), .ZN(n8001) );
  NOR2_X1 U8104 ( .A1(n8004), .A2(n8005), .ZN(n7991) );
  NOR2_X1 U8105 ( .A1(n8006), .A2(n8007), .ZN(n8005) );
  NOR2_X1 U8106 ( .A1(n8008), .A2(n8009), .ZN(n8006) );
  NAND2_X1 U8107 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  NAND2_X1 U8108 ( .A1(n7954), .A2(n7984), .ZN(n8011) );
  INV_X1 U8109 ( .A(n8012), .ZN(n7984) );
  NAND2_X1 U8110 ( .A1(n7996), .A2(n7955), .ZN(n8010) );
  INV_X1 U8111 ( .A(n7990), .ZN(n7996) );
  NOR2_X1 U8112 ( .A1(n8013), .A2(n7989), .ZN(n8008) );
  NOR2_X1 U8113 ( .A1(n8014), .A2(n8015), .ZN(n8004) );
  NOR2_X1 U8114 ( .A1(n8016), .A2(n8017), .ZN(n8015) );
  NAND2_X1 U8115 ( .A1(n8018), .A2(n8019), .ZN(n8017) );
  NAND2_X1 U8116 ( .A1(n7954), .A2(n8012), .ZN(n8019) );
  NAND2_X1 U8117 ( .A1(n7955), .A2(n7990), .ZN(n8018) );
  AND2_X1 U8118 ( .A1(n7989), .A2(n7988), .ZN(n8016) );
  INV_X1 U8119 ( .A(n8007), .ZN(n8014) );
  NAND2_X1 U8120 ( .A1(n8000), .A2(n8020), .ZN(n8007) );
  NAND2_X1 U8121 ( .A1(n8021), .A2(n8022), .ZN(Result_61_) );
  NAND2_X1 U8122 ( .A1(n8023), .A2(n7959), .ZN(n8022) );
  XOR2_X1 U8123 ( .A(n8024), .B(n8025), .Z(n8023) );
  XOR2_X1 U8124 ( .A(n8026), .B(n8027), .Z(n8024) );
  NOR2_X1 U8125 ( .A1(n8028), .A2(n8029), .ZN(n8021) );
  NOR2_X1 U8126 ( .A1(n8030), .A2(n8031), .ZN(n8029) );
  NOR2_X1 U8127 ( .A1(n8032), .A2(n8033), .ZN(n8030) );
  NAND2_X1 U8128 ( .A1(n8034), .A2(n8035), .ZN(n8033) );
  NAND2_X1 U8129 ( .A1(n7954), .A2(n8036), .ZN(n8035) );
  NAND2_X1 U8130 ( .A1(n7955), .A2(n8037), .ZN(n8034) );
  NOR2_X1 U8131 ( .A1(n8038), .A2(n8013), .ZN(n8032) );
  NOR2_X1 U8132 ( .A1(n8039), .A2(n8040), .ZN(n8028) );
  INV_X1 U8133 ( .A(n8031), .ZN(n8040) );
  XNOR2_X1 U8134 ( .A(n8041), .B(b_29_), .ZN(n8031) );
  NOR2_X1 U8135 ( .A1(n8042), .A2(n8043), .ZN(n8039) );
  NAND2_X1 U8136 ( .A1(n8044), .A2(n8045), .ZN(n8043) );
  OR2_X1 U8137 ( .A1(n8036), .A2(n7951), .ZN(n8045) );
  NAND2_X1 U8138 ( .A1(n7955), .A2(n8046), .ZN(n8044) );
  NOR2_X1 U8139 ( .A1(n8047), .A2(n8013), .ZN(n8042) );
  NAND2_X1 U8140 ( .A1(n8048), .A2(n8049), .ZN(Result_60_) );
  NAND2_X1 U8141 ( .A1(n7959), .A2(n8050), .ZN(n8049) );
  XNOR2_X1 U8142 ( .A(n8051), .B(n8052), .ZN(n8050) );
  XNOR2_X1 U8143 ( .A(n8053), .B(n8054), .ZN(n8052) );
  NOR2_X1 U8144 ( .A1(n7999), .A2(n8055), .ZN(n8054) );
  NOR2_X1 U8145 ( .A1(n8056), .A2(n8057), .ZN(n8048) );
  NOR2_X1 U8146 ( .A1(n8058), .A2(n8059), .ZN(n8057) );
  NOR2_X1 U8147 ( .A1(n8060), .A2(n8061), .ZN(n8058) );
  NAND2_X1 U8148 ( .A1(n8062), .A2(n8063), .ZN(n8061) );
  NAND2_X1 U8149 ( .A1(n7954), .A2(n8064), .ZN(n8063) );
  NAND2_X1 U8150 ( .A1(n7955), .A2(n8065), .ZN(n8062) );
  NOR2_X1 U8151 ( .A1(n8066), .A2(n8013), .ZN(n8060) );
  NOR2_X1 U8152 ( .A1(n8067), .A2(n8068), .ZN(n8056) );
  INV_X1 U8153 ( .A(n8059), .ZN(n8068) );
  XNOR2_X1 U8154 ( .A(n8069), .B(a_28_), .ZN(n8059) );
  NOR2_X1 U8155 ( .A1(n8070), .A2(n8071), .ZN(n8067) );
  NAND2_X1 U8156 ( .A1(n8072), .A2(n8073), .ZN(n8071) );
  OR2_X1 U8157 ( .A1(n8064), .A2(n7951), .ZN(n8073) );
  NAND2_X1 U8158 ( .A1(n7955), .A2(n8074), .ZN(n8072) );
  NOR2_X1 U8159 ( .A1(n8075), .A2(n8013), .ZN(n8070) );
  NAND2_X1 U8160 ( .A1(n7956), .A2(n8076), .ZN(Result_5_) );
  NAND2_X1 U8161 ( .A1(n8077), .A2(n7959), .ZN(n8076) );
  XOR2_X1 U8162 ( .A(n8078), .B(n8079), .Z(n8077) );
  AND2_X1 U8163 ( .A1(n8080), .A2(n8081), .ZN(n8079) );
  NAND2_X1 U8164 ( .A1(n8082), .A2(n8083), .ZN(Result_59_) );
  NAND2_X1 U8165 ( .A1(n8084), .A2(n7959), .ZN(n8083) );
  XNOR2_X1 U8166 ( .A(n8085), .B(n8086), .ZN(n8084) );
  XOR2_X1 U8167 ( .A(n8087), .B(n8088), .Z(n8086) );
  NAND2_X1 U8168 ( .A1(a_27_), .A2(b_31_), .ZN(n8088) );
  NOR2_X1 U8169 ( .A1(n8089), .A2(n8090), .ZN(n8082) );
  NOR2_X1 U8170 ( .A1(n8091), .A2(n8092), .ZN(n8090) );
  NOR2_X1 U8171 ( .A1(n8093), .A2(n8094), .ZN(n8091) );
  NAND2_X1 U8172 ( .A1(n8095), .A2(n8096), .ZN(n8094) );
  NAND2_X1 U8173 ( .A1(n7954), .A2(n8097), .ZN(n8096) );
  NAND2_X1 U8174 ( .A1(n7955), .A2(n8098), .ZN(n8095) );
  NOR2_X1 U8175 ( .A1(n8099), .A2(n8013), .ZN(n8093) );
  NOR2_X1 U8176 ( .A1(n8100), .A2(n8101), .ZN(n8089) );
  INV_X1 U8177 ( .A(n8092), .ZN(n8101) );
  XNOR2_X1 U8178 ( .A(n8102), .B(a_27_), .ZN(n8092) );
  NOR2_X1 U8179 ( .A1(n8103), .A2(n8104), .ZN(n8100) );
  NAND2_X1 U8180 ( .A1(n8105), .A2(n8106), .ZN(n8104) );
  OR2_X1 U8181 ( .A1(n8097), .A2(n7951), .ZN(n8106) );
  NAND2_X1 U8182 ( .A1(n7955), .A2(n8107), .ZN(n8105) );
  NOR2_X1 U8183 ( .A1(n8108), .A2(n8013), .ZN(n8103) );
  NAND2_X1 U8184 ( .A1(n8109), .A2(n8110), .ZN(Result_58_) );
  NAND2_X1 U8185 ( .A1(n8111), .A2(n7959), .ZN(n8110) );
  XOR2_X1 U8186 ( .A(n8112), .B(n8113), .Z(n8111) );
  XOR2_X1 U8187 ( .A(n8114), .B(n8115), .Z(n8112) );
  NOR2_X1 U8188 ( .A1(n7999), .A2(n8116), .ZN(n8115) );
  NOR2_X1 U8189 ( .A1(n8117), .A2(n8118), .ZN(n8109) );
  NOR2_X1 U8190 ( .A1(n8119), .A2(n8120), .ZN(n8118) );
  NOR2_X1 U8191 ( .A1(n8121), .A2(n8122), .ZN(n8119) );
  NAND2_X1 U8192 ( .A1(n8123), .A2(n8124), .ZN(n8122) );
  NAND2_X1 U8193 ( .A1(n7954), .A2(n8125), .ZN(n8124) );
  NAND2_X1 U8194 ( .A1(n7955), .A2(n8126), .ZN(n8123) );
  NOR2_X1 U8195 ( .A1(n8127), .A2(n8013), .ZN(n8121) );
  NOR2_X1 U8196 ( .A1(n8128), .A2(n8129), .ZN(n8117) );
  INV_X1 U8197 ( .A(n8120), .ZN(n8129) );
  XNOR2_X1 U8198 ( .A(n8130), .B(a_26_), .ZN(n8120) );
  NOR2_X1 U8199 ( .A1(n8131), .A2(n8132), .ZN(n8128) );
  NAND2_X1 U8200 ( .A1(n8133), .A2(n8134), .ZN(n8132) );
  NAND2_X1 U8201 ( .A1(n8135), .A2(n7954), .ZN(n8134) );
  NAND2_X1 U8202 ( .A1(n7955), .A2(n8136), .ZN(n8133) );
  NOR2_X1 U8203 ( .A1(n8137), .A2(n8013), .ZN(n8131) );
  NAND2_X1 U8204 ( .A1(n8138), .A2(n8139), .ZN(Result_57_) );
  NAND2_X1 U8205 ( .A1(n7959), .A2(n8140), .ZN(n8139) );
  XNOR2_X1 U8206 ( .A(n8141), .B(n8142), .ZN(n8140) );
  NAND2_X1 U8207 ( .A1(n8143), .A2(n8144), .ZN(n8141) );
  NOR2_X1 U8208 ( .A1(n8145), .A2(n8146), .ZN(n8138) );
  NOR2_X1 U8209 ( .A1(n8147), .A2(n8148), .ZN(n8146) );
  NOR2_X1 U8210 ( .A1(n8149), .A2(n8150), .ZN(n8147) );
  NAND2_X1 U8211 ( .A1(n8151), .A2(n8152), .ZN(n8150) );
  NAND2_X1 U8212 ( .A1(n7954), .A2(n8153), .ZN(n8152) );
  NAND2_X1 U8213 ( .A1(n7955), .A2(n8154), .ZN(n8151) );
  NOR2_X1 U8214 ( .A1(n8155), .A2(n8013), .ZN(n8149) );
  NOR2_X1 U8215 ( .A1(n8156), .A2(n8157), .ZN(n8145) );
  INV_X1 U8216 ( .A(n8148), .ZN(n8157) );
  XNOR2_X1 U8217 ( .A(n8158), .B(b_25_), .ZN(n8148) );
  NOR2_X1 U8218 ( .A1(n8159), .A2(n8160), .ZN(n8156) );
  NAND2_X1 U8219 ( .A1(n8161), .A2(n8162), .ZN(n8160) );
  OR2_X1 U8220 ( .A1(n8153), .A2(n7951), .ZN(n8162) );
  NAND2_X1 U8221 ( .A1(n7955), .A2(n8163), .ZN(n8161) );
  NOR2_X1 U8222 ( .A1(n8164), .A2(n8013), .ZN(n8159) );
  NAND2_X1 U8223 ( .A1(n8165), .A2(n8166), .ZN(Result_56_) );
  NAND2_X1 U8224 ( .A1(n7959), .A2(n8167), .ZN(n8166) );
  XOR2_X1 U8225 ( .A(n8168), .B(n8169), .Z(n8167) );
  XNOR2_X1 U8226 ( .A(n8170), .B(n8171), .ZN(n8169) );
  NAND2_X1 U8227 ( .A1(a_24_), .A2(b_31_), .ZN(n8170) );
  NOR2_X1 U8228 ( .A1(n8172), .A2(n8173), .ZN(n8165) );
  NOR2_X1 U8229 ( .A1(n8174), .A2(n8175), .ZN(n8173) );
  NOR2_X1 U8230 ( .A1(n8176), .A2(n8177), .ZN(n8174) );
  NAND2_X1 U8231 ( .A1(n8178), .A2(n8179), .ZN(n8177) );
  NAND2_X1 U8232 ( .A1(n7954), .A2(n8180), .ZN(n8179) );
  NAND2_X1 U8233 ( .A1(n7955), .A2(n8181), .ZN(n8178) );
  NOR2_X1 U8234 ( .A1(n8182), .A2(n8013), .ZN(n8176) );
  NOR2_X1 U8235 ( .A1(n8183), .A2(n8184), .ZN(n8172) );
  INV_X1 U8236 ( .A(n8175), .ZN(n8184) );
  XNOR2_X1 U8237 ( .A(n8185), .B(a_24_), .ZN(n8175) );
  NOR2_X1 U8238 ( .A1(n8186), .A2(n8187), .ZN(n8183) );
  NAND2_X1 U8239 ( .A1(n8188), .A2(n8189), .ZN(n8187) );
  NAND2_X1 U8240 ( .A1(n8190), .A2(n7954), .ZN(n8189) );
  NAND2_X1 U8241 ( .A1(n7955), .A2(n8191), .ZN(n8188) );
  NOR2_X1 U8242 ( .A1(n8192), .A2(n8013), .ZN(n8186) );
  NAND2_X1 U8243 ( .A1(n8193), .A2(n8194), .ZN(Result_55_) );
  NAND2_X1 U8244 ( .A1(n8195), .A2(n7959), .ZN(n8194) );
  XNOR2_X1 U8245 ( .A(n8196), .B(n8197), .ZN(n8195) );
  NAND2_X1 U8246 ( .A1(n8198), .A2(n8199), .ZN(n8196) );
  NOR2_X1 U8247 ( .A1(n8200), .A2(n8201), .ZN(n8193) );
  NOR2_X1 U8248 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  NOR2_X1 U8249 ( .A1(n8204), .A2(n8205), .ZN(n8202) );
  NAND2_X1 U8250 ( .A1(n8206), .A2(n8207), .ZN(n8205) );
  NAND2_X1 U8251 ( .A1(n7954), .A2(n8208), .ZN(n8207) );
  NAND2_X1 U8252 ( .A1(n7955), .A2(n8209), .ZN(n8206) );
  NOR2_X1 U8253 ( .A1(n8210), .A2(n8013), .ZN(n8204) );
  NOR2_X1 U8254 ( .A1(n8211), .A2(n8212), .ZN(n8200) );
  INV_X1 U8255 ( .A(n8203), .ZN(n8212) );
  XNOR2_X1 U8256 ( .A(n8213), .B(b_23_), .ZN(n8203) );
  NOR2_X1 U8257 ( .A1(n8214), .A2(n8215), .ZN(n8211) );
  NAND2_X1 U8258 ( .A1(n8216), .A2(n8217), .ZN(n8215) );
  OR2_X1 U8259 ( .A1(n8208), .A2(n7951), .ZN(n8217) );
  NAND2_X1 U8260 ( .A1(n7955), .A2(n8218), .ZN(n8216) );
  NOR2_X1 U8261 ( .A1(n8219), .A2(n8013), .ZN(n8214) );
  NAND2_X1 U8262 ( .A1(n8220), .A2(n8221), .ZN(Result_54_) );
  NAND2_X1 U8263 ( .A1(n7959), .A2(n8222), .ZN(n8221) );
  XNOR2_X1 U8264 ( .A(n8223), .B(n8224), .ZN(n8222) );
  XOR2_X1 U8265 ( .A(n8225), .B(n8226), .Z(n8224) );
  NAND2_X1 U8266 ( .A1(a_22_), .A2(b_31_), .ZN(n8226) );
  NOR2_X1 U8267 ( .A1(n8227), .A2(n8228), .ZN(n8220) );
  NOR2_X1 U8268 ( .A1(n8229), .A2(n8230), .ZN(n8228) );
  NOR2_X1 U8269 ( .A1(n8231), .A2(n8232), .ZN(n8229) );
  NAND2_X1 U8270 ( .A1(n8233), .A2(n8234), .ZN(n8232) );
  NAND2_X1 U8271 ( .A1(n7954), .A2(n8235), .ZN(n8234) );
  NAND2_X1 U8272 ( .A1(n7955), .A2(n8236), .ZN(n8233) );
  NOR2_X1 U8273 ( .A1(n8237), .A2(n8013), .ZN(n8231) );
  NOR2_X1 U8274 ( .A1(n8238), .A2(n8239), .ZN(n8227) );
  INV_X1 U8275 ( .A(n8230), .ZN(n8239) );
  XNOR2_X1 U8276 ( .A(n8240), .B(a_22_), .ZN(n8230) );
  NOR2_X1 U8277 ( .A1(n8241), .A2(n8242), .ZN(n8238) );
  NAND2_X1 U8278 ( .A1(n8243), .A2(n8244), .ZN(n8242) );
  NAND2_X1 U8279 ( .A1(n8245), .A2(n7954), .ZN(n8244) );
  NAND2_X1 U8280 ( .A1(n7955), .A2(n8246), .ZN(n8243) );
  NOR2_X1 U8281 ( .A1(n8247), .A2(n8013), .ZN(n8241) );
  NAND2_X1 U8282 ( .A1(n8248), .A2(n8249), .ZN(Result_53_) );
  NAND2_X1 U8283 ( .A1(n7959), .A2(n8250), .ZN(n8249) );
  XNOR2_X1 U8284 ( .A(n8251), .B(n8252), .ZN(n8250) );
  XOR2_X1 U8285 ( .A(n8253), .B(n8254), .Z(n8252) );
  NAND2_X1 U8286 ( .A1(a_21_), .A2(b_31_), .ZN(n8254) );
  NOR2_X1 U8287 ( .A1(n8255), .A2(n8256), .ZN(n8248) );
  NOR2_X1 U8288 ( .A1(n8257), .A2(n8258), .ZN(n8256) );
  NOR2_X1 U8289 ( .A1(n8259), .A2(n8260), .ZN(n8257) );
  NAND2_X1 U8290 ( .A1(n8261), .A2(n8262), .ZN(n8260) );
  NAND2_X1 U8291 ( .A1(n7954), .A2(n8263), .ZN(n8262) );
  NAND2_X1 U8292 ( .A1(n7955), .A2(n8264), .ZN(n8261) );
  NOR2_X1 U8293 ( .A1(n8265), .A2(n8013), .ZN(n8259) );
  NOR2_X1 U8294 ( .A1(n8266), .A2(n8267), .ZN(n8255) );
  INV_X1 U8295 ( .A(n8258), .ZN(n8267) );
  XNOR2_X1 U8296 ( .A(n8268), .B(b_21_), .ZN(n8258) );
  NOR2_X1 U8297 ( .A1(n8269), .A2(n8270), .ZN(n8266) );
  NAND2_X1 U8298 ( .A1(n8271), .A2(n8272), .ZN(n8270) );
  OR2_X1 U8299 ( .A1(n8263), .A2(n7951), .ZN(n8272) );
  NAND2_X1 U8300 ( .A1(n7955), .A2(n8273), .ZN(n8271) );
  NOR2_X1 U8301 ( .A1(n8274), .A2(n8013), .ZN(n8269) );
  NAND2_X1 U8302 ( .A1(n8275), .A2(n8276), .ZN(Result_52_) );
  NAND2_X1 U8303 ( .A1(n7959), .A2(n8277), .ZN(n8276) );
  XNOR2_X1 U8304 ( .A(n8278), .B(n8279), .ZN(n8277) );
  XOR2_X1 U8305 ( .A(n8280), .B(n8281), .Z(n8279) );
  NAND2_X1 U8306 ( .A1(a_20_), .A2(b_31_), .ZN(n8281) );
  NOR2_X1 U8307 ( .A1(n8282), .A2(n8283), .ZN(n8275) );
  NOR2_X1 U8308 ( .A1(n8284), .A2(n8285), .ZN(n8283) );
  NOR2_X1 U8309 ( .A1(n8286), .A2(n8287), .ZN(n8284) );
  NAND2_X1 U8310 ( .A1(n8288), .A2(n8289), .ZN(n8287) );
  NAND2_X1 U8311 ( .A1(n8290), .A2(n7954), .ZN(n8289) );
  NAND2_X1 U8312 ( .A1(n7955), .A2(n8291), .ZN(n8288) );
  NOR2_X1 U8313 ( .A1(n8292), .A2(n8013), .ZN(n8286) );
  NOR2_X1 U8314 ( .A1(n8293), .A2(n8294), .ZN(n8282) );
  NOR2_X1 U8315 ( .A1(n8295), .A2(n8296), .ZN(n8294) );
  NAND2_X1 U8316 ( .A1(n8297), .A2(n8298), .ZN(n8296) );
  NAND2_X1 U8317 ( .A1(n7954), .A2(n8299), .ZN(n8298) );
  NAND2_X1 U8318 ( .A1(n7955), .A2(n8300), .ZN(n8297) );
  NOR2_X1 U8319 ( .A1(n8301), .A2(n8013), .ZN(n8295) );
  INV_X1 U8320 ( .A(n8285), .ZN(n8293) );
  NAND2_X1 U8321 ( .A1(n8302), .A2(n8303), .ZN(n8285) );
  NAND2_X1 U8322 ( .A1(n8304), .A2(n8305), .ZN(Result_51_) );
  NAND2_X1 U8323 ( .A1(n8306), .A2(n7959), .ZN(n8305) );
  XNOR2_X1 U8324 ( .A(n8307), .B(n8308), .ZN(n8306) );
  XNOR2_X1 U8325 ( .A(n8309), .B(n8310), .ZN(n8308) );
  NOR2_X1 U8326 ( .A1(n8311), .A2(n8312), .ZN(n8304) );
  NOR2_X1 U8327 ( .A1(n8313), .A2(n8314), .ZN(n8312) );
  NOR2_X1 U8328 ( .A1(n8315), .A2(n8316), .ZN(n8313) );
  NAND2_X1 U8329 ( .A1(n8317), .A2(n8318), .ZN(n8316) );
  NAND2_X1 U8330 ( .A1(n7954), .A2(n8319), .ZN(n8318) );
  NAND2_X1 U8331 ( .A1(n7955), .A2(n8320), .ZN(n8317) );
  NOR2_X1 U8332 ( .A1(n8321), .A2(n8013), .ZN(n8315) );
  NOR2_X1 U8333 ( .A1(n8322), .A2(n8323), .ZN(n8311) );
  INV_X1 U8334 ( .A(n8314), .ZN(n8323) );
  XNOR2_X1 U8335 ( .A(n8324), .B(b_19_), .ZN(n8314) );
  NOR2_X1 U8336 ( .A1(n8325), .A2(n8326), .ZN(n8322) );
  NAND2_X1 U8337 ( .A1(n8327), .A2(n8328), .ZN(n8326) );
  OR2_X1 U8338 ( .A1(n8319), .A2(n7951), .ZN(n8328) );
  NAND2_X1 U8339 ( .A1(n7955), .A2(n8329), .ZN(n8327) );
  NOR2_X1 U8340 ( .A1(n8330), .A2(n8013), .ZN(n8325) );
  NAND2_X1 U8341 ( .A1(n8331), .A2(n8332), .ZN(Result_50_) );
  NAND2_X1 U8342 ( .A1(n7959), .A2(n8333), .ZN(n8332) );
  XOR2_X1 U8343 ( .A(n8334), .B(n8335), .Z(n8333) );
  XNOR2_X1 U8344 ( .A(n8336), .B(n8337), .ZN(n8335) );
  NAND2_X1 U8345 ( .A1(a_18_), .A2(b_31_), .ZN(n8336) );
  NOR2_X1 U8346 ( .A1(n8338), .A2(n8339), .ZN(n8331) );
  NOR2_X1 U8347 ( .A1(n8340), .A2(n8341), .ZN(n8339) );
  NOR2_X1 U8348 ( .A1(n8342), .A2(n8343), .ZN(n8340) );
  NAND2_X1 U8349 ( .A1(n8344), .A2(n8345), .ZN(n8343) );
  OR2_X1 U8350 ( .A1(n8346), .A2(n7951), .ZN(n8345) );
  NAND2_X1 U8351 ( .A1(n7955), .A2(n8347), .ZN(n8344) );
  NOR2_X1 U8352 ( .A1(n8348), .A2(n8013), .ZN(n8342) );
  NOR2_X1 U8353 ( .A1(n8349), .A2(n8350), .ZN(n8338) );
  NOR2_X1 U8354 ( .A1(n8351), .A2(n8352), .ZN(n8350) );
  NAND2_X1 U8355 ( .A1(n8353), .A2(n8354), .ZN(n8352) );
  NAND2_X1 U8356 ( .A1(n7954), .A2(n8346), .ZN(n8354) );
  NAND2_X1 U8357 ( .A1(n7955), .A2(n8355), .ZN(n8353) );
  NOR2_X1 U8358 ( .A1(n8356), .A2(n8013), .ZN(n8351) );
  INV_X1 U8359 ( .A(n8341), .ZN(n8349) );
  NAND2_X1 U8360 ( .A1(n8357), .A2(n8358), .ZN(n8341) );
  NAND2_X1 U8361 ( .A1(n7956), .A2(n8359), .ZN(Result_4_) );
  NAND2_X1 U8362 ( .A1(n8360), .A2(n7959), .ZN(n8359) );
  XOR2_X1 U8363 ( .A(n8361), .B(n8362), .Z(n8360) );
  AND2_X1 U8364 ( .A1(n8363), .A2(n8364), .ZN(n8362) );
  NAND2_X1 U8365 ( .A1(n8365), .A2(n8366), .ZN(Result_49_) );
  NAND2_X1 U8366 ( .A1(n8367), .A2(n7959), .ZN(n8366) );
  XNOR2_X1 U8367 ( .A(n8368), .B(n8369), .ZN(n8367) );
  XNOR2_X1 U8368 ( .A(n8370), .B(n8371), .ZN(n8369) );
  NOR2_X1 U8369 ( .A1(n8372), .A2(n8373), .ZN(n8365) );
  NOR2_X1 U8370 ( .A1(n8374), .A2(n8375), .ZN(n8373) );
  NOR2_X1 U8371 ( .A1(n8376), .A2(n8377), .ZN(n8374) );
  NAND2_X1 U8372 ( .A1(n8378), .A2(n8379), .ZN(n8377) );
  NAND2_X1 U8373 ( .A1(n7954), .A2(n8380), .ZN(n8379) );
  NAND2_X1 U8374 ( .A1(n7955), .A2(n8381), .ZN(n8378) );
  NOR2_X1 U8375 ( .A1(n8382), .A2(n8013), .ZN(n8376) );
  NOR2_X1 U8376 ( .A1(n8383), .A2(n8384), .ZN(n8372) );
  INV_X1 U8377 ( .A(n8375), .ZN(n8384) );
  XNOR2_X1 U8378 ( .A(n8385), .B(b_17_), .ZN(n8375) );
  NOR2_X1 U8379 ( .A1(n8386), .A2(n8387), .ZN(n8383) );
  NAND2_X1 U8380 ( .A1(n8388), .A2(n8389), .ZN(n8387) );
  OR2_X1 U8381 ( .A1(n8380), .A2(n7951), .ZN(n8389) );
  NAND2_X1 U8382 ( .A1(n7955), .A2(n8390), .ZN(n8388) );
  NOR2_X1 U8383 ( .A1(n8391), .A2(n8013), .ZN(n8386) );
  NAND2_X1 U8384 ( .A1(n8392), .A2(n8393), .ZN(Result_48_) );
  NAND2_X1 U8385 ( .A1(n7959), .A2(n8394), .ZN(n8393) );
  XNOR2_X1 U8386 ( .A(n8395), .B(n8396), .ZN(n8394) );
  XOR2_X1 U8387 ( .A(n8397), .B(n8398), .Z(n8396) );
  NAND2_X1 U8388 ( .A1(a_16_), .A2(b_31_), .ZN(n8398) );
  NOR2_X1 U8389 ( .A1(n8399), .A2(n8400), .ZN(n8392) );
  NOR2_X1 U8390 ( .A1(n8401), .A2(n8402), .ZN(n8400) );
  NOR2_X1 U8391 ( .A1(n8403), .A2(n8404), .ZN(n8401) );
  NAND2_X1 U8392 ( .A1(n8405), .A2(n8406), .ZN(n8404) );
  OR2_X1 U8393 ( .A1(n8407), .A2(n7951), .ZN(n8406) );
  NAND2_X1 U8394 ( .A1(n7955), .A2(n8408), .ZN(n8405) );
  NOR2_X1 U8395 ( .A1(n8409), .A2(n8013), .ZN(n8403) );
  NOR2_X1 U8396 ( .A1(n8410), .A2(n8411), .ZN(n8399) );
  NOR2_X1 U8397 ( .A1(n8412), .A2(n8413), .ZN(n8411) );
  NAND2_X1 U8398 ( .A1(n8414), .A2(n8415), .ZN(n8413) );
  NAND2_X1 U8399 ( .A1(n7954), .A2(n8407), .ZN(n8415) );
  NAND2_X1 U8400 ( .A1(n7955), .A2(n8416), .ZN(n8414) );
  NOR2_X1 U8401 ( .A1(n8417), .A2(n8013), .ZN(n8412) );
  INV_X1 U8402 ( .A(n8402), .ZN(n8410) );
  NAND2_X1 U8403 ( .A1(n8418), .A2(n8419), .ZN(n8402) );
  NAND2_X1 U8404 ( .A1(n8420), .A2(n8421), .ZN(Result_47_) );
  NAND2_X1 U8405 ( .A1(n8422), .A2(n7959), .ZN(n8421) );
  XOR2_X1 U8406 ( .A(n8423), .B(n8424), .Z(n8422) );
  XOR2_X1 U8407 ( .A(n8425), .B(n8426), .Z(n8423) );
  NOR2_X1 U8408 ( .A1(n8427), .A2(n8428), .ZN(n8420) );
  NOR2_X1 U8409 ( .A1(n8429), .A2(n8430), .ZN(n8428) );
  NOR2_X1 U8410 ( .A1(n8431), .A2(n8432), .ZN(n8429) );
  NAND2_X1 U8411 ( .A1(n8433), .A2(n8434), .ZN(n8432) );
  NAND2_X1 U8412 ( .A1(n7954), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U8413 ( .A1(n7955), .A2(n8436), .ZN(n8433) );
  NOR2_X1 U8414 ( .A1(n8437), .A2(n8013), .ZN(n8431) );
  NOR2_X1 U8415 ( .A1(n8438), .A2(n8439), .ZN(n8427) );
  INV_X1 U8416 ( .A(n8430), .ZN(n8439) );
  XNOR2_X1 U8417 ( .A(n8440), .B(b_15_), .ZN(n8430) );
  NOR2_X1 U8418 ( .A1(n8441), .A2(n8442), .ZN(n8438) );
  NAND2_X1 U8419 ( .A1(n8443), .A2(n8444), .ZN(n8442) );
  OR2_X1 U8420 ( .A1(n8435), .A2(n7951), .ZN(n8444) );
  NAND2_X1 U8421 ( .A1(n7955), .A2(n8445), .ZN(n8443) );
  NOR2_X1 U8422 ( .A1(n8446), .A2(n8013), .ZN(n8441) );
  NAND2_X1 U8423 ( .A1(n8447), .A2(n8448), .ZN(Result_46_) );
  NAND2_X1 U8424 ( .A1(n7959), .A2(n8449), .ZN(n8448) );
  XNOR2_X1 U8425 ( .A(n8450), .B(n8451), .ZN(n8449) );
  XOR2_X1 U8426 ( .A(n8452), .B(n8453), .Z(n8451) );
  NAND2_X1 U8427 ( .A1(a_14_), .A2(b_31_), .ZN(n8453) );
  NOR2_X1 U8428 ( .A1(n8454), .A2(n8455), .ZN(n8447) );
  NOR2_X1 U8429 ( .A1(n8456), .A2(n8457), .ZN(n8455) );
  NOR2_X1 U8430 ( .A1(n8458), .A2(n8459), .ZN(n8456) );
  NAND2_X1 U8431 ( .A1(n8460), .A2(n8461), .ZN(n8459) );
  OR2_X1 U8432 ( .A1(n8462), .A2(n7951), .ZN(n8461) );
  NAND2_X1 U8433 ( .A1(n7955), .A2(n8463), .ZN(n8460) );
  NOR2_X1 U8434 ( .A1(n8464), .A2(n8013), .ZN(n8458) );
  NOR2_X1 U8435 ( .A1(n8465), .A2(n8466), .ZN(n8454) );
  NOR2_X1 U8436 ( .A1(n8467), .A2(n8468), .ZN(n8466) );
  NAND2_X1 U8437 ( .A1(n8469), .A2(n8470), .ZN(n8468) );
  NAND2_X1 U8438 ( .A1(n7954), .A2(n8462), .ZN(n8470) );
  NAND2_X1 U8439 ( .A1(n7955), .A2(n8471), .ZN(n8469) );
  NOR2_X1 U8440 ( .A1(n8472), .A2(n8013), .ZN(n8467) );
  INV_X1 U8441 ( .A(n8457), .ZN(n8465) );
  NAND2_X1 U8442 ( .A1(n8473), .A2(n8474), .ZN(n8457) );
  NAND2_X1 U8443 ( .A1(n8475), .A2(n8476), .ZN(Result_45_) );
  NAND2_X1 U8444 ( .A1(n8477), .A2(n7959), .ZN(n8476) );
  XOR2_X1 U8445 ( .A(n8478), .B(n8479), .Z(n8477) );
  XOR2_X1 U8446 ( .A(n8480), .B(n8481), .Z(n8478) );
  NOR2_X1 U8447 ( .A1(n8482), .A2(n8483), .ZN(n8475) );
  NOR2_X1 U8448 ( .A1(n8484), .A2(n8485), .ZN(n8483) );
  NOR2_X1 U8449 ( .A1(n8486), .A2(n8487), .ZN(n8484) );
  NAND2_X1 U8450 ( .A1(n8488), .A2(n8489), .ZN(n8487) );
  NAND2_X1 U8451 ( .A1(n7954), .A2(n8490), .ZN(n8489) );
  NAND2_X1 U8452 ( .A1(n7955), .A2(n8491), .ZN(n8488) );
  NOR2_X1 U8453 ( .A1(n8492), .A2(n8013), .ZN(n8486) );
  NOR2_X1 U8454 ( .A1(n8493), .A2(n8494), .ZN(n8482) );
  INV_X1 U8455 ( .A(n8485), .ZN(n8494) );
  XNOR2_X1 U8456 ( .A(n8495), .B(b_13_), .ZN(n8485) );
  NOR2_X1 U8457 ( .A1(n8496), .A2(n8497), .ZN(n8493) );
  NAND2_X1 U8458 ( .A1(n8498), .A2(n8499), .ZN(n8497) );
  OR2_X1 U8459 ( .A1(n8490), .A2(n7951), .ZN(n8499) );
  NAND2_X1 U8460 ( .A1(n7955), .A2(n8500), .ZN(n8498) );
  NOR2_X1 U8461 ( .A1(n8501), .A2(n8013), .ZN(n8496) );
  NAND2_X1 U8462 ( .A1(n8502), .A2(n8503), .ZN(Result_44_) );
  NAND2_X1 U8463 ( .A1(n7959), .A2(n8504), .ZN(n8503) );
  XNOR2_X1 U8464 ( .A(n8505), .B(n8506), .ZN(n8504) );
  XOR2_X1 U8465 ( .A(n8507), .B(n8508), .Z(n8506) );
  NAND2_X1 U8466 ( .A1(a_12_), .A2(b_31_), .ZN(n8508) );
  NOR2_X1 U8467 ( .A1(n8509), .A2(n8510), .ZN(n8502) );
  NOR2_X1 U8468 ( .A1(n8511), .A2(n8512), .ZN(n8510) );
  NOR2_X1 U8469 ( .A1(n8513), .A2(n8514), .ZN(n8511) );
  NAND2_X1 U8470 ( .A1(n8515), .A2(n8516), .ZN(n8514) );
  OR2_X1 U8471 ( .A1(n8517), .A2(n7951), .ZN(n8516) );
  NAND2_X1 U8472 ( .A1(n7955), .A2(n8518), .ZN(n8515) );
  NOR2_X1 U8473 ( .A1(n8519), .A2(n8013), .ZN(n8513) );
  NOR2_X1 U8474 ( .A1(n8520), .A2(n8521), .ZN(n8509) );
  NOR2_X1 U8475 ( .A1(n8522), .A2(n8523), .ZN(n8521) );
  NAND2_X1 U8476 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  NAND2_X1 U8477 ( .A1(n7954), .A2(n8517), .ZN(n8525) );
  NAND2_X1 U8478 ( .A1(n7955), .A2(n8526), .ZN(n8524) );
  NOR2_X1 U8479 ( .A1(n8527), .A2(n8013), .ZN(n8522) );
  INV_X1 U8480 ( .A(n8512), .ZN(n8520) );
  NAND2_X1 U8481 ( .A1(n8528), .A2(n8529), .ZN(n8512) );
  NAND2_X1 U8482 ( .A1(n8530), .A2(n8531), .ZN(Result_43_) );
  NAND2_X1 U8483 ( .A1(n8532), .A2(n7959), .ZN(n8531) );
  XOR2_X1 U8484 ( .A(n8533), .B(n8534), .Z(n8532) );
  XOR2_X1 U8485 ( .A(n8535), .B(n8536), .Z(n8533) );
  NOR2_X1 U8486 ( .A1(n8537), .A2(n8538), .ZN(n8530) );
  NOR2_X1 U8487 ( .A1(n8539), .A2(n8540), .ZN(n8538) );
  NOR2_X1 U8488 ( .A1(n8541), .A2(n8542), .ZN(n8539) );
  NAND2_X1 U8489 ( .A1(n8543), .A2(n8544), .ZN(n8542) );
  NAND2_X1 U8490 ( .A1(n7954), .A2(n8545), .ZN(n8544) );
  NAND2_X1 U8491 ( .A1(n7955), .A2(n8546), .ZN(n8543) );
  NOR2_X1 U8492 ( .A1(n8547), .A2(n8013), .ZN(n8541) );
  NOR2_X1 U8493 ( .A1(n8548), .A2(n8549), .ZN(n8537) );
  INV_X1 U8494 ( .A(n8540), .ZN(n8549) );
  XNOR2_X1 U8495 ( .A(n8550), .B(b_11_), .ZN(n8540) );
  NOR2_X1 U8496 ( .A1(n8551), .A2(n8552), .ZN(n8548) );
  NAND2_X1 U8497 ( .A1(n8553), .A2(n8554), .ZN(n8552) );
  OR2_X1 U8498 ( .A1(n8545), .A2(n7951), .ZN(n8554) );
  NAND2_X1 U8499 ( .A1(n7955), .A2(n8555), .ZN(n8553) );
  NOR2_X1 U8500 ( .A1(n8556), .A2(n8013), .ZN(n8551) );
  NAND2_X1 U8501 ( .A1(n8557), .A2(n8558), .ZN(Result_42_) );
  NAND2_X1 U8502 ( .A1(n7959), .A2(n8559), .ZN(n8558) );
  XNOR2_X1 U8503 ( .A(n8560), .B(n8561), .ZN(n8559) );
  XOR2_X1 U8504 ( .A(n8562), .B(n8563), .Z(n8561) );
  NAND2_X1 U8505 ( .A1(a_10_), .A2(b_31_), .ZN(n8563) );
  NOR2_X1 U8506 ( .A1(n8564), .A2(n8565), .ZN(n8557) );
  NOR2_X1 U8507 ( .A1(n8566), .A2(n8567), .ZN(n8565) );
  NOR2_X1 U8508 ( .A1(n8568), .A2(n8569), .ZN(n8566) );
  NAND2_X1 U8509 ( .A1(n8570), .A2(n8571), .ZN(n8569) );
  OR2_X1 U8510 ( .A1(n8572), .A2(n7951), .ZN(n8571) );
  NAND2_X1 U8511 ( .A1(n7955), .A2(n8573), .ZN(n8570) );
  NOR2_X1 U8512 ( .A1(n8574), .A2(n8013), .ZN(n8568) );
  NOR2_X1 U8513 ( .A1(n8575), .A2(n8576), .ZN(n8564) );
  NOR2_X1 U8514 ( .A1(n8577), .A2(n8578), .ZN(n8576) );
  NAND2_X1 U8515 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
  NAND2_X1 U8516 ( .A1(n7954), .A2(n8572), .ZN(n8580) );
  NAND2_X1 U8517 ( .A1(n7955), .A2(n8581), .ZN(n8579) );
  NOR2_X1 U8518 ( .A1(n8582), .A2(n8013), .ZN(n8577) );
  INV_X1 U8519 ( .A(n8567), .ZN(n8575) );
  NAND2_X1 U8520 ( .A1(n8583), .A2(n8584), .ZN(n8567) );
  NAND2_X1 U8521 ( .A1(n8585), .A2(n8586), .ZN(Result_41_) );
  NAND2_X1 U8522 ( .A1(n7959), .A2(n8587), .ZN(n8586) );
  XOR2_X1 U8523 ( .A(n8588), .B(n8589), .Z(n8587) );
  XOR2_X1 U8524 ( .A(n8590), .B(n8591), .Z(n8589) );
  NOR2_X1 U8525 ( .A1(n8592), .A2(n8593), .ZN(n8585) );
  NOR2_X1 U8526 ( .A1(n8594), .A2(n8595), .ZN(n8593) );
  NOR2_X1 U8527 ( .A1(n8596), .A2(n8597), .ZN(n8594) );
  NAND2_X1 U8528 ( .A1(n8598), .A2(n8599), .ZN(n8597) );
  NAND2_X1 U8529 ( .A1(n7954), .A2(n8600), .ZN(n8599) );
  NAND2_X1 U8530 ( .A1(n7955), .A2(n8601), .ZN(n8598) );
  NOR2_X1 U8531 ( .A1(n8602), .A2(n8013), .ZN(n8596) );
  NOR2_X1 U8532 ( .A1(n8603), .A2(n8604), .ZN(n8592) );
  INV_X1 U8533 ( .A(n8595), .ZN(n8604) );
  XNOR2_X1 U8534 ( .A(n8605), .B(b_9_), .ZN(n8595) );
  NOR2_X1 U8535 ( .A1(n8606), .A2(n8607), .ZN(n8603) );
  NAND2_X1 U8536 ( .A1(n8608), .A2(n8609), .ZN(n8607) );
  OR2_X1 U8537 ( .A1(n8600), .A2(n7951), .ZN(n8609) );
  NAND2_X1 U8538 ( .A1(n7955), .A2(n8610), .ZN(n8608) );
  NOR2_X1 U8539 ( .A1(n8611), .A2(n8013), .ZN(n8606) );
  NAND2_X1 U8540 ( .A1(n8612), .A2(n8613), .ZN(Result_40_) );
  NAND2_X1 U8541 ( .A1(n7959), .A2(n8614), .ZN(n8613) );
  XOR2_X1 U8542 ( .A(n8615), .B(n8616), .Z(n8614) );
  XOR2_X1 U8543 ( .A(n8617), .B(n8618), .Z(n8616) );
  NOR2_X1 U8544 ( .A1(n7999), .A2(n8619), .ZN(n8618) );
  NOR2_X1 U8545 ( .A1(n8620), .A2(n8621), .ZN(n8612) );
  NOR2_X1 U8546 ( .A1(n8622), .A2(n8623), .ZN(n8621) );
  NOR2_X1 U8547 ( .A1(n8624), .A2(n8625), .ZN(n8622) );
  NAND2_X1 U8548 ( .A1(n8626), .A2(n8627), .ZN(n8625) );
  OR2_X1 U8549 ( .A1(n8628), .A2(n7951), .ZN(n8627) );
  NAND2_X1 U8550 ( .A1(n7955), .A2(n8629), .ZN(n8626) );
  NOR2_X1 U8551 ( .A1(n8630), .A2(n8013), .ZN(n8624) );
  NOR2_X1 U8552 ( .A1(n8631), .A2(n8632), .ZN(n8620) );
  NOR2_X1 U8553 ( .A1(n8633), .A2(n8634), .ZN(n8632) );
  NAND2_X1 U8554 ( .A1(n8635), .A2(n8636), .ZN(n8634) );
  NAND2_X1 U8555 ( .A1(n7954), .A2(n8628), .ZN(n8636) );
  NAND2_X1 U8556 ( .A1(n7955), .A2(n8637), .ZN(n8635) );
  NOR2_X1 U8557 ( .A1(n8638), .A2(n8013), .ZN(n8633) );
  INV_X1 U8558 ( .A(n8623), .ZN(n8631) );
  NAND2_X1 U8559 ( .A1(n8639), .A2(n8640), .ZN(n8623) );
  NAND2_X1 U8560 ( .A1(n7956), .A2(n8641), .ZN(Result_3_) );
  NAND2_X1 U8561 ( .A1(n8642), .A2(n7959), .ZN(n8641) );
  XOR2_X1 U8562 ( .A(n8643), .B(n8644), .Z(n8642) );
  AND2_X1 U8563 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  NAND2_X1 U8564 ( .A1(n8647), .A2(n8648), .ZN(Result_39_) );
  NAND2_X1 U8565 ( .A1(n8649), .A2(n7959), .ZN(n8648) );
  XOR2_X1 U8566 ( .A(n8650), .B(n8651), .Z(n8649) );
  XOR2_X1 U8567 ( .A(n8652), .B(n8653), .Z(n8650) );
  NOR2_X1 U8568 ( .A1(n8654), .A2(n8655), .ZN(n8647) );
  NOR2_X1 U8569 ( .A1(n8656), .A2(n8657), .ZN(n8655) );
  NOR2_X1 U8570 ( .A1(n8658), .A2(n8659), .ZN(n8656) );
  NAND2_X1 U8571 ( .A1(n8660), .A2(n8661), .ZN(n8659) );
  NAND2_X1 U8572 ( .A1(n7954), .A2(n8662), .ZN(n8661) );
  NAND2_X1 U8573 ( .A1(n7955), .A2(n8663), .ZN(n8660) );
  NOR2_X1 U8574 ( .A1(n8664), .A2(n8013), .ZN(n8658) );
  NOR2_X1 U8575 ( .A1(n8665), .A2(n8666), .ZN(n8654) );
  INV_X1 U8576 ( .A(n8657), .ZN(n8666) );
  XNOR2_X1 U8577 ( .A(n8667), .B(a_7_), .ZN(n8657) );
  NOR2_X1 U8578 ( .A1(n8668), .A2(n8669), .ZN(n8665) );
  NAND2_X1 U8579 ( .A1(n8670), .A2(n8671), .ZN(n8669) );
  OR2_X1 U8580 ( .A1(n8662), .A2(n7951), .ZN(n8671) );
  NAND2_X1 U8581 ( .A1(n7955), .A2(n8672), .ZN(n8670) );
  NOR2_X1 U8582 ( .A1(n8673), .A2(n8013), .ZN(n8668) );
  NAND2_X1 U8583 ( .A1(n8674), .A2(n8675), .ZN(Result_38_) );
  NAND2_X1 U8584 ( .A1(n8676), .A2(n7959), .ZN(n8675) );
  XOR2_X1 U8585 ( .A(n8677), .B(n8678), .Z(n8676) );
  XOR2_X1 U8586 ( .A(n8679), .B(n8680), .Z(n8677) );
  NOR2_X1 U8587 ( .A1(n7999), .A2(n8681), .ZN(n8680) );
  NOR2_X1 U8588 ( .A1(n8682), .A2(n8683), .ZN(n8674) );
  NOR2_X1 U8589 ( .A1(n8684), .A2(n8685), .ZN(n8683) );
  NOR2_X1 U8590 ( .A1(n8686), .A2(n8687), .ZN(n8684) );
  NAND2_X1 U8591 ( .A1(n8688), .A2(n8689), .ZN(n8687) );
  OR2_X1 U8592 ( .A1(n8690), .A2(n7951), .ZN(n8689) );
  NAND2_X1 U8593 ( .A1(n7955), .A2(n8691), .ZN(n8688) );
  NOR2_X1 U8594 ( .A1(n8692), .A2(n8013), .ZN(n8686) );
  NOR2_X1 U8595 ( .A1(n8693), .A2(n8694), .ZN(n8682) );
  NOR2_X1 U8596 ( .A1(n8695), .A2(n8696), .ZN(n8694) );
  NAND2_X1 U8597 ( .A1(n8697), .A2(n8698), .ZN(n8696) );
  NAND2_X1 U8598 ( .A1(n7954), .A2(n8690), .ZN(n8698) );
  NAND2_X1 U8599 ( .A1(n7955), .A2(n8699), .ZN(n8697) );
  NOR2_X1 U8600 ( .A1(n8700), .A2(n8013), .ZN(n8695) );
  INV_X1 U8601 ( .A(n8685), .ZN(n8693) );
  NAND2_X1 U8602 ( .A1(n8701), .A2(n8702), .ZN(n8685) );
  NAND2_X1 U8603 ( .A1(n8703), .A2(n8704), .ZN(Result_37_) );
  NAND2_X1 U8604 ( .A1(n8705), .A2(n7959), .ZN(n8704) );
  XOR2_X1 U8605 ( .A(n8706), .B(n8707), .Z(n8705) );
  XOR2_X1 U8606 ( .A(n8708), .B(n8709), .Z(n8706) );
  NOR2_X1 U8607 ( .A1(n8710), .A2(n8711), .ZN(n8703) );
  NOR2_X1 U8608 ( .A1(n8712), .A2(n8713), .ZN(n8711) );
  NOR2_X1 U8609 ( .A1(n8714), .A2(n8715), .ZN(n8712) );
  NAND2_X1 U8610 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
  NAND2_X1 U8611 ( .A1(n7954), .A2(n8718), .ZN(n8717) );
  NAND2_X1 U8612 ( .A1(n7955), .A2(n8719), .ZN(n8716) );
  NOR2_X1 U8613 ( .A1(n8720), .A2(n8013), .ZN(n8714) );
  NOR2_X1 U8614 ( .A1(n8721), .A2(n8722), .ZN(n8710) );
  INV_X1 U8615 ( .A(n8713), .ZN(n8722) );
  XNOR2_X1 U8616 ( .A(n8723), .B(b_5_), .ZN(n8713) );
  NOR2_X1 U8617 ( .A1(n8724), .A2(n8725), .ZN(n8721) );
  NAND2_X1 U8618 ( .A1(n8726), .A2(n8727), .ZN(n8725) );
  OR2_X1 U8619 ( .A1(n8718), .A2(n7951), .ZN(n8727) );
  NAND2_X1 U8620 ( .A1(n7955), .A2(n8728), .ZN(n8726) );
  NOR2_X1 U8621 ( .A1(n8729), .A2(n8013), .ZN(n8724) );
  NAND2_X1 U8622 ( .A1(n8730), .A2(n8731), .ZN(Result_36_) );
  NAND2_X1 U8623 ( .A1(n7959), .A2(n8732), .ZN(n8731) );
  XNOR2_X1 U8624 ( .A(n8733), .B(n8734), .ZN(n8732) );
  XOR2_X1 U8625 ( .A(n8735), .B(n8736), .Z(n8734) );
  NAND2_X1 U8626 ( .A1(a_4_), .A2(b_31_), .ZN(n8736) );
  NOR2_X1 U8627 ( .A1(n8737), .A2(n8738), .ZN(n8730) );
  NOR2_X1 U8628 ( .A1(n8739), .A2(n8740), .ZN(n8738) );
  NOR2_X1 U8629 ( .A1(n8741), .A2(n8742), .ZN(n8739) );
  NAND2_X1 U8630 ( .A1(n8743), .A2(n8744), .ZN(n8742) );
  OR2_X1 U8631 ( .A1(n8745), .A2(n7951), .ZN(n8744) );
  NAND2_X1 U8632 ( .A1(n7955), .A2(n8746), .ZN(n8743) );
  NOR2_X1 U8633 ( .A1(n8747), .A2(n8013), .ZN(n8741) );
  NOR2_X1 U8634 ( .A1(n8748), .A2(n8749), .ZN(n8737) );
  NOR2_X1 U8635 ( .A1(n8750), .A2(n8751), .ZN(n8749) );
  NAND2_X1 U8636 ( .A1(n8752), .A2(n8753), .ZN(n8751) );
  NAND2_X1 U8637 ( .A1(n7954), .A2(n8745), .ZN(n8753) );
  NAND2_X1 U8638 ( .A1(n7955), .A2(n8754), .ZN(n8752) );
  NOR2_X1 U8639 ( .A1(n8755), .A2(n8013), .ZN(n8750) );
  INV_X1 U8640 ( .A(n8740), .ZN(n8748) );
  NAND2_X1 U8641 ( .A1(n8756), .A2(n8757), .ZN(n8740) );
  NAND2_X1 U8642 ( .A1(n8758), .A2(n8759), .ZN(Result_35_) );
  NAND2_X1 U8643 ( .A1(n8760), .A2(n7959), .ZN(n8759) );
  XOR2_X1 U8644 ( .A(n8761), .B(n8762), .Z(n8760) );
  XOR2_X1 U8645 ( .A(n8763), .B(n8764), .Z(n8761) );
  NOR2_X1 U8646 ( .A1(n8765), .A2(n8766), .ZN(n8758) );
  NOR2_X1 U8647 ( .A1(n8767), .A2(n8768), .ZN(n8766) );
  NOR2_X1 U8648 ( .A1(n8769), .A2(n8770), .ZN(n8767) );
  NAND2_X1 U8649 ( .A1(n8771), .A2(n8772), .ZN(n8770) );
  NAND2_X1 U8650 ( .A1(n7954), .A2(n8773), .ZN(n8772) );
  NAND2_X1 U8651 ( .A1(n7955), .A2(n8774), .ZN(n8771) );
  NOR2_X1 U8652 ( .A1(n8775), .A2(n8013), .ZN(n8769) );
  NOR2_X1 U8653 ( .A1(n8776), .A2(n8777), .ZN(n8765) );
  INV_X1 U8654 ( .A(n8768), .ZN(n8777) );
  XNOR2_X1 U8655 ( .A(n8778), .B(b_3_), .ZN(n8768) );
  NOR2_X1 U8656 ( .A1(n8779), .A2(n8780), .ZN(n8776) );
  NAND2_X1 U8657 ( .A1(n8781), .A2(n8782), .ZN(n8780) );
  OR2_X1 U8658 ( .A1(n8773), .A2(n7951), .ZN(n8782) );
  NAND2_X1 U8659 ( .A1(n7955), .A2(n8783), .ZN(n8781) );
  NOR2_X1 U8660 ( .A1(n8784), .A2(n8013), .ZN(n8779) );
  NAND2_X1 U8661 ( .A1(n8785), .A2(n8786), .ZN(Result_34_) );
  NAND2_X1 U8662 ( .A1(n7959), .A2(n8787), .ZN(n8786) );
  XOR2_X1 U8663 ( .A(n8788), .B(n8789), .Z(n8787) );
  XOR2_X1 U8664 ( .A(n8790), .B(n8791), .Z(n8789) );
  NOR2_X1 U8665 ( .A1(n7999), .A2(n8792), .ZN(n8791) );
  NOR2_X1 U8666 ( .A1(n8793), .A2(n8794), .ZN(n8785) );
  NOR2_X1 U8667 ( .A1(n8795), .A2(n8796), .ZN(n8794) );
  NOR2_X1 U8668 ( .A1(n8797), .A2(n8798), .ZN(n8795) );
  NAND2_X1 U8669 ( .A1(n8799), .A2(n8800), .ZN(n8798) );
  OR2_X1 U8670 ( .A1(n8801), .A2(n7951), .ZN(n8800) );
  NAND2_X1 U8671 ( .A1(n7955), .A2(n8802), .ZN(n8799) );
  NOR2_X1 U8672 ( .A1(n8803), .A2(n8013), .ZN(n8797) );
  NOR2_X1 U8673 ( .A1(n8804), .A2(n8805), .ZN(n8793) );
  NOR2_X1 U8674 ( .A1(n8806), .A2(n8807), .ZN(n8805) );
  NAND2_X1 U8675 ( .A1(n8808), .A2(n8809), .ZN(n8807) );
  NAND2_X1 U8676 ( .A1(n7954), .A2(n8801), .ZN(n8809) );
  NAND2_X1 U8677 ( .A1(n7955), .A2(n8810), .ZN(n8808) );
  NOR2_X1 U8678 ( .A1(n8811), .A2(n8013), .ZN(n8806) );
  INV_X1 U8679 ( .A(n8796), .ZN(n8804) );
  NAND2_X1 U8680 ( .A1(n8812), .A2(n8813), .ZN(n8796) );
  NAND2_X1 U8681 ( .A1(n8814), .A2(n8815), .ZN(Result_33_) );
  NAND2_X1 U8682 ( .A1(n7959), .A2(n8816), .ZN(n8815) );
  XOR2_X1 U8683 ( .A(n8817), .B(n8818), .Z(n8816) );
  XOR2_X1 U8684 ( .A(n8819), .B(n8820), .Z(n8818) );
  NOR2_X1 U8685 ( .A1(n8821), .A2(n8822), .ZN(n8814) );
  NOR2_X1 U8686 ( .A1(n8823), .A2(n8824), .ZN(n8822) );
  NOR2_X1 U8687 ( .A1(n8825), .A2(n8826), .ZN(n8823) );
  NAND2_X1 U8688 ( .A1(n8827), .A2(n8828), .ZN(n8826) );
  NAND2_X1 U8689 ( .A1(n7954), .A2(n8829), .ZN(n8828) );
  NAND2_X1 U8690 ( .A1(n7955), .A2(n8830), .ZN(n8827) );
  NOR2_X1 U8691 ( .A1(n8831), .A2(n8013), .ZN(n8825) );
  NOR2_X1 U8692 ( .A1(n8832), .A2(n8833), .ZN(n8821) );
  INV_X1 U8693 ( .A(n8824), .ZN(n8833) );
  XNOR2_X1 U8694 ( .A(n8834), .B(a_1_), .ZN(n8824) );
  NOR2_X1 U8695 ( .A1(n8835), .A2(n8836), .ZN(n8832) );
  NAND2_X1 U8696 ( .A1(n8837), .A2(n8838), .ZN(n8836) );
  OR2_X1 U8697 ( .A1(n8829), .A2(n7951), .ZN(n8838) );
  NAND2_X1 U8698 ( .A1(n7955), .A2(n8839), .ZN(n8837) );
  NOR2_X1 U8699 ( .A1(n8840), .A2(n8013), .ZN(n8835) );
  NAND2_X1 U8700 ( .A1(n8841), .A2(n8842), .ZN(Result_32_) );
  NAND2_X1 U8701 ( .A1(n7959), .A2(n8843), .ZN(n8842) );
  XNOR2_X1 U8702 ( .A(n8844), .B(n8845), .ZN(n8843) );
  XOR2_X1 U8703 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND2_X1 U8704 ( .A1(a_0_), .A2(b_31_), .ZN(n8847) );
  NOR2_X1 U8705 ( .A1(n8848), .A2(n8849), .ZN(n8841) );
  NOR2_X1 U8706 ( .A1(n8850), .A2(n8851), .ZN(n8849) );
  NOR2_X1 U8707 ( .A1(n8852), .A2(n8853), .ZN(n8850) );
  NAND2_X1 U8708 ( .A1(n8854), .A2(n8855), .ZN(n8853) );
  NAND2_X1 U8709 ( .A1(n7954), .A2(n8856), .ZN(n8855) );
  NAND2_X1 U8710 ( .A1(n7955), .A2(n8857), .ZN(n8854) );
  NOR2_X1 U8711 ( .A1(n8858), .A2(n8013), .ZN(n8852) );
  NOR2_X1 U8712 ( .A1(n8859), .A2(n8860), .ZN(n8848) );
  NOR2_X1 U8713 ( .A1(n8861), .A2(n8862), .ZN(n8860) );
  NAND2_X1 U8714 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  OR2_X1 U8715 ( .A1(n8856), .A2(n7951), .ZN(n8864) );
  NAND2_X1 U8716 ( .A1(n8865), .A2(n8866), .ZN(n8856) );
  OR2_X1 U8717 ( .A1(n8829), .A2(n8867), .ZN(n8866) );
  NAND2_X1 U8718 ( .A1(n8812), .A2(n8868), .ZN(n8829) );
  NAND2_X1 U8719 ( .A1(n8813), .A2(n8801), .ZN(n8868) );
  NAND2_X1 U8720 ( .A1(n8869), .A2(n8870), .ZN(n8801) );
  NAND2_X1 U8721 ( .A1(n8871), .A2(n8773), .ZN(n8870) );
  NAND2_X1 U8722 ( .A1(n8756), .A2(n8872), .ZN(n8773) );
  NAND2_X1 U8723 ( .A1(n8757), .A2(n8745), .ZN(n8872) );
  NAND2_X1 U8724 ( .A1(n8873), .A2(n8874), .ZN(n8745) );
  NAND2_X1 U8725 ( .A1(n8875), .A2(n8718), .ZN(n8874) );
  NAND2_X1 U8726 ( .A1(n8701), .A2(n8876), .ZN(n8718) );
  NAND2_X1 U8727 ( .A1(n8702), .A2(n8690), .ZN(n8876) );
  NAND2_X1 U8728 ( .A1(n8877), .A2(n8878), .ZN(n8690) );
  NAND2_X1 U8729 ( .A1(n8879), .A2(n8662), .ZN(n8878) );
  NAND2_X1 U8730 ( .A1(n8639), .A2(n8880), .ZN(n8662) );
  NAND2_X1 U8731 ( .A1(n8640), .A2(n8628), .ZN(n8880) );
  NAND2_X1 U8732 ( .A1(n8881), .A2(n8882), .ZN(n8628) );
  NAND2_X1 U8733 ( .A1(n8883), .A2(n8600), .ZN(n8882) );
  NAND2_X1 U8734 ( .A1(n8583), .A2(n8884), .ZN(n8600) );
  NAND2_X1 U8735 ( .A1(n8584), .A2(n8572), .ZN(n8884) );
  NAND2_X1 U8736 ( .A1(n8885), .A2(n8886), .ZN(n8572) );
  NAND2_X1 U8737 ( .A1(n8887), .A2(n8545), .ZN(n8886) );
  NAND2_X1 U8738 ( .A1(n8528), .A2(n8888), .ZN(n8545) );
  NAND2_X1 U8739 ( .A1(n8529), .A2(n8517), .ZN(n8888) );
  NAND2_X1 U8740 ( .A1(n8889), .A2(n8890), .ZN(n8517) );
  NAND2_X1 U8741 ( .A1(n8891), .A2(n8490), .ZN(n8890) );
  NAND2_X1 U8742 ( .A1(n8473), .A2(n8892), .ZN(n8490) );
  NAND2_X1 U8743 ( .A1(n8474), .A2(n8462), .ZN(n8892) );
  NAND2_X1 U8744 ( .A1(n8893), .A2(n8894), .ZN(n8462) );
  NAND2_X1 U8745 ( .A1(n8895), .A2(n8435), .ZN(n8894) );
  NAND2_X1 U8746 ( .A1(n8418), .A2(n8896), .ZN(n8435) );
  NAND2_X1 U8747 ( .A1(n8419), .A2(n8407), .ZN(n8896) );
  NAND2_X1 U8748 ( .A1(n8897), .A2(n8898), .ZN(n8407) );
  NAND2_X1 U8749 ( .A1(n8899), .A2(n8380), .ZN(n8898) );
  NAND2_X1 U8750 ( .A1(n8357), .A2(n8900), .ZN(n8380) );
  NAND2_X1 U8751 ( .A1(n8358), .A2(n8346), .ZN(n8900) );
  NAND2_X1 U8752 ( .A1(n8901), .A2(n8902), .ZN(n8346) );
  NAND2_X1 U8753 ( .A1(n8903), .A2(n8319), .ZN(n8902) );
  NAND2_X1 U8754 ( .A1(n8302), .A2(n8904), .ZN(n8319) );
  NAND2_X1 U8755 ( .A1(n8303), .A2(n8299), .ZN(n8904) );
  INV_X1 U8756 ( .A(n8290), .ZN(n8299) );
  NOR2_X1 U8757 ( .A1(n8905), .A2(n8906), .ZN(n8290) );
  AND2_X1 U8758 ( .A1(n8907), .A2(n8263), .ZN(n8906) );
  NAND2_X1 U8759 ( .A1(n8908), .A2(n8909), .ZN(n8263) );
  NAND2_X1 U8760 ( .A1(n8910), .A2(n8235), .ZN(n8909) );
  INV_X1 U8761 ( .A(n8245), .ZN(n8235) );
  NOR2_X1 U8762 ( .A1(n8911), .A2(n8912), .ZN(n8245) );
  AND2_X1 U8763 ( .A1(n8913), .A2(n8208), .ZN(n8912) );
  NAND2_X1 U8764 ( .A1(n8914), .A2(n8915), .ZN(n8208) );
  NAND2_X1 U8765 ( .A1(n8916), .A2(n8180), .ZN(n8915) );
  INV_X1 U8766 ( .A(n8190), .ZN(n8180) );
  NOR2_X1 U8767 ( .A1(n8917), .A2(n8918), .ZN(n8190) );
  AND2_X1 U8768 ( .A1(n8919), .A2(n8153), .ZN(n8918) );
  NAND2_X1 U8769 ( .A1(n8920), .A2(n8921), .ZN(n8153) );
  NAND2_X1 U8770 ( .A1(n8922), .A2(n8125), .ZN(n8921) );
  INV_X1 U8771 ( .A(n8135), .ZN(n8125) );
  NOR2_X1 U8772 ( .A1(n8923), .A2(n8924), .ZN(n8135) );
  AND2_X1 U8773 ( .A1(n8925), .A2(n8097), .ZN(n8924) );
  NAND2_X1 U8774 ( .A1(n8926), .A2(n8927), .ZN(n8097) );
  NAND2_X1 U8775 ( .A1(n8928), .A2(n8064), .ZN(n8927) );
  NAND2_X1 U8776 ( .A1(n8929), .A2(n8930), .ZN(n8064) );
  NAND2_X1 U8777 ( .A1(n8931), .A2(n8036), .ZN(n8930) );
  NAND2_X1 U8778 ( .A1(n8932), .A2(n8933), .ZN(n8036) );
  NAND2_X1 U8779 ( .A1(b_30_), .A2(n8934), .ZN(n8933) );
  NAND2_X1 U8780 ( .A1(n8935), .A2(n8012), .ZN(n8934) );
  NAND2_X1 U8781 ( .A1(a_31_), .A2(b_31_), .ZN(n8012) );
  NAND2_X1 U8782 ( .A1(n7953), .A2(b_31_), .ZN(n8932) );
  NAND2_X1 U8783 ( .A1(n8936), .A2(n8041), .ZN(n8931) );
  NAND2_X1 U8784 ( .A1(n8069), .A2(n8055), .ZN(n8928) );
  NAND2_X1 U8785 ( .A1(n8102), .A2(n8937), .ZN(n8925) );
  NAND2_X1 U8786 ( .A1(n8130), .A2(n8116), .ZN(n8922) );
  NAND2_X1 U8787 ( .A1(n8938), .A2(n8158), .ZN(n8919) );
  NAND2_X1 U8788 ( .A1(n8185), .A2(n8939), .ZN(n8916) );
  NAND2_X1 U8789 ( .A1(n8940), .A2(n8213), .ZN(n8913) );
  NAND2_X1 U8790 ( .A1(n8240), .A2(n8941), .ZN(n8910) );
  NAND2_X1 U8791 ( .A1(n8942), .A2(n8268), .ZN(n8907) );
  NAND2_X1 U8792 ( .A1(n8943), .A2(n8944), .ZN(n8303) );
  NAND2_X1 U8793 ( .A1(n8945), .A2(n8324), .ZN(n8903) );
  NAND2_X1 U8794 ( .A1(n8946), .A2(n8947), .ZN(n8358) );
  NAND2_X1 U8795 ( .A1(n8948), .A2(n8385), .ZN(n8899) );
  NAND2_X1 U8796 ( .A1(n8949), .A2(n8950), .ZN(n8419) );
  NAND2_X1 U8797 ( .A1(n8951), .A2(n8440), .ZN(n8895) );
  NAND2_X1 U8798 ( .A1(n8952), .A2(n8953), .ZN(n8474) );
  NAND2_X1 U8799 ( .A1(n8954), .A2(n8495), .ZN(n8891) );
  NAND2_X1 U8800 ( .A1(n8955), .A2(n8956), .ZN(n8529) );
  NAND2_X1 U8801 ( .A1(n8957), .A2(n8550), .ZN(n8887) );
  NAND2_X1 U8802 ( .A1(n8958), .A2(n8959), .ZN(n8584) );
  NAND2_X1 U8803 ( .A1(n8960), .A2(n8605), .ZN(n8883) );
  NAND2_X1 U8804 ( .A1(n8961), .A2(n8619), .ZN(n8640) );
  NAND2_X1 U8805 ( .A1(n8667), .A2(n8962), .ZN(n8879) );
  NAND2_X1 U8806 ( .A1(n8963), .A2(n8681), .ZN(n8702) );
  NAND2_X1 U8807 ( .A1(n8964), .A2(n8723), .ZN(n8875) );
  NAND2_X1 U8808 ( .A1(n8965), .A2(n8966), .ZN(n8757) );
  NAND2_X1 U8809 ( .A1(n8967), .A2(n8778), .ZN(n8871) );
  NAND2_X1 U8810 ( .A1(n8968), .A2(n8792), .ZN(n8813) );
  NAND2_X1 U8811 ( .A1(n8834), .A2(n8969), .ZN(n8865) );
  NAND2_X1 U8812 ( .A1(n7955), .A2(n8970), .ZN(n8863) );
  NOR2_X1 U8813 ( .A1(n8971), .A2(n8013), .ZN(n8861) );
  INV_X1 U8814 ( .A(n8851), .ZN(n8859) );
  NAND2_X1 U8815 ( .A1(n8972), .A2(n8973), .ZN(n8851) );
  NAND2_X1 U8816 ( .A1(n8974), .A2(n8975), .ZN(n8973) );
  NAND2_X1 U8817 ( .A1(n7956), .A2(n8976), .ZN(Result_31_) );
  NAND2_X1 U8818 ( .A1(n7959), .A2(n8977), .ZN(n8976) );
  XOR2_X1 U8819 ( .A(n8978), .B(n8979), .Z(n8977) );
  NAND2_X1 U8820 ( .A1(n7956), .A2(n8980), .ZN(Result_30_) );
  NAND2_X1 U8821 ( .A1(n8981), .A2(n7959), .ZN(n8980) );
  NOR2_X1 U8822 ( .A1(n8982), .A2(n8983), .ZN(n8981) );
  NOR2_X1 U8823 ( .A1(n8984), .A2(n8985), .ZN(n8983) );
  NAND2_X1 U8824 ( .A1(n7956), .A2(n8986), .ZN(Result_2_) );
  NAND2_X1 U8825 ( .A1(n8987), .A2(n7959), .ZN(n8986) );
  XOR2_X1 U8826 ( .A(n8988), .B(n8989), .Z(n8987) );
  AND2_X1 U8827 ( .A1(n8990), .A2(n8991), .ZN(n8989) );
  NAND2_X1 U8828 ( .A1(n7956), .A2(n8992), .ZN(Result_29_) );
  NAND2_X1 U8829 ( .A1(n7959), .A2(n8993), .ZN(n8992) );
  XNOR2_X1 U8830 ( .A(n8982), .B(n8994), .ZN(n8993) );
  NAND2_X1 U8831 ( .A1(n8995), .A2(n8996), .ZN(n8994) );
  NAND2_X1 U8832 ( .A1(n7956), .A2(n8997), .ZN(Result_28_) );
  NAND2_X1 U8833 ( .A1(n8998), .A2(n7959), .ZN(n8997) );
  XNOR2_X1 U8834 ( .A(n8999), .B(n9000), .ZN(n8998) );
  NAND2_X1 U8835 ( .A1(n9001), .A2(n9002), .ZN(n8999) );
  NAND2_X1 U8836 ( .A1(n7956), .A2(n9003), .ZN(Result_27_) );
  NAND2_X1 U8837 ( .A1(n9004), .A2(n7959), .ZN(n9003) );
  XOR2_X1 U8838 ( .A(n9005), .B(n9006), .Z(n9004) );
  AND2_X1 U8839 ( .A1(n9007), .A2(n9008), .ZN(n9006) );
  NAND2_X1 U8840 ( .A1(n7956), .A2(n9009), .ZN(Result_26_) );
  NAND2_X1 U8841 ( .A1(n9010), .A2(n7959), .ZN(n9009) );
  XOR2_X1 U8842 ( .A(n9011), .B(n9012), .Z(n9010) );
  AND2_X1 U8843 ( .A1(n9013), .A2(n9014), .ZN(n9012) );
  NAND2_X1 U8844 ( .A1(n7956), .A2(n9015), .ZN(Result_25_) );
  NAND2_X1 U8845 ( .A1(n9016), .A2(n7959), .ZN(n9015) );
  XOR2_X1 U8846 ( .A(n9017), .B(n9018), .Z(n9016) );
  AND2_X1 U8847 ( .A1(n9019), .A2(n9020), .ZN(n9018) );
  NAND2_X1 U8848 ( .A1(n7956), .A2(n9021), .ZN(Result_24_) );
  NAND2_X1 U8849 ( .A1(n9022), .A2(n7959), .ZN(n9021) );
  XOR2_X1 U8850 ( .A(n9023), .B(n9024), .Z(n9022) );
  AND2_X1 U8851 ( .A1(n9025), .A2(n9026), .ZN(n9024) );
  NAND2_X1 U8852 ( .A1(n7956), .A2(n9027), .ZN(Result_23_) );
  NAND2_X1 U8853 ( .A1(n9028), .A2(n7959), .ZN(n9027) );
  XOR2_X1 U8854 ( .A(n9029), .B(n9030), .Z(n9028) );
  AND2_X1 U8855 ( .A1(n9031), .A2(n9032), .ZN(n9030) );
  NAND2_X1 U8856 ( .A1(n7956), .A2(n9033), .ZN(Result_22_) );
  NAND2_X1 U8857 ( .A1(n9034), .A2(n7959), .ZN(n9033) );
  XOR2_X1 U8858 ( .A(n9035), .B(n9036), .Z(n9034) );
  AND2_X1 U8859 ( .A1(n9037), .A2(n9038), .ZN(n9036) );
  NAND2_X1 U8860 ( .A1(n7956), .A2(n9039), .ZN(Result_21_) );
  NAND2_X1 U8861 ( .A1(n9040), .A2(n7959), .ZN(n9039) );
  XOR2_X1 U8862 ( .A(n9041), .B(n9042), .Z(n9040) );
  AND2_X1 U8863 ( .A1(n9043), .A2(n9044), .ZN(n9042) );
  NAND2_X1 U8864 ( .A1(n7956), .A2(n9045), .ZN(Result_20_) );
  NAND2_X1 U8865 ( .A1(n9046), .A2(n7959), .ZN(n9045) );
  XOR2_X1 U8866 ( .A(n9047), .B(n9048), .Z(n9046) );
  AND2_X1 U8867 ( .A1(n9049), .A2(n9050), .ZN(n9048) );
  NAND2_X1 U8868 ( .A1(n7956), .A2(n9051), .ZN(Result_1_) );
  NAND2_X1 U8869 ( .A1(n9052), .A2(n7959), .ZN(n9051) );
  XNOR2_X1 U8870 ( .A(n9053), .B(n9054), .ZN(n9052) );
  NOR2_X1 U8871 ( .A1(n9055), .A2(n9056), .ZN(n9054) );
  NAND2_X1 U8872 ( .A1(n7956), .A2(n9057), .ZN(Result_19_) );
  NAND2_X1 U8873 ( .A1(n9058), .A2(n7959), .ZN(n9057) );
  XOR2_X1 U8874 ( .A(n9059), .B(n9060), .Z(n9058) );
  AND2_X1 U8875 ( .A1(n9061), .A2(n9062), .ZN(n9060) );
  NAND2_X1 U8876 ( .A1(n7956), .A2(n9063), .ZN(Result_18_) );
  NAND2_X1 U8877 ( .A1(n9064), .A2(n7959), .ZN(n9063) );
  XOR2_X1 U8878 ( .A(n9065), .B(n9066), .Z(n9064) );
  AND2_X1 U8879 ( .A1(n9067), .A2(n9068), .ZN(n9066) );
  NAND2_X1 U8880 ( .A1(n7956), .A2(n9069), .ZN(Result_17_) );
  NAND2_X1 U8881 ( .A1(n9070), .A2(n7959), .ZN(n9069) );
  XOR2_X1 U8882 ( .A(n9071), .B(n9072), .Z(n9070) );
  AND2_X1 U8883 ( .A1(n9073), .A2(n9074), .ZN(n9072) );
  NAND2_X1 U8884 ( .A1(n7956), .A2(n9075), .ZN(Result_16_) );
  NAND2_X1 U8885 ( .A1(n9076), .A2(n7959), .ZN(n9075) );
  XOR2_X1 U8886 ( .A(n9077), .B(n9078), .Z(n9076) );
  AND2_X1 U8887 ( .A1(n9079), .A2(n9080), .ZN(n9078) );
  NAND2_X1 U8888 ( .A1(n7956), .A2(n9081), .ZN(Result_15_) );
  NAND2_X1 U8889 ( .A1(n9082), .A2(n7959), .ZN(n9081) );
  XOR2_X1 U8890 ( .A(n9083), .B(n9084), .Z(n9082) );
  AND2_X1 U8891 ( .A1(n9085), .A2(n9086), .ZN(n9084) );
  NAND2_X1 U8892 ( .A1(n7956), .A2(n9087), .ZN(Result_14_) );
  NAND2_X1 U8893 ( .A1(n9088), .A2(n7959), .ZN(n9087) );
  XOR2_X1 U8894 ( .A(n9089), .B(n9090), .Z(n9088) );
  AND2_X1 U8895 ( .A1(n9091), .A2(n9092), .ZN(n9090) );
  NAND2_X1 U8896 ( .A1(n7956), .A2(n9093), .ZN(Result_13_) );
  NAND2_X1 U8897 ( .A1(n9094), .A2(n7959), .ZN(n9093) );
  XOR2_X1 U8898 ( .A(n9095), .B(n9096), .Z(n9094) );
  AND2_X1 U8899 ( .A1(n9097), .A2(n9098), .ZN(n9096) );
  NAND2_X1 U8900 ( .A1(n7956), .A2(n9099), .ZN(Result_12_) );
  NAND2_X1 U8901 ( .A1(n9100), .A2(n7959), .ZN(n9099) );
  XOR2_X1 U8902 ( .A(n9101), .B(n9102), .Z(n9100) );
  AND2_X1 U8903 ( .A1(n9103), .A2(n9104), .ZN(n9102) );
  NAND2_X1 U8904 ( .A1(n7956), .A2(n9105), .ZN(Result_11_) );
  NAND2_X1 U8905 ( .A1(n9106), .A2(n7959), .ZN(n9105) );
  XOR2_X1 U8906 ( .A(n9107), .B(n9108), .Z(n9106) );
  AND2_X1 U8907 ( .A1(n9109), .A2(n9110), .ZN(n9108) );
  NAND2_X1 U8908 ( .A1(n7956), .A2(n9111), .ZN(Result_10_) );
  NAND2_X1 U8909 ( .A1(n9112), .A2(n7959), .ZN(n9111) );
  XOR2_X1 U8910 ( .A(n9113), .B(n9114), .Z(n9112) );
  AND2_X1 U8911 ( .A1(n9115), .A2(n9116), .ZN(n9114) );
  NAND2_X1 U8912 ( .A1(n7956), .A2(n9117), .ZN(Result_0_) );
  NAND2_X1 U8913 ( .A1(n7959), .A2(n9118), .ZN(n9117) );
  NAND2_X1 U8914 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  NAND2_X1 U8915 ( .A1(a_0_), .A2(n9121), .ZN(n9120) );
  NOR2_X1 U8916 ( .A1(n9056), .A2(n9122), .ZN(n9119) );
  NOR2_X1 U8917 ( .A1(n9053), .A2(n9055), .ZN(n9122) );
  AND2_X1 U8918 ( .A1(n9123), .A2(n9124), .ZN(n9055) );
  XOR2_X1 U8919 ( .A(n8972), .B(n9121), .Z(n9123) );
  AND2_X1 U8920 ( .A1(n8991), .A2(n9125), .ZN(n9053) );
  NAND2_X1 U8921 ( .A1(n8990), .A2(n8988), .ZN(n9125) );
  NAND2_X1 U8922 ( .A1(n8645), .A2(n9126), .ZN(n8988) );
  NAND2_X1 U8923 ( .A1(n8646), .A2(n8643), .ZN(n9126) );
  NAND2_X1 U8924 ( .A1(n8364), .A2(n9127), .ZN(n8643) );
  NAND2_X1 U8925 ( .A1(n8363), .A2(n8361), .ZN(n9127) );
  NAND2_X1 U8926 ( .A1(n8080), .A2(n9128), .ZN(n8361) );
  NAND2_X1 U8927 ( .A1(n8081), .A2(n8078), .ZN(n9128) );
  NAND2_X1 U8928 ( .A1(n7981), .A2(n9129), .ZN(n8078) );
  NAND2_X1 U8929 ( .A1(n7980), .A2(n7978), .ZN(n9129) );
  NAND2_X1 U8930 ( .A1(n7974), .A2(n9130), .ZN(n7978) );
  NAND2_X1 U8931 ( .A1(n7975), .A2(n7972), .ZN(n9130) );
  NAND2_X1 U8932 ( .A1(n7969), .A2(n9131), .ZN(n7972) );
  NAND2_X1 U8933 ( .A1(n7968), .A2(n7966), .ZN(n9131) );
  NAND2_X1 U8934 ( .A1(n7962), .A2(n9132), .ZN(n7966) );
  NAND2_X1 U8935 ( .A1(n7963), .A2(n7960), .ZN(n9132) );
  NAND2_X1 U8936 ( .A1(n9116), .A2(n9133), .ZN(n7960) );
  NAND2_X1 U8937 ( .A1(n9113), .A2(n9115), .ZN(n9133) );
  NAND2_X1 U8938 ( .A1(n9134), .A2(n9135), .ZN(n9115) );
  NAND2_X1 U8939 ( .A1(n9109), .A2(n9136), .ZN(n9113) );
  NAND2_X1 U8940 ( .A1(n9107), .A2(n9110), .ZN(n9136) );
  NAND2_X1 U8941 ( .A1(n9137), .A2(n9138), .ZN(n9110) );
  NAND2_X1 U8942 ( .A1(n9104), .A2(n9139), .ZN(n9107) );
  NAND2_X1 U8943 ( .A1(n9101), .A2(n9103), .ZN(n9139) );
  NAND2_X1 U8944 ( .A1(n9140), .A2(n9141), .ZN(n9103) );
  XNOR2_X1 U8945 ( .A(n9142), .B(n9143), .ZN(n9140) );
  NAND2_X1 U8946 ( .A1(n9097), .A2(n9144), .ZN(n9101) );
  NAND2_X1 U8947 ( .A1(n9095), .A2(n9098), .ZN(n9144) );
  NAND2_X1 U8948 ( .A1(n9145), .A2(n9146), .ZN(n9098) );
  NAND2_X1 U8949 ( .A1(n9092), .A2(n9147), .ZN(n9095) );
  NAND2_X1 U8950 ( .A1(n9091), .A2(n9089), .ZN(n9147) );
  NAND2_X1 U8951 ( .A1(n9086), .A2(n9148), .ZN(n9089) );
  NAND2_X1 U8952 ( .A1(n9085), .A2(n9083), .ZN(n9148) );
  NAND2_X1 U8953 ( .A1(n9080), .A2(n9149), .ZN(n9083) );
  NAND2_X1 U8954 ( .A1(n9077), .A2(n9079), .ZN(n9149) );
  NAND2_X1 U8955 ( .A1(n9150), .A2(n9151), .ZN(n9079) );
  NAND2_X1 U8956 ( .A1(n9152), .A2(n9153), .ZN(n9151) );
  XOR2_X1 U8957 ( .A(n9154), .B(n9155), .Z(n9150) );
  NAND2_X1 U8958 ( .A1(n9074), .A2(n9156), .ZN(n9077) );
  NAND2_X1 U8959 ( .A1(n9073), .A2(n9071), .ZN(n9156) );
  NAND2_X1 U8960 ( .A1(n9067), .A2(n9157), .ZN(n9071) );
  NAND2_X1 U8961 ( .A1(n9065), .A2(n9068), .ZN(n9157) );
  NAND2_X1 U8962 ( .A1(n9158), .A2(n9159), .ZN(n9068) );
  NAND2_X1 U8963 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  XOR2_X1 U8964 ( .A(n9162), .B(n9163), .Z(n9158) );
  NAND2_X1 U8965 ( .A1(n9062), .A2(n9164), .ZN(n9065) );
  NAND2_X1 U8966 ( .A1(n9059), .A2(n9061), .ZN(n9164) );
  NAND2_X1 U8967 ( .A1(n9165), .A2(n9166), .ZN(n9061) );
  NAND2_X1 U8968 ( .A1(n9167), .A2(n9168), .ZN(n9166) );
  XNOR2_X1 U8969 ( .A(n9161), .B(n9160), .ZN(n9165) );
  NAND2_X1 U8970 ( .A1(n9050), .A2(n9169), .ZN(n9059) );
  NAND2_X1 U8971 ( .A1(n9047), .A2(n9049), .ZN(n9169) );
  NAND2_X1 U8972 ( .A1(n9170), .A2(n9171), .ZN(n9049) );
  NAND2_X1 U8973 ( .A1(n9043), .A2(n9172), .ZN(n9047) );
  NAND2_X1 U8974 ( .A1(n9044), .A2(n9041), .ZN(n9172) );
  NAND2_X1 U8975 ( .A1(n9037), .A2(n9173), .ZN(n9041) );
  NAND2_X1 U8976 ( .A1(n9035), .A2(n9038), .ZN(n9173) );
  NAND2_X1 U8977 ( .A1(n9174), .A2(n9175), .ZN(n9038) );
  NAND2_X1 U8978 ( .A1(n9176), .A2(n9177), .ZN(n9175) );
  XNOR2_X1 U8979 ( .A(n9178), .B(n9179), .ZN(n9174) );
  NAND2_X1 U8980 ( .A1(n9032), .A2(n9180), .ZN(n9035) );
  NAND2_X1 U8981 ( .A1(n9029), .A2(n9031), .ZN(n9180) );
  NAND2_X1 U8982 ( .A1(n9181), .A2(n9182), .ZN(n9031) );
  NAND2_X1 U8983 ( .A1(n9183), .A2(n9184), .ZN(n9182) );
  XOR2_X1 U8984 ( .A(n9177), .B(n9185), .Z(n9181) );
  NAND2_X1 U8985 ( .A1(n9026), .A2(n9186), .ZN(n9029) );
  NAND2_X1 U8986 ( .A1(n9023), .A2(n9025), .ZN(n9186) );
  NAND2_X1 U8987 ( .A1(n9187), .A2(n9188), .ZN(n9025) );
  NAND2_X1 U8988 ( .A1(n9019), .A2(n9189), .ZN(n9023) );
  NAND2_X1 U8989 ( .A1(n9020), .A2(n9017), .ZN(n9189) );
  NAND2_X1 U8990 ( .A1(n9190), .A2(n9013), .ZN(n9017) );
  NAND2_X1 U8991 ( .A1(n9191), .A2(n9192), .ZN(n9013) );
  XOR2_X1 U8992 ( .A(n9193), .B(n9194), .Z(n9191) );
  NAND2_X1 U8993 ( .A1(n9014), .A2(n9011), .ZN(n9190) );
  NAND2_X1 U8994 ( .A1(n9008), .A2(n9195), .ZN(n9011) );
  NAND2_X1 U8995 ( .A1(n9005), .A2(n9007), .ZN(n9195) );
  NAND2_X1 U8996 ( .A1(n9196), .A2(n9197), .ZN(n9007) );
  NAND2_X1 U8997 ( .A1(n9001), .A2(n9198), .ZN(n9005) );
  NAND2_X1 U8998 ( .A1(n9000), .A2(n9002), .ZN(n9198) );
  NAND2_X1 U8999 ( .A1(n9199), .A2(n9200), .ZN(n9002) );
  NAND2_X1 U9000 ( .A1(n9201), .A2(n9202), .ZN(n9200) );
  XNOR2_X1 U9001 ( .A(n9203), .B(n9204), .ZN(n9199) );
  NAND2_X1 U9002 ( .A1(n8996), .A2(n9205), .ZN(n9000) );
  NAND2_X1 U9003 ( .A1(n8982), .A2(n8995), .ZN(n9205) );
  NAND2_X1 U9004 ( .A1(n9206), .A2(n9207), .ZN(n8995) );
  NAND2_X1 U9005 ( .A1(n9208), .A2(n9209), .ZN(n9207) );
  XNOR2_X1 U9006 ( .A(n9202), .B(n9201), .ZN(n9206) );
  AND2_X1 U9007 ( .A1(n8984), .A2(n8985), .ZN(n8982) );
  XOR2_X1 U9008 ( .A(n9209), .B(n9208), .Z(n8985) );
  NOR2_X1 U9009 ( .A1(n8978), .A2(n8979), .ZN(n8984) );
  XNOR2_X1 U9010 ( .A(n9210), .B(n9211), .ZN(n8979) );
  XOR2_X1 U9011 ( .A(n9212), .B(n9213), .Z(n9210) );
  NOR2_X1 U9012 ( .A1(n8002), .A2(n8974), .ZN(n9213) );
  AND2_X1 U9013 ( .A1(n9214), .A2(n9215), .ZN(n8978) );
  NAND2_X1 U9014 ( .A1(n9216), .A2(a_0_), .ZN(n9215) );
  NOR2_X1 U9015 ( .A1(n9217), .A2(n7999), .ZN(n9216) );
  NOR2_X1 U9016 ( .A1(n8844), .A2(n8846), .ZN(n9217) );
  NAND2_X1 U9017 ( .A1(n8844), .A2(n8846), .ZN(n9214) );
  NAND2_X1 U9018 ( .A1(n9218), .A2(n9219), .ZN(n8846) );
  NAND2_X1 U9019 ( .A1(n8820), .A2(n9220), .ZN(n9219) );
  NAND2_X1 U9020 ( .A1(n8819), .A2(n8817), .ZN(n9220) );
  NOR2_X1 U9021 ( .A1(n8969), .A2(n7999), .ZN(n8820) );
  OR2_X1 U9022 ( .A1(n8817), .A2(n8819), .ZN(n9218) );
  AND2_X1 U9023 ( .A1(n9221), .A2(n9222), .ZN(n8819) );
  NAND2_X1 U9024 ( .A1(n9223), .A2(a_2_), .ZN(n9222) );
  NOR2_X1 U9025 ( .A1(n9224), .A2(n7999), .ZN(n9223) );
  NOR2_X1 U9026 ( .A1(n8788), .A2(n8790), .ZN(n9224) );
  NAND2_X1 U9027 ( .A1(n8788), .A2(n8790), .ZN(n9221) );
  NAND2_X1 U9028 ( .A1(n9225), .A2(n9226), .ZN(n8790) );
  NAND2_X1 U9029 ( .A1(n8764), .A2(n9227), .ZN(n9226) );
  OR2_X1 U9030 ( .A1(n8763), .A2(n8762), .ZN(n9227) );
  NOR2_X1 U9031 ( .A1(n8778), .A2(n7999), .ZN(n8764) );
  NAND2_X1 U9032 ( .A1(n8762), .A2(n8763), .ZN(n9225) );
  NAND2_X1 U9033 ( .A1(n9228), .A2(n9229), .ZN(n8763) );
  NAND2_X1 U9034 ( .A1(n9230), .A2(a_4_), .ZN(n9229) );
  NOR2_X1 U9035 ( .A1(n9231), .A2(n7999), .ZN(n9230) );
  NOR2_X1 U9036 ( .A1(n8733), .A2(n8735), .ZN(n9231) );
  NAND2_X1 U9037 ( .A1(n8733), .A2(n8735), .ZN(n9228) );
  NAND2_X1 U9038 ( .A1(n9232), .A2(n9233), .ZN(n8735) );
  NAND2_X1 U9039 ( .A1(n8709), .A2(n9234), .ZN(n9233) );
  OR2_X1 U9040 ( .A1(n8708), .A2(n8707), .ZN(n9234) );
  NOR2_X1 U9041 ( .A1(n8723), .A2(n7999), .ZN(n8709) );
  NAND2_X1 U9042 ( .A1(n8707), .A2(n8708), .ZN(n9232) );
  NAND2_X1 U9043 ( .A1(n9235), .A2(n9236), .ZN(n8708) );
  NAND2_X1 U9044 ( .A1(n9237), .A2(a_6_), .ZN(n9236) );
  NOR2_X1 U9045 ( .A1(n9238), .A2(n7999), .ZN(n9237) );
  NOR2_X1 U9046 ( .A1(n8678), .A2(n8679), .ZN(n9238) );
  NAND2_X1 U9047 ( .A1(n8678), .A2(n8679), .ZN(n9235) );
  NAND2_X1 U9048 ( .A1(n9239), .A2(n9240), .ZN(n8679) );
  NAND2_X1 U9049 ( .A1(n8653), .A2(n9241), .ZN(n9240) );
  OR2_X1 U9050 ( .A1(n8652), .A2(n8651), .ZN(n9241) );
  NOR2_X1 U9051 ( .A1(n8962), .A2(n7999), .ZN(n8653) );
  NAND2_X1 U9052 ( .A1(n8651), .A2(n8652), .ZN(n9239) );
  NAND2_X1 U9053 ( .A1(n9242), .A2(n9243), .ZN(n8652) );
  NAND2_X1 U9054 ( .A1(n9244), .A2(a_8_), .ZN(n9243) );
  NOR2_X1 U9055 ( .A1(n9245), .A2(n7999), .ZN(n9244) );
  NOR2_X1 U9056 ( .A1(n8615), .A2(n8617), .ZN(n9245) );
  NAND2_X1 U9057 ( .A1(n8615), .A2(n8617), .ZN(n9242) );
  NAND2_X1 U9058 ( .A1(n9246), .A2(n9247), .ZN(n8617) );
  NAND2_X1 U9059 ( .A1(n8591), .A2(n9248), .ZN(n9247) );
  NAND2_X1 U9060 ( .A1(n8590), .A2(n8588), .ZN(n9248) );
  NOR2_X1 U9061 ( .A1(n8605), .A2(n7999), .ZN(n8591) );
  OR2_X1 U9062 ( .A1(n8588), .A2(n8590), .ZN(n9246) );
  AND2_X1 U9063 ( .A1(n9249), .A2(n9250), .ZN(n8590) );
  NAND2_X1 U9064 ( .A1(n9251), .A2(a_10_), .ZN(n9250) );
  NOR2_X1 U9065 ( .A1(n9252), .A2(n7999), .ZN(n9251) );
  NOR2_X1 U9066 ( .A1(n8560), .A2(n8562), .ZN(n9252) );
  NAND2_X1 U9067 ( .A1(n8560), .A2(n8562), .ZN(n9249) );
  NAND2_X1 U9068 ( .A1(n9253), .A2(n9254), .ZN(n8562) );
  NAND2_X1 U9069 ( .A1(n8536), .A2(n9255), .ZN(n9254) );
  OR2_X1 U9070 ( .A1(n8535), .A2(n8534), .ZN(n9255) );
  NOR2_X1 U9071 ( .A1(n8550), .A2(n7999), .ZN(n8536) );
  NAND2_X1 U9072 ( .A1(n8534), .A2(n8535), .ZN(n9253) );
  NAND2_X1 U9073 ( .A1(n9256), .A2(n9257), .ZN(n8535) );
  NAND2_X1 U9074 ( .A1(n9258), .A2(a_12_), .ZN(n9257) );
  NOR2_X1 U9075 ( .A1(n9259), .A2(n7999), .ZN(n9258) );
  NOR2_X1 U9076 ( .A1(n8505), .A2(n8507), .ZN(n9259) );
  NAND2_X1 U9077 ( .A1(n8505), .A2(n8507), .ZN(n9256) );
  NAND2_X1 U9078 ( .A1(n9260), .A2(n9261), .ZN(n8507) );
  NAND2_X1 U9079 ( .A1(n8481), .A2(n9262), .ZN(n9261) );
  OR2_X1 U9080 ( .A1(n8480), .A2(n8479), .ZN(n9262) );
  NOR2_X1 U9081 ( .A1(n8495), .A2(n7999), .ZN(n8481) );
  NAND2_X1 U9082 ( .A1(n8479), .A2(n8480), .ZN(n9260) );
  NAND2_X1 U9083 ( .A1(n9263), .A2(n9264), .ZN(n8480) );
  NAND2_X1 U9084 ( .A1(n9265), .A2(a_14_), .ZN(n9264) );
  NOR2_X1 U9085 ( .A1(n9266), .A2(n7999), .ZN(n9265) );
  NOR2_X1 U9086 ( .A1(n8450), .A2(n8452), .ZN(n9266) );
  NAND2_X1 U9087 ( .A1(n8450), .A2(n8452), .ZN(n9263) );
  NAND2_X1 U9088 ( .A1(n9267), .A2(n9268), .ZN(n8452) );
  NAND2_X1 U9089 ( .A1(n8426), .A2(n9269), .ZN(n9268) );
  OR2_X1 U9090 ( .A1(n8425), .A2(n8424), .ZN(n9269) );
  NOR2_X1 U9091 ( .A1(n8440), .A2(n7999), .ZN(n8426) );
  NAND2_X1 U9092 ( .A1(n8424), .A2(n8425), .ZN(n9267) );
  NAND2_X1 U9093 ( .A1(n9270), .A2(n9271), .ZN(n8425) );
  NAND2_X1 U9094 ( .A1(n9272), .A2(a_16_), .ZN(n9271) );
  NOR2_X1 U9095 ( .A1(n9273), .A2(n7999), .ZN(n9272) );
  NOR2_X1 U9096 ( .A1(n8395), .A2(n8397), .ZN(n9273) );
  NAND2_X1 U9097 ( .A1(n8395), .A2(n8397), .ZN(n9270) );
  NAND2_X1 U9098 ( .A1(n9274), .A2(n9275), .ZN(n8397) );
  NAND2_X1 U9099 ( .A1(n8371), .A2(n9276), .ZN(n9275) );
  OR2_X1 U9100 ( .A1(n8370), .A2(n8368), .ZN(n9276) );
  NOR2_X1 U9101 ( .A1(n8385), .A2(n7999), .ZN(n8371) );
  NAND2_X1 U9102 ( .A1(n8368), .A2(n8370), .ZN(n9274) );
  NAND2_X1 U9103 ( .A1(n9277), .A2(n9278), .ZN(n8370) );
  NAND2_X1 U9104 ( .A1(n9279), .A2(a_18_), .ZN(n9278) );
  NOR2_X1 U9105 ( .A1(n9280), .A2(n7999), .ZN(n9279) );
  NOR2_X1 U9106 ( .A1(n8334), .A2(n8337), .ZN(n9280) );
  NAND2_X1 U9107 ( .A1(n8334), .A2(n8337), .ZN(n9277) );
  NAND2_X1 U9108 ( .A1(n9281), .A2(n9282), .ZN(n8337) );
  NAND2_X1 U9109 ( .A1(n8307), .A2(n9283), .ZN(n9282) );
  OR2_X1 U9110 ( .A1(n8309), .A2(n8310), .ZN(n9283) );
  XOR2_X1 U9111 ( .A(n9284), .B(n9285), .Z(n8307) );
  XNOR2_X1 U9112 ( .A(n9286), .B(n9287), .ZN(n9284) );
  NAND2_X1 U9113 ( .A1(a_20_), .A2(b_30_), .ZN(n9286) );
  NAND2_X1 U9114 ( .A1(n8310), .A2(n8309), .ZN(n9281) );
  NAND2_X1 U9115 ( .A1(n9288), .A2(n9289), .ZN(n8309) );
  NAND2_X1 U9116 ( .A1(n9290), .A2(a_20_), .ZN(n9289) );
  NOR2_X1 U9117 ( .A1(n9291), .A2(n7999), .ZN(n9290) );
  NOR2_X1 U9118 ( .A1(n8278), .A2(n8280), .ZN(n9291) );
  NAND2_X1 U9119 ( .A1(n8278), .A2(n8280), .ZN(n9288) );
  NAND2_X1 U9120 ( .A1(n9292), .A2(n9293), .ZN(n8280) );
  NAND2_X1 U9121 ( .A1(n9294), .A2(a_21_), .ZN(n9293) );
  NOR2_X1 U9122 ( .A1(n9295), .A2(n7999), .ZN(n9294) );
  NOR2_X1 U9123 ( .A1(n8251), .A2(n8253), .ZN(n9295) );
  NAND2_X1 U9124 ( .A1(n8251), .A2(n8253), .ZN(n9292) );
  NAND2_X1 U9125 ( .A1(n9296), .A2(n9297), .ZN(n8253) );
  NAND2_X1 U9126 ( .A1(n9298), .A2(a_22_), .ZN(n9297) );
  NOR2_X1 U9127 ( .A1(n9299), .A2(n7999), .ZN(n9298) );
  NOR2_X1 U9128 ( .A1(n8223), .A2(n8225), .ZN(n9299) );
  NAND2_X1 U9129 ( .A1(n8223), .A2(n8225), .ZN(n9296) );
  NAND2_X1 U9130 ( .A1(n8198), .A2(n9300), .ZN(n8225) );
  NAND2_X1 U9131 ( .A1(n8197), .A2(n8199), .ZN(n9300) );
  NAND2_X1 U9132 ( .A1(n9301), .A2(n9302), .ZN(n8199) );
  NAND2_X1 U9133 ( .A1(a_23_), .A2(b_31_), .ZN(n9302) );
  INV_X1 U9134 ( .A(n9303), .ZN(n9301) );
  XOR2_X1 U9135 ( .A(n9304), .B(n9305), .Z(n8197) );
  XOR2_X1 U9136 ( .A(n9306), .B(n9307), .Z(n9304) );
  NOR2_X1 U9137 ( .A1(n8002), .A2(n8939), .ZN(n9307) );
  NAND2_X1 U9138 ( .A1(a_23_), .A2(n9303), .ZN(n8198) );
  NAND2_X1 U9139 ( .A1(n9308), .A2(n9309), .ZN(n9303) );
  NAND2_X1 U9140 ( .A1(n9310), .A2(a_24_), .ZN(n9309) );
  NOR2_X1 U9141 ( .A1(n9311), .A2(n7999), .ZN(n9310) );
  NOR2_X1 U9142 ( .A1(n8168), .A2(n8171), .ZN(n9311) );
  NAND2_X1 U9143 ( .A1(n8168), .A2(n8171), .ZN(n9308) );
  NAND2_X1 U9144 ( .A1(n8143), .A2(n9312), .ZN(n8171) );
  NAND2_X1 U9145 ( .A1(n8142), .A2(n8144), .ZN(n9312) );
  NAND2_X1 U9146 ( .A1(n9313), .A2(n9314), .ZN(n8144) );
  NAND2_X1 U9147 ( .A1(a_25_), .A2(b_31_), .ZN(n9314) );
  INV_X1 U9148 ( .A(n9315), .ZN(n9313) );
  XNOR2_X1 U9149 ( .A(n9316), .B(n9317), .ZN(n8142) );
  NAND2_X1 U9150 ( .A1(n9318), .A2(n9319), .ZN(n9316) );
  NAND2_X1 U9151 ( .A1(a_25_), .A2(n9315), .ZN(n8143) );
  NAND2_X1 U9152 ( .A1(n9320), .A2(n9321), .ZN(n9315) );
  NAND2_X1 U9153 ( .A1(n9322), .A2(a_26_), .ZN(n9321) );
  NOR2_X1 U9154 ( .A1(n9323), .A2(n7999), .ZN(n9322) );
  NOR2_X1 U9155 ( .A1(n8113), .A2(n8114), .ZN(n9323) );
  NAND2_X1 U9156 ( .A1(n8113), .A2(n8114), .ZN(n9320) );
  NAND2_X1 U9157 ( .A1(n9324), .A2(n9325), .ZN(n8114) );
  NAND2_X1 U9158 ( .A1(n9326), .A2(a_27_), .ZN(n9325) );
  NOR2_X1 U9159 ( .A1(n9327), .A2(n7999), .ZN(n9326) );
  NOR2_X1 U9160 ( .A1(n8085), .A2(n8087), .ZN(n9327) );
  NAND2_X1 U9161 ( .A1(n8085), .A2(n8087), .ZN(n9324) );
  NAND2_X1 U9162 ( .A1(n9328), .A2(n9329), .ZN(n8087) );
  NAND2_X1 U9163 ( .A1(n9330), .A2(a_28_), .ZN(n9329) );
  NOR2_X1 U9164 ( .A1(n9331), .A2(n7999), .ZN(n9330) );
  NOR2_X1 U9165 ( .A1(n8051), .A2(n8053), .ZN(n9331) );
  NAND2_X1 U9166 ( .A1(n8051), .A2(n8053), .ZN(n9328) );
  NAND2_X1 U9167 ( .A1(n9332), .A2(n9333), .ZN(n8053) );
  NAND2_X1 U9168 ( .A1(n8027), .A2(n9334), .ZN(n9333) );
  OR2_X1 U9169 ( .A1(n8026), .A2(n8025), .ZN(n9334) );
  AND2_X1 U9170 ( .A1(n9335), .A2(n7953), .ZN(n8027) );
  NOR2_X1 U9171 ( .A1(n7999), .A2(n8002), .ZN(n9335) );
  NAND2_X1 U9172 ( .A1(n8025), .A2(n8026), .ZN(n9332) );
  NAND2_X1 U9173 ( .A1(n9336), .A2(n9337), .ZN(n8026) );
  NAND2_X1 U9174 ( .A1(b_29_), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U9175 ( .A1(n8003), .A2(n9339), .ZN(n9338) );
  NAND2_X1 U9176 ( .A1(a_31_), .A2(n8002), .ZN(n9339) );
  NAND2_X1 U9177 ( .A1(b_30_), .A2(n9340), .ZN(n9336) );
  NAND2_X1 U9178 ( .A1(n9341), .A2(n9342), .ZN(n9340) );
  NAND2_X1 U9179 ( .A1(a_30_), .A2(n8936), .ZN(n9342) );
  NOR2_X1 U9180 ( .A1(n8041), .A2(n7999), .ZN(n8025) );
  XOR2_X1 U9181 ( .A(n9343), .B(n9344), .Z(n8051) );
  XOR2_X1 U9182 ( .A(n9345), .B(n9346), .Z(n9343) );
  XOR2_X1 U9183 ( .A(n9347), .B(n9348), .Z(n8085) );
  XNOR2_X1 U9184 ( .A(n9349), .B(n9350), .ZN(n9347) );
  NAND2_X1 U9185 ( .A1(a_28_), .A2(b_30_), .ZN(n9349) );
  XNOR2_X1 U9186 ( .A(n9351), .B(n9352), .ZN(n8113) );
  NAND2_X1 U9187 ( .A1(n9353), .A2(n9354), .ZN(n9351) );
  XNOR2_X1 U9188 ( .A(n9355), .B(n9356), .ZN(n8168) );
  XNOR2_X1 U9189 ( .A(n9357), .B(n9358), .ZN(n9356) );
  XOR2_X1 U9190 ( .A(n9359), .B(n9360), .Z(n8223) );
  XOR2_X1 U9191 ( .A(n9361), .B(n9362), .Z(n9359) );
  XOR2_X1 U9192 ( .A(n9363), .B(n9364), .Z(n8251) );
  XOR2_X1 U9193 ( .A(n9365), .B(n9366), .Z(n9363) );
  NOR2_X1 U9194 ( .A1(n8002), .A2(n8941), .ZN(n9366) );
  XNOR2_X1 U9195 ( .A(n9367), .B(n9368), .ZN(n8278) );
  XNOR2_X1 U9196 ( .A(n9369), .B(n9370), .ZN(n9368) );
  NOR2_X1 U9197 ( .A1(n8324), .A2(n7999), .ZN(n8310) );
  XNOR2_X1 U9198 ( .A(n9371), .B(n9372), .ZN(n8334) );
  XNOR2_X1 U9199 ( .A(n9373), .B(n9374), .ZN(n9372) );
  XOR2_X1 U9200 ( .A(n9375), .B(n9376), .Z(n8368) );
  XNOR2_X1 U9201 ( .A(n9377), .B(n9378), .ZN(n9375) );
  NAND2_X1 U9202 ( .A1(a_18_), .A2(b_30_), .ZN(n9377) );
  XOR2_X1 U9203 ( .A(n9379), .B(n9380), .Z(n8395) );
  XOR2_X1 U9204 ( .A(n9381), .B(n9382), .Z(n9379) );
  XOR2_X1 U9205 ( .A(n9383), .B(n9384), .Z(n8424) );
  XOR2_X1 U9206 ( .A(n9385), .B(n9386), .Z(n9383) );
  NOR2_X1 U9207 ( .A1(n8002), .A2(n8950), .ZN(n9386) );
  XOR2_X1 U9208 ( .A(n9387), .B(n9388), .Z(n8450) );
  XOR2_X1 U9209 ( .A(n9389), .B(n9390), .Z(n9387) );
  XOR2_X1 U9210 ( .A(n9391), .B(n9392), .Z(n8479) );
  XOR2_X1 U9211 ( .A(n9393), .B(n9394), .Z(n9391) );
  NOR2_X1 U9212 ( .A1(n8002), .A2(n8953), .ZN(n9394) );
  XOR2_X1 U9213 ( .A(n9395), .B(n9396), .Z(n8505) );
  XOR2_X1 U9214 ( .A(n9397), .B(n9398), .Z(n9395) );
  XOR2_X1 U9215 ( .A(n9399), .B(n9400), .Z(n8534) );
  XOR2_X1 U9216 ( .A(n9401), .B(n9402), .Z(n9399) );
  NOR2_X1 U9217 ( .A1(n8002), .A2(n8956), .ZN(n9402) );
  XOR2_X1 U9218 ( .A(n9403), .B(n9404), .Z(n8560) );
  XOR2_X1 U9219 ( .A(n9405), .B(n9406), .Z(n9403) );
  XOR2_X1 U9220 ( .A(n9407), .B(n9408), .Z(n8588) );
  XOR2_X1 U9221 ( .A(n9409), .B(n9410), .Z(n9408) );
  NAND2_X1 U9222 ( .A1(a_10_), .A2(b_30_), .ZN(n9410) );
  XOR2_X1 U9223 ( .A(n9411), .B(n9412), .Z(n8615) );
  XOR2_X1 U9224 ( .A(n9413), .B(n9414), .Z(n9411) );
  XOR2_X1 U9225 ( .A(n9415), .B(n9416), .Z(n8651) );
  XOR2_X1 U9226 ( .A(n9417), .B(n9418), .Z(n9415) );
  NOR2_X1 U9227 ( .A1(n8002), .A2(n8619), .ZN(n9418) );
  XNOR2_X1 U9228 ( .A(n9419), .B(n9420), .ZN(n8678) );
  XNOR2_X1 U9229 ( .A(n9421), .B(n9422), .ZN(n9419) );
  XOR2_X1 U9230 ( .A(n9423), .B(n9424), .Z(n8707) );
  XOR2_X1 U9231 ( .A(n9425), .B(n9426), .Z(n9423) );
  NOR2_X1 U9232 ( .A1(n8002), .A2(n8681), .ZN(n9426) );
  XOR2_X1 U9233 ( .A(n9427), .B(n9428), .Z(n8733) );
  XOR2_X1 U9234 ( .A(n9429), .B(n9430), .Z(n9427) );
  XNOR2_X1 U9235 ( .A(n9431), .B(n9432), .ZN(n8762) );
  XOR2_X1 U9236 ( .A(n9433), .B(n9434), .Z(n9432) );
  NAND2_X1 U9237 ( .A1(a_4_), .A2(b_30_), .ZN(n9434) );
  XOR2_X1 U9238 ( .A(n9435), .B(n9436), .Z(n8788) );
  XOR2_X1 U9239 ( .A(n9437), .B(n9438), .Z(n9435) );
  XNOR2_X1 U9240 ( .A(n9439), .B(n9440), .ZN(n8817) );
  XOR2_X1 U9241 ( .A(n9441), .B(n9442), .Z(n9439) );
  NOR2_X1 U9242 ( .A1(n8002), .A2(n8792), .ZN(n9442) );
  XOR2_X1 U9243 ( .A(n9443), .B(n9444), .Z(n8844) );
  XNOR2_X1 U9244 ( .A(n9445), .B(n9446), .ZN(n9443) );
  NAND2_X1 U9245 ( .A1(a_1_), .A2(b_30_), .ZN(n9445) );
  NAND2_X1 U9246 ( .A1(n9447), .A2(n9448), .ZN(n8996) );
  XOR2_X1 U9247 ( .A(n9202), .B(n9201), .Z(n9448) );
  AND2_X1 U9248 ( .A1(n9209), .A2(n9208), .ZN(n9447) );
  XOR2_X1 U9249 ( .A(n9449), .B(n9450), .Z(n9208) );
  XOR2_X1 U9250 ( .A(n9451), .B(n9452), .Z(n9449) );
  NOR2_X1 U9251 ( .A1(n8974), .A2(n8936), .ZN(n9452) );
  NAND2_X1 U9252 ( .A1(n9453), .A2(n9454), .ZN(n9209) );
  NAND2_X1 U9253 ( .A1(n9455), .A2(a_0_), .ZN(n9454) );
  NOR2_X1 U9254 ( .A1(n9456), .A2(n8002), .ZN(n9455) );
  NOR2_X1 U9255 ( .A1(n9211), .A2(n9212), .ZN(n9456) );
  NAND2_X1 U9256 ( .A1(n9211), .A2(n9212), .ZN(n9453) );
  NAND2_X1 U9257 ( .A1(n9457), .A2(n9458), .ZN(n9212) );
  NAND2_X1 U9258 ( .A1(n9459), .A2(a_1_), .ZN(n9458) );
  NOR2_X1 U9259 ( .A1(n9460), .A2(n8002), .ZN(n9459) );
  NOR2_X1 U9260 ( .A1(n9446), .A2(n9444), .ZN(n9460) );
  NAND2_X1 U9261 ( .A1(n9444), .A2(n9446), .ZN(n9457) );
  NAND2_X1 U9262 ( .A1(n9461), .A2(n9462), .ZN(n9446) );
  NAND2_X1 U9263 ( .A1(n9463), .A2(a_2_), .ZN(n9462) );
  NOR2_X1 U9264 ( .A1(n9464), .A2(n8002), .ZN(n9463) );
  NOR2_X1 U9265 ( .A1(n9441), .A2(n9440), .ZN(n9464) );
  NAND2_X1 U9266 ( .A1(n9440), .A2(n9441), .ZN(n9461) );
  NAND2_X1 U9267 ( .A1(n9465), .A2(n9466), .ZN(n9441) );
  NAND2_X1 U9268 ( .A1(n9438), .A2(n9467), .ZN(n9466) );
  OR2_X1 U9269 ( .A1(n9436), .A2(n9437), .ZN(n9467) );
  NOR2_X1 U9270 ( .A1(n8778), .A2(n8002), .ZN(n9438) );
  NAND2_X1 U9271 ( .A1(n9436), .A2(n9437), .ZN(n9465) );
  NAND2_X1 U9272 ( .A1(n9468), .A2(n9469), .ZN(n9437) );
  NAND2_X1 U9273 ( .A1(n9470), .A2(a_4_), .ZN(n9469) );
  NOR2_X1 U9274 ( .A1(n9471), .A2(n8002), .ZN(n9470) );
  NOR2_X1 U9275 ( .A1(n9431), .A2(n9433), .ZN(n9471) );
  NAND2_X1 U9276 ( .A1(n9431), .A2(n9433), .ZN(n9468) );
  NAND2_X1 U9277 ( .A1(n9472), .A2(n9473), .ZN(n9433) );
  NAND2_X1 U9278 ( .A1(n9430), .A2(n9474), .ZN(n9473) );
  OR2_X1 U9279 ( .A1(n9428), .A2(n9429), .ZN(n9474) );
  NOR2_X1 U9280 ( .A1(n8723), .A2(n8002), .ZN(n9430) );
  NAND2_X1 U9281 ( .A1(n9428), .A2(n9429), .ZN(n9472) );
  NAND2_X1 U9282 ( .A1(n9475), .A2(n9476), .ZN(n9429) );
  NAND2_X1 U9283 ( .A1(n9477), .A2(a_6_), .ZN(n9476) );
  NOR2_X1 U9284 ( .A1(n9478), .A2(n8002), .ZN(n9477) );
  NOR2_X1 U9285 ( .A1(n9424), .A2(n9425), .ZN(n9478) );
  NAND2_X1 U9286 ( .A1(n9424), .A2(n9425), .ZN(n9475) );
  NAND2_X1 U9287 ( .A1(n9479), .A2(n9480), .ZN(n9425) );
  NAND2_X1 U9288 ( .A1(n9422), .A2(n9481), .ZN(n9480) );
  NAND2_X1 U9289 ( .A1(n9421), .A2(n9420), .ZN(n9481) );
  NOR2_X1 U9290 ( .A1(n8962), .A2(n8002), .ZN(n9422) );
  OR2_X1 U9291 ( .A1(n9420), .A2(n9421), .ZN(n9479) );
  AND2_X1 U9292 ( .A1(n9482), .A2(n9483), .ZN(n9421) );
  NAND2_X1 U9293 ( .A1(n9484), .A2(a_8_), .ZN(n9483) );
  NOR2_X1 U9294 ( .A1(n9485), .A2(n8002), .ZN(n9484) );
  NOR2_X1 U9295 ( .A1(n9416), .A2(n9417), .ZN(n9485) );
  NAND2_X1 U9296 ( .A1(n9416), .A2(n9417), .ZN(n9482) );
  NAND2_X1 U9297 ( .A1(n9486), .A2(n9487), .ZN(n9417) );
  NAND2_X1 U9298 ( .A1(n9414), .A2(n9488), .ZN(n9487) );
  OR2_X1 U9299 ( .A1(n9412), .A2(n9413), .ZN(n9488) );
  NOR2_X1 U9300 ( .A1(n8605), .A2(n8002), .ZN(n9414) );
  NAND2_X1 U9301 ( .A1(n9412), .A2(n9413), .ZN(n9486) );
  NAND2_X1 U9302 ( .A1(n9489), .A2(n9490), .ZN(n9413) );
  NAND2_X1 U9303 ( .A1(n9491), .A2(a_10_), .ZN(n9490) );
  NOR2_X1 U9304 ( .A1(n9492), .A2(n8002), .ZN(n9491) );
  NOR2_X1 U9305 ( .A1(n9409), .A2(n9407), .ZN(n9492) );
  NAND2_X1 U9306 ( .A1(n9407), .A2(n9409), .ZN(n9489) );
  NAND2_X1 U9307 ( .A1(n9493), .A2(n9494), .ZN(n9409) );
  NAND2_X1 U9308 ( .A1(n9406), .A2(n9495), .ZN(n9494) );
  OR2_X1 U9309 ( .A1(n9404), .A2(n9405), .ZN(n9495) );
  NOR2_X1 U9310 ( .A1(n8550), .A2(n8002), .ZN(n9406) );
  NAND2_X1 U9311 ( .A1(n9404), .A2(n9405), .ZN(n9493) );
  NAND2_X1 U9312 ( .A1(n9496), .A2(n9497), .ZN(n9405) );
  NAND2_X1 U9313 ( .A1(n9498), .A2(a_12_), .ZN(n9497) );
  NOR2_X1 U9314 ( .A1(n9499), .A2(n8002), .ZN(n9498) );
  NOR2_X1 U9315 ( .A1(n9400), .A2(n9401), .ZN(n9499) );
  NAND2_X1 U9316 ( .A1(n9400), .A2(n9401), .ZN(n9496) );
  NAND2_X1 U9317 ( .A1(n9500), .A2(n9501), .ZN(n9401) );
  NAND2_X1 U9318 ( .A1(n9398), .A2(n9502), .ZN(n9501) );
  OR2_X1 U9319 ( .A1(n9396), .A2(n9397), .ZN(n9502) );
  NOR2_X1 U9320 ( .A1(n8495), .A2(n8002), .ZN(n9398) );
  NAND2_X1 U9321 ( .A1(n9396), .A2(n9397), .ZN(n9500) );
  NAND2_X1 U9322 ( .A1(n9503), .A2(n9504), .ZN(n9397) );
  NAND2_X1 U9323 ( .A1(n9505), .A2(a_14_), .ZN(n9504) );
  NOR2_X1 U9324 ( .A1(n9506), .A2(n8002), .ZN(n9505) );
  NOR2_X1 U9325 ( .A1(n9392), .A2(n9393), .ZN(n9506) );
  NAND2_X1 U9326 ( .A1(n9392), .A2(n9393), .ZN(n9503) );
  NAND2_X1 U9327 ( .A1(n9507), .A2(n9508), .ZN(n9393) );
  NAND2_X1 U9328 ( .A1(n9390), .A2(n9509), .ZN(n9508) );
  OR2_X1 U9329 ( .A1(n9388), .A2(n9389), .ZN(n9509) );
  NOR2_X1 U9330 ( .A1(n8440), .A2(n8002), .ZN(n9390) );
  NAND2_X1 U9331 ( .A1(n9388), .A2(n9389), .ZN(n9507) );
  NAND2_X1 U9332 ( .A1(n9510), .A2(n9511), .ZN(n9389) );
  NAND2_X1 U9333 ( .A1(n9512), .A2(a_16_), .ZN(n9511) );
  NOR2_X1 U9334 ( .A1(n9513), .A2(n8002), .ZN(n9512) );
  NOR2_X1 U9335 ( .A1(n9384), .A2(n9385), .ZN(n9513) );
  NAND2_X1 U9336 ( .A1(n9384), .A2(n9385), .ZN(n9510) );
  NAND2_X1 U9337 ( .A1(n9514), .A2(n9515), .ZN(n9385) );
  NAND2_X1 U9338 ( .A1(n9382), .A2(n9516), .ZN(n9515) );
  OR2_X1 U9339 ( .A1(n9380), .A2(n9381), .ZN(n9516) );
  NOR2_X1 U9340 ( .A1(n8385), .A2(n8002), .ZN(n9382) );
  NAND2_X1 U9341 ( .A1(n9380), .A2(n9381), .ZN(n9514) );
  NAND2_X1 U9342 ( .A1(n9517), .A2(n9518), .ZN(n9381) );
  NAND2_X1 U9343 ( .A1(n9519), .A2(a_18_), .ZN(n9518) );
  NOR2_X1 U9344 ( .A1(n9520), .A2(n8002), .ZN(n9519) );
  NOR2_X1 U9345 ( .A1(n9376), .A2(n9378), .ZN(n9520) );
  NAND2_X1 U9346 ( .A1(n9376), .A2(n9378), .ZN(n9517) );
  NAND2_X1 U9347 ( .A1(n9521), .A2(n9522), .ZN(n9378) );
  NAND2_X1 U9348 ( .A1(n9374), .A2(n9523), .ZN(n9522) );
  OR2_X1 U9349 ( .A1(n9371), .A2(n9373), .ZN(n9523) );
  NOR2_X1 U9350 ( .A1(n8324), .A2(n8002), .ZN(n9374) );
  NAND2_X1 U9351 ( .A1(n9371), .A2(n9373), .ZN(n9521) );
  NAND2_X1 U9352 ( .A1(n9524), .A2(n9525), .ZN(n9373) );
  NAND2_X1 U9353 ( .A1(n9526), .A2(a_20_), .ZN(n9525) );
  NOR2_X1 U9354 ( .A1(n9527), .A2(n8002), .ZN(n9526) );
  NOR2_X1 U9355 ( .A1(n9285), .A2(n9287), .ZN(n9527) );
  NAND2_X1 U9356 ( .A1(n9285), .A2(n9287), .ZN(n9524) );
  NAND2_X1 U9357 ( .A1(n9528), .A2(n9529), .ZN(n9287) );
  NAND2_X1 U9358 ( .A1(n9370), .A2(n9530), .ZN(n9529) );
  OR2_X1 U9359 ( .A1(n9367), .A2(n9369), .ZN(n9530) );
  NOR2_X1 U9360 ( .A1(n8268), .A2(n8002), .ZN(n9370) );
  NAND2_X1 U9361 ( .A1(n9367), .A2(n9369), .ZN(n9528) );
  NAND2_X1 U9362 ( .A1(n9531), .A2(n9532), .ZN(n9369) );
  NAND2_X1 U9363 ( .A1(n9533), .A2(a_22_), .ZN(n9532) );
  NOR2_X1 U9364 ( .A1(n9534), .A2(n8002), .ZN(n9533) );
  NOR2_X1 U9365 ( .A1(n9365), .A2(n9364), .ZN(n9534) );
  NAND2_X1 U9366 ( .A1(n9364), .A2(n9365), .ZN(n9531) );
  NAND2_X1 U9367 ( .A1(n9535), .A2(n9536), .ZN(n9365) );
  NAND2_X1 U9368 ( .A1(n9362), .A2(n9537), .ZN(n9536) );
  OR2_X1 U9369 ( .A1(n9360), .A2(n9361), .ZN(n9537) );
  NOR2_X1 U9370 ( .A1(n8213), .A2(n8002), .ZN(n9362) );
  NAND2_X1 U9371 ( .A1(n9360), .A2(n9361), .ZN(n9535) );
  NAND2_X1 U9372 ( .A1(n9538), .A2(n9539), .ZN(n9361) );
  NAND2_X1 U9373 ( .A1(n9540), .A2(a_24_), .ZN(n9539) );
  NOR2_X1 U9374 ( .A1(n9541), .A2(n8002), .ZN(n9540) );
  NOR2_X1 U9375 ( .A1(n9306), .A2(n9305), .ZN(n9541) );
  NAND2_X1 U9376 ( .A1(n9305), .A2(n9306), .ZN(n9538) );
  NAND2_X1 U9377 ( .A1(n9542), .A2(n9543), .ZN(n9306) );
  NAND2_X1 U9378 ( .A1(n9358), .A2(n9544), .ZN(n9543) );
  OR2_X1 U9379 ( .A1(n9355), .A2(n9357), .ZN(n9544) );
  NOR2_X1 U9380 ( .A1(n8158), .A2(n8002), .ZN(n9358) );
  NAND2_X1 U9381 ( .A1(n9355), .A2(n9357), .ZN(n9542) );
  NAND2_X1 U9382 ( .A1(n9318), .A2(n9545), .ZN(n9357) );
  NAND2_X1 U9383 ( .A1(n9317), .A2(n9319), .ZN(n9545) );
  NAND2_X1 U9384 ( .A1(n9546), .A2(n9547), .ZN(n9319) );
  NAND2_X1 U9385 ( .A1(a_26_), .A2(b_30_), .ZN(n9547) );
  INV_X1 U9386 ( .A(n9548), .ZN(n9546) );
  XNOR2_X1 U9387 ( .A(n9549), .B(n9550), .ZN(n9317) );
  NAND2_X1 U9388 ( .A1(n9551), .A2(n9552), .ZN(n9549) );
  NAND2_X1 U9389 ( .A1(a_26_), .A2(n9548), .ZN(n9318) );
  NAND2_X1 U9390 ( .A1(n9353), .A2(n9553), .ZN(n9548) );
  NAND2_X1 U9391 ( .A1(n9352), .A2(n9354), .ZN(n9553) );
  NAND2_X1 U9392 ( .A1(n9554), .A2(n9555), .ZN(n9354) );
  NAND2_X1 U9393 ( .A1(a_27_), .A2(b_30_), .ZN(n9555) );
  INV_X1 U9394 ( .A(n9556), .ZN(n9554) );
  XOR2_X1 U9395 ( .A(n9557), .B(n9558), .Z(n9352) );
  XNOR2_X1 U9396 ( .A(n9559), .B(n9560), .ZN(n9557) );
  NAND2_X1 U9397 ( .A1(b_29_), .A2(a_28_), .ZN(n9559) );
  NAND2_X1 U9398 ( .A1(a_27_), .A2(n9556), .ZN(n9353) );
  NAND2_X1 U9399 ( .A1(n9561), .A2(n9562), .ZN(n9556) );
  NAND2_X1 U9400 ( .A1(n9563), .A2(a_28_), .ZN(n9562) );
  NOR2_X1 U9401 ( .A1(n9564), .A2(n8002), .ZN(n9563) );
  NOR2_X1 U9402 ( .A1(n9348), .A2(n9350), .ZN(n9564) );
  NAND2_X1 U9403 ( .A1(n9348), .A2(n9350), .ZN(n9561) );
  NAND2_X1 U9404 ( .A1(n9565), .A2(n9566), .ZN(n9350) );
  NAND2_X1 U9405 ( .A1(n9344), .A2(n9567), .ZN(n9566) );
  OR2_X1 U9406 ( .A1(n9345), .A2(n9346), .ZN(n9567) );
  NOR2_X1 U9407 ( .A1(n8041), .A2(n8002), .ZN(n9344) );
  NAND2_X1 U9408 ( .A1(n9346), .A2(n9345), .ZN(n9565) );
  NAND2_X1 U9409 ( .A1(n9568), .A2(n9569), .ZN(n9345) );
  NAND2_X1 U9410 ( .A1(b_28_), .A2(n9570), .ZN(n9569) );
  NAND2_X1 U9411 ( .A1(n8003), .A2(n9571), .ZN(n9570) );
  NAND2_X1 U9412 ( .A1(a_31_), .A2(n8936), .ZN(n9571) );
  NAND2_X1 U9413 ( .A1(b_29_), .A2(n9572), .ZN(n9568) );
  NAND2_X1 U9414 ( .A1(n9341), .A2(n9573), .ZN(n9572) );
  NAND2_X1 U9415 ( .A1(a_30_), .A2(n8069), .ZN(n9573) );
  AND2_X1 U9416 ( .A1(n9574), .A2(n7953), .ZN(n9346) );
  NOR2_X1 U9417 ( .A1(n8002), .A2(n8936), .ZN(n9574) );
  XNOR2_X1 U9418 ( .A(n9575), .B(n8929), .ZN(n9348) );
  XOR2_X1 U9419 ( .A(n9576), .B(n9577), .Z(n9575) );
  XNOR2_X1 U9420 ( .A(n9578), .B(n9579), .ZN(n9355) );
  NAND2_X1 U9421 ( .A1(n9580), .A2(n9581), .ZN(n9578) );
  XNOR2_X1 U9422 ( .A(n9582), .B(n9583), .ZN(n9305) );
  XNOR2_X1 U9423 ( .A(n9584), .B(n9585), .ZN(n9582) );
  XOR2_X1 U9424 ( .A(n9586), .B(n9587), .Z(n9360) );
  XOR2_X1 U9425 ( .A(n9588), .B(n9589), .Z(n9586) );
  NOR2_X1 U9426 ( .A1(n8939), .A2(n8936), .ZN(n9589) );
  XNOR2_X1 U9427 ( .A(n9590), .B(n9591), .ZN(n9364) );
  XNOR2_X1 U9428 ( .A(n9592), .B(n9593), .ZN(n9591) );
  XOR2_X1 U9429 ( .A(n9594), .B(n9595), .Z(n9367) );
  XNOR2_X1 U9430 ( .A(n9596), .B(n9597), .ZN(n9594) );
  NAND2_X1 U9431 ( .A1(b_29_), .A2(a_22_), .ZN(n9596) );
  XNOR2_X1 U9432 ( .A(n9598), .B(n9599), .ZN(n9285) );
  XNOR2_X1 U9433 ( .A(n9600), .B(n9601), .ZN(n9599) );
  XOR2_X1 U9434 ( .A(n9602), .B(n9603), .Z(n9371) );
  XNOR2_X1 U9435 ( .A(n9604), .B(n9605), .ZN(n9602) );
  NAND2_X1 U9436 ( .A1(b_29_), .A2(a_20_), .ZN(n9604) );
  XNOR2_X1 U9437 ( .A(n9606), .B(n9607), .ZN(n9376) );
  XNOR2_X1 U9438 ( .A(n9608), .B(n9609), .ZN(n9607) );
  XOR2_X1 U9439 ( .A(n9610), .B(n9611), .Z(n9380) );
  XOR2_X1 U9440 ( .A(n9612), .B(n9613), .Z(n9610) );
  NOR2_X1 U9441 ( .A1(n8947), .A2(n8936), .ZN(n9613) );
  XOR2_X1 U9442 ( .A(n9614), .B(n9615), .Z(n9384) );
  XOR2_X1 U9443 ( .A(n9616), .B(n9617), .Z(n9614) );
  XOR2_X1 U9444 ( .A(n9618), .B(n9619), .Z(n9388) );
  XOR2_X1 U9445 ( .A(n9620), .B(n9621), .Z(n9618) );
  NOR2_X1 U9446 ( .A1(n8950), .A2(n8936), .ZN(n9621) );
  XOR2_X1 U9447 ( .A(n9622), .B(n9623), .Z(n9392) );
  XOR2_X1 U9448 ( .A(n9624), .B(n9625), .Z(n9622) );
  XOR2_X1 U9449 ( .A(n9626), .B(n9627), .Z(n9396) );
  XOR2_X1 U9450 ( .A(n9628), .B(n9629), .Z(n9626) );
  NOR2_X1 U9451 ( .A1(n8953), .A2(n8936), .ZN(n9629) );
  XOR2_X1 U9452 ( .A(n9630), .B(n9631), .Z(n9400) );
  XOR2_X1 U9453 ( .A(n9632), .B(n9633), .Z(n9630) );
  XNOR2_X1 U9454 ( .A(n9634), .B(n9635), .ZN(n9404) );
  XOR2_X1 U9455 ( .A(n9636), .B(n9637), .Z(n9635) );
  NAND2_X1 U9456 ( .A1(b_29_), .A2(a_12_), .ZN(n9637) );
  XNOR2_X1 U9457 ( .A(n9638), .B(n9639), .ZN(n9407) );
  XNOR2_X1 U9458 ( .A(n9640), .B(n9641), .ZN(n9638) );
  XOR2_X1 U9459 ( .A(n9642), .B(n9643), .Z(n9412) );
  XOR2_X1 U9460 ( .A(n9644), .B(n9645), .Z(n9642) );
  NOR2_X1 U9461 ( .A1(n8959), .A2(n8936), .ZN(n9645) );
  XOR2_X1 U9462 ( .A(n9646), .B(n9647), .Z(n9416) );
  XOR2_X1 U9463 ( .A(n9648), .B(n9649), .Z(n9646) );
  XNOR2_X1 U9464 ( .A(n9650), .B(n9651), .ZN(n9420) );
  XOR2_X1 U9465 ( .A(n9652), .B(n9653), .Z(n9650) );
  NOR2_X1 U9466 ( .A1(n8619), .A2(n8936), .ZN(n9653) );
  XOR2_X1 U9467 ( .A(n9654), .B(n9655), .Z(n9424) );
  XOR2_X1 U9468 ( .A(n9656), .B(n9657), .Z(n9654) );
  XNOR2_X1 U9469 ( .A(n9658), .B(n9659), .ZN(n9428) );
  XOR2_X1 U9470 ( .A(n9660), .B(n9661), .Z(n9659) );
  NAND2_X1 U9471 ( .A1(b_29_), .A2(a_6_), .ZN(n9661) );
  XOR2_X1 U9472 ( .A(n9662), .B(n9663), .Z(n9431) );
  XOR2_X1 U9473 ( .A(n9664), .B(n9665), .Z(n9662) );
  XOR2_X1 U9474 ( .A(n9666), .B(n9667), .Z(n9436) );
  XOR2_X1 U9475 ( .A(n9668), .B(n9669), .Z(n9666) );
  NOR2_X1 U9476 ( .A1(n8966), .A2(n8936), .ZN(n9669) );
  XOR2_X1 U9477 ( .A(n9670), .B(n9671), .Z(n9440) );
  XOR2_X1 U9478 ( .A(n9672), .B(n9673), .Z(n9670) );
  NOR2_X1 U9479 ( .A1(n8778), .A2(n8936), .ZN(n9673) );
  XNOR2_X1 U9480 ( .A(n9674), .B(n9675), .ZN(n9444) );
  XNOR2_X1 U9481 ( .A(n9676), .B(n9677), .ZN(n9674) );
  XOR2_X1 U9482 ( .A(n9678), .B(n9679), .Z(n9211) );
  XOR2_X1 U9483 ( .A(n9680), .B(n9681), .Z(n9678) );
  NOR2_X1 U9484 ( .A1(n8969), .A2(n8936), .ZN(n9681) );
  NAND2_X1 U9485 ( .A1(n9682), .A2(n9683), .ZN(n9001) );
  XOR2_X1 U9486 ( .A(n9203), .B(n9204), .Z(n9683) );
  AND2_X1 U9487 ( .A1(n9202), .A2(n9201), .ZN(n9682) );
  XOR2_X1 U9488 ( .A(n9684), .B(n9685), .Z(n9201) );
  XOR2_X1 U9489 ( .A(n9686), .B(n9687), .Z(n9684) );
  NAND2_X1 U9490 ( .A1(n9688), .A2(n9689), .ZN(n9202) );
  NAND2_X1 U9491 ( .A1(n9690), .A2(b_29_), .ZN(n9689) );
  NOR2_X1 U9492 ( .A1(n9691), .A2(n8974), .ZN(n9690) );
  NOR2_X1 U9493 ( .A1(n9450), .A2(n9451), .ZN(n9691) );
  NAND2_X1 U9494 ( .A1(n9450), .A2(n9451), .ZN(n9688) );
  NAND2_X1 U9495 ( .A1(n9692), .A2(n9693), .ZN(n9451) );
  NAND2_X1 U9496 ( .A1(n9694), .A2(b_29_), .ZN(n9693) );
  NOR2_X1 U9497 ( .A1(n9695), .A2(n8969), .ZN(n9694) );
  NOR2_X1 U9498 ( .A1(n9679), .A2(n9680), .ZN(n9695) );
  NAND2_X1 U9499 ( .A1(n9679), .A2(n9680), .ZN(n9692) );
  NAND2_X1 U9500 ( .A1(n9696), .A2(n9697), .ZN(n9680) );
  NAND2_X1 U9501 ( .A1(n9676), .A2(n9698), .ZN(n9697) );
  NAND2_X1 U9502 ( .A1(n9675), .A2(n9677), .ZN(n9698) );
  NAND2_X1 U9503 ( .A1(n9699), .A2(n9700), .ZN(n9676) );
  NAND2_X1 U9504 ( .A1(n9701), .A2(b_29_), .ZN(n9700) );
  NOR2_X1 U9505 ( .A1(n9702), .A2(n8778), .ZN(n9701) );
  NOR2_X1 U9506 ( .A1(n9671), .A2(n9672), .ZN(n9702) );
  NAND2_X1 U9507 ( .A1(n9671), .A2(n9672), .ZN(n9699) );
  NAND2_X1 U9508 ( .A1(n9703), .A2(n9704), .ZN(n9672) );
  NAND2_X1 U9509 ( .A1(n9705), .A2(b_29_), .ZN(n9704) );
  NOR2_X1 U9510 ( .A1(n9706), .A2(n8966), .ZN(n9705) );
  NOR2_X1 U9511 ( .A1(n9667), .A2(n9668), .ZN(n9706) );
  NAND2_X1 U9512 ( .A1(n9667), .A2(n9668), .ZN(n9703) );
  NAND2_X1 U9513 ( .A1(n9707), .A2(n9708), .ZN(n9668) );
  NAND2_X1 U9514 ( .A1(n9665), .A2(n9709), .ZN(n9708) );
  OR2_X1 U9515 ( .A1(n9664), .A2(n9663), .ZN(n9709) );
  NOR2_X1 U9516 ( .A1(n8936), .A2(n8723), .ZN(n9665) );
  NAND2_X1 U9517 ( .A1(n9663), .A2(n9664), .ZN(n9707) );
  NAND2_X1 U9518 ( .A1(n9710), .A2(n9711), .ZN(n9664) );
  NAND2_X1 U9519 ( .A1(n9712), .A2(b_29_), .ZN(n9711) );
  NOR2_X1 U9520 ( .A1(n9713), .A2(n8681), .ZN(n9712) );
  NOR2_X1 U9521 ( .A1(n9658), .A2(n9660), .ZN(n9713) );
  NAND2_X1 U9522 ( .A1(n9658), .A2(n9660), .ZN(n9710) );
  NAND2_X1 U9523 ( .A1(n9714), .A2(n9715), .ZN(n9660) );
  NAND2_X1 U9524 ( .A1(n9657), .A2(n9716), .ZN(n9715) );
  OR2_X1 U9525 ( .A1(n9656), .A2(n9655), .ZN(n9716) );
  NOR2_X1 U9526 ( .A1(n8936), .A2(n8962), .ZN(n9657) );
  NAND2_X1 U9527 ( .A1(n9655), .A2(n9656), .ZN(n9714) );
  NAND2_X1 U9528 ( .A1(n9717), .A2(n9718), .ZN(n9656) );
  NAND2_X1 U9529 ( .A1(n9719), .A2(b_29_), .ZN(n9718) );
  NOR2_X1 U9530 ( .A1(n9720), .A2(n8619), .ZN(n9719) );
  NOR2_X1 U9531 ( .A1(n9651), .A2(n9652), .ZN(n9720) );
  NAND2_X1 U9532 ( .A1(n9651), .A2(n9652), .ZN(n9717) );
  NAND2_X1 U9533 ( .A1(n9721), .A2(n9722), .ZN(n9652) );
  NAND2_X1 U9534 ( .A1(n9649), .A2(n9723), .ZN(n9722) );
  OR2_X1 U9535 ( .A1(n9648), .A2(n9647), .ZN(n9723) );
  NOR2_X1 U9536 ( .A1(n8936), .A2(n8605), .ZN(n9649) );
  NAND2_X1 U9537 ( .A1(n9647), .A2(n9648), .ZN(n9721) );
  NAND2_X1 U9538 ( .A1(n9724), .A2(n9725), .ZN(n9648) );
  NAND2_X1 U9539 ( .A1(n9726), .A2(b_29_), .ZN(n9725) );
  NOR2_X1 U9540 ( .A1(n9727), .A2(n8959), .ZN(n9726) );
  NOR2_X1 U9541 ( .A1(n9643), .A2(n9644), .ZN(n9727) );
  NAND2_X1 U9542 ( .A1(n9643), .A2(n9644), .ZN(n9724) );
  NAND2_X1 U9543 ( .A1(n9728), .A2(n9729), .ZN(n9644) );
  NAND2_X1 U9544 ( .A1(n9641), .A2(n9730), .ZN(n9729) );
  NAND2_X1 U9545 ( .A1(n9640), .A2(n9639), .ZN(n9730) );
  NOR2_X1 U9546 ( .A1(n8936), .A2(n8550), .ZN(n9641) );
  OR2_X1 U9547 ( .A1(n9639), .A2(n9640), .ZN(n9728) );
  AND2_X1 U9548 ( .A1(n9731), .A2(n9732), .ZN(n9640) );
  NAND2_X1 U9549 ( .A1(n9733), .A2(b_29_), .ZN(n9732) );
  NOR2_X1 U9550 ( .A1(n9734), .A2(n8956), .ZN(n9733) );
  NOR2_X1 U9551 ( .A1(n9634), .A2(n9636), .ZN(n9734) );
  NAND2_X1 U9552 ( .A1(n9634), .A2(n9636), .ZN(n9731) );
  NAND2_X1 U9553 ( .A1(n9735), .A2(n9736), .ZN(n9636) );
  NAND2_X1 U9554 ( .A1(n9633), .A2(n9737), .ZN(n9736) );
  OR2_X1 U9555 ( .A1(n9632), .A2(n9631), .ZN(n9737) );
  NOR2_X1 U9556 ( .A1(n8936), .A2(n8495), .ZN(n9633) );
  NAND2_X1 U9557 ( .A1(n9631), .A2(n9632), .ZN(n9735) );
  NAND2_X1 U9558 ( .A1(n9738), .A2(n9739), .ZN(n9632) );
  NAND2_X1 U9559 ( .A1(n9740), .A2(b_29_), .ZN(n9739) );
  NOR2_X1 U9560 ( .A1(n9741), .A2(n8953), .ZN(n9740) );
  NOR2_X1 U9561 ( .A1(n9627), .A2(n9628), .ZN(n9741) );
  NAND2_X1 U9562 ( .A1(n9627), .A2(n9628), .ZN(n9738) );
  NAND2_X1 U9563 ( .A1(n9742), .A2(n9743), .ZN(n9628) );
  NAND2_X1 U9564 ( .A1(n9625), .A2(n9744), .ZN(n9743) );
  OR2_X1 U9565 ( .A1(n9624), .A2(n9623), .ZN(n9744) );
  NOR2_X1 U9566 ( .A1(n8936), .A2(n8440), .ZN(n9625) );
  NAND2_X1 U9567 ( .A1(n9623), .A2(n9624), .ZN(n9742) );
  NAND2_X1 U9568 ( .A1(n9745), .A2(n9746), .ZN(n9624) );
  NAND2_X1 U9569 ( .A1(n9747), .A2(b_29_), .ZN(n9746) );
  NOR2_X1 U9570 ( .A1(n9748), .A2(n8950), .ZN(n9747) );
  NOR2_X1 U9571 ( .A1(n9619), .A2(n9620), .ZN(n9748) );
  NAND2_X1 U9572 ( .A1(n9619), .A2(n9620), .ZN(n9745) );
  NAND2_X1 U9573 ( .A1(n9749), .A2(n9750), .ZN(n9620) );
  NAND2_X1 U9574 ( .A1(n9617), .A2(n9751), .ZN(n9750) );
  OR2_X1 U9575 ( .A1(n9616), .A2(n9615), .ZN(n9751) );
  NOR2_X1 U9576 ( .A1(n8936), .A2(n8385), .ZN(n9617) );
  NAND2_X1 U9577 ( .A1(n9615), .A2(n9616), .ZN(n9749) );
  NAND2_X1 U9578 ( .A1(n9752), .A2(n9753), .ZN(n9616) );
  NAND2_X1 U9579 ( .A1(n9754), .A2(b_29_), .ZN(n9753) );
  NOR2_X1 U9580 ( .A1(n9755), .A2(n8947), .ZN(n9754) );
  NOR2_X1 U9581 ( .A1(n9611), .A2(n9612), .ZN(n9755) );
  NAND2_X1 U9582 ( .A1(n9611), .A2(n9612), .ZN(n9752) );
  NAND2_X1 U9583 ( .A1(n9756), .A2(n9757), .ZN(n9612) );
  NAND2_X1 U9584 ( .A1(n9609), .A2(n9758), .ZN(n9757) );
  OR2_X1 U9585 ( .A1(n9608), .A2(n9606), .ZN(n9758) );
  NOR2_X1 U9586 ( .A1(n8936), .A2(n8324), .ZN(n9609) );
  NAND2_X1 U9587 ( .A1(n9606), .A2(n9608), .ZN(n9756) );
  NAND2_X1 U9588 ( .A1(n9759), .A2(n9760), .ZN(n9608) );
  NAND2_X1 U9589 ( .A1(n9761), .A2(b_29_), .ZN(n9760) );
  NOR2_X1 U9590 ( .A1(n9762), .A2(n8944), .ZN(n9761) );
  NOR2_X1 U9591 ( .A1(n9603), .A2(n9605), .ZN(n9762) );
  NAND2_X1 U9592 ( .A1(n9603), .A2(n9605), .ZN(n9759) );
  NAND2_X1 U9593 ( .A1(n9763), .A2(n9764), .ZN(n9605) );
  NAND2_X1 U9594 ( .A1(n9601), .A2(n9765), .ZN(n9764) );
  OR2_X1 U9595 ( .A1(n9600), .A2(n9598), .ZN(n9765) );
  NOR2_X1 U9596 ( .A1(n8936), .A2(n8268), .ZN(n9601) );
  NAND2_X1 U9597 ( .A1(n9598), .A2(n9600), .ZN(n9763) );
  NAND2_X1 U9598 ( .A1(n9766), .A2(n9767), .ZN(n9600) );
  NAND2_X1 U9599 ( .A1(n9768), .A2(b_29_), .ZN(n9767) );
  NOR2_X1 U9600 ( .A1(n9769), .A2(n8941), .ZN(n9768) );
  NOR2_X1 U9601 ( .A1(n9595), .A2(n9597), .ZN(n9769) );
  NAND2_X1 U9602 ( .A1(n9595), .A2(n9597), .ZN(n9766) );
  NAND2_X1 U9603 ( .A1(n9770), .A2(n9771), .ZN(n9597) );
  NAND2_X1 U9604 ( .A1(n9593), .A2(n9772), .ZN(n9771) );
  OR2_X1 U9605 ( .A1(n9592), .A2(n9590), .ZN(n9772) );
  NOR2_X1 U9606 ( .A1(n8936), .A2(n8213), .ZN(n9593) );
  NAND2_X1 U9607 ( .A1(n9590), .A2(n9592), .ZN(n9770) );
  NAND2_X1 U9608 ( .A1(n9773), .A2(n9774), .ZN(n9592) );
  NAND2_X1 U9609 ( .A1(n9775), .A2(b_29_), .ZN(n9774) );
  NOR2_X1 U9610 ( .A1(n9776), .A2(n8939), .ZN(n9775) );
  NOR2_X1 U9611 ( .A1(n9587), .A2(n9588), .ZN(n9776) );
  NAND2_X1 U9612 ( .A1(n9587), .A2(n9588), .ZN(n9773) );
  NAND2_X1 U9613 ( .A1(n9777), .A2(n9778), .ZN(n9588) );
  NAND2_X1 U9614 ( .A1(n9585), .A2(n9779), .ZN(n9778) );
  NAND2_X1 U9615 ( .A1(n9584), .A2(n9583), .ZN(n9779) );
  NOR2_X1 U9616 ( .A1(n8936), .A2(n8158), .ZN(n9585) );
  OR2_X1 U9617 ( .A1(n9583), .A2(n9584), .ZN(n9777) );
  AND2_X1 U9618 ( .A1(n9580), .A2(n9780), .ZN(n9584) );
  NAND2_X1 U9619 ( .A1(n9579), .A2(n9581), .ZN(n9780) );
  NAND2_X1 U9620 ( .A1(n9781), .A2(n9782), .ZN(n9581) );
  NAND2_X1 U9621 ( .A1(b_29_), .A2(a_26_), .ZN(n9782) );
  INV_X1 U9622 ( .A(n9783), .ZN(n9781) );
  XNOR2_X1 U9623 ( .A(n9784), .B(n9785), .ZN(n9579) );
  NAND2_X1 U9624 ( .A1(n9786), .A2(n9787), .ZN(n9784) );
  NAND2_X1 U9625 ( .A1(a_26_), .A2(n9783), .ZN(n9580) );
  NAND2_X1 U9626 ( .A1(n9551), .A2(n9788), .ZN(n9783) );
  NAND2_X1 U9627 ( .A1(n9550), .A2(n9552), .ZN(n9788) );
  NAND2_X1 U9628 ( .A1(n9789), .A2(n9790), .ZN(n9552) );
  NAND2_X1 U9629 ( .A1(b_29_), .A2(a_27_), .ZN(n9790) );
  INV_X1 U9630 ( .A(n9791), .ZN(n9789) );
  XOR2_X1 U9631 ( .A(n9792), .B(n9793), .Z(n9550) );
  XOR2_X1 U9632 ( .A(n8926), .B(n9794), .Z(n9792) );
  NAND2_X1 U9633 ( .A1(a_27_), .A2(n9791), .ZN(n9551) );
  NAND2_X1 U9634 ( .A1(n9795), .A2(n9796), .ZN(n9791) );
  NAND2_X1 U9635 ( .A1(n9797), .A2(b_29_), .ZN(n9796) );
  NOR2_X1 U9636 ( .A1(n9798), .A2(n8055), .ZN(n9797) );
  NOR2_X1 U9637 ( .A1(n9558), .A2(n9560), .ZN(n9798) );
  NAND2_X1 U9638 ( .A1(n9558), .A2(n9560), .ZN(n9795) );
  NAND2_X1 U9639 ( .A1(n9799), .A2(n9800), .ZN(n9560) );
  NAND2_X1 U9640 ( .A1(n9801), .A2(n9802), .ZN(n9800) );
  OR2_X1 U9641 ( .A1(n9576), .A2(n9577), .ZN(n9802) );
  INV_X1 U9642 ( .A(n8929), .ZN(n9801) );
  NAND2_X1 U9643 ( .A1(b_29_), .A2(a_29_), .ZN(n8929) );
  NAND2_X1 U9644 ( .A1(n9577), .A2(n9576), .ZN(n9799) );
  NAND2_X1 U9645 ( .A1(n9803), .A2(n9804), .ZN(n9576) );
  NAND2_X1 U9646 ( .A1(b_27_), .A2(n9805), .ZN(n9804) );
  NAND2_X1 U9647 ( .A1(n8003), .A2(n9806), .ZN(n9805) );
  NAND2_X1 U9648 ( .A1(a_31_), .A2(n8069), .ZN(n9806) );
  NAND2_X1 U9649 ( .A1(b_28_), .A2(n9807), .ZN(n9803) );
  NAND2_X1 U9650 ( .A1(n9341), .A2(n9808), .ZN(n9807) );
  NAND2_X1 U9651 ( .A1(a_30_), .A2(n8102), .ZN(n9808) );
  AND2_X1 U9652 ( .A1(n9809), .A2(n7953), .ZN(n9577) );
  NOR2_X1 U9653 ( .A1(n8936), .A2(n8069), .ZN(n9809) );
  XOR2_X1 U9654 ( .A(n9810), .B(n9811), .Z(n9558) );
  XOR2_X1 U9655 ( .A(n9812), .B(n9813), .Z(n9810) );
  XOR2_X1 U9656 ( .A(n9814), .B(n9815), .Z(n9583) );
  NAND2_X1 U9657 ( .A1(n9816), .A2(n9817), .ZN(n9814) );
  XNOR2_X1 U9658 ( .A(n9818), .B(n9819), .ZN(n9587) );
  XNOR2_X1 U9659 ( .A(n9820), .B(n9821), .ZN(n9819) );
  XOR2_X1 U9660 ( .A(n9822), .B(n9823), .Z(n9590) );
  XOR2_X1 U9661 ( .A(n9824), .B(n9825), .Z(n9822) );
  NOR2_X1 U9662 ( .A1(n8939), .A2(n8069), .ZN(n9825) );
  XNOR2_X1 U9663 ( .A(n9826), .B(n9827), .ZN(n9595) );
  XNOR2_X1 U9664 ( .A(n9828), .B(n9829), .ZN(n9827) );
  XOR2_X1 U9665 ( .A(n9830), .B(n9831), .Z(n9598) );
  XOR2_X1 U9666 ( .A(n9832), .B(n9833), .Z(n9830) );
  NOR2_X1 U9667 ( .A1(n8941), .A2(n8069), .ZN(n9833) );
  XNOR2_X1 U9668 ( .A(n9834), .B(n9835), .ZN(n9603) );
  XNOR2_X1 U9669 ( .A(n9836), .B(n9837), .ZN(n9835) );
  XOR2_X1 U9670 ( .A(n9838), .B(n9839), .Z(n9606) );
  XOR2_X1 U9671 ( .A(n9840), .B(n9841), .Z(n9838) );
  NOR2_X1 U9672 ( .A1(n8944), .A2(n8069), .ZN(n9841) );
  XNOR2_X1 U9673 ( .A(n9842), .B(n9843), .ZN(n9611) );
  XNOR2_X1 U9674 ( .A(n9844), .B(n9845), .ZN(n9843) );
  XOR2_X1 U9675 ( .A(n9846), .B(n9847), .Z(n9615) );
  XOR2_X1 U9676 ( .A(n9848), .B(n9849), .Z(n9846) );
  NOR2_X1 U9677 ( .A1(n8947), .A2(n8069), .ZN(n9849) );
  XOR2_X1 U9678 ( .A(n9850), .B(n9851), .Z(n9619) );
  XOR2_X1 U9679 ( .A(n9852), .B(n9853), .Z(n9850) );
  XOR2_X1 U9680 ( .A(n9854), .B(n9855), .Z(n9623) );
  XOR2_X1 U9681 ( .A(n9856), .B(n9857), .Z(n9854) );
  NOR2_X1 U9682 ( .A1(n8950), .A2(n8069), .ZN(n9857) );
  XOR2_X1 U9683 ( .A(n9858), .B(n9859), .Z(n9627) );
  XOR2_X1 U9684 ( .A(n9860), .B(n9861), .Z(n9858) );
  XNOR2_X1 U9685 ( .A(n9862), .B(n9863), .ZN(n9631) );
  XOR2_X1 U9686 ( .A(n9864), .B(n9865), .Z(n9863) );
  NAND2_X1 U9687 ( .A1(b_28_), .A2(a_14_), .ZN(n9865) );
  XOR2_X1 U9688 ( .A(n9866), .B(n9867), .Z(n9634) );
  XOR2_X1 U9689 ( .A(n9868), .B(n9869), .Z(n9866) );
  XNOR2_X1 U9690 ( .A(n9870), .B(n9871), .ZN(n9639) );
  XOR2_X1 U9691 ( .A(n9872), .B(n9873), .Z(n9870) );
  NOR2_X1 U9692 ( .A1(n8956), .A2(n8069), .ZN(n9873) );
  XOR2_X1 U9693 ( .A(n9874), .B(n9875), .Z(n9643) );
  XOR2_X1 U9694 ( .A(n9876), .B(n9877), .Z(n9874) );
  XOR2_X1 U9695 ( .A(n9878), .B(n9879), .Z(n9647) );
  XOR2_X1 U9696 ( .A(n9880), .B(n9881), .Z(n9878) );
  NOR2_X1 U9697 ( .A1(n8959), .A2(n8069), .ZN(n9881) );
  XNOR2_X1 U9698 ( .A(n9882), .B(n9883), .ZN(n9651) );
  XNOR2_X1 U9699 ( .A(n9884), .B(n9885), .ZN(n9882) );
  XOR2_X1 U9700 ( .A(n9886), .B(n9887), .Z(n9655) );
  XOR2_X1 U9701 ( .A(n9888), .B(n9889), .Z(n9886) );
  NOR2_X1 U9702 ( .A1(n8619), .A2(n8069), .ZN(n9889) );
  XNOR2_X1 U9703 ( .A(n9890), .B(n9891), .ZN(n9658) );
  XNOR2_X1 U9704 ( .A(n9892), .B(n9893), .ZN(n9891) );
  XOR2_X1 U9705 ( .A(n9894), .B(n9895), .Z(n9663) );
  XOR2_X1 U9706 ( .A(n9896), .B(n9897), .Z(n9894) );
  NOR2_X1 U9707 ( .A1(n8681), .A2(n8069), .ZN(n9897) );
  XOR2_X1 U9708 ( .A(n9898), .B(n9899), .Z(n9667) );
  XOR2_X1 U9709 ( .A(n9900), .B(n9901), .Z(n9898) );
  XNOR2_X1 U9710 ( .A(n9902), .B(n9903), .ZN(n9671) );
  XOR2_X1 U9711 ( .A(n9904), .B(n9905), .Z(n9903) );
  NAND2_X1 U9712 ( .A1(b_28_), .A2(a_4_), .ZN(n9905) );
  OR2_X1 U9713 ( .A1(n9677), .A2(n9675), .ZN(n9696) );
  XNOR2_X1 U9714 ( .A(n9906), .B(n9907), .ZN(n9675) );
  XNOR2_X1 U9715 ( .A(n9908), .B(n9909), .ZN(n9906) );
  NAND2_X1 U9716 ( .A1(b_28_), .A2(a_3_), .ZN(n9908) );
  NAND2_X1 U9717 ( .A1(b_29_), .A2(a_2_), .ZN(n9677) );
  XOR2_X1 U9718 ( .A(n9910), .B(n9911), .Z(n9679) );
  XOR2_X1 U9719 ( .A(n9912), .B(n9913), .Z(n9910) );
  XOR2_X1 U9720 ( .A(n9914), .B(n9915), .Z(n9450) );
  XOR2_X1 U9721 ( .A(n9916), .B(n9917), .Z(n9914) );
  OR2_X1 U9722 ( .A1(n9197), .A2(n9196), .ZN(n9008) );
  NAND2_X1 U9723 ( .A1(n9918), .A2(n9919), .ZN(n9196) );
  NAND2_X1 U9724 ( .A1(n9920), .A2(n9921), .ZN(n9919) );
  NAND2_X1 U9725 ( .A1(n9204), .A2(n9203), .ZN(n9197) );
  NAND2_X1 U9726 ( .A1(n9922), .A2(n9923), .ZN(n9203) );
  NAND2_X1 U9727 ( .A1(n9687), .A2(n9924), .ZN(n9923) );
  OR2_X1 U9728 ( .A1(n9686), .A2(n9685), .ZN(n9924) );
  NOR2_X1 U9729 ( .A1(n8069), .A2(n8974), .ZN(n9687) );
  NAND2_X1 U9730 ( .A1(n9685), .A2(n9686), .ZN(n9922) );
  NAND2_X1 U9731 ( .A1(n9925), .A2(n9926), .ZN(n9686) );
  NAND2_X1 U9732 ( .A1(n9917), .A2(n9927), .ZN(n9926) );
  OR2_X1 U9733 ( .A1(n9916), .A2(n9915), .ZN(n9927) );
  NOR2_X1 U9734 ( .A1(n8069), .A2(n8969), .ZN(n9917) );
  NAND2_X1 U9735 ( .A1(n9915), .A2(n9916), .ZN(n9925) );
  NAND2_X1 U9736 ( .A1(n9928), .A2(n9929), .ZN(n9916) );
  NAND2_X1 U9737 ( .A1(n9912), .A2(n9930), .ZN(n9929) );
  OR2_X1 U9738 ( .A1(n9911), .A2(n9913), .ZN(n9930) );
  NAND2_X1 U9739 ( .A1(n9931), .A2(n9932), .ZN(n9912) );
  NAND2_X1 U9740 ( .A1(n9933), .A2(b_28_), .ZN(n9932) );
  NOR2_X1 U9741 ( .A1(n9934), .A2(n8778), .ZN(n9933) );
  NOR2_X1 U9742 ( .A1(n9907), .A2(n9909), .ZN(n9934) );
  NAND2_X1 U9743 ( .A1(n9907), .A2(n9909), .ZN(n9931) );
  NAND2_X1 U9744 ( .A1(n9935), .A2(n9936), .ZN(n9909) );
  NAND2_X1 U9745 ( .A1(n9937), .A2(b_28_), .ZN(n9936) );
  NOR2_X1 U9746 ( .A1(n9938), .A2(n8966), .ZN(n9937) );
  NOR2_X1 U9747 ( .A1(n9902), .A2(n9904), .ZN(n9938) );
  NAND2_X1 U9748 ( .A1(n9902), .A2(n9904), .ZN(n9935) );
  NAND2_X1 U9749 ( .A1(n9939), .A2(n9940), .ZN(n9904) );
  NAND2_X1 U9750 ( .A1(n9901), .A2(n9941), .ZN(n9940) );
  OR2_X1 U9751 ( .A1(n9900), .A2(n9899), .ZN(n9941) );
  NOR2_X1 U9752 ( .A1(n8069), .A2(n8723), .ZN(n9901) );
  NAND2_X1 U9753 ( .A1(n9899), .A2(n9900), .ZN(n9939) );
  NAND2_X1 U9754 ( .A1(n9942), .A2(n9943), .ZN(n9900) );
  NAND2_X1 U9755 ( .A1(n9944), .A2(b_28_), .ZN(n9943) );
  NOR2_X1 U9756 ( .A1(n9945), .A2(n8681), .ZN(n9944) );
  NOR2_X1 U9757 ( .A1(n9895), .A2(n9896), .ZN(n9945) );
  NAND2_X1 U9758 ( .A1(n9895), .A2(n9896), .ZN(n9942) );
  NAND2_X1 U9759 ( .A1(n9946), .A2(n9947), .ZN(n9896) );
  NAND2_X1 U9760 ( .A1(n9893), .A2(n9948), .ZN(n9947) );
  OR2_X1 U9761 ( .A1(n9892), .A2(n9890), .ZN(n9948) );
  NOR2_X1 U9762 ( .A1(n8069), .A2(n8962), .ZN(n9893) );
  NAND2_X1 U9763 ( .A1(n9890), .A2(n9892), .ZN(n9946) );
  NAND2_X1 U9764 ( .A1(n9949), .A2(n9950), .ZN(n9892) );
  NAND2_X1 U9765 ( .A1(n9951), .A2(b_28_), .ZN(n9950) );
  NOR2_X1 U9766 ( .A1(n9952), .A2(n8619), .ZN(n9951) );
  NOR2_X1 U9767 ( .A1(n9887), .A2(n9888), .ZN(n9952) );
  NAND2_X1 U9768 ( .A1(n9887), .A2(n9888), .ZN(n9949) );
  NAND2_X1 U9769 ( .A1(n9953), .A2(n9954), .ZN(n9888) );
  NAND2_X1 U9770 ( .A1(n9885), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U9771 ( .A1(n9884), .A2(n9883), .ZN(n9955) );
  NOR2_X1 U9772 ( .A1(n8069), .A2(n8605), .ZN(n9885) );
  OR2_X1 U9773 ( .A1(n9883), .A2(n9884), .ZN(n9953) );
  AND2_X1 U9774 ( .A1(n9956), .A2(n9957), .ZN(n9884) );
  NAND2_X1 U9775 ( .A1(n9958), .A2(b_28_), .ZN(n9957) );
  NOR2_X1 U9776 ( .A1(n9959), .A2(n8959), .ZN(n9958) );
  NOR2_X1 U9777 ( .A1(n9879), .A2(n9880), .ZN(n9959) );
  NAND2_X1 U9778 ( .A1(n9879), .A2(n9880), .ZN(n9956) );
  NAND2_X1 U9779 ( .A1(n9960), .A2(n9961), .ZN(n9880) );
  NAND2_X1 U9780 ( .A1(n9877), .A2(n9962), .ZN(n9961) );
  OR2_X1 U9781 ( .A1(n9876), .A2(n9875), .ZN(n9962) );
  NOR2_X1 U9782 ( .A1(n8069), .A2(n8550), .ZN(n9877) );
  NAND2_X1 U9783 ( .A1(n9875), .A2(n9876), .ZN(n9960) );
  NAND2_X1 U9784 ( .A1(n9963), .A2(n9964), .ZN(n9876) );
  NAND2_X1 U9785 ( .A1(n9965), .A2(b_28_), .ZN(n9964) );
  NOR2_X1 U9786 ( .A1(n9966), .A2(n8956), .ZN(n9965) );
  NOR2_X1 U9787 ( .A1(n9871), .A2(n9872), .ZN(n9966) );
  NAND2_X1 U9788 ( .A1(n9871), .A2(n9872), .ZN(n9963) );
  NAND2_X1 U9789 ( .A1(n9967), .A2(n9968), .ZN(n9872) );
  NAND2_X1 U9790 ( .A1(n9869), .A2(n9969), .ZN(n9968) );
  OR2_X1 U9791 ( .A1(n9868), .A2(n9867), .ZN(n9969) );
  NOR2_X1 U9792 ( .A1(n8069), .A2(n8495), .ZN(n9869) );
  NAND2_X1 U9793 ( .A1(n9867), .A2(n9868), .ZN(n9967) );
  NAND2_X1 U9794 ( .A1(n9970), .A2(n9971), .ZN(n9868) );
  NAND2_X1 U9795 ( .A1(n9972), .A2(b_28_), .ZN(n9971) );
  NOR2_X1 U9796 ( .A1(n9973), .A2(n8953), .ZN(n9972) );
  NOR2_X1 U9797 ( .A1(n9862), .A2(n9864), .ZN(n9973) );
  NAND2_X1 U9798 ( .A1(n9862), .A2(n9864), .ZN(n9970) );
  NAND2_X1 U9799 ( .A1(n9974), .A2(n9975), .ZN(n9864) );
  NAND2_X1 U9800 ( .A1(n9861), .A2(n9976), .ZN(n9975) );
  OR2_X1 U9801 ( .A1(n9860), .A2(n9859), .ZN(n9976) );
  NOR2_X1 U9802 ( .A1(n8069), .A2(n8440), .ZN(n9861) );
  NAND2_X1 U9803 ( .A1(n9859), .A2(n9860), .ZN(n9974) );
  NAND2_X1 U9804 ( .A1(n9977), .A2(n9978), .ZN(n9860) );
  NAND2_X1 U9805 ( .A1(n9979), .A2(b_28_), .ZN(n9978) );
  NOR2_X1 U9806 ( .A1(n9980), .A2(n8950), .ZN(n9979) );
  NOR2_X1 U9807 ( .A1(n9855), .A2(n9856), .ZN(n9980) );
  NAND2_X1 U9808 ( .A1(n9855), .A2(n9856), .ZN(n9977) );
  NAND2_X1 U9809 ( .A1(n9981), .A2(n9982), .ZN(n9856) );
  NAND2_X1 U9810 ( .A1(n9853), .A2(n9983), .ZN(n9982) );
  OR2_X1 U9811 ( .A1(n9852), .A2(n9851), .ZN(n9983) );
  NOR2_X1 U9812 ( .A1(n8069), .A2(n8385), .ZN(n9853) );
  NAND2_X1 U9813 ( .A1(n9851), .A2(n9852), .ZN(n9981) );
  NAND2_X1 U9814 ( .A1(n9984), .A2(n9985), .ZN(n9852) );
  NAND2_X1 U9815 ( .A1(n9986), .A2(b_28_), .ZN(n9985) );
  NOR2_X1 U9816 ( .A1(n9987), .A2(n8947), .ZN(n9986) );
  NOR2_X1 U9817 ( .A1(n9847), .A2(n9848), .ZN(n9987) );
  NAND2_X1 U9818 ( .A1(n9847), .A2(n9848), .ZN(n9984) );
  NAND2_X1 U9819 ( .A1(n9988), .A2(n9989), .ZN(n9848) );
  NAND2_X1 U9820 ( .A1(n9845), .A2(n9990), .ZN(n9989) );
  OR2_X1 U9821 ( .A1(n9844), .A2(n9842), .ZN(n9990) );
  NOR2_X1 U9822 ( .A1(n8069), .A2(n8324), .ZN(n9845) );
  NAND2_X1 U9823 ( .A1(n9842), .A2(n9844), .ZN(n9988) );
  NAND2_X1 U9824 ( .A1(n9991), .A2(n9992), .ZN(n9844) );
  NAND2_X1 U9825 ( .A1(n9993), .A2(b_28_), .ZN(n9992) );
  NOR2_X1 U9826 ( .A1(n9994), .A2(n8944), .ZN(n9993) );
  NOR2_X1 U9827 ( .A1(n9839), .A2(n9840), .ZN(n9994) );
  NAND2_X1 U9828 ( .A1(n9839), .A2(n9840), .ZN(n9991) );
  NAND2_X1 U9829 ( .A1(n9995), .A2(n9996), .ZN(n9840) );
  NAND2_X1 U9830 ( .A1(n9837), .A2(n9997), .ZN(n9996) );
  OR2_X1 U9831 ( .A1(n9836), .A2(n9834), .ZN(n9997) );
  NOR2_X1 U9832 ( .A1(n8069), .A2(n8268), .ZN(n9837) );
  NAND2_X1 U9833 ( .A1(n9834), .A2(n9836), .ZN(n9995) );
  NAND2_X1 U9834 ( .A1(n9998), .A2(n9999), .ZN(n9836) );
  NAND2_X1 U9835 ( .A1(n10000), .A2(b_28_), .ZN(n9999) );
  NOR2_X1 U9836 ( .A1(n10001), .A2(n8941), .ZN(n10000) );
  NOR2_X1 U9837 ( .A1(n9831), .A2(n9832), .ZN(n10001) );
  NAND2_X1 U9838 ( .A1(n9831), .A2(n9832), .ZN(n9998) );
  NAND2_X1 U9839 ( .A1(n10002), .A2(n10003), .ZN(n9832) );
  NAND2_X1 U9840 ( .A1(n9829), .A2(n10004), .ZN(n10003) );
  OR2_X1 U9841 ( .A1(n9828), .A2(n9826), .ZN(n10004) );
  NOR2_X1 U9842 ( .A1(n8069), .A2(n8213), .ZN(n9829) );
  NAND2_X1 U9843 ( .A1(n9826), .A2(n9828), .ZN(n10002) );
  NAND2_X1 U9844 ( .A1(n10005), .A2(n10006), .ZN(n9828) );
  NAND2_X1 U9845 ( .A1(n10007), .A2(b_28_), .ZN(n10006) );
  NOR2_X1 U9846 ( .A1(n10008), .A2(n8939), .ZN(n10007) );
  NOR2_X1 U9847 ( .A1(n9823), .A2(n9824), .ZN(n10008) );
  NAND2_X1 U9848 ( .A1(n9823), .A2(n9824), .ZN(n10005) );
  NAND2_X1 U9849 ( .A1(n10009), .A2(n10010), .ZN(n9824) );
  NAND2_X1 U9850 ( .A1(n9821), .A2(n10011), .ZN(n10010) );
  OR2_X1 U9851 ( .A1(n9820), .A2(n9818), .ZN(n10011) );
  NOR2_X1 U9852 ( .A1(n8069), .A2(n8158), .ZN(n9821) );
  NAND2_X1 U9853 ( .A1(n9818), .A2(n9820), .ZN(n10009) );
  NAND2_X1 U9854 ( .A1(n9816), .A2(n10012), .ZN(n9820) );
  NAND2_X1 U9855 ( .A1(n9815), .A2(n9817), .ZN(n10012) );
  NAND2_X1 U9856 ( .A1(n10013), .A2(n10014), .ZN(n9817) );
  NAND2_X1 U9857 ( .A1(b_28_), .A2(a_26_), .ZN(n10014) );
  INV_X1 U9858 ( .A(n10015), .ZN(n10013) );
  XNOR2_X1 U9859 ( .A(n10016), .B(n10017), .ZN(n9815) );
  XNOR2_X1 U9860 ( .A(n8923), .B(n10018), .ZN(n10017) );
  NAND2_X1 U9861 ( .A1(a_26_), .A2(n10015), .ZN(n9816) );
  NAND2_X1 U9862 ( .A1(n9786), .A2(n10019), .ZN(n10015) );
  NAND2_X1 U9863 ( .A1(n9785), .A2(n9787), .ZN(n10019) );
  NAND2_X1 U9864 ( .A1(n10020), .A2(n10021), .ZN(n9787) );
  NAND2_X1 U9865 ( .A1(b_28_), .A2(a_27_), .ZN(n10021) );
  INV_X1 U9866 ( .A(n10022), .ZN(n10020) );
  XOR2_X1 U9867 ( .A(n10023), .B(n10024), .Z(n9785) );
  XNOR2_X1 U9868 ( .A(n10025), .B(n10026), .ZN(n10023) );
  NAND2_X1 U9869 ( .A1(b_27_), .A2(a_28_), .ZN(n10025) );
  NAND2_X1 U9870 ( .A1(a_27_), .A2(n10022), .ZN(n9786) );
  NAND2_X1 U9871 ( .A1(n10027), .A2(n10028), .ZN(n10022) );
  NAND2_X1 U9872 ( .A1(n9793), .A2(n10029), .ZN(n10028) );
  NAND2_X1 U9873 ( .A1(n9794), .A2(n8926), .ZN(n10029) );
  INV_X1 U9874 ( .A(n10030), .ZN(n9794) );
  XOR2_X1 U9875 ( .A(n10031), .B(n10032), .Z(n9793) );
  XOR2_X1 U9876 ( .A(n10033), .B(n10034), .Z(n10031) );
  NAND2_X1 U9877 ( .A1(n10035), .A2(n10030), .ZN(n10027) );
  NAND2_X1 U9878 ( .A1(n10036), .A2(n10037), .ZN(n10030) );
  NAND2_X1 U9879 ( .A1(n9811), .A2(n10038), .ZN(n10037) );
  OR2_X1 U9880 ( .A1(n9812), .A2(n9813), .ZN(n10038) );
  NOR2_X1 U9881 ( .A1(n8069), .A2(n8041), .ZN(n9811) );
  NAND2_X1 U9882 ( .A1(n9813), .A2(n9812), .ZN(n10036) );
  NAND2_X1 U9883 ( .A1(n10039), .A2(n10040), .ZN(n9812) );
  NAND2_X1 U9884 ( .A1(b_26_), .A2(n10041), .ZN(n10040) );
  NAND2_X1 U9885 ( .A1(n8003), .A2(n10042), .ZN(n10041) );
  NAND2_X1 U9886 ( .A1(a_31_), .A2(n8102), .ZN(n10042) );
  NAND2_X1 U9887 ( .A1(b_27_), .A2(n10043), .ZN(n10039) );
  NAND2_X1 U9888 ( .A1(n9341), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U9889 ( .A1(a_30_), .A2(n8130), .ZN(n10044) );
  AND2_X1 U9890 ( .A1(n10045), .A2(n7953), .ZN(n9813) );
  NOR2_X1 U9891 ( .A1(n8069), .A2(n8102), .ZN(n10045) );
  INV_X1 U9892 ( .A(n8926), .ZN(n10035) );
  NAND2_X1 U9893 ( .A1(b_28_), .A2(a_28_), .ZN(n8926) );
  XNOR2_X1 U9894 ( .A(n10046), .B(n10047), .ZN(n9818) );
  NAND2_X1 U9895 ( .A1(n10048), .A2(n10049), .ZN(n10046) );
  XNOR2_X1 U9896 ( .A(n10050), .B(n10051), .ZN(n9823) );
  XNOR2_X1 U9897 ( .A(n10052), .B(n10053), .ZN(n10051) );
  XNOR2_X1 U9898 ( .A(n10054), .B(n10055), .ZN(n9826) );
  XOR2_X1 U9899 ( .A(n10056), .B(n10057), .Z(n10055) );
  NAND2_X1 U9900 ( .A1(b_27_), .A2(a_24_), .ZN(n10057) );
  XNOR2_X1 U9901 ( .A(n10058), .B(n10059), .ZN(n9831) );
  XNOR2_X1 U9902 ( .A(n10060), .B(n10061), .ZN(n10059) );
  XOR2_X1 U9903 ( .A(n10062), .B(n10063), .Z(n9834) );
  XOR2_X1 U9904 ( .A(n10064), .B(n10065), .Z(n10062) );
  NOR2_X1 U9905 ( .A1(n8941), .A2(n8102), .ZN(n10065) );
  XNOR2_X1 U9906 ( .A(n10066), .B(n10067), .ZN(n9839) );
  XNOR2_X1 U9907 ( .A(n10068), .B(n10069), .ZN(n10067) );
  XOR2_X1 U9908 ( .A(n10070), .B(n10071), .Z(n9842) );
  XOR2_X1 U9909 ( .A(n10072), .B(n10073), .Z(n10070) );
  NOR2_X1 U9910 ( .A1(n8944), .A2(n8102), .ZN(n10073) );
  XNOR2_X1 U9911 ( .A(n10074), .B(n10075), .ZN(n9847) );
  XNOR2_X1 U9912 ( .A(n10076), .B(n10077), .ZN(n10075) );
  XOR2_X1 U9913 ( .A(n10078), .B(n10079), .Z(n9851) );
  XOR2_X1 U9914 ( .A(n10080), .B(n10081), .Z(n10078) );
  NOR2_X1 U9915 ( .A1(n8947), .A2(n8102), .ZN(n10081) );
  XOR2_X1 U9916 ( .A(n10082), .B(n10083), .Z(n9855) );
  XOR2_X1 U9917 ( .A(n10084), .B(n10085), .Z(n10082) );
  XNOR2_X1 U9918 ( .A(n10086), .B(n10087), .ZN(n9859) );
  XOR2_X1 U9919 ( .A(n10088), .B(n10089), .Z(n10087) );
  NAND2_X1 U9920 ( .A1(b_27_), .A2(a_16_), .ZN(n10089) );
  XOR2_X1 U9921 ( .A(n10090), .B(n10091), .Z(n9862) );
  XOR2_X1 U9922 ( .A(n10092), .B(n10093), .Z(n10090) );
  XOR2_X1 U9923 ( .A(n10094), .B(n10095), .Z(n9867) );
  XOR2_X1 U9924 ( .A(n10096), .B(n10097), .Z(n10094) );
  NOR2_X1 U9925 ( .A1(n8953), .A2(n8102), .ZN(n10097) );
  XNOR2_X1 U9926 ( .A(n10098), .B(n10099), .ZN(n9871) );
  XNOR2_X1 U9927 ( .A(n10100), .B(n10101), .ZN(n10098) );
  XOR2_X1 U9928 ( .A(n10102), .B(n10103), .Z(n9875) );
  XOR2_X1 U9929 ( .A(n10104), .B(n10105), .Z(n10102) );
  NOR2_X1 U9930 ( .A1(n8956), .A2(n8102), .ZN(n10105) );
  XOR2_X1 U9931 ( .A(n10106), .B(n10107), .Z(n9879) );
  XOR2_X1 U9932 ( .A(n10108), .B(n10109), .Z(n10106) );
  XOR2_X1 U9933 ( .A(n10110), .B(n10111), .Z(n9883) );
  XOR2_X1 U9934 ( .A(n10112), .B(n10113), .Z(n10111) );
  NAND2_X1 U9935 ( .A1(b_27_), .A2(a_10_), .ZN(n10113) );
  XOR2_X1 U9936 ( .A(n10114), .B(n10115), .Z(n9887) );
  XOR2_X1 U9937 ( .A(n10116), .B(n10117), .Z(n10114) );
  XNOR2_X1 U9938 ( .A(n10118), .B(n10119), .ZN(n9890) );
  XOR2_X1 U9939 ( .A(n10120), .B(n10121), .Z(n10119) );
  NAND2_X1 U9940 ( .A1(b_27_), .A2(a_8_), .ZN(n10121) );
  XOR2_X1 U9941 ( .A(n10122), .B(n10123), .Z(n9895) );
  XOR2_X1 U9942 ( .A(n10124), .B(n10125), .Z(n10122) );
  NOR2_X1 U9943 ( .A1(n8962), .A2(n8102), .ZN(n10125) );
  XOR2_X1 U9944 ( .A(n10126), .B(n10127), .Z(n9899) );
  XOR2_X1 U9945 ( .A(n10128), .B(n10129), .Z(n10126) );
  NOR2_X1 U9946 ( .A1(n8681), .A2(n8102), .ZN(n10129) );
  XNOR2_X1 U9947 ( .A(n10130), .B(n10131), .ZN(n9902) );
  XNOR2_X1 U9948 ( .A(n10132), .B(n10133), .ZN(n10130) );
  XOR2_X1 U9949 ( .A(n10134), .B(n10135), .Z(n9907) );
  XOR2_X1 U9950 ( .A(n10136), .B(n10137), .Z(n10134) );
  NOR2_X1 U9951 ( .A1(n8966), .A2(n8102), .ZN(n10137) );
  NAND2_X1 U9952 ( .A1(n9913), .A2(n9911), .ZN(n9928) );
  XNOR2_X1 U9953 ( .A(n10138), .B(n10139), .ZN(n9911) );
  NAND2_X1 U9954 ( .A1(n10140), .A2(n10141), .ZN(n10138) );
  NOR2_X1 U9955 ( .A1(n8069), .A2(n8792), .ZN(n9913) );
  XNOR2_X1 U9956 ( .A(n10142), .B(n10143), .ZN(n9915) );
  NAND2_X1 U9957 ( .A1(n10144), .A2(n10145), .ZN(n10142) );
  XOR2_X1 U9958 ( .A(n10146), .B(n10147), .Z(n9685) );
  XOR2_X1 U9959 ( .A(n10148), .B(n10149), .Z(n10146) );
  NOR2_X1 U9960 ( .A1(n8969), .A2(n8102), .ZN(n10149) );
  XOR2_X1 U9961 ( .A(n10150), .B(n10151), .Z(n9204) );
  XNOR2_X1 U9962 ( .A(n10152), .B(n10153), .ZN(n10151) );
  NAND2_X1 U9963 ( .A1(n10154), .A2(n9918), .ZN(n9014) );
  INV_X1 U9964 ( .A(n9192), .ZN(n9918) );
  NOR2_X1 U9965 ( .A1(n9921), .A2(n9920), .ZN(n9192) );
  XOR2_X1 U9966 ( .A(n10155), .B(n10156), .Z(n9920) );
  XNOR2_X1 U9967 ( .A(n10157), .B(n10158), .ZN(n10155) );
  NAND2_X1 U9968 ( .A1(n10159), .A2(n10160), .ZN(n9921) );
  NAND2_X1 U9969 ( .A1(n10152), .A2(n10161), .ZN(n10160) );
  OR2_X1 U9970 ( .A1(n10153), .A2(n10150), .ZN(n10161) );
  AND2_X1 U9971 ( .A1(n10162), .A2(n10163), .ZN(n10152) );
  NAND2_X1 U9972 ( .A1(n10164), .A2(b_27_), .ZN(n10163) );
  NOR2_X1 U9973 ( .A1(n10165), .A2(n8969), .ZN(n10164) );
  NOR2_X1 U9974 ( .A1(n10147), .A2(n10148), .ZN(n10165) );
  NAND2_X1 U9975 ( .A1(n10147), .A2(n10148), .ZN(n10162) );
  NAND2_X1 U9976 ( .A1(n10144), .A2(n10166), .ZN(n10148) );
  NAND2_X1 U9977 ( .A1(n10143), .A2(n10145), .ZN(n10166) );
  NAND2_X1 U9978 ( .A1(n10167), .A2(n10168), .ZN(n10145) );
  NAND2_X1 U9979 ( .A1(b_27_), .A2(a_2_), .ZN(n10168) );
  INV_X1 U9980 ( .A(n10169), .ZN(n10167) );
  XNOR2_X1 U9981 ( .A(n10170), .B(n10171), .ZN(n10143) );
  XNOR2_X1 U9982 ( .A(n10172), .B(n10173), .ZN(n10170) );
  NAND2_X1 U9983 ( .A1(a_2_), .A2(n10169), .ZN(n10144) );
  NAND2_X1 U9984 ( .A1(n10140), .A2(n10174), .ZN(n10169) );
  NAND2_X1 U9985 ( .A1(n10139), .A2(n10141), .ZN(n10174) );
  NAND2_X1 U9986 ( .A1(n10175), .A2(n10176), .ZN(n10141) );
  NAND2_X1 U9987 ( .A1(b_27_), .A2(a_3_), .ZN(n10176) );
  INV_X1 U9988 ( .A(n10177), .ZN(n10175) );
  XNOR2_X1 U9989 ( .A(n10178), .B(n10179), .ZN(n10139) );
  XNOR2_X1 U9990 ( .A(n10180), .B(n10181), .ZN(n10178) );
  NAND2_X1 U9991 ( .A1(a_3_), .A2(n10177), .ZN(n10140) );
  NAND2_X1 U9992 ( .A1(n10182), .A2(n10183), .ZN(n10177) );
  NAND2_X1 U9993 ( .A1(n10184), .A2(b_27_), .ZN(n10183) );
  NOR2_X1 U9994 ( .A1(n10185), .A2(n8966), .ZN(n10184) );
  NOR2_X1 U9995 ( .A1(n10135), .A2(n10136), .ZN(n10185) );
  NAND2_X1 U9996 ( .A1(n10135), .A2(n10136), .ZN(n10182) );
  NAND2_X1 U9997 ( .A1(n10186), .A2(n10187), .ZN(n10136) );
  NAND2_X1 U9998 ( .A1(n10133), .A2(n10188), .ZN(n10187) );
  NAND2_X1 U9999 ( .A1(n10132), .A2(n10131), .ZN(n10188) );
  NOR2_X1 U10000 ( .A1(n8102), .A2(n8723), .ZN(n10133) );
  OR2_X1 U10001 ( .A1(n10131), .A2(n10132), .ZN(n10186) );
  AND2_X1 U10002 ( .A1(n10189), .A2(n10190), .ZN(n10132) );
  NAND2_X1 U10003 ( .A1(n10191), .A2(b_27_), .ZN(n10190) );
  NOR2_X1 U10004 ( .A1(n10192), .A2(n8681), .ZN(n10191) );
  NOR2_X1 U10005 ( .A1(n10127), .A2(n10128), .ZN(n10192) );
  NAND2_X1 U10006 ( .A1(n10127), .A2(n10128), .ZN(n10189) );
  NAND2_X1 U10007 ( .A1(n10193), .A2(n10194), .ZN(n10128) );
  NAND2_X1 U10008 ( .A1(n10195), .A2(b_27_), .ZN(n10194) );
  NOR2_X1 U10009 ( .A1(n10196), .A2(n8962), .ZN(n10195) );
  NOR2_X1 U10010 ( .A1(n10123), .A2(n10124), .ZN(n10196) );
  NAND2_X1 U10011 ( .A1(n10123), .A2(n10124), .ZN(n10193) );
  NAND2_X1 U10012 ( .A1(n10197), .A2(n10198), .ZN(n10124) );
  NAND2_X1 U10013 ( .A1(n10199), .A2(b_27_), .ZN(n10198) );
  NOR2_X1 U10014 ( .A1(n10200), .A2(n8619), .ZN(n10199) );
  NOR2_X1 U10015 ( .A1(n10118), .A2(n10120), .ZN(n10200) );
  NAND2_X1 U10016 ( .A1(n10118), .A2(n10120), .ZN(n10197) );
  NAND2_X1 U10017 ( .A1(n10201), .A2(n10202), .ZN(n10120) );
  NAND2_X1 U10018 ( .A1(n10116), .A2(n10203), .ZN(n10202) );
  OR2_X1 U10019 ( .A1(n10117), .A2(n10115), .ZN(n10203) );
  NOR2_X1 U10020 ( .A1(n8102), .A2(n8605), .ZN(n10116) );
  NAND2_X1 U10021 ( .A1(n10115), .A2(n10117), .ZN(n10201) );
  NAND2_X1 U10022 ( .A1(n10204), .A2(n10205), .ZN(n10117) );
  NAND2_X1 U10023 ( .A1(n10206), .A2(b_27_), .ZN(n10205) );
  NOR2_X1 U10024 ( .A1(n10207), .A2(n8959), .ZN(n10206) );
  NOR2_X1 U10025 ( .A1(n10110), .A2(n10112), .ZN(n10207) );
  NAND2_X1 U10026 ( .A1(n10110), .A2(n10112), .ZN(n10204) );
  NAND2_X1 U10027 ( .A1(n10208), .A2(n10209), .ZN(n10112) );
  NAND2_X1 U10028 ( .A1(n10109), .A2(n10210), .ZN(n10209) );
  OR2_X1 U10029 ( .A1(n10108), .A2(n10107), .ZN(n10210) );
  NOR2_X1 U10030 ( .A1(n8102), .A2(n8550), .ZN(n10109) );
  NAND2_X1 U10031 ( .A1(n10107), .A2(n10108), .ZN(n10208) );
  NAND2_X1 U10032 ( .A1(n10211), .A2(n10212), .ZN(n10108) );
  NAND2_X1 U10033 ( .A1(n10213), .A2(b_27_), .ZN(n10212) );
  NOR2_X1 U10034 ( .A1(n10214), .A2(n8956), .ZN(n10213) );
  NOR2_X1 U10035 ( .A1(n10103), .A2(n10104), .ZN(n10214) );
  NAND2_X1 U10036 ( .A1(n10103), .A2(n10104), .ZN(n10211) );
  NAND2_X1 U10037 ( .A1(n10215), .A2(n10216), .ZN(n10104) );
  NAND2_X1 U10038 ( .A1(n10101), .A2(n10217), .ZN(n10216) );
  NAND2_X1 U10039 ( .A1(n10100), .A2(n10099), .ZN(n10217) );
  NOR2_X1 U10040 ( .A1(n8102), .A2(n8495), .ZN(n10101) );
  OR2_X1 U10041 ( .A1(n10099), .A2(n10100), .ZN(n10215) );
  AND2_X1 U10042 ( .A1(n10218), .A2(n10219), .ZN(n10100) );
  NAND2_X1 U10043 ( .A1(n10220), .A2(b_27_), .ZN(n10219) );
  NOR2_X1 U10044 ( .A1(n10221), .A2(n8953), .ZN(n10220) );
  NOR2_X1 U10045 ( .A1(n10095), .A2(n10096), .ZN(n10221) );
  NAND2_X1 U10046 ( .A1(n10095), .A2(n10096), .ZN(n10218) );
  NAND2_X1 U10047 ( .A1(n10222), .A2(n10223), .ZN(n10096) );
  NAND2_X1 U10048 ( .A1(n10093), .A2(n10224), .ZN(n10223) );
  OR2_X1 U10049 ( .A1(n10092), .A2(n10091), .ZN(n10224) );
  NOR2_X1 U10050 ( .A1(n8102), .A2(n8440), .ZN(n10093) );
  NAND2_X1 U10051 ( .A1(n10091), .A2(n10092), .ZN(n10222) );
  NAND2_X1 U10052 ( .A1(n10225), .A2(n10226), .ZN(n10092) );
  NAND2_X1 U10053 ( .A1(n10227), .A2(b_27_), .ZN(n10226) );
  NOR2_X1 U10054 ( .A1(n10228), .A2(n8950), .ZN(n10227) );
  NOR2_X1 U10055 ( .A1(n10086), .A2(n10088), .ZN(n10228) );
  NAND2_X1 U10056 ( .A1(n10086), .A2(n10088), .ZN(n10225) );
  NAND2_X1 U10057 ( .A1(n10229), .A2(n10230), .ZN(n10088) );
  NAND2_X1 U10058 ( .A1(n10085), .A2(n10231), .ZN(n10230) );
  OR2_X1 U10059 ( .A1(n10084), .A2(n10083), .ZN(n10231) );
  NOR2_X1 U10060 ( .A1(n8102), .A2(n8385), .ZN(n10085) );
  NAND2_X1 U10061 ( .A1(n10083), .A2(n10084), .ZN(n10229) );
  NAND2_X1 U10062 ( .A1(n10232), .A2(n10233), .ZN(n10084) );
  NAND2_X1 U10063 ( .A1(n10234), .A2(b_27_), .ZN(n10233) );
  NOR2_X1 U10064 ( .A1(n10235), .A2(n8947), .ZN(n10234) );
  NOR2_X1 U10065 ( .A1(n10079), .A2(n10080), .ZN(n10235) );
  NAND2_X1 U10066 ( .A1(n10079), .A2(n10080), .ZN(n10232) );
  NAND2_X1 U10067 ( .A1(n10236), .A2(n10237), .ZN(n10080) );
  NAND2_X1 U10068 ( .A1(n10077), .A2(n10238), .ZN(n10237) );
  OR2_X1 U10069 ( .A1(n10076), .A2(n10074), .ZN(n10238) );
  NOR2_X1 U10070 ( .A1(n8102), .A2(n8324), .ZN(n10077) );
  NAND2_X1 U10071 ( .A1(n10074), .A2(n10076), .ZN(n10236) );
  NAND2_X1 U10072 ( .A1(n10239), .A2(n10240), .ZN(n10076) );
  NAND2_X1 U10073 ( .A1(n10241), .A2(b_27_), .ZN(n10240) );
  NOR2_X1 U10074 ( .A1(n10242), .A2(n8944), .ZN(n10241) );
  NOR2_X1 U10075 ( .A1(n10071), .A2(n10072), .ZN(n10242) );
  NAND2_X1 U10076 ( .A1(n10071), .A2(n10072), .ZN(n10239) );
  NAND2_X1 U10077 ( .A1(n10243), .A2(n10244), .ZN(n10072) );
  NAND2_X1 U10078 ( .A1(n10069), .A2(n10245), .ZN(n10244) );
  OR2_X1 U10079 ( .A1(n10068), .A2(n10066), .ZN(n10245) );
  NOR2_X1 U10080 ( .A1(n8102), .A2(n8268), .ZN(n10069) );
  NAND2_X1 U10081 ( .A1(n10066), .A2(n10068), .ZN(n10243) );
  NAND2_X1 U10082 ( .A1(n10246), .A2(n10247), .ZN(n10068) );
  NAND2_X1 U10083 ( .A1(n10248), .A2(b_27_), .ZN(n10247) );
  NOR2_X1 U10084 ( .A1(n10249), .A2(n8941), .ZN(n10248) );
  NOR2_X1 U10085 ( .A1(n10063), .A2(n10064), .ZN(n10249) );
  NAND2_X1 U10086 ( .A1(n10063), .A2(n10064), .ZN(n10246) );
  NAND2_X1 U10087 ( .A1(n10250), .A2(n10251), .ZN(n10064) );
  NAND2_X1 U10088 ( .A1(n10061), .A2(n10252), .ZN(n10251) );
  OR2_X1 U10089 ( .A1(n10060), .A2(n10058), .ZN(n10252) );
  NOR2_X1 U10090 ( .A1(n8102), .A2(n8213), .ZN(n10061) );
  NAND2_X1 U10091 ( .A1(n10058), .A2(n10060), .ZN(n10250) );
  NAND2_X1 U10092 ( .A1(n10253), .A2(n10254), .ZN(n10060) );
  NAND2_X1 U10093 ( .A1(n10255), .A2(b_27_), .ZN(n10254) );
  NOR2_X1 U10094 ( .A1(n10256), .A2(n8939), .ZN(n10255) );
  NOR2_X1 U10095 ( .A1(n10054), .A2(n10056), .ZN(n10256) );
  NAND2_X1 U10096 ( .A1(n10054), .A2(n10056), .ZN(n10253) );
  NAND2_X1 U10097 ( .A1(n10257), .A2(n10258), .ZN(n10056) );
  NAND2_X1 U10098 ( .A1(n10053), .A2(n10259), .ZN(n10258) );
  OR2_X1 U10099 ( .A1(n10052), .A2(n10050), .ZN(n10259) );
  NOR2_X1 U10100 ( .A1(n8102), .A2(n8158), .ZN(n10053) );
  NAND2_X1 U10101 ( .A1(n10050), .A2(n10052), .ZN(n10257) );
  NAND2_X1 U10102 ( .A1(n10048), .A2(n10260), .ZN(n10052) );
  NAND2_X1 U10103 ( .A1(n10047), .A2(n10049), .ZN(n10260) );
  NAND2_X1 U10104 ( .A1(n10261), .A2(n10262), .ZN(n10049) );
  NAND2_X1 U10105 ( .A1(b_27_), .A2(a_26_), .ZN(n10262) );
  INV_X1 U10106 ( .A(n10263), .ZN(n10261) );
  XNOR2_X1 U10107 ( .A(n10264), .B(n10265), .ZN(n10047) );
  NAND2_X1 U10108 ( .A1(n10266), .A2(n10267), .ZN(n10264) );
  NAND2_X1 U10109 ( .A1(a_26_), .A2(n10263), .ZN(n10048) );
  NAND2_X1 U10110 ( .A1(n10268), .A2(n10269), .ZN(n10263) );
  NAND2_X1 U10111 ( .A1(n10016), .A2(n10270), .ZN(n10269) );
  OR2_X1 U10112 ( .A1(n10018), .A2(n8923), .ZN(n10270) );
  XOR2_X1 U10113 ( .A(n10271), .B(n10272), .Z(n10016) );
  XNOR2_X1 U10114 ( .A(n10273), .B(n10274), .ZN(n10271) );
  NAND2_X1 U10115 ( .A1(b_26_), .A2(a_28_), .ZN(n10273) );
  NAND2_X1 U10116 ( .A1(n8923), .A2(n10018), .ZN(n10268) );
  NAND2_X1 U10117 ( .A1(n10275), .A2(n10276), .ZN(n10018) );
  NAND2_X1 U10118 ( .A1(n10277), .A2(b_27_), .ZN(n10276) );
  NOR2_X1 U10119 ( .A1(n10278), .A2(n8055), .ZN(n10277) );
  NOR2_X1 U10120 ( .A1(n10024), .A2(n10026), .ZN(n10278) );
  NAND2_X1 U10121 ( .A1(n10024), .A2(n10026), .ZN(n10275) );
  NAND2_X1 U10122 ( .A1(n10279), .A2(n10280), .ZN(n10026) );
  NAND2_X1 U10123 ( .A1(n10032), .A2(n10281), .ZN(n10280) );
  OR2_X1 U10124 ( .A1(n10033), .A2(n10034), .ZN(n10281) );
  NOR2_X1 U10125 ( .A1(n8102), .A2(n8041), .ZN(n10032) );
  NAND2_X1 U10126 ( .A1(n10034), .A2(n10033), .ZN(n10279) );
  NAND2_X1 U10127 ( .A1(n10282), .A2(n10283), .ZN(n10033) );
  NAND2_X1 U10128 ( .A1(b_25_), .A2(n10284), .ZN(n10283) );
  NAND2_X1 U10129 ( .A1(n8003), .A2(n10285), .ZN(n10284) );
  NAND2_X1 U10130 ( .A1(a_31_), .A2(n8130), .ZN(n10285) );
  NAND2_X1 U10131 ( .A1(b_26_), .A2(n10286), .ZN(n10282) );
  NAND2_X1 U10132 ( .A1(n9341), .A2(n10287), .ZN(n10286) );
  NAND2_X1 U10133 ( .A1(a_30_), .A2(n8938), .ZN(n10287) );
  AND2_X1 U10134 ( .A1(n10288), .A2(n7953), .ZN(n10034) );
  NOR2_X1 U10135 ( .A1(n8102), .A2(n8130), .ZN(n10288) );
  XOR2_X1 U10136 ( .A(n10289), .B(n10290), .Z(n10024) );
  XOR2_X1 U10137 ( .A(n10291), .B(n10292), .Z(n10289) );
  NOR2_X1 U10138 ( .A1(n8102), .A2(n8937), .ZN(n8923) );
  XOR2_X1 U10139 ( .A(n10293), .B(n10294), .Z(n10050) );
  XOR2_X1 U10140 ( .A(n10295), .B(n10296), .Z(n10293) );
  XNOR2_X1 U10141 ( .A(n10297), .B(n10298), .ZN(n10054) );
  XNOR2_X1 U10142 ( .A(n10299), .B(n10300), .ZN(n10298) );
  XOR2_X1 U10143 ( .A(n10301), .B(n10302), .Z(n10058) );
  XOR2_X1 U10144 ( .A(n10303), .B(n10304), .Z(n10301) );
  NOR2_X1 U10145 ( .A1(n8939), .A2(n8130), .ZN(n10304) );
  XNOR2_X1 U10146 ( .A(n10305), .B(n10306), .ZN(n10063) );
  XNOR2_X1 U10147 ( .A(n10307), .B(n10308), .ZN(n10306) );
  XOR2_X1 U10148 ( .A(n10309), .B(n10310), .Z(n10066) );
  XOR2_X1 U10149 ( .A(n10311), .B(n10312), .Z(n10309) );
  NOR2_X1 U10150 ( .A1(n8941), .A2(n8130), .ZN(n10312) );
  XNOR2_X1 U10151 ( .A(n10313), .B(n10314), .ZN(n10071) );
  XNOR2_X1 U10152 ( .A(n10315), .B(n10316), .ZN(n10314) );
  XOR2_X1 U10153 ( .A(n10317), .B(n10318), .Z(n10074) );
  XOR2_X1 U10154 ( .A(n10319), .B(n10320), .Z(n10317) );
  NOR2_X1 U10155 ( .A1(n8944), .A2(n8130), .ZN(n10320) );
  XOR2_X1 U10156 ( .A(n10321), .B(n10322), .Z(n10079) );
  XOR2_X1 U10157 ( .A(n10323), .B(n10324), .Z(n10321) );
  XOR2_X1 U10158 ( .A(n10325), .B(n10326), .Z(n10083) );
  XOR2_X1 U10159 ( .A(n10327), .B(n10328), .Z(n10325) );
  NOR2_X1 U10160 ( .A1(n8947), .A2(n8130), .ZN(n10328) );
  XOR2_X1 U10161 ( .A(n10329), .B(n10330), .Z(n10086) );
  XOR2_X1 U10162 ( .A(n10331), .B(n10332), .Z(n10329) );
  XOR2_X1 U10163 ( .A(n10333), .B(n10334), .Z(n10091) );
  XOR2_X1 U10164 ( .A(n10335), .B(n10336), .Z(n10333) );
  NOR2_X1 U10165 ( .A1(n8950), .A2(n8130), .ZN(n10336) );
  XOR2_X1 U10166 ( .A(n10337), .B(n10338), .Z(n10095) );
  XOR2_X1 U10167 ( .A(n10339), .B(n10340), .Z(n10337) );
  XNOR2_X1 U10168 ( .A(n10341), .B(n10342), .ZN(n10099) );
  XOR2_X1 U10169 ( .A(n10343), .B(n10344), .Z(n10341) );
  NOR2_X1 U10170 ( .A1(n8953), .A2(n8130), .ZN(n10344) );
  XOR2_X1 U10171 ( .A(n10345), .B(n10346), .Z(n10103) );
  XOR2_X1 U10172 ( .A(n10347), .B(n10348), .Z(n10345) );
  XNOR2_X1 U10173 ( .A(n10349), .B(n10350), .ZN(n10107) );
  XOR2_X1 U10174 ( .A(n10351), .B(n10352), .Z(n10350) );
  NAND2_X1 U10175 ( .A1(b_26_), .A2(a_12_), .ZN(n10352) );
  XNOR2_X1 U10176 ( .A(n10353), .B(n10354), .ZN(n10110) );
  XNOR2_X1 U10177 ( .A(n10355), .B(n10356), .ZN(n10353) );
  XNOR2_X1 U10178 ( .A(n10357), .B(n10358), .ZN(n10115) );
  XOR2_X1 U10179 ( .A(n10359), .B(n10360), .Z(n10358) );
  NAND2_X1 U10180 ( .A1(b_26_), .A2(a_10_), .ZN(n10360) );
  XOR2_X1 U10181 ( .A(n10361), .B(n10362), .Z(n10118) );
  XOR2_X1 U10182 ( .A(n10363), .B(n10364), .Z(n10361) );
  XOR2_X1 U10183 ( .A(n10365), .B(n10366), .Z(n10123) );
  XOR2_X1 U10184 ( .A(n10367), .B(n10368), .Z(n10365) );
  NOR2_X1 U10185 ( .A1(n8619), .A2(n8130), .ZN(n10368) );
  XNOR2_X1 U10186 ( .A(n10369), .B(n10370), .ZN(n10127) );
  NAND2_X1 U10187 ( .A1(n10371), .A2(n10372), .ZN(n10369) );
  XNOR2_X1 U10188 ( .A(n10373), .B(n10374), .ZN(n10131) );
  XOR2_X1 U10189 ( .A(n10375), .B(n10376), .Z(n10373) );
  NOR2_X1 U10190 ( .A1(n8681), .A2(n8130), .ZN(n10376) );
  XOR2_X1 U10191 ( .A(n10377), .B(n10378), .Z(n10135) );
  XOR2_X1 U10192 ( .A(n10379), .B(n10380), .Z(n10377) );
  NOR2_X1 U10193 ( .A1(n8723), .A2(n8130), .ZN(n10380) );
  XNOR2_X1 U10194 ( .A(n10381), .B(n10382), .ZN(n10147) );
  NAND2_X1 U10195 ( .A1(n10383), .A2(n10384), .ZN(n10381) );
  NAND2_X1 U10196 ( .A1(n10150), .A2(n10153), .ZN(n10159) );
  NAND2_X1 U10197 ( .A1(b_27_), .A2(a_0_), .ZN(n10153) );
  XNOR2_X1 U10198 ( .A(n10385), .B(n10386), .ZN(n10150) );
  XOR2_X1 U10199 ( .A(n10387), .B(n10388), .Z(n10385) );
  NOR2_X1 U10200 ( .A1(n8969), .A2(n8130), .ZN(n10388) );
  NAND2_X1 U10201 ( .A1(n10389), .A2(n10390), .ZN(n10154) );
  NAND2_X1 U10202 ( .A1(n9194), .A2(n9193), .ZN(n10390) );
  NAND2_X1 U10203 ( .A1(n10389), .A2(n10391), .ZN(n9020) );
  NAND2_X1 U10204 ( .A1(n10392), .A2(n9188), .ZN(n10391) );
  INV_X1 U10205 ( .A(n10393), .ZN(n10389) );
  NAND2_X1 U10206 ( .A1(n10394), .A2(n10393), .ZN(n9019) );
  NOR2_X1 U10207 ( .A1(n9193), .A2(n9194), .ZN(n10393) );
  AND2_X1 U10208 ( .A1(n10395), .A2(n10396), .ZN(n9194) );
  NAND2_X1 U10209 ( .A1(n10158), .A2(n10397), .ZN(n10396) );
  NAND2_X1 U10210 ( .A1(n10157), .A2(n10156), .ZN(n10397) );
  NOR2_X1 U10211 ( .A1(n8130), .A2(n8974), .ZN(n10158) );
  OR2_X1 U10212 ( .A1(n10156), .A2(n10157), .ZN(n10395) );
  AND2_X1 U10213 ( .A1(n10398), .A2(n10399), .ZN(n10157) );
  NAND2_X1 U10214 ( .A1(n10400), .A2(b_26_), .ZN(n10399) );
  NOR2_X1 U10215 ( .A1(n10401), .A2(n8969), .ZN(n10400) );
  NOR2_X1 U10216 ( .A1(n10387), .A2(n10386), .ZN(n10401) );
  NAND2_X1 U10217 ( .A1(n10386), .A2(n10387), .ZN(n10398) );
  NAND2_X1 U10218 ( .A1(n10383), .A2(n10402), .ZN(n10387) );
  NAND2_X1 U10219 ( .A1(n10382), .A2(n10384), .ZN(n10402) );
  NAND2_X1 U10220 ( .A1(n10403), .A2(n10404), .ZN(n10384) );
  NAND2_X1 U10221 ( .A1(b_26_), .A2(a_2_), .ZN(n10404) );
  INV_X1 U10222 ( .A(n10405), .ZN(n10403) );
  XOR2_X1 U10223 ( .A(n10406), .B(n10407), .Z(n10382) );
  XOR2_X1 U10224 ( .A(n10408), .B(n10409), .Z(n10406) );
  NOR2_X1 U10225 ( .A1(n8778), .A2(n8938), .ZN(n10409) );
  NAND2_X1 U10226 ( .A1(a_2_), .A2(n10405), .ZN(n10383) );
  NAND2_X1 U10227 ( .A1(n10410), .A2(n10411), .ZN(n10405) );
  NAND2_X1 U10228 ( .A1(n10173), .A2(n10412), .ZN(n10411) );
  NAND2_X1 U10229 ( .A1(n10172), .A2(n10171), .ZN(n10412) );
  NOR2_X1 U10230 ( .A1(n8130), .A2(n8778), .ZN(n10173) );
  OR2_X1 U10231 ( .A1(n10171), .A2(n10172), .ZN(n10410) );
  AND2_X1 U10232 ( .A1(n10413), .A2(n10414), .ZN(n10172) );
  NAND2_X1 U10233 ( .A1(n10181), .A2(n10415), .ZN(n10414) );
  NAND2_X1 U10234 ( .A1(n10180), .A2(n10179), .ZN(n10415) );
  NOR2_X1 U10235 ( .A1(n8130), .A2(n8966), .ZN(n10181) );
  OR2_X1 U10236 ( .A1(n10179), .A2(n10180), .ZN(n10413) );
  AND2_X1 U10237 ( .A1(n10416), .A2(n10417), .ZN(n10180) );
  NAND2_X1 U10238 ( .A1(n10418), .A2(b_26_), .ZN(n10417) );
  NOR2_X1 U10239 ( .A1(n10419), .A2(n8723), .ZN(n10418) );
  NOR2_X1 U10240 ( .A1(n10379), .A2(n10378), .ZN(n10419) );
  NAND2_X1 U10241 ( .A1(n10378), .A2(n10379), .ZN(n10416) );
  NAND2_X1 U10242 ( .A1(n10420), .A2(n10421), .ZN(n10379) );
  NAND2_X1 U10243 ( .A1(n10422), .A2(b_26_), .ZN(n10421) );
  NOR2_X1 U10244 ( .A1(n10423), .A2(n8681), .ZN(n10422) );
  NOR2_X1 U10245 ( .A1(n10375), .A2(n10374), .ZN(n10423) );
  NAND2_X1 U10246 ( .A1(n10374), .A2(n10375), .ZN(n10420) );
  NAND2_X1 U10247 ( .A1(n10371), .A2(n10424), .ZN(n10375) );
  NAND2_X1 U10248 ( .A1(n10370), .A2(n10372), .ZN(n10424) );
  NAND2_X1 U10249 ( .A1(n10425), .A2(n10426), .ZN(n10372) );
  NAND2_X1 U10250 ( .A1(b_26_), .A2(a_7_), .ZN(n10426) );
  INV_X1 U10251 ( .A(n10427), .ZN(n10425) );
  XOR2_X1 U10252 ( .A(n10428), .B(n10429), .Z(n10370) );
  XOR2_X1 U10253 ( .A(n10430), .B(n10431), .Z(n10428) );
  NOR2_X1 U10254 ( .A1(n8619), .A2(n8938), .ZN(n10431) );
  NAND2_X1 U10255 ( .A1(a_7_), .A2(n10427), .ZN(n10371) );
  NAND2_X1 U10256 ( .A1(n10432), .A2(n10433), .ZN(n10427) );
  NAND2_X1 U10257 ( .A1(n10434), .A2(b_26_), .ZN(n10433) );
  NOR2_X1 U10258 ( .A1(n10435), .A2(n8619), .ZN(n10434) );
  NOR2_X1 U10259 ( .A1(n10366), .A2(n10367), .ZN(n10435) );
  NAND2_X1 U10260 ( .A1(n10366), .A2(n10367), .ZN(n10432) );
  NAND2_X1 U10261 ( .A1(n10436), .A2(n10437), .ZN(n10367) );
  NAND2_X1 U10262 ( .A1(n10364), .A2(n10438), .ZN(n10437) );
  OR2_X1 U10263 ( .A1(n10362), .A2(n10363), .ZN(n10438) );
  NOR2_X1 U10264 ( .A1(n8130), .A2(n8605), .ZN(n10364) );
  NAND2_X1 U10265 ( .A1(n10362), .A2(n10363), .ZN(n10436) );
  NAND2_X1 U10266 ( .A1(n10439), .A2(n10440), .ZN(n10363) );
  NAND2_X1 U10267 ( .A1(n10441), .A2(b_26_), .ZN(n10440) );
  NOR2_X1 U10268 ( .A1(n10442), .A2(n8959), .ZN(n10441) );
  NOR2_X1 U10269 ( .A1(n10357), .A2(n10359), .ZN(n10442) );
  NAND2_X1 U10270 ( .A1(n10357), .A2(n10359), .ZN(n10439) );
  NAND2_X1 U10271 ( .A1(n10443), .A2(n10444), .ZN(n10359) );
  NAND2_X1 U10272 ( .A1(n10356), .A2(n10445), .ZN(n10444) );
  NAND2_X1 U10273 ( .A1(n10355), .A2(n10354), .ZN(n10445) );
  NOR2_X1 U10274 ( .A1(n8130), .A2(n8550), .ZN(n10356) );
  OR2_X1 U10275 ( .A1(n10354), .A2(n10355), .ZN(n10443) );
  AND2_X1 U10276 ( .A1(n10446), .A2(n10447), .ZN(n10355) );
  NAND2_X1 U10277 ( .A1(n10448), .A2(b_26_), .ZN(n10447) );
  NOR2_X1 U10278 ( .A1(n10449), .A2(n8956), .ZN(n10448) );
  NOR2_X1 U10279 ( .A1(n10349), .A2(n10351), .ZN(n10449) );
  NAND2_X1 U10280 ( .A1(n10349), .A2(n10351), .ZN(n10446) );
  NAND2_X1 U10281 ( .A1(n10450), .A2(n10451), .ZN(n10351) );
  NAND2_X1 U10282 ( .A1(n10348), .A2(n10452), .ZN(n10451) );
  OR2_X1 U10283 ( .A1(n10346), .A2(n10347), .ZN(n10452) );
  NOR2_X1 U10284 ( .A1(n8130), .A2(n8495), .ZN(n10348) );
  NAND2_X1 U10285 ( .A1(n10346), .A2(n10347), .ZN(n10450) );
  NAND2_X1 U10286 ( .A1(n10453), .A2(n10454), .ZN(n10347) );
  NAND2_X1 U10287 ( .A1(n10455), .A2(b_26_), .ZN(n10454) );
  NOR2_X1 U10288 ( .A1(n10456), .A2(n8953), .ZN(n10455) );
  NOR2_X1 U10289 ( .A1(n10343), .A2(n10342), .ZN(n10456) );
  NAND2_X1 U10290 ( .A1(n10342), .A2(n10343), .ZN(n10453) );
  NAND2_X1 U10291 ( .A1(n10457), .A2(n10458), .ZN(n10343) );
  NAND2_X1 U10292 ( .A1(n10340), .A2(n10459), .ZN(n10458) );
  OR2_X1 U10293 ( .A1(n10338), .A2(n10339), .ZN(n10459) );
  NOR2_X1 U10294 ( .A1(n8130), .A2(n8440), .ZN(n10340) );
  NAND2_X1 U10295 ( .A1(n10338), .A2(n10339), .ZN(n10457) );
  NAND2_X1 U10296 ( .A1(n10460), .A2(n10461), .ZN(n10339) );
  NAND2_X1 U10297 ( .A1(n10462), .A2(b_26_), .ZN(n10461) );
  NOR2_X1 U10298 ( .A1(n10463), .A2(n8950), .ZN(n10462) );
  NOR2_X1 U10299 ( .A1(n10334), .A2(n10335), .ZN(n10463) );
  NAND2_X1 U10300 ( .A1(n10334), .A2(n10335), .ZN(n10460) );
  NAND2_X1 U10301 ( .A1(n10464), .A2(n10465), .ZN(n10335) );
  NAND2_X1 U10302 ( .A1(n10332), .A2(n10466), .ZN(n10465) );
  OR2_X1 U10303 ( .A1(n10330), .A2(n10331), .ZN(n10466) );
  NOR2_X1 U10304 ( .A1(n8130), .A2(n8385), .ZN(n10332) );
  NAND2_X1 U10305 ( .A1(n10330), .A2(n10331), .ZN(n10464) );
  NAND2_X1 U10306 ( .A1(n10467), .A2(n10468), .ZN(n10331) );
  NAND2_X1 U10307 ( .A1(n10469), .A2(b_26_), .ZN(n10468) );
  NOR2_X1 U10308 ( .A1(n10470), .A2(n8947), .ZN(n10469) );
  NOR2_X1 U10309 ( .A1(n10326), .A2(n10327), .ZN(n10470) );
  NAND2_X1 U10310 ( .A1(n10326), .A2(n10327), .ZN(n10467) );
  NAND2_X1 U10311 ( .A1(n10471), .A2(n10472), .ZN(n10327) );
  NAND2_X1 U10312 ( .A1(n10324), .A2(n10473), .ZN(n10472) );
  OR2_X1 U10313 ( .A1(n10322), .A2(n10323), .ZN(n10473) );
  NOR2_X1 U10314 ( .A1(n8130), .A2(n8324), .ZN(n10324) );
  NAND2_X1 U10315 ( .A1(n10322), .A2(n10323), .ZN(n10471) );
  NAND2_X1 U10316 ( .A1(n10474), .A2(n10475), .ZN(n10323) );
  NAND2_X1 U10317 ( .A1(n10476), .A2(b_26_), .ZN(n10475) );
  NOR2_X1 U10318 ( .A1(n10477), .A2(n8944), .ZN(n10476) );
  NOR2_X1 U10319 ( .A1(n10318), .A2(n10319), .ZN(n10477) );
  NAND2_X1 U10320 ( .A1(n10318), .A2(n10319), .ZN(n10474) );
  NAND2_X1 U10321 ( .A1(n10478), .A2(n10479), .ZN(n10319) );
  NAND2_X1 U10322 ( .A1(n10316), .A2(n10480), .ZN(n10479) );
  OR2_X1 U10323 ( .A1(n10313), .A2(n10315), .ZN(n10480) );
  NOR2_X1 U10324 ( .A1(n8130), .A2(n8268), .ZN(n10316) );
  NAND2_X1 U10325 ( .A1(n10313), .A2(n10315), .ZN(n10478) );
  NAND2_X1 U10326 ( .A1(n10481), .A2(n10482), .ZN(n10315) );
  NAND2_X1 U10327 ( .A1(n10483), .A2(b_26_), .ZN(n10482) );
  NOR2_X1 U10328 ( .A1(n10484), .A2(n8941), .ZN(n10483) );
  NOR2_X1 U10329 ( .A1(n10310), .A2(n10311), .ZN(n10484) );
  NAND2_X1 U10330 ( .A1(n10310), .A2(n10311), .ZN(n10481) );
  NAND2_X1 U10331 ( .A1(n10485), .A2(n10486), .ZN(n10311) );
  NAND2_X1 U10332 ( .A1(n10308), .A2(n10487), .ZN(n10486) );
  OR2_X1 U10333 ( .A1(n10305), .A2(n10307), .ZN(n10487) );
  NOR2_X1 U10334 ( .A1(n8130), .A2(n8213), .ZN(n10308) );
  NAND2_X1 U10335 ( .A1(n10305), .A2(n10307), .ZN(n10485) );
  NAND2_X1 U10336 ( .A1(n10488), .A2(n10489), .ZN(n10307) );
  NAND2_X1 U10337 ( .A1(n10490), .A2(b_26_), .ZN(n10489) );
  NOR2_X1 U10338 ( .A1(n10491), .A2(n8939), .ZN(n10490) );
  NOR2_X1 U10339 ( .A1(n10302), .A2(n10303), .ZN(n10491) );
  NAND2_X1 U10340 ( .A1(n10302), .A2(n10303), .ZN(n10488) );
  NAND2_X1 U10341 ( .A1(n10492), .A2(n10493), .ZN(n10303) );
  NAND2_X1 U10342 ( .A1(n10300), .A2(n10494), .ZN(n10493) );
  OR2_X1 U10343 ( .A1(n10297), .A2(n10299), .ZN(n10494) );
  NOR2_X1 U10344 ( .A1(n8130), .A2(n8158), .ZN(n10300) );
  NAND2_X1 U10345 ( .A1(n10297), .A2(n10299), .ZN(n10492) );
  NAND2_X1 U10346 ( .A1(n10495), .A2(n10496), .ZN(n10299) );
  NAND2_X1 U10347 ( .A1(n10294), .A2(n10497), .ZN(n10496) );
  OR2_X1 U10348 ( .A1(n10295), .A2(n10296), .ZN(n10497) );
  XNOR2_X1 U10349 ( .A(n10498), .B(n10499), .ZN(n10294) );
  NAND2_X1 U10350 ( .A1(n10500), .A2(n10501), .ZN(n10498) );
  NAND2_X1 U10351 ( .A1(n10296), .A2(n10295), .ZN(n10495) );
  NAND2_X1 U10352 ( .A1(n10266), .A2(n10502), .ZN(n10295) );
  NAND2_X1 U10353 ( .A1(n10265), .A2(n10267), .ZN(n10502) );
  NAND2_X1 U10354 ( .A1(n10503), .A2(n10504), .ZN(n10267) );
  NAND2_X1 U10355 ( .A1(b_26_), .A2(a_27_), .ZN(n10504) );
  INV_X1 U10356 ( .A(n10505), .ZN(n10503) );
  XOR2_X1 U10357 ( .A(n10506), .B(n10507), .Z(n10265) );
  XNOR2_X1 U10358 ( .A(n10508), .B(n10509), .ZN(n10506) );
  NAND2_X1 U10359 ( .A1(b_25_), .A2(a_28_), .ZN(n10508) );
  NAND2_X1 U10360 ( .A1(a_27_), .A2(n10505), .ZN(n10266) );
  NAND2_X1 U10361 ( .A1(n10510), .A2(n10511), .ZN(n10505) );
  NAND2_X1 U10362 ( .A1(n10512), .A2(b_26_), .ZN(n10511) );
  NOR2_X1 U10363 ( .A1(n10513), .A2(n8055), .ZN(n10512) );
  NOR2_X1 U10364 ( .A1(n10272), .A2(n10274), .ZN(n10513) );
  NAND2_X1 U10365 ( .A1(n10272), .A2(n10274), .ZN(n10510) );
  NAND2_X1 U10366 ( .A1(n10514), .A2(n10515), .ZN(n10274) );
  NAND2_X1 U10367 ( .A1(n10290), .A2(n10516), .ZN(n10515) );
  OR2_X1 U10368 ( .A1(n10291), .A2(n10292), .ZN(n10516) );
  NOR2_X1 U10369 ( .A1(n8130), .A2(n8041), .ZN(n10290) );
  NAND2_X1 U10370 ( .A1(n10292), .A2(n10291), .ZN(n10514) );
  NAND2_X1 U10371 ( .A1(n10517), .A2(n10518), .ZN(n10291) );
  NAND2_X1 U10372 ( .A1(b_24_), .A2(n10519), .ZN(n10518) );
  NAND2_X1 U10373 ( .A1(n8003), .A2(n10520), .ZN(n10519) );
  NAND2_X1 U10374 ( .A1(a_31_), .A2(n8938), .ZN(n10520) );
  NAND2_X1 U10375 ( .A1(b_25_), .A2(n10521), .ZN(n10517) );
  NAND2_X1 U10376 ( .A1(n9341), .A2(n10522), .ZN(n10521) );
  NAND2_X1 U10377 ( .A1(a_30_), .A2(n8185), .ZN(n10522) );
  AND2_X1 U10378 ( .A1(n10523), .A2(n7953), .ZN(n10292) );
  NOR2_X1 U10379 ( .A1(n8130), .A2(n8938), .ZN(n10523) );
  XOR2_X1 U10380 ( .A(n10524), .B(n10525), .Z(n10272) );
  XOR2_X1 U10381 ( .A(n10526), .B(n10527), .Z(n10524) );
  INV_X1 U10382 ( .A(n8920), .ZN(n10296) );
  NAND2_X1 U10383 ( .A1(b_26_), .A2(a_26_), .ZN(n8920) );
  XNOR2_X1 U10384 ( .A(n10528), .B(n10529), .ZN(n10297) );
  NAND2_X1 U10385 ( .A1(n10530), .A2(n10531), .ZN(n10528) );
  XNOR2_X1 U10386 ( .A(n10532), .B(n10533), .ZN(n10302) );
  XNOR2_X1 U10387 ( .A(n10534), .B(n8917), .ZN(n10533) );
  XOR2_X1 U10388 ( .A(n10535), .B(n10536), .Z(n10305) );
  XOR2_X1 U10389 ( .A(n10537), .B(n10538), .Z(n10535) );
  NOR2_X1 U10390 ( .A1(n8939), .A2(n8938), .ZN(n10538) );
  XNOR2_X1 U10391 ( .A(n10539), .B(n10540), .ZN(n10310) );
  XNOR2_X1 U10392 ( .A(n10541), .B(n10542), .ZN(n10540) );
  XOR2_X1 U10393 ( .A(n10543), .B(n10544), .Z(n10313) );
  XOR2_X1 U10394 ( .A(n10545), .B(n10546), .Z(n10543) );
  NOR2_X1 U10395 ( .A1(n8941), .A2(n8938), .ZN(n10546) );
  XOR2_X1 U10396 ( .A(n10547), .B(n10548), .Z(n10318) );
  XOR2_X1 U10397 ( .A(n10549), .B(n10550), .Z(n10547) );
  XOR2_X1 U10398 ( .A(n10551), .B(n10552), .Z(n10322) );
  XOR2_X1 U10399 ( .A(n10553), .B(n10554), .Z(n10551) );
  NOR2_X1 U10400 ( .A1(n8944), .A2(n8938), .ZN(n10554) );
  XNOR2_X1 U10401 ( .A(n10555), .B(n10556), .ZN(n10326) );
  XNOR2_X1 U10402 ( .A(n10557), .B(n10558), .ZN(n10556) );
  XOR2_X1 U10403 ( .A(n10559), .B(n10560), .Z(n10330) );
  XOR2_X1 U10404 ( .A(n10561), .B(n10562), .Z(n10559) );
  NOR2_X1 U10405 ( .A1(n8947), .A2(n8938), .ZN(n10562) );
  XOR2_X1 U10406 ( .A(n10563), .B(n10564), .Z(n10334) );
  XOR2_X1 U10407 ( .A(n10565), .B(n10566), .Z(n10563) );
  XOR2_X1 U10408 ( .A(n10567), .B(n10568), .Z(n10338) );
  XOR2_X1 U10409 ( .A(n10569), .B(n10570), .Z(n10567) );
  NOR2_X1 U10410 ( .A1(n8950), .A2(n8938), .ZN(n10570) );
  XNOR2_X1 U10411 ( .A(n10571), .B(n10572), .ZN(n10342) );
  XNOR2_X1 U10412 ( .A(n10573), .B(n10574), .ZN(n10571) );
  XNOR2_X1 U10413 ( .A(n10575), .B(n10576), .ZN(n10346) );
  XOR2_X1 U10414 ( .A(n10577), .B(n10578), .Z(n10576) );
  NAND2_X1 U10415 ( .A1(b_25_), .A2(a_14_), .ZN(n10578) );
  XOR2_X1 U10416 ( .A(n10579), .B(n10580), .Z(n10349) );
  XOR2_X1 U10417 ( .A(n10581), .B(n10582), .Z(n10579) );
  XNOR2_X1 U10418 ( .A(n10583), .B(n10584), .ZN(n10354) );
  XOR2_X1 U10419 ( .A(n10585), .B(n10586), .Z(n10583) );
  NOR2_X1 U10420 ( .A1(n8956), .A2(n8938), .ZN(n10586) );
  XOR2_X1 U10421 ( .A(n10587), .B(n10588), .Z(n10357) );
  XOR2_X1 U10422 ( .A(n10589), .B(n10590), .Z(n10587) );
  NOR2_X1 U10423 ( .A1(n8550), .A2(n8938), .ZN(n10590) );
  XOR2_X1 U10424 ( .A(n10591), .B(n10592), .Z(n10362) );
  XOR2_X1 U10425 ( .A(n10593), .B(n10594), .Z(n10591) );
  NOR2_X1 U10426 ( .A1(n8959), .A2(n8938), .ZN(n10594) );
  XOR2_X1 U10427 ( .A(n10595), .B(n10596), .Z(n10366) );
  XOR2_X1 U10428 ( .A(n10597), .B(n10598), .Z(n10595) );
  XNOR2_X1 U10429 ( .A(n10599), .B(n10600), .ZN(n10374) );
  NAND2_X1 U10430 ( .A1(n10601), .A2(n10602), .ZN(n10599) );
  XNOR2_X1 U10431 ( .A(n10603), .B(n10604), .ZN(n10378) );
  XNOR2_X1 U10432 ( .A(n10605), .B(n10606), .ZN(n10603) );
  XNOR2_X1 U10433 ( .A(n10607), .B(n10608), .ZN(n10179) );
  XOR2_X1 U10434 ( .A(n10609), .B(n10610), .Z(n10607) );
  NOR2_X1 U10435 ( .A1(n8723), .A2(n8938), .ZN(n10610) );
  XNOR2_X1 U10436 ( .A(n10611), .B(n10612), .ZN(n10171) );
  XOR2_X1 U10437 ( .A(n10613), .B(n10614), .Z(n10611) );
  NOR2_X1 U10438 ( .A1(n8966), .A2(n8938), .ZN(n10614) );
  XNOR2_X1 U10439 ( .A(n10615), .B(n10616), .ZN(n10386) );
  NAND2_X1 U10440 ( .A1(n10617), .A2(n10618), .ZN(n10615) );
  XNOR2_X1 U10441 ( .A(n10619), .B(n10620), .ZN(n10156) );
  XOR2_X1 U10442 ( .A(n10621), .B(n10622), .Z(n10619) );
  NOR2_X1 U10443 ( .A1(n8969), .A2(n8938), .ZN(n10622) );
  XOR2_X1 U10444 ( .A(n10623), .B(n10624), .Z(n9193) );
  XNOR2_X1 U10445 ( .A(n10625), .B(n10626), .ZN(n10623) );
  AND2_X1 U10446 ( .A1(n9188), .A2(n10392), .ZN(n10394) );
  NAND2_X1 U10447 ( .A1(n10627), .A2(n10628), .ZN(n10392) );
  XOR2_X1 U10448 ( .A(n10629), .B(n10630), .Z(n10628) );
  NOR2_X1 U10449 ( .A1(n10631), .A2(n10632), .ZN(n10627) );
  NOR2_X1 U10450 ( .A1(n10625), .A2(n10624), .ZN(n10632) );
  INV_X1 U10451 ( .A(n10633), .ZN(n10631) );
  OR2_X1 U10452 ( .A1(n9188), .A2(n9187), .ZN(n9026) );
  XNOR2_X1 U10453 ( .A(n9184), .B(n9183), .ZN(n9187) );
  NAND2_X1 U10454 ( .A1(n10634), .A2(n10635), .ZN(n9188) );
  NAND2_X1 U10455 ( .A1(n10636), .A2(n10633), .ZN(n10635) );
  NAND2_X1 U10456 ( .A1(n10626), .A2(n10637), .ZN(n10633) );
  NAND2_X1 U10457 ( .A1(n10625), .A2(n10624), .ZN(n10637) );
  NOR2_X1 U10458 ( .A1(n8938), .A2(n8974), .ZN(n10626) );
  OR2_X1 U10459 ( .A1(n10624), .A2(n10625), .ZN(n10636) );
  AND2_X1 U10460 ( .A1(n10638), .A2(n10639), .ZN(n10625) );
  NAND2_X1 U10461 ( .A1(n10640), .A2(b_25_), .ZN(n10639) );
  NOR2_X1 U10462 ( .A1(n10641), .A2(n8969), .ZN(n10640) );
  NOR2_X1 U10463 ( .A1(n10620), .A2(n10621), .ZN(n10641) );
  NAND2_X1 U10464 ( .A1(n10620), .A2(n10621), .ZN(n10638) );
  NAND2_X1 U10465 ( .A1(n10617), .A2(n10642), .ZN(n10621) );
  NAND2_X1 U10466 ( .A1(n10616), .A2(n10618), .ZN(n10642) );
  NAND2_X1 U10467 ( .A1(n10643), .A2(n10644), .ZN(n10618) );
  NAND2_X1 U10468 ( .A1(b_25_), .A2(a_2_), .ZN(n10644) );
  INV_X1 U10469 ( .A(n10645), .ZN(n10643) );
  XNOR2_X1 U10470 ( .A(n10646), .B(n10647), .ZN(n10616) );
  NAND2_X1 U10471 ( .A1(n10648), .A2(n10649), .ZN(n10646) );
  NAND2_X1 U10472 ( .A1(a_2_), .A2(n10645), .ZN(n10617) );
  NAND2_X1 U10473 ( .A1(n10650), .A2(n10651), .ZN(n10645) );
  NAND2_X1 U10474 ( .A1(n10652), .A2(b_25_), .ZN(n10651) );
  NOR2_X1 U10475 ( .A1(n10653), .A2(n8778), .ZN(n10652) );
  NOR2_X1 U10476 ( .A1(n10407), .A2(n10408), .ZN(n10653) );
  NAND2_X1 U10477 ( .A1(n10407), .A2(n10408), .ZN(n10650) );
  NAND2_X1 U10478 ( .A1(n10654), .A2(n10655), .ZN(n10408) );
  NAND2_X1 U10479 ( .A1(n10656), .A2(b_25_), .ZN(n10655) );
  NOR2_X1 U10480 ( .A1(n10657), .A2(n8966), .ZN(n10656) );
  NOR2_X1 U10481 ( .A1(n10612), .A2(n10613), .ZN(n10657) );
  NAND2_X1 U10482 ( .A1(n10612), .A2(n10613), .ZN(n10654) );
  NAND2_X1 U10483 ( .A1(n10658), .A2(n10659), .ZN(n10613) );
  NAND2_X1 U10484 ( .A1(n10660), .A2(b_25_), .ZN(n10659) );
  NOR2_X1 U10485 ( .A1(n10661), .A2(n8723), .ZN(n10660) );
  NOR2_X1 U10486 ( .A1(n10608), .A2(n10609), .ZN(n10661) );
  NAND2_X1 U10487 ( .A1(n10608), .A2(n10609), .ZN(n10658) );
  NAND2_X1 U10488 ( .A1(n10662), .A2(n10663), .ZN(n10609) );
  NAND2_X1 U10489 ( .A1(n10605), .A2(n10664), .ZN(n10663) );
  NAND2_X1 U10490 ( .A1(n10604), .A2(n10606), .ZN(n10664) );
  NAND2_X1 U10491 ( .A1(n10601), .A2(n10665), .ZN(n10605) );
  NAND2_X1 U10492 ( .A1(n10600), .A2(n10602), .ZN(n10665) );
  NAND2_X1 U10493 ( .A1(n10666), .A2(n10667), .ZN(n10602) );
  NAND2_X1 U10494 ( .A1(b_25_), .A2(a_7_), .ZN(n10667) );
  INV_X1 U10495 ( .A(n10668), .ZN(n10666) );
  XOR2_X1 U10496 ( .A(n10669), .B(n10670), .Z(n10600) );
  XOR2_X1 U10497 ( .A(n10671), .B(n10672), .Z(n10669) );
  NOR2_X1 U10498 ( .A1(n8619), .A2(n8185), .ZN(n10672) );
  NAND2_X1 U10499 ( .A1(a_7_), .A2(n10668), .ZN(n10601) );
  NAND2_X1 U10500 ( .A1(n10673), .A2(n10674), .ZN(n10668) );
  NAND2_X1 U10501 ( .A1(n10675), .A2(b_25_), .ZN(n10674) );
  NOR2_X1 U10502 ( .A1(n10676), .A2(n8619), .ZN(n10675) );
  NOR2_X1 U10503 ( .A1(n10429), .A2(n10430), .ZN(n10676) );
  NAND2_X1 U10504 ( .A1(n10429), .A2(n10430), .ZN(n10673) );
  NAND2_X1 U10505 ( .A1(n10677), .A2(n10678), .ZN(n10430) );
  NAND2_X1 U10506 ( .A1(n10598), .A2(n10679), .ZN(n10678) );
  OR2_X1 U10507 ( .A1(n10597), .A2(n10596), .ZN(n10679) );
  NOR2_X1 U10508 ( .A1(n8938), .A2(n8605), .ZN(n10598) );
  NAND2_X1 U10509 ( .A1(n10596), .A2(n10597), .ZN(n10677) );
  NAND2_X1 U10510 ( .A1(n10680), .A2(n10681), .ZN(n10597) );
  NAND2_X1 U10511 ( .A1(n10682), .A2(b_25_), .ZN(n10681) );
  NOR2_X1 U10512 ( .A1(n10683), .A2(n8959), .ZN(n10682) );
  NOR2_X1 U10513 ( .A1(n10592), .A2(n10593), .ZN(n10683) );
  NAND2_X1 U10514 ( .A1(n10592), .A2(n10593), .ZN(n10680) );
  NAND2_X1 U10515 ( .A1(n10684), .A2(n10685), .ZN(n10593) );
  NAND2_X1 U10516 ( .A1(n10686), .A2(b_25_), .ZN(n10685) );
  NOR2_X1 U10517 ( .A1(n10687), .A2(n8550), .ZN(n10686) );
  NOR2_X1 U10518 ( .A1(n10588), .A2(n10589), .ZN(n10687) );
  NAND2_X1 U10519 ( .A1(n10588), .A2(n10589), .ZN(n10684) );
  NAND2_X1 U10520 ( .A1(n10688), .A2(n10689), .ZN(n10589) );
  NAND2_X1 U10521 ( .A1(n10690), .A2(b_25_), .ZN(n10689) );
  NOR2_X1 U10522 ( .A1(n10691), .A2(n8956), .ZN(n10690) );
  NOR2_X1 U10523 ( .A1(n10584), .A2(n10585), .ZN(n10691) );
  NAND2_X1 U10524 ( .A1(n10584), .A2(n10585), .ZN(n10688) );
  NAND2_X1 U10525 ( .A1(n10692), .A2(n10693), .ZN(n10585) );
  NAND2_X1 U10526 ( .A1(n10582), .A2(n10694), .ZN(n10693) );
  OR2_X1 U10527 ( .A1(n10581), .A2(n10580), .ZN(n10694) );
  NOR2_X1 U10528 ( .A1(n8938), .A2(n8495), .ZN(n10582) );
  NAND2_X1 U10529 ( .A1(n10580), .A2(n10581), .ZN(n10692) );
  NAND2_X1 U10530 ( .A1(n10695), .A2(n10696), .ZN(n10581) );
  NAND2_X1 U10531 ( .A1(n10697), .A2(b_25_), .ZN(n10696) );
  NOR2_X1 U10532 ( .A1(n10698), .A2(n8953), .ZN(n10697) );
  NOR2_X1 U10533 ( .A1(n10575), .A2(n10577), .ZN(n10698) );
  NAND2_X1 U10534 ( .A1(n10575), .A2(n10577), .ZN(n10695) );
  NAND2_X1 U10535 ( .A1(n10699), .A2(n10700), .ZN(n10577) );
  NAND2_X1 U10536 ( .A1(n10574), .A2(n10701), .ZN(n10700) );
  NAND2_X1 U10537 ( .A1(n10573), .A2(n10572), .ZN(n10701) );
  NOR2_X1 U10538 ( .A1(n8938), .A2(n8440), .ZN(n10574) );
  OR2_X1 U10539 ( .A1(n10572), .A2(n10573), .ZN(n10699) );
  AND2_X1 U10540 ( .A1(n10702), .A2(n10703), .ZN(n10573) );
  NAND2_X1 U10541 ( .A1(n10704), .A2(b_25_), .ZN(n10703) );
  NOR2_X1 U10542 ( .A1(n10705), .A2(n8950), .ZN(n10704) );
  NOR2_X1 U10543 ( .A1(n10568), .A2(n10569), .ZN(n10705) );
  NAND2_X1 U10544 ( .A1(n10568), .A2(n10569), .ZN(n10702) );
  NAND2_X1 U10545 ( .A1(n10706), .A2(n10707), .ZN(n10569) );
  NAND2_X1 U10546 ( .A1(n10566), .A2(n10708), .ZN(n10707) );
  OR2_X1 U10547 ( .A1(n10565), .A2(n10564), .ZN(n10708) );
  NOR2_X1 U10548 ( .A1(n8938), .A2(n8385), .ZN(n10566) );
  NAND2_X1 U10549 ( .A1(n10564), .A2(n10565), .ZN(n10706) );
  NAND2_X1 U10550 ( .A1(n10709), .A2(n10710), .ZN(n10565) );
  NAND2_X1 U10551 ( .A1(n10711), .A2(b_25_), .ZN(n10710) );
  NOR2_X1 U10552 ( .A1(n10712), .A2(n8947), .ZN(n10711) );
  NOR2_X1 U10553 ( .A1(n10560), .A2(n10561), .ZN(n10712) );
  NAND2_X1 U10554 ( .A1(n10560), .A2(n10561), .ZN(n10709) );
  NAND2_X1 U10555 ( .A1(n10713), .A2(n10714), .ZN(n10561) );
  NAND2_X1 U10556 ( .A1(n10558), .A2(n10715), .ZN(n10714) );
  OR2_X1 U10557 ( .A1(n10557), .A2(n10555), .ZN(n10715) );
  NOR2_X1 U10558 ( .A1(n8938), .A2(n8324), .ZN(n10558) );
  NAND2_X1 U10559 ( .A1(n10555), .A2(n10557), .ZN(n10713) );
  NAND2_X1 U10560 ( .A1(n10716), .A2(n10717), .ZN(n10557) );
  NAND2_X1 U10561 ( .A1(n10718), .A2(b_25_), .ZN(n10717) );
  NOR2_X1 U10562 ( .A1(n10719), .A2(n8944), .ZN(n10718) );
  NOR2_X1 U10563 ( .A1(n10552), .A2(n10553), .ZN(n10719) );
  NAND2_X1 U10564 ( .A1(n10552), .A2(n10553), .ZN(n10716) );
  NAND2_X1 U10565 ( .A1(n10720), .A2(n10721), .ZN(n10553) );
  NAND2_X1 U10566 ( .A1(n10550), .A2(n10722), .ZN(n10721) );
  OR2_X1 U10567 ( .A1(n10549), .A2(n10548), .ZN(n10722) );
  NOR2_X1 U10568 ( .A1(n8938), .A2(n8268), .ZN(n10550) );
  NAND2_X1 U10569 ( .A1(n10548), .A2(n10549), .ZN(n10720) );
  NAND2_X1 U10570 ( .A1(n10723), .A2(n10724), .ZN(n10549) );
  NAND2_X1 U10571 ( .A1(n10725), .A2(b_25_), .ZN(n10724) );
  NOR2_X1 U10572 ( .A1(n10726), .A2(n8941), .ZN(n10725) );
  NOR2_X1 U10573 ( .A1(n10544), .A2(n10545), .ZN(n10726) );
  NAND2_X1 U10574 ( .A1(n10544), .A2(n10545), .ZN(n10723) );
  NAND2_X1 U10575 ( .A1(n10727), .A2(n10728), .ZN(n10545) );
  NAND2_X1 U10576 ( .A1(n10542), .A2(n10729), .ZN(n10728) );
  OR2_X1 U10577 ( .A1(n10541), .A2(n10539), .ZN(n10729) );
  NOR2_X1 U10578 ( .A1(n8938), .A2(n8213), .ZN(n10542) );
  NAND2_X1 U10579 ( .A1(n10539), .A2(n10541), .ZN(n10727) );
  NAND2_X1 U10580 ( .A1(n10730), .A2(n10731), .ZN(n10541) );
  NAND2_X1 U10581 ( .A1(n10732), .A2(b_25_), .ZN(n10731) );
  NOR2_X1 U10582 ( .A1(n10733), .A2(n8939), .ZN(n10732) );
  NOR2_X1 U10583 ( .A1(n10536), .A2(n10537), .ZN(n10733) );
  NAND2_X1 U10584 ( .A1(n10536), .A2(n10537), .ZN(n10730) );
  NAND2_X1 U10585 ( .A1(n10734), .A2(n10735), .ZN(n10537) );
  NAND2_X1 U10586 ( .A1(n8917), .A2(n10736), .ZN(n10735) );
  OR2_X1 U10587 ( .A1(n10534), .A2(n10532), .ZN(n10736) );
  NOR2_X1 U10588 ( .A1(n8938), .A2(n8158), .ZN(n8917) );
  NAND2_X1 U10589 ( .A1(n10532), .A2(n10534), .ZN(n10734) );
  NAND2_X1 U10590 ( .A1(n10530), .A2(n10737), .ZN(n10534) );
  NAND2_X1 U10591 ( .A1(n10529), .A2(n10531), .ZN(n10737) );
  NAND2_X1 U10592 ( .A1(n10738), .A2(n10739), .ZN(n10531) );
  NAND2_X1 U10593 ( .A1(b_25_), .A2(a_26_), .ZN(n10739) );
  INV_X1 U10594 ( .A(n10740), .ZN(n10738) );
  XNOR2_X1 U10595 ( .A(n10741), .B(n10742), .ZN(n10529) );
  NAND2_X1 U10596 ( .A1(n10743), .A2(n10744), .ZN(n10741) );
  NAND2_X1 U10597 ( .A1(a_26_), .A2(n10740), .ZN(n10530) );
  NAND2_X1 U10598 ( .A1(n10500), .A2(n10745), .ZN(n10740) );
  NAND2_X1 U10599 ( .A1(n10499), .A2(n10501), .ZN(n10745) );
  NAND2_X1 U10600 ( .A1(n10746), .A2(n10747), .ZN(n10501) );
  NAND2_X1 U10601 ( .A1(b_25_), .A2(a_27_), .ZN(n10747) );
  INV_X1 U10602 ( .A(n10748), .ZN(n10746) );
  XOR2_X1 U10603 ( .A(n10749), .B(n10750), .Z(n10499) );
  XNOR2_X1 U10604 ( .A(n10751), .B(n10752), .ZN(n10749) );
  NAND2_X1 U10605 ( .A1(b_24_), .A2(a_28_), .ZN(n10751) );
  NAND2_X1 U10606 ( .A1(a_27_), .A2(n10748), .ZN(n10500) );
  NAND2_X1 U10607 ( .A1(n10753), .A2(n10754), .ZN(n10748) );
  NAND2_X1 U10608 ( .A1(n10755), .A2(b_25_), .ZN(n10754) );
  NOR2_X1 U10609 ( .A1(n10756), .A2(n8055), .ZN(n10755) );
  NOR2_X1 U10610 ( .A1(n10507), .A2(n10509), .ZN(n10756) );
  NAND2_X1 U10611 ( .A1(n10507), .A2(n10509), .ZN(n10753) );
  NAND2_X1 U10612 ( .A1(n10757), .A2(n10758), .ZN(n10509) );
  NAND2_X1 U10613 ( .A1(n10525), .A2(n10759), .ZN(n10758) );
  OR2_X1 U10614 ( .A1(n10526), .A2(n10527), .ZN(n10759) );
  NOR2_X1 U10615 ( .A1(n8938), .A2(n8041), .ZN(n10525) );
  NAND2_X1 U10616 ( .A1(n10527), .A2(n10526), .ZN(n10757) );
  NAND2_X1 U10617 ( .A1(n10760), .A2(n10761), .ZN(n10526) );
  NAND2_X1 U10618 ( .A1(b_23_), .A2(n10762), .ZN(n10761) );
  NAND2_X1 U10619 ( .A1(n8003), .A2(n10763), .ZN(n10762) );
  NAND2_X1 U10620 ( .A1(a_31_), .A2(n8185), .ZN(n10763) );
  NAND2_X1 U10621 ( .A1(b_24_), .A2(n10764), .ZN(n10760) );
  NAND2_X1 U10622 ( .A1(n9341), .A2(n10765), .ZN(n10764) );
  NAND2_X1 U10623 ( .A1(a_30_), .A2(n8940), .ZN(n10765) );
  AND2_X1 U10624 ( .A1(n10766), .A2(n7953), .ZN(n10527) );
  NOR2_X1 U10625 ( .A1(n8938), .A2(n8185), .ZN(n10766) );
  XOR2_X1 U10626 ( .A(n10767), .B(n10768), .Z(n10507) );
  XOR2_X1 U10627 ( .A(n10769), .B(n10770), .Z(n10767) );
  XNOR2_X1 U10628 ( .A(n10771), .B(n10772), .ZN(n10532) );
  NAND2_X1 U10629 ( .A1(n10773), .A2(n10774), .ZN(n10771) );
  XNOR2_X1 U10630 ( .A(n10775), .B(n10776), .ZN(n10536) );
  XNOR2_X1 U10631 ( .A(n10777), .B(n10778), .ZN(n10776) );
  XOR2_X1 U10632 ( .A(n10779), .B(n10780), .Z(n10539) );
  XOR2_X1 U10633 ( .A(n10781), .B(n10782), .Z(n10779) );
  XNOR2_X1 U10634 ( .A(n10783), .B(n10784), .ZN(n10544) );
  XNOR2_X1 U10635 ( .A(n10785), .B(n10786), .ZN(n10784) );
  XOR2_X1 U10636 ( .A(n10787), .B(n10788), .Z(n10548) );
  XOR2_X1 U10637 ( .A(n10789), .B(n10790), .Z(n10787) );
  NOR2_X1 U10638 ( .A1(n8941), .A2(n8185), .ZN(n10790) );
  XNOR2_X1 U10639 ( .A(n10791), .B(n10792), .ZN(n10552) );
  XNOR2_X1 U10640 ( .A(n10793), .B(n10794), .ZN(n10792) );
  XOR2_X1 U10641 ( .A(n10795), .B(n10796), .Z(n10555) );
  XOR2_X1 U10642 ( .A(n10797), .B(n10798), .Z(n10795) );
  NOR2_X1 U10643 ( .A1(n8944), .A2(n8185), .ZN(n10798) );
  XNOR2_X1 U10644 ( .A(n10799), .B(n10800), .ZN(n10560) );
  XNOR2_X1 U10645 ( .A(n10801), .B(n10802), .ZN(n10800) );
  XOR2_X1 U10646 ( .A(n10803), .B(n10804), .Z(n10564) );
  XOR2_X1 U10647 ( .A(n10805), .B(n10806), .Z(n10803) );
  NOR2_X1 U10648 ( .A1(n8947), .A2(n8185), .ZN(n10806) );
  XOR2_X1 U10649 ( .A(n10807), .B(n10808), .Z(n10568) );
  XOR2_X1 U10650 ( .A(n10809), .B(n10810), .Z(n10807) );
  XOR2_X1 U10651 ( .A(n10811), .B(n10812), .Z(n10572) );
  XOR2_X1 U10652 ( .A(n10813), .B(n10814), .Z(n10812) );
  NAND2_X1 U10653 ( .A1(b_24_), .A2(a_16_), .ZN(n10814) );
  XOR2_X1 U10654 ( .A(n10815), .B(n10816), .Z(n10575) );
  XOR2_X1 U10655 ( .A(n10817), .B(n10818), .Z(n10815) );
  XOR2_X1 U10656 ( .A(n10819), .B(n10820), .Z(n10580) );
  XOR2_X1 U10657 ( .A(n10821), .B(n10822), .Z(n10819) );
  NOR2_X1 U10658 ( .A1(n8953), .A2(n8185), .ZN(n10822) );
  XNOR2_X1 U10659 ( .A(n10823), .B(n10824), .ZN(n10584) );
  XNOR2_X1 U10660 ( .A(n10825), .B(n10826), .ZN(n10823) );
  XOR2_X1 U10661 ( .A(n10827), .B(n10828), .Z(n10588) );
  XOR2_X1 U10662 ( .A(n10829), .B(n10830), .Z(n10827) );
  NOR2_X1 U10663 ( .A1(n8956), .A2(n8185), .ZN(n10830) );
  XOR2_X1 U10664 ( .A(n10831), .B(n10832), .Z(n10592) );
  XOR2_X1 U10665 ( .A(n10833), .B(n10834), .Z(n10831) );
  NOR2_X1 U10666 ( .A1(n8550), .A2(n8185), .ZN(n10834) );
  XOR2_X1 U10667 ( .A(n10835), .B(n10836), .Z(n10596) );
  XOR2_X1 U10668 ( .A(n10837), .B(n10838), .Z(n10835) );
  NOR2_X1 U10669 ( .A1(n8959), .A2(n8185), .ZN(n10838) );
  XNOR2_X1 U10670 ( .A(n10839), .B(n10840), .ZN(n10429) );
  XNOR2_X1 U10671 ( .A(n10841), .B(n10842), .ZN(n10839) );
  OR2_X1 U10672 ( .A1(n10606), .A2(n10604), .ZN(n10662) );
  XOR2_X1 U10673 ( .A(n10843), .B(n10844), .Z(n10604) );
  NAND2_X1 U10674 ( .A1(n10845), .A2(n10846), .ZN(n10843) );
  NAND2_X1 U10675 ( .A1(b_25_), .A2(a_6_), .ZN(n10606) );
  XNOR2_X1 U10676 ( .A(n10847), .B(n10848), .ZN(n10608) );
  XNOR2_X1 U10677 ( .A(n10849), .B(n10850), .ZN(n10847) );
  XNOR2_X1 U10678 ( .A(n10851), .B(n10852), .ZN(n10612) );
  XNOR2_X1 U10679 ( .A(n10853), .B(n10854), .ZN(n10851) );
  XOR2_X1 U10680 ( .A(n10855), .B(n10856), .Z(n10407) );
  XOR2_X1 U10681 ( .A(n10857), .B(n10858), .Z(n10855) );
  NOR2_X1 U10682 ( .A1(n8966), .A2(n8185), .ZN(n10858) );
  XNOR2_X1 U10683 ( .A(n10859), .B(n10860), .ZN(n10620) );
  NAND2_X1 U10684 ( .A1(n10861), .A2(n10862), .ZN(n10859) );
  XNOR2_X1 U10685 ( .A(n10863), .B(n10864), .ZN(n10624) );
  XOR2_X1 U10686 ( .A(n10865), .B(n10866), .Z(n10863) );
  XOR2_X1 U10687 ( .A(n10867), .B(n10629), .Z(n10634) );
  XNOR2_X1 U10688 ( .A(n10868), .B(n10869), .ZN(n10629) );
  NOR2_X1 U10689 ( .A1(n8974), .A2(n8185), .ZN(n10869) );
  INV_X1 U10690 ( .A(n10630), .ZN(n10867) );
  NAND2_X1 U10691 ( .A1(n10870), .A2(n10871), .ZN(n9032) );
  XOR2_X1 U10692 ( .A(n9177), .B(n9176), .Z(n10871) );
  INV_X1 U10693 ( .A(n9185), .ZN(n9176) );
  AND2_X1 U10694 ( .A1(n9184), .A2(n9183), .ZN(n10870) );
  XOR2_X1 U10695 ( .A(n10872), .B(n10873), .Z(n9183) );
  XOR2_X1 U10696 ( .A(n10874), .B(n10875), .Z(n10872) );
  NOR2_X1 U10697 ( .A1(n8974), .A2(n8940), .ZN(n10875) );
  NAND2_X1 U10698 ( .A1(n10876), .A2(n10877), .ZN(n9184) );
  NAND2_X1 U10699 ( .A1(n10878), .A2(b_24_), .ZN(n10877) );
  NOR2_X1 U10700 ( .A1(n10879), .A2(n8974), .ZN(n10878) );
  NOR2_X1 U10701 ( .A1(n10630), .A2(n10868), .ZN(n10879) );
  NAND2_X1 U10702 ( .A1(n10630), .A2(n10868), .ZN(n10876) );
  NAND2_X1 U10703 ( .A1(n10880), .A2(n10881), .ZN(n10868) );
  NAND2_X1 U10704 ( .A1(n10865), .A2(n10882), .ZN(n10881) );
  OR2_X1 U10705 ( .A1(n10864), .A2(n10866), .ZN(n10882) );
  NAND2_X1 U10706 ( .A1(n10861), .A2(n10883), .ZN(n10865) );
  NAND2_X1 U10707 ( .A1(n10860), .A2(n10862), .ZN(n10883) );
  NAND2_X1 U10708 ( .A1(n10884), .A2(n10885), .ZN(n10862) );
  NAND2_X1 U10709 ( .A1(b_24_), .A2(a_2_), .ZN(n10885) );
  INV_X1 U10710 ( .A(n10886), .ZN(n10884) );
  XNOR2_X1 U10711 ( .A(n10887), .B(n10888), .ZN(n10860) );
  XOR2_X1 U10712 ( .A(n10889), .B(n10890), .Z(n10888) );
  NAND2_X1 U10713 ( .A1(b_23_), .A2(a_3_), .ZN(n10890) );
  NAND2_X1 U10714 ( .A1(a_2_), .A2(n10886), .ZN(n10861) );
  NAND2_X1 U10715 ( .A1(n10648), .A2(n10891), .ZN(n10886) );
  NAND2_X1 U10716 ( .A1(n10647), .A2(n10649), .ZN(n10891) );
  NAND2_X1 U10717 ( .A1(n10892), .A2(n10893), .ZN(n10649) );
  NAND2_X1 U10718 ( .A1(b_24_), .A2(a_3_), .ZN(n10893) );
  INV_X1 U10719 ( .A(n10894), .ZN(n10892) );
  XOR2_X1 U10720 ( .A(n10895), .B(n10896), .Z(n10647) );
  XOR2_X1 U10721 ( .A(n10897), .B(n10898), .Z(n10895) );
  NOR2_X1 U10722 ( .A1(n8966), .A2(n8940), .ZN(n10898) );
  NAND2_X1 U10723 ( .A1(a_3_), .A2(n10894), .ZN(n10648) );
  NAND2_X1 U10724 ( .A1(n10899), .A2(n10900), .ZN(n10894) );
  NAND2_X1 U10725 ( .A1(n10901), .A2(b_24_), .ZN(n10900) );
  NOR2_X1 U10726 ( .A1(n10902), .A2(n8966), .ZN(n10901) );
  NOR2_X1 U10727 ( .A1(n10856), .A2(n10857), .ZN(n10902) );
  NAND2_X1 U10728 ( .A1(n10856), .A2(n10857), .ZN(n10899) );
  NAND2_X1 U10729 ( .A1(n10903), .A2(n10904), .ZN(n10857) );
  NAND2_X1 U10730 ( .A1(n10854), .A2(n10905), .ZN(n10904) );
  NAND2_X1 U10731 ( .A1(n10853), .A2(n10852), .ZN(n10905) );
  NOR2_X1 U10732 ( .A1(n8185), .A2(n8723), .ZN(n10854) );
  OR2_X1 U10733 ( .A1(n10852), .A2(n10853), .ZN(n10903) );
  AND2_X1 U10734 ( .A1(n10906), .A2(n10907), .ZN(n10853) );
  NAND2_X1 U10735 ( .A1(n10849), .A2(n10908), .ZN(n10907) );
  NAND2_X1 U10736 ( .A1(n10848), .A2(n10850), .ZN(n10908) );
  NAND2_X1 U10737 ( .A1(n10845), .A2(n10909), .ZN(n10849) );
  NAND2_X1 U10738 ( .A1(n10844), .A2(n10846), .ZN(n10909) );
  NAND2_X1 U10739 ( .A1(n10910), .A2(n10911), .ZN(n10846) );
  NAND2_X1 U10740 ( .A1(b_24_), .A2(a_7_), .ZN(n10911) );
  INV_X1 U10741 ( .A(n10912), .ZN(n10910) );
  XNOR2_X1 U10742 ( .A(n10913), .B(n10914), .ZN(n10844) );
  XNOR2_X1 U10743 ( .A(n10915), .B(n10916), .ZN(n10914) );
  NAND2_X1 U10744 ( .A1(a_7_), .A2(n10912), .ZN(n10845) );
  NAND2_X1 U10745 ( .A1(n10917), .A2(n10918), .ZN(n10912) );
  NAND2_X1 U10746 ( .A1(n10919), .A2(b_24_), .ZN(n10918) );
  NOR2_X1 U10747 ( .A1(n10920), .A2(n8619), .ZN(n10919) );
  NOR2_X1 U10748 ( .A1(n10670), .A2(n10671), .ZN(n10920) );
  NAND2_X1 U10749 ( .A1(n10670), .A2(n10671), .ZN(n10917) );
  NAND2_X1 U10750 ( .A1(n10921), .A2(n10922), .ZN(n10671) );
  NAND2_X1 U10751 ( .A1(n10842), .A2(n10923), .ZN(n10922) );
  NAND2_X1 U10752 ( .A1(n10841), .A2(n10840), .ZN(n10923) );
  NOR2_X1 U10753 ( .A1(n8185), .A2(n8605), .ZN(n10842) );
  OR2_X1 U10754 ( .A1(n10840), .A2(n10841), .ZN(n10921) );
  AND2_X1 U10755 ( .A1(n10924), .A2(n10925), .ZN(n10841) );
  NAND2_X1 U10756 ( .A1(n10926), .A2(b_24_), .ZN(n10925) );
  NOR2_X1 U10757 ( .A1(n10927), .A2(n8959), .ZN(n10926) );
  NOR2_X1 U10758 ( .A1(n10836), .A2(n10837), .ZN(n10927) );
  NAND2_X1 U10759 ( .A1(n10836), .A2(n10837), .ZN(n10924) );
  NAND2_X1 U10760 ( .A1(n10928), .A2(n10929), .ZN(n10837) );
  NAND2_X1 U10761 ( .A1(n10930), .A2(b_24_), .ZN(n10929) );
  NOR2_X1 U10762 ( .A1(n10931), .A2(n8550), .ZN(n10930) );
  NOR2_X1 U10763 ( .A1(n10832), .A2(n10833), .ZN(n10931) );
  NAND2_X1 U10764 ( .A1(n10832), .A2(n10833), .ZN(n10928) );
  NAND2_X1 U10765 ( .A1(n10932), .A2(n10933), .ZN(n10833) );
  NAND2_X1 U10766 ( .A1(n10934), .A2(b_24_), .ZN(n10933) );
  NOR2_X1 U10767 ( .A1(n10935), .A2(n8956), .ZN(n10934) );
  NOR2_X1 U10768 ( .A1(n10828), .A2(n10829), .ZN(n10935) );
  NAND2_X1 U10769 ( .A1(n10828), .A2(n10829), .ZN(n10932) );
  NAND2_X1 U10770 ( .A1(n10936), .A2(n10937), .ZN(n10829) );
  NAND2_X1 U10771 ( .A1(n10826), .A2(n10938), .ZN(n10937) );
  NAND2_X1 U10772 ( .A1(n10825), .A2(n10824), .ZN(n10938) );
  NOR2_X1 U10773 ( .A1(n8185), .A2(n8495), .ZN(n10826) );
  OR2_X1 U10774 ( .A1(n10824), .A2(n10825), .ZN(n10936) );
  AND2_X1 U10775 ( .A1(n10939), .A2(n10940), .ZN(n10825) );
  NAND2_X1 U10776 ( .A1(n10941), .A2(b_24_), .ZN(n10940) );
  NOR2_X1 U10777 ( .A1(n10942), .A2(n8953), .ZN(n10941) );
  NOR2_X1 U10778 ( .A1(n10820), .A2(n10821), .ZN(n10942) );
  NAND2_X1 U10779 ( .A1(n10820), .A2(n10821), .ZN(n10939) );
  NAND2_X1 U10780 ( .A1(n10943), .A2(n10944), .ZN(n10821) );
  NAND2_X1 U10781 ( .A1(n10818), .A2(n10945), .ZN(n10944) );
  OR2_X1 U10782 ( .A1(n10817), .A2(n10816), .ZN(n10945) );
  NOR2_X1 U10783 ( .A1(n8185), .A2(n8440), .ZN(n10818) );
  NAND2_X1 U10784 ( .A1(n10816), .A2(n10817), .ZN(n10943) );
  NAND2_X1 U10785 ( .A1(n10946), .A2(n10947), .ZN(n10817) );
  NAND2_X1 U10786 ( .A1(n10948), .A2(b_24_), .ZN(n10947) );
  NOR2_X1 U10787 ( .A1(n10949), .A2(n8950), .ZN(n10948) );
  NOR2_X1 U10788 ( .A1(n10811), .A2(n10813), .ZN(n10949) );
  NAND2_X1 U10789 ( .A1(n10811), .A2(n10813), .ZN(n10946) );
  NAND2_X1 U10790 ( .A1(n10950), .A2(n10951), .ZN(n10813) );
  NAND2_X1 U10791 ( .A1(n10810), .A2(n10952), .ZN(n10951) );
  OR2_X1 U10792 ( .A1(n10809), .A2(n10808), .ZN(n10952) );
  NOR2_X1 U10793 ( .A1(n8185), .A2(n8385), .ZN(n10810) );
  NAND2_X1 U10794 ( .A1(n10808), .A2(n10809), .ZN(n10950) );
  NAND2_X1 U10795 ( .A1(n10953), .A2(n10954), .ZN(n10809) );
  NAND2_X1 U10796 ( .A1(n10955), .A2(b_24_), .ZN(n10954) );
  NOR2_X1 U10797 ( .A1(n10956), .A2(n8947), .ZN(n10955) );
  NOR2_X1 U10798 ( .A1(n10804), .A2(n10805), .ZN(n10956) );
  NAND2_X1 U10799 ( .A1(n10804), .A2(n10805), .ZN(n10953) );
  NAND2_X1 U10800 ( .A1(n10957), .A2(n10958), .ZN(n10805) );
  NAND2_X1 U10801 ( .A1(n10802), .A2(n10959), .ZN(n10958) );
  OR2_X1 U10802 ( .A1(n10801), .A2(n10799), .ZN(n10959) );
  NOR2_X1 U10803 ( .A1(n8185), .A2(n8324), .ZN(n10802) );
  NAND2_X1 U10804 ( .A1(n10799), .A2(n10801), .ZN(n10957) );
  NAND2_X1 U10805 ( .A1(n10960), .A2(n10961), .ZN(n10801) );
  NAND2_X1 U10806 ( .A1(n10962), .A2(b_24_), .ZN(n10961) );
  NOR2_X1 U10807 ( .A1(n10963), .A2(n8944), .ZN(n10962) );
  NOR2_X1 U10808 ( .A1(n10796), .A2(n10797), .ZN(n10963) );
  NAND2_X1 U10809 ( .A1(n10796), .A2(n10797), .ZN(n10960) );
  NAND2_X1 U10810 ( .A1(n10964), .A2(n10965), .ZN(n10797) );
  NAND2_X1 U10811 ( .A1(n10794), .A2(n10966), .ZN(n10965) );
  OR2_X1 U10812 ( .A1(n10793), .A2(n10791), .ZN(n10966) );
  NOR2_X1 U10813 ( .A1(n8185), .A2(n8268), .ZN(n10794) );
  NAND2_X1 U10814 ( .A1(n10791), .A2(n10793), .ZN(n10964) );
  NAND2_X1 U10815 ( .A1(n10967), .A2(n10968), .ZN(n10793) );
  NAND2_X1 U10816 ( .A1(n10969), .A2(b_24_), .ZN(n10968) );
  NOR2_X1 U10817 ( .A1(n10970), .A2(n8941), .ZN(n10969) );
  NOR2_X1 U10818 ( .A1(n10788), .A2(n10789), .ZN(n10970) );
  NAND2_X1 U10819 ( .A1(n10788), .A2(n10789), .ZN(n10967) );
  NAND2_X1 U10820 ( .A1(n10971), .A2(n10972), .ZN(n10789) );
  NAND2_X1 U10821 ( .A1(n10786), .A2(n10973), .ZN(n10972) );
  OR2_X1 U10822 ( .A1(n10785), .A2(n10783), .ZN(n10973) );
  NOR2_X1 U10823 ( .A1(n8185), .A2(n8213), .ZN(n10786) );
  NAND2_X1 U10824 ( .A1(n10783), .A2(n10785), .ZN(n10971) );
  NAND2_X1 U10825 ( .A1(n10974), .A2(n10975), .ZN(n10785) );
  NAND2_X1 U10826 ( .A1(n10780), .A2(n10976), .ZN(n10975) );
  OR2_X1 U10827 ( .A1(n10781), .A2(n10782), .ZN(n10976) );
  XNOR2_X1 U10828 ( .A(n10977), .B(n10978), .ZN(n10780) );
  XNOR2_X1 U10829 ( .A(n10979), .B(n10980), .ZN(n10978) );
  NAND2_X1 U10830 ( .A1(n10782), .A2(n10781), .ZN(n10974) );
  NAND2_X1 U10831 ( .A1(n10981), .A2(n10982), .ZN(n10781) );
  NAND2_X1 U10832 ( .A1(n10778), .A2(n10983), .ZN(n10982) );
  OR2_X1 U10833 ( .A1(n10777), .A2(n10775), .ZN(n10983) );
  NOR2_X1 U10834 ( .A1(n8185), .A2(n8158), .ZN(n10778) );
  NAND2_X1 U10835 ( .A1(n10775), .A2(n10777), .ZN(n10981) );
  NAND2_X1 U10836 ( .A1(n10773), .A2(n10984), .ZN(n10777) );
  NAND2_X1 U10837 ( .A1(n10772), .A2(n10774), .ZN(n10984) );
  NAND2_X1 U10838 ( .A1(n10985), .A2(n10986), .ZN(n10774) );
  NAND2_X1 U10839 ( .A1(b_24_), .A2(a_26_), .ZN(n10986) );
  INV_X1 U10840 ( .A(n10987), .ZN(n10985) );
  XNOR2_X1 U10841 ( .A(n10988), .B(n10989), .ZN(n10772) );
  NAND2_X1 U10842 ( .A1(n10990), .A2(n10991), .ZN(n10988) );
  NAND2_X1 U10843 ( .A1(a_26_), .A2(n10987), .ZN(n10773) );
  NAND2_X1 U10844 ( .A1(n10743), .A2(n10992), .ZN(n10987) );
  NAND2_X1 U10845 ( .A1(n10742), .A2(n10744), .ZN(n10992) );
  NAND2_X1 U10846 ( .A1(n10993), .A2(n10994), .ZN(n10744) );
  NAND2_X1 U10847 ( .A1(b_24_), .A2(a_27_), .ZN(n10994) );
  INV_X1 U10848 ( .A(n10995), .ZN(n10993) );
  XOR2_X1 U10849 ( .A(n10996), .B(n10997), .Z(n10742) );
  XNOR2_X1 U10850 ( .A(n10998), .B(n10999), .ZN(n10996) );
  NAND2_X1 U10851 ( .A1(b_23_), .A2(a_28_), .ZN(n10998) );
  NAND2_X1 U10852 ( .A1(a_27_), .A2(n10995), .ZN(n10743) );
  NAND2_X1 U10853 ( .A1(n11000), .A2(n11001), .ZN(n10995) );
  NAND2_X1 U10854 ( .A1(n11002), .A2(b_24_), .ZN(n11001) );
  NOR2_X1 U10855 ( .A1(n11003), .A2(n8055), .ZN(n11002) );
  NOR2_X1 U10856 ( .A1(n10750), .A2(n10752), .ZN(n11003) );
  NAND2_X1 U10857 ( .A1(n10750), .A2(n10752), .ZN(n11000) );
  NAND2_X1 U10858 ( .A1(n11004), .A2(n11005), .ZN(n10752) );
  NAND2_X1 U10859 ( .A1(n10768), .A2(n11006), .ZN(n11005) );
  OR2_X1 U10860 ( .A1(n10769), .A2(n10770), .ZN(n11006) );
  NOR2_X1 U10861 ( .A1(n8185), .A2(n8041), .ZN(n10768) );
  NAND2_X1 U10862 ( .A1(n10770), .A2(n10769), .ZN(n11004) );
  NAND2_X1 U10863 ( .A1(n11007), .A2(n11008), .ZN(n10769) );
  NAND2_X1 U10864 ( .A1(b_22_), .A2(n11009), .ZN(n11008) );
  NAND2_X1 U10865 ( .A1(n8003), .A2(n11010), .ZN(n11009) );
  NAND2_X1 U10866 ( .A1(a_31_), .A2(n8940), .ZN(n11010) );
  NAND2_X1 U10867 ( .A1(b_23_), .A2(n11011), .ZN(n11007) );
  NAND2_X1 U10868 ( .A1(n9341), .A2(n11012), .ZN(n11011) );
  NAND2_X1 U10869 ( .A1(a_30_), .A2(n8240), .ZN(n11012) );
  AND2_X1 U10870 ( .A1(n11013), .A2(n7953), .ZN(n10770) );
  NOR2_X1 U10871 ( .A1(n8185), .A2(n8940), .ZN(n11013) );
  XOR2_X1 U10872 ( .A(n11014), .B(n11015), .Z(n10750) );
  XOR2_X1 U10873 ( .A(n11016), .B(n11017), .Z(n11014) );
  XNOR2_X1 U10874 ( .A(n11018), .B(n11019), .ZN(n10775) );
  NAND2_X1 U10875 ( .A1(n11020), .A2(n11021), .ZN(n11018) );
  INV_X1 U10876 ( .A(n8914), .ZN(n10782) );
  NAND2_X1 U10877 ( .A1(b_24_), .A2(a_24_), .ZN(n8914) );
  XOR2_X1 U10878 ( .A(n11022), .B(n11023), .Z(n10783) );
  XOR2_X1 U10879 ( .A(n11024), .B(n11025), .Z(n11022) );
  NOR2_X1 U10880 ( .A1(n8939), .A2(n8940), .ZN(n11025) );
  XNOR2_X1 U10881 ( .A(n11026), .B(n11027), .ZN(n10788) );
  XNOR2_X1 U10882 ( .A(n11028), .B(n8911), .ZN(n11027) );
  XOR2_X1 U10883 ( .A(n11029), .B(n11030), .Z(n10791) );
  XOR2_X1 U10884 ( .A(n11031), .B(n11032), .Z(n11029) );
  NOR2_X1 U10885 ( .A1(n8941), .A2(n8940), .ZN(n11032) );
  XNOR2_X1 U10886 ( .A(n11033), .B(n11034), .ZN(n10796) );
  XNOR2_X1 U10887 ( .A(n11035), .B(n11036), .ZN(n11034) );
  XOR2_X1 U10888 ( .A(n11037), .B(n11038), .Z(n10799) );
  XOR2_X1 U10889 ( .A(n11039), .B(n11040), .Z(n11037) );
  NOR2_X1 U10890 ( .A1(n8944), .A2(n8940), .ZN(n11040) );
  XOR2_X1 U10891 ( .A(n11041), .B(n11042), .Z(n10804) );
  XOR2_X1 U10892 ( .A(n11043), .B(n11044), .Z(n11041) );
  XNOR2_X1 U10893 ( .A(n11045), .B(n11046), .ZN(n10808) );
  XOR2_X1 U10894 ( .A(n11047), .B(n11048), .Z(n11046) );
  NAND2_X1 U10895 ( .A1(b_23_), .A2(a_18_), .ZN(n11048) );
  XNOR2_X1 U10896 ( .A(n11049), .B(n11050), .ZN(n10811) );
  XNOR2_X1 U10897 ( .A(n11051), .B(n11052), .ZN(n11049) );
  XOR2_X1 U10898 ( .A(n11053), .B(n11054), .Z(n10816) );
  XOR2_X1 U10899 ( .A(n11055), .B(n11056), .Z(n11053) );
  NOR2_X1 U10900 ( .A1(n8950), .A2(n8940), .ZN(n11056) );
  XOR2_X1 U10901 ( .A(n11057), .B(n11058), .Z(n10820) );
  XOR2_X1 U10902 ( .A(n11059), .B(n11060), .Z(n11057) );
  NOR2_X1 U10903 ( .A1(n8440), .A2(n8940), .ZN(n11060) );
  XOR2_X1 U10904 ( .A(n11061), .B(n11062), .Z(n10824) );
  NAND2_X1 U10905 ( .A1(n11063), .A2(n11064), .ZN(n11061) );
  XOR2_X1 U10906 ( .A(n11065), .B(n11066), .Z(n10828) );
  XOR2_X1 U10907 ( .A(n11067), .B(n11068), .Z(n11065) );
  XOR2_X1 U10908 ( .A(n11069), .B(n11070), .Z(n10832) );
  XOR2_X1 U10909 ( .A(n11071), .B(n11072), .Z(n11069) );
  NOR2_X1 U10910 ( .A1(n8956), .A2(n8940), .ZN(n11072) );
  XOR2_X1 U10911 ( .A(n11073), .B(n11074), .Z(n10836) );
  XOR2_X1 U10912 ( .A(n11075), .B(n11076), .Z(n11073) );
  NOR2_X1 U10913 ( .A1(n8550), .A2(n8940), .ZN(n11076) );
  XOR2_X1 U10914 ( .A(n11077), .B(n11078), .Z(n10840) );
  NAND2_X1 U10915 ( .A1(n11079), .A2(n11080), .ZN(n11077) );
  XNOR2_X1 U10916 ( .A(n11081), .B(n11082), .ZN(n10670) );
  XNOR2_X1 U10917 ( .A(n11083), .B(n11084), .ZN(n11082) );
  OR2_X1 U10918 ( .A1(n10850), .A2(n10848), .ZN(n10906) );
  XOR2_X1 U10919 ( .A(n11085), .B(n11086), .Z(n10848) );
  XOR2_X1 U10920 ( .A(n11087), .B(n11088), .Z(n11086) );
  NAND2_X1 U10921 ( .A1(b_23_), .A2(a_7_), .ZN(n11088) );
  NAND2_X1 U10922 ( .A1(b_24_), .A2(a_6_), .ZN(n10850) );
  XOR2_X1 U10923 ( .A(n11089), .B(n11090), .Z(n10852) );
  NAND2_X1 U10924 ( .A1(n11091), .A2(n11092), .ZN(n11089) );
  XOR2_X1 U10925 ( .A(n11093), .B(n11094), .Z(n10856) );
  XOR2_X1 U10926 ( .A(n11095), .B(n11096), .Z(n11093) );
  NOR2_X1 U10927 ( .A1(n8723), .A2(n8940), .ZN(n11096) );
  NAND2_X1 U10928 ( .A1(n10866), .A2(n10864), .ZN(n10880) );
  XOR2_X1 U10929 ( .A(n11097), .B(n11098), .Z(n10864) );
  XOR2_X1 U10930 ( .A(n11099), .B(n11100), .Z(n11097) );
  NOR2_X1 U10931 ( .A1(n8792), .A2(n8940), .ZN(n11100) );
  NOR2_X1 U10932 ( .A1(n8185), .A2(n8969), .ZN(n10866) );
  XOR2_X1 U10933 ( .A(n11101), .B(n11102), .Z(n10630) );
  XOR2_X1 U10934 ( .A(n11103), .B(n11104), .Z(n11101) );
  NOR2_X1 U10935 ( .A1(n8969), .A2(n8940), .ZN(n11104) );
  NAND2_X1 U10936 ( .A1(n11105), .A2(n11106), .ZN(n9037) );
  AND2_X1 U10937 ( .A1(n11107), .A2(n9177), .ZN(n11106) );
  NAND2_X1 U10938 ( .A1(n11108), .A2(n11109), .ZN(n9177) );
  NAND2_X1 U10939 ( .A1(n11110), .A2(b_23_), .ZN(n11109) );
  NOR2_X1 U10940 ( .A1(n11111), .A2(n8974), .ZN(n11110) );
  NOR2_X1 U10941 ( .A1(n10873), .A2(n10874), .ZN(n11111) );
  NAND2_X1 U10942 ( .A1(n10873), .A2(n10874), .ZN(n11108) );
  NAND2_X1 U10943 ( .A1(n11112), .A2(n11113), .ZN(n10874) );
  NAND2_X1 U10944 ( .A1(n11114), .A2(b_23_), .ZN(n11113) );
  NOR2_X1 U10945 ( .A1(n11115), .A2(n8969), .ZN(n11114) );
  NOR2_X1 U10946 ( .A1(n11102), .A2(n11103), .ZN(n11115) );
  NAND2_X1 U10947 ( .A1(n11102), .A2(n11103), .ZN(n11112) );
  NAND2_X1 U10948 ( .A1(n11116), .A2(n11117), .ZN(n11103) );
  NAND2_X1 U10949 ( .A1(n11118), .A2(b_23_), .ZN(n11117) );
  NOR2_X1 U10950 ( .A1(n11119), .A2(n8792), .ZN(n11118) );
  NOR2_X1 U10951 ( .A1(n11098), .A2(n11099), .ZN(n11119) );
  NAND2_X1 U10952 ( .A1(n11098), .A2(n11099), .ZN(n11116) );
  NAND2_X1 U10953 ( .A1(n11120), .A2(n11121), .ZN(n11099) );
  NAND2_X1 U10954 ( .A1(n11122), .A2(b_23_), .ZN(n11121) );
  NOR2_X1 U10955 ( .A1(n11123), .A2(n8778), .ZN(n11122) );
  NOR2_X1 U10956 ( .A1(n10887), .A2(n10889), .ZN(n11123) );
  NAND2_X1 U10957 ( .A1(n10887), .A2(n10889), .ZN(n11120) );
  NAND2_X1 U10958 ( .A1(n11124), .A2(n11125), .ZN(n10889) );
  NAND2_X1 U10959 ( .A1(n11126), .A2(b_23_), .ZN(n11125) );
  NOR2_X1 U10960 ( .A1(n11127), .A2(n8966), .ZN(n11126) );
  NOR2_X1 U10961 ( .A1(n10896), .A2(n10897), .ZN(n11127) );
  NAND2_X1 U10962 ( .A1(n10896), .A2(n10897), .ZN(n11124) );
  NAND2_X1 U10963 ( .A1(n11128), .A2(n11129), .ZN(n10897) );
  NAND2_X1 U10964 ( .A1(n11130), .A2(b_23_), .ZN(n11129) );
  NOR2_X1 U10965 ( .A1(n11131), .A2(n8723), .ZN(n11130) );
  NOR2_X1 U10966 ( .A1(n11094), .A2(n11095), .ZN(n11131) );
  NAND2_X1 U10967 ( .A1(n11094), .A2(n11095), .ZN(n11128) );
  NAND2_X1 U10968 ( .A1(n11091), .A2(n11132), .ZN(n11095) );
  NAND2_X1 U10969 ( .A1(n11090), .A2(n11092), .ZN(n11132) );
  NAND2_X1 U10970 ( .A1(n11133), .A2(n11134), .ZN(n11092) );
  NAND2_X1 U10971 ( .A1(b_23_), .A2(a_6_), .ZN(n11134) );
  INV_X1 U10972 ( .A(n11135), .ZN(n11133) );
  XNOR2_X1 U10973 ( .A(n11136), .B(n11137), .ZN(n11090) );
  XNOR2_X1 U10974 ( .A(n11138), .B(n11139), .ZN(n11137) );
  NAND2_X1 U10975 ( .A1(a_6_), .A2(n11135), .ZN(n11091) );
  NAND2_X1 U10976 ( .A1(n11140), .A2(n11141), .ZN(n11135) );
  NAND2_X1 U10977 ( .A1(n11142), .A2(b_23_), .ZN(n11141) );
  NOR2_X1 U10978 ( .A1(n11143), .A2(n8962), .ZN(n11142) );
  NOR2_X1 U10979 ( .A1(n11085), .A2(n11087), .ZN(n11143) );
  NAND2_X1 U10980 ( .A1(n11085), .A2(n11087), .ZN(n11140) );
  NAND2_X1 U10981 ( .A1(n11144), .A2(n11145), .ZN(n11087) );
  NAND2_X1 U10982 ( .A1(n10916), .A2(n11146), .ZN(n11145) );
  OR2_X1 U10983 ( .A1(n10915), .A2(n10913), .ZN(n11146) );
  NOR2_X1 U10984 ( .A1(n8940), .A2(n8619), .ZN(n10916) );
  NAND2_X1 U10985 ( .A1(n10913), .A2(n10915), .ZN(n11144) );
  NAND2_X1 U10986 ( .A1(n11147), .A2(n11148), .ZN(n10915) );
  NAND2_X1 U10987 ( .A1(n11084), .A2(n11149), .ZN(n11148) );
  OR2_X1 U10988 ( .A1(n11083), .A2(n11081), .ZN(n11149) );
  NOR2_X1 U10989 ( .A1(n8940), .A2(n8605), .ZN(n11084) );
  NAND2_X1 U10990 ( .A1(n11081), .A2(n11083), .ZN(n11147) );
  NAND2_X1 U10991 ( .A1(n11079), .A2(n11150), .ZN(n11083) );
  NAND2_X1 U10992 ( .A1(n11078), .A2(n11080), .ZN(n11150) );
  NAND2_X1 U10993 ( .A1(n11151), .A2(n11152), .ZN(n11080) );
  NAND2_X1 U10994 ( .A1(b_23_), .A2(a_10_), .ZN(n11152) );
  INV_X1 U10995 ( .A(n11153), .ZN(n11151) );
  XOR2_X1 U10996 ( .A(n11154), .B(n11155), .Z(n11078) );
  XOR2_X1 U10997 ( .A(n11156), .B(n11157), .Z(n11154) );
  NAND2_X1 U10998 ( .A1(a_10_), .A2(n11153), .ZN(n11079) );
  NAND2_X1 U10999 ( .A1(n11158), .A2(n11159), .ZN(n11153) );
  NAND2_X1 U11000 ( .A1(n11160), .A2(b_23_), .ZN(n11159) );
  NOR2_X1 U11001 ( .A1(n11161), .A2(n8550), .ZN(n11160) );
  NOR2_X1 U11002 ( .A1(n11074), .A2(n11075), .ZN(n11161) );
  NAND2_X1 U11003 ( .A1(n11074), .A2(n11075), .ZN(n11158) );
  NAND2_X1 U11004 ( .A1(n11162), .A2(n11163), .ZN(n11075) );
  NAND2_X1 U11005 ( .A1(n11164), .A2(b_23_), .ZN(n11163) );
  NOR2_X1 U11006 ( .A1(n11165), .A2(n8956), .ZN(n11164) );
  NOR2_X1 U11007 ( .A1(n11070), .A2(n11071), .ZN(n11165) );
  NAND2_X1 U11008 ( .A1(n11070), .A2(n11071), .ZN(n11162) );
  NAND2_X1 U11009 ( .A1(n11166), .A2(n11167), .ZN(n11071) );
  NAND2_X1 U11010 ( .A1(n11068), .A2(n11168), .ZN(n11167) );
  OR2_X1 U11011 ( .A1(n11067), .A2(n11066), .ZN(n11168) );
  NOR2_X1 U11012 ( .A1(n8940), .A2(n8495), .ZN(n11068) );
  NAND2_X1 U11013 ( .A1(n11066), .A2(n11067), .ZN(n11166) );
  NAND2_X1 U11014 ( .A1(n11063), .A2(n11169), .ZN(n11067) );
  NAND2_X1 U11015 ( .A1(n11062), .A2(n11064), .ZN(n11169) );
  NAND2_X1 U11016 ( .A1(n11170), .A2(n11171), .ZN(n11064) );
  NAND2_X1 U11017 ( .A1(b_23_), .A2(a_14_), .ZN(n11171) );
  INV_X1 U11018 ( .A(n11172), .ZN(n11170) );
  XOR2_X1 U11019 ( .A(n11173), .B(n11174), .Z(n11062) );
  XOR2_X1 U11020 ( .A(n11175), .B(n11176), .Z(n11173) );
  NAND2_X1 U11021 ( .A1(a_14_), .A2(n11172), .ZN(n11063) );
  NAND2_X1 U11022 ( .A1(n11177), .A2(n11178), .ZN(n11172) );
  NAND2_X1 U11023 ( .A1(n11179), .A2(b_23_), .ZN(n11178) );
  NOR2_X1 U11024 ( .A1(n11180), .A2(n8440), .ZN(n11179) );
  NOR2_X1 U11025 ( .A1(n11058), .A2(n11059), .ZN(n11180) );
  NAND2_X1 U11026 ( .A1(n11058), .A2(n11059), .ZN(n11177) );
  NAND2_X1 U11027 ( .A1(n11181), .A2(n11182), .ZN(n11059) );
  NAND2_X1 U11028 ( .A1(n11183), .A2(b_23_), .ZN(n11182) );
  NOR2_X1 U11029 ( .A1(n11184), .A2(n8950), .ZN(n11183) );
  NOR2_X1 U11030 ( .A1(n11054), .A2(n11055), .ZN(n11184) );
  NAND2_X1 U11031 ( .A1(n11054), .A2(n11055), .ZN(n11181) );
  NAND2_X1 U11032 ( .A1(n11185), .A2(n11186), .ZN(n11055) );
  NAND2_X1 U11033 ( .A1(n11052), .A2(n11187), .ZN(n11186) );
  NAND2_X1 U11034 ( .A1(n11051), .A2(n11050), .ZN(n11187) );
  NOR2_X1 U11035 ( .A1(n8940), .A2(n8385), .ZN(n11052) );
  OR2_X1 U11036 ( .A1(n11050), .A2(n11051), .ZN(n11185) );
  AND2_X1 U11037 ( .A1(n11188), .A2(n11189), .ZN(n11051) );
  NAND2_X1 U11038 ( .A1(n11190), .A2(b_23_), .ZN(n11189) );
  NOR2_X1 U11039 ( .A1(n11191), .A2(n8947), .ZN(n11190) );
  NOR2_X1 U11040 ( .A1(n11045), .A2(n11047), .ZN(n11191) );
  NAND2_X1 U11041 ( .A1(n11045), .A2(n11047), .ZN(n11188) );
  NAND2_X1 U11042 ( .A1(n11192), .A2(n11193), .ZN(n11047) );
  NAND2_X1 U11043 ( .A1(n11044), .A2(n11194), .ZN(n11193) );
  OR2_X1 U11044 ( .A1(n11043), .A2(n11042), .ZN(n11194) );
  NOR2_X1 U11045 ( .A1(n8940), .A2(n8324), .ZN(n11044) );
  NAND2_X1 U11046 ( .A1(n11042), .A2(n11043), .ZN(n11192) );
  NAND2_X1 U11047 ( .A1(n11195), .A2(n11196), .ZN(n11043) );
  NAND2_X1 U11048 ( .A1(n11197), .A2(b_23_), .ZN(n11196) );
  NOR2_X1 U11049 ( .A1(n11198), .A2(n8944), .ZN(n11197) );
  NOR2_X1 U11050 ( .A1(n11038), .A2(n11039), .ZN(n11198) );
  NAND2_X1 U11051 ( .A1(n11038), .A2(n11039), .ZN(n11195) );
  NAND2_X1 U11052 ( .A1(n11199), .A2(n11200), .ZN(n11039) );
  NAND2_X1 U11053 ( .A1(n11036), .A2(n11201), .ZN(n11200) );
  OR2_X1 U11054 ( .A1(n11035), .A2(n11033), .ZN(n11201) );
  NOR2_X1 U11055 ( .A1(n8940), .A2(n8268), .ZN(n11036) );
  NAND2_X1 U11056 ( .A1(n11033), .A2(n11035), .ZN(n11199) );
  NAND2_X1 U11057 ( .A1(n11202), .A2(n11203), .ZN(n11035) );
  NAND2_X1 U11058 ( .A1(n11204), .A2(b_23_), .ZN(n11203) );
  NOR2_X1 U11059 ( .A1(n11205), .A2(n8941), .ZN(n11204) );
  NOR2_X1 U11060 ( .A1(n11030), .A2(n11031), .ZN(n11205) );
  NAND2_X1 U11061 ( .A1(n11030), .A2(n11031), .ZN(n11202) );
  NAND2_X1 U11062 ( .A1(n11206), .A2(n11207), .ZN(n11031) );
  NAND2_X1 U11063 ( .A1(n8911), .A2(n11208), .ZN(n11207) );
  OR2_X1 U11064 ( .A1(n11028), .A2(n11026), .ZN(n11208) );
  NOR2_X1 U11065 ( .A1(n8940), .A2(n8213), .ZN(n8911) );
  NAND2_X1 U11066 ( .A1(n11026), .A2(n11028), .ZN(n11206) );
  NAND2_X1 U11067 ( .A1(n11209), .A2(n11210), .ZN(n11028) );
  NAND2_X1 U11068 ( .A1(n11211), .A2(b_23_), .ZN(n11210) );
  NOR2_X1 U11069 ( .A1(n11212), .A2(n8939), .ZN(n11211) );
  NOR2_X1 U11070 ( .A1(n11023), .A2(n11024), .ZN(n11212) );
  NAND2_X1 U11071 ( .A1(n11023), .A2(n11024), .ZN(n11209) );
  NAND2_X1 U11072 ( .A1(n11213), .A2(n11214), .ZN(n11024) );
  NAND2_X1 U11073 ( .A1(n10980), .A2(n11215), .ZN(n11214) );
  OR2_X1 U11074 ( .A1(n10979), .A2(n10977), .ZN(n11215) );
  NOR2_X1 U11075 ( .A1(n8940), .A2(n8158), .ZN(n10980) );
  NAND2_X1 U11076 ( .A1(n10977), .A2(n10979), .ZN(n11213) );
  NAND2_X1 U11077 ( .A1(n11020), .A2(n11216), .ZN(n10979) );
  NAND2_X1 U11078 ( .A1(n11019), .A2(n11021), .ZN(n11216) );
  NAND2_X1 U11079 ( .A1(n11217), .A2(n11218), .ZN(n11021) );
  NAND2_X1 U11080 ( .A1(b_23_), .A2(a_26_), .ZN(n11218) );
  INV_X1 U11081 ( .A(n11219), .ZN(n11217) );
  XNOR2_X1 U11082 ( .A(n11220), .B(n11221), .ZN(n11019) );
  NAND2_X1 U11083 ( .A1(n11222), .A2(n11223), .ZN(n11220) );
  NAND2_X1 U11084 ( .A1(a_26_), .A2(n11219), .ZN(n11020) );
  NAND2_X1 U11085 ( .A1(n10990), .A2(n11224), .ZN(n11219) );
  NAND2_X1 U11086 ( .A1(n10989), .A2(n10991), .ZN(n11224) );
  NAND2_X1 U11087 ( .A1(n11225), .A2(n11226), .ZN(n10991) );
  NAND2_X1 U11088 ( .A1(b_23_), .A2(a_27_), .ZN(n11226) );
  INV_X1 U11089 ( .A(n11227), .ZN(n11225) );
  XOR2_X1 U11090 ( .A(n11228), .B(n11229), .Z(n10989) );
  XNOR2_X1 U11091 ( .A(n11230), .B(n11231), .ZN(n11228) );
  NAND2_X1 U11092 ( .A1(b_22_), .A2(a_28_), .ZN(n11230) );
  NAND2_X1 U11093 ( .A1(a_27_), .A2(n11227), .ZN(n10990) );
  NAND2_X1 U11094 ( .A1(n11232), .A2(n11233), .ZN(n11227) );
  NAND2_X1 U11095 ( .A1(n11234), .A2(b_23_), .ZN(n11233) );
  NOR2_X1 U11096 ( .A1(n11235), .A2(n8055), .ZN(n11234) );
  NOR2_X1 U11097 ( .A1(n10997), .A2(n10999), .ZN(n11235) );
  NAND2_X1 U11098 ( .A1(n10997), .A2(n10999), .ZN(n11232) );
  NAND2_X1 U11099 ( .A1(n11236), .A2(n11237), .ZN(n10999) );
  NAND2_X1 U11100 ( .A1(n11015), .A2(n11238), .ZN(n11237) );
  OR2_X1 U11101 ( .A1(n11016), .A2(n11017), .ZN(n11238) );
  NOR2_X1 U11102 ( .A1(n8940), .A2(n8041), .ZN(n11015) );
  NAND2_X1 U11103 ( .A1(n11017), .A2(n11016), .ZN(n11236) );
  NAND2_X1 U11104 ( .A1(n11239), .A2(n11240), .ZN(n11016) );
  NAND2_X1 U11105 ( .A1(b_21_), .A2(n11241), .ZN(n11240) );
  NAND2_X1 U11106 ( .A1(n8003), .A2(n11242), .ZN(n11241) );
  NAND2_X1 U11107 ( .A1(a_31_), .A2(n8240), .ZN(n11242) );
  NAND2_X1 U11108 ( .A1(b_22_), .A2(n11243), .ZN(n11239) );
  NAND2_X1 U11109 ( .A1(n9341), .A2(n11244), .ZN(n11243) );
  NAND2_X1 U11110 ( .A1(a_30_), .A2(n8942), .ZN(n11244) );
  AND2_X1 U11111 ( .A1(n11245), .A2(n7953), .ZN(n11017) );
  NOR2_X1 U11112 ( .A1(n8940), .A2(n8240), .ZN(n11245) );
  XOR2_X1 U11113 ( .A(n11246), .B(n11247), .Z(n10997) );
  XOR2_X1 U11114 ( .A(n11248), .B(n11249), .Z(n11246) );
  XNOR2_X1 U11115 ( .A(n11250), .B(n11251), .ZN(n10977) );
  NAND2_X1 U11116 ( .A1(n11252), .A2(n11253), .ZN(n11250) );
  XNOR2_X1 U11117 ( .A(n11254), .B(n11255), .ZN(n11023) );
  XNOR2_X1 U11118 ( .A(n11256), .B(n11257), .ZN(n11255) );
  XOR2_X1 U11119 ( .A(n11258), .B(n11259), .Z(n11026) );
  XOR2_X1 U11120 ( .A(n11260), .B(n11261), .Z(n11258) );
  NOR2_X1 U11121 ( .A1(n8939), .A2(n8240), .ZN(n11261) );
  XNOR2_X1 U11122 ( .A(n11262), .B(n11263), .ZN(n11030) );
  XNOR2_X1 U11123 ( .A(n11264), .B(n11265), .ZN(n11263) );
  XOR2_X1 U11124 ( .A(n11266), .B(n11267), .Z(n11033) );
  XOR2_X1 U11125 ( .A(n11268), .B(n11269), .Z(n11266) );
  XNOR2_X1 U11126 ( .A(n11270), .B(n11271), .ZN(n11038) );
  XNOR2_X1 U11127 ( .A(n11272), .B(n11273), .ZN(n11271) );
  XOR2_X1 U11128 ( .A(n11274), .B(n11275), .Z(n11042) );
  XOR2_X1 U11129 ( .A(n11276), .B(n11277), .Z(n11274) );
  NOR2_X1 U11130 ( .A1(n8944), .A2(n8240), .ZN(n11277) );
  XNOR2_X1 U11131 ( .A(n11278), .B(n11279), .ZN(n11045) );
  XNOR2_X1 U11132 ( .A(n11280), .B(n11281), .ZN(n11279) );
  XNOR2_X1 U11133 ( .A(n11282), .B(n11283), .ZN(n11050) );
  XOR2_X1 U11134 ( .A(n11284), .B(n11285), .Z(n11282) );
  NOR2_X1 U11135 ( .A1(n8947), .A2(n8240), .ZN(n11285) );
  XOR2_X1 U11136 ( .A(n11286), .B(n11287), .Z(n11054) );
  XOR2_X1 U11137 ( .A(n11288), .B(n11289), .Z(n11286) );
  XOR2_X1 U11138 ( .A(n11290), .B(n11291), .Z(n11058) );
  XOR2_X1 U11139 ( .A(n11292), .B(n11293), .Z(n11290) );
  NOR2_X1 U11140 ( .A1(n8950), .A2(n8240), .ZN(n11293) );
  XNOR2_X1 U11141 ( .A(n11294), .B(n11295), .ZN(n11066) );
  XOR2_X1 U11142 ( .A(n11296), .B(n11297), .Z(n11295) );
  NAND2_X1 U11143 ( .A1(b_22_), .A2(a_14_), .ZN(n11297) );
  XOR2_X1 U11144 ( .A(n11298), .B(n11299), .Z(n11070) );
  XOR2_X1 U11145 ( .A(n11300), .B(n11301), .Z(n11298) );
  XNOR2_X1 U11146 ( .A(n11302), .B(n11303), .ZN(n11074) );
  XOR2_X1 U11147 ( .A(n11304), .B(n11305), .Z(n11303) );
  NAND2_X1 U11148 ( .A1(b_22_), .A2(a_12_), .ZN(n11305) );
  XOR2_X1 U11149 ( .A(n11306), .B(n11307), .Z(n11081) );
  XOR2_X1 U11150 ( .A(n11308), .B(n11309), .Z(n11306) );
  NOR2_X1 U11151 ( .A1(n8959), .A2(n8240), .ZN(n11309) );
  XOR2_X1 U11152 ( .A(n11310), .B(n11311), .Z(n10913) );
  XOR2_X1 U11153 ( .A(n11312), .B(n11313), .Z(n11310) );
  NOR2_X1 U11154 ( .A1(n8605), .A2(n8240), .ZN(n11313) );
  XNOR2_X1 U11155 ( .A(n11314), .B(n11315), .ZN(n11085) );
  XNOR2_X1 U11156 ( .A(n11316), .B(n11317), .ZN(n11315) );
  XNOR2_X1 U11157 ( .A(n11318), .B(n11319), .ZN(n11094) );
  XNOR2_X1 U11158 ( .A(n11320), .B(n11321), .ZN(n11319) );
  XNOR2_X1 U11159 ( .A(n11322), .B(n11323), .ZN(n10896) );
  XOR2_X1 U11160 ( .A(n11324), .B(n11325), .Z(n11323) );
  NAND2_X1 U11161 ( .A1(b_22_), .A2(a_5_), .ZN(n11325) );
  XNOR2_X1 U11162 ( .A(n11326), .B(n11327), .ZN(n10887) );
  NAND2_X1 U11163 ( .A1(n11328), .A2(n11329), .ZN(n11326) );
  XOR2_X1 U11164 ( .A(n11330), .B(n11331), .Z(n11098) );
  XOR2_X1 U11165 ( .A(n11332), .B(n11333), .Z(n11330) );
  XNOR2_X1 U11166 ( .A(n11334), .B(n11335), .ZN(n11102) );
  XNOR2_X1 U11167 ( .A(n11336), .B(n11337), .ZN(n11334) );
  XNOR2_X1 U11168 ( .A(n11338), .B(n11339), .ZN(n10873) );
  XOR2_X1 U11169 ( .A(n11340), .B(n11341), .Z(n11339) );
  NAND2_X1 U11170 ( .A1(b_22_), .A2(a_1_), .ZN(n11341) );
  NOR2_X1 U11171 ( .A1(n11342), .A2(n9185), .ZN(n11105) );
  XOR2_X1 U11172 ( .A(n11343), .B(n11344), .Z(n9185) );
  XNOR2_X1 U11173 ( .A(n11345), .B(n11346), .ZN(n11343) );
  NOR2_X1 U11174 ( .A1(n9178), .A2(n9179), .ZN(n11342) );
  NAND2_X1 U11175 ( .A1(n11107), .A2(n11347), .ZN(n9044) );
  NAND2_X1 U11176 ( .A1(n11348), .A2(n9171), .ZN(n11347) );
  NAND2_X1 U11177 ( .A1(n11349), .A2(n11350), .ZN(n9043) );
  INV_X1 U11178 ( .A(n11107), .ZN(n11350) );
  NAND2_X1 U11179 ( .A1(n9178), .A2(n9179), .ZN(n11107) );
  NAND2_X1 U11180 ( .A1(n11351), .A2(n11352), .ZN(n9179) );
  NAND2_X1 U11181 ( .A1(n11346), .A2(n11353), .ZN(n11352) );
  NAND2_X1 U11182 ( .A1(n11345), .A2(n11344), .ZN(n11353) );
  NOR2_X1 U11183 ( .A1(n8240), .A2(n8974), .ZN(n11346) );
  OR2_X1 U11184 ( .A1(n11344), .A2(n11345), .ZN(n11351) );
  AND2_X1 U11185 ( .A1(n11354), .A2(n11355), .ZN(n11345) );
  NAND2_X1 U11186 ( .A1(n11356), .A2(b_22_), .ZN(n11355) );
  NOR2_X1 U11187 ( .A1(n11357), .A2(n8969), .ZN(n11356) );
  NOR2_X1 U11188 ( .A1(n11338), .A2(n11340), .ZN(n11357) );
  NAND2_X1 U11189 ( .A1(n11338), .A2(n11340), .ZN(n11354) );
  NAND2_X1 U11190 ( .A1(n11358), .A2(n11359), .ZN(n11340) );
  NAND2_X1 U11191 ( .A1(n11337), .A2(n11360), .ZN(n11359) );
  NAND2_X1 U11192 ( .A1(n11336), .A2(n11335), .ZN(n11360) );
  NOR2_X1 U11193 ( .A1(n8240), .A2(n8792), .ZN(n11337) );
  OR2_X1 U11194 ( .A1(n11335), .A2(n11336), .ZN(n11358) );
  AND2_X1 U11195 ( .A1(n11361), .A2(n11362), .ZN(n11336) );
  NAND2_X1 U11196 ( .A1(n11333), .A2(n11363), .ZN(n11362) );
  OR2_X1 U11197 ( .A1(n11331), .A2(n11332), .ZN(n11363) );
  NOR2_X1 U11198 ( .A1(n8240), .A2(n8778), .ZN(n11333) );
  NAND2_X1 U11199 ( .A1(n11331), .A2(n11332), .ZN(n11361) );
  NAND2_X1 U11200 ( .A1(n11328), .A2(n11364), .ZN(n11332) );
  NAND2_X1 U11201 ( .A1(n11327), .A2(n11329), .ZN(n11364) );
  NAND2_X1 U11202 ( .A1(n11365), .A2(n11366), .ZN(n11329) );
  NAND2_X1 U11203 ( .A1(b_22_), .A2(a_4_), .ZN(n11366) );
  INV_X1 U11204 ( .A(n11367), .ZN(n11365) );
  XOR2_X1 U11205 ( .A(n11368), .B(n11369), .Z(n11327) );
  XOR2_X1 U11206 ( .A(n11370), .B(n11371), .Z(n11368) );
  NOR2_X1 U11207 ( .A1(n8723), .A2(n8942), .ZN(n11371) );
  NAND2_X1 U11208 ( .A1(a_4_), .A2(n11367), .ZN(n11328) );
  NAND2_X1 U11209 ( .A1(n11372), .A2(n11373), .ZN(n11367) );
  NAND2_X1 U11210 ( .A1(n11374), .A2(b_22_), .ZN(n11373) );
  NOR2_X1 U11211 ( .A1(n11375), .A2(n8723), .ZN(n11374) );
  NOR2_X1 U11212 ( .A1(n11324), .A2(n11322), .ZN(n11375) );
  NAND2_X1 U11213 ( .A1(n11322), .A2(n11324), .ZN(n11372) );
  NAND2_X1 U11214 ( .A1(n11376), .A2(n11377), .ZN(n11324) );
  NAND2_X1 U11215 ( .A1(n11321), .A2(n11378), .ZN(n11377) );
  OR2_X1 U11216 ( .A1(n11320), .A2(n11318), .ZN(n11378) );
  NOR2_X1 U11217 ( .A1(n8240), .A2(n8681), .ZN(n11321) );
  NAND2_X1 U11218 ( .A1(n11318), .A2(n11320), .ZN(n11376) );
  NAND2_X1 U11219 ( .A1(n11379), .A2(n11380), .ZN(n11320) );
  NAND2_X1 U11220 ( .A1(n11139), .A2(n11381), .ZN(n11380) );
  OR2_X1 U11221 ( .A1(n11136), .A2(n11138), .ZN(n11381) );
  NOR2_X1 U11222 ( .A1(n8240), .A2(n8962), .ZN(n11139) );
  NAND2_X1 U11223 ( .A1(n11136), .A2(n11138), .ZN(n11379) );
  NAND2_X1 U11224 ( .A1(n11382), .A2(n11383), .ZN(n11138) );
  NAND2_X1 U11225 ( .A1(n11317), .A2(n11384), .ZN(n11383) );
  OR2_X1 U11226 ( .A1(n11316), .A2(n11314), .ZN(n11384) );
  NOR2_X1 U11227 ( .A1(n8240), .A2(n8619), .ZN(n11317) );
  NAND2_X1 U11228 ( .A1(n11314), .A2(n11316), .ZN(n11382) );
  NAND2_X1 U11229 ( .A1(n11385), .A2(n11386), .ZN(n11316) );
  NAND2_X1 U11230 ( .A1(n11387), .A2(b_22_), .ZN(n11386) );
  NOR2_X1 U11231 ( .A1(n11388), .A2(n8605), .ZN(n11387) );
  NOR2_X1 U11232 ( .A1(n11311), .A2(n11312), .ZN(n11388) );
  NAND2_X1 U11233 ( .A1(n11311), .A2(n11312), .ZN(n11385) );
  NAND2_X1 U11234 ( .A1(n11389), .A2(n11390), .ZN(n11312) );
  NAND2_X1 U11235 ( .A1(n11391), .A2(b_22_), .ZN(n11390) );
  NOR2_X1 U11236 ( .A1(n11392), .A2(n8959), .ZN(n11391) );
  NOR2_X1 U11237 ( .A1(n11307), .A2(n11308), .ZN(n11392) );
  NAND2_X1 U11238 ( .A1(n11307), .A2(n11308), .ZN(n11389) );
  NAND2_X1 U11239 ( .A1(n11393), .A2(n11394), .ZN(n11308) );
  NAND2_X1 U11240 ( .A1(n11157), .A2(n11395), .ZN(n11394) );
  OR2_X1 U11241 ( .A1(n11155), .A2(n11156), .ZN(n11395) );
  NOR2_X1 U11242 ( .A1(n8240), .A2(n8550), .ZN(n11157) );
  NAND2_X1 U11243 ( .A1(n11155), .A2(n11156), .ZN(n11393) );
  NAND2_X1 U11244 ( .A1(n11396), .A2(n11397), .ZN(n11156) );
  NAND2_X1 U11245 ( .A1(n11398), .A2(b_22_), .ZN(n11397) );
  NOR2_X1 U11246 ( .A1(n11399), .A2(n8956), .ZN(n11398) );
  NOR2_X1 U11247 ( .A1(n11302), .A2(n11304), .ZN(n11399) );
  NAND2_X1 U11248 ( .A1(n11302), .A2(n11304), .ZN(n11396) );
  NAND2_X1 U11249 ( .A1(n11400), .A2(n11401), .ZN(n11304) );
  NAND2_X1 U11250 ( .A1(n11301), .A2(n11402), .ZN(n11401) );
  OR2_X1 U11251 ( .A1(n11299), .A2(n11300), .ZN(n11402) );
  NOR2_X1 U11252 ( .A1(n8240), .A2(n8495), .ZN(n11301) );
  NAND2_X1 U11253 ( .A1(n11299), .A2(n11300), .ZN(n11400) );
  NAND2_X1 U11254 ( .A1(n11403), .A2(n11404), .ZN(n11300) );
  NAND2_X1 U11255 ( .A1(n11405), .A2(b_22_), .ZN(n11404) );
  NOR2_X1 U11256 ( .A1(n11406), .A2(n8953), .ZN(n11405) );
  NOR2_X1 U11257 ( .A1(n11294), .A2(n11296), .ZN(n11406) );
  NAND2_X1 U11258 ( .A1(n11294), .A2(n11296), .ZN(n11403) );
  NAND2_X1 U11259 ( .A1(n11407), .A2(n11408), .ZN(n11296) );
  NAND2_X1 U11260 ( .A1(n11176), .A2(n11409), .ZN(n11408) );
  OR2_X1 U11261 ( .A1(n11174), .A2(n11175), .ZN(n11409) );
  NOR2_X1 U11262 ( .A1(n8240), .A2(n8440), .ZN(n11176) );
  NAND2_X1 U11263 ( .A1(n11174), .A2(n11175), .ZN(n11407) );
  NAND2_X1 U11264 ( .A1(n11410), .A2(n11411), .ZN(n11175) );
  NAND2_X1 U11265 ( .A1(n11412), .A2(b_22_), .ZN(n11411) );
  NOR2_X1 U11266 ( .A1(n11413), .A2(n8950), .ZN(n11412) );
  NOR2_X1 U11267 ( .A1(n11291), .A2(n11292), .ZN(n11413) );
  NAND2_X1 U11268 ( .A1(n11291), .A2(n11292), .ZN(n11410) );
  NAND2_X1 U11269 ( .A1(n11414), .A2(n11415), .ZN(n11292) );
  NAND2_X1 U11270 ( .A1(n11289), .A2(n11416), .ZN(n11415) );
  OR2_X1 U11271 ( .A1(n11287), .A2(n11288), .ZN(n11416) );
  NOR2_X1 U11272 ( .A1(n8240), .A2(n8385), .ZN(n11289) );
  NAND2_X1 U11273 ( .A1(n11287), .A2(n11288), .ZN(n11414) );
  NAND2_X1 U11274 ( .A1(n11417), .A2(n11418), .ZN(n11288) );
  NAND2_X1 U11275 ( .A1(n11419), .A2(b_22_), .ZN(n11418) );
  NOR2_X1 U11276 ( .A1(n11420), .A2(n8947), .ZN(n11419) );
  NOR2_X1 U11277 ( .A1(n11284), .A2(n11283), .ZN(n11420) );
  NAND2_X1 U11278 ( .A1(n11283), .A2(n11284), .ZN(n11417) );
  NAND2_X1 U11279 ( .A1(n11421), .A2(n11422), .ZN(n11284) );
  NAND2_X1 U11280 ( .A1(n11281), .A2(n11423), .ZN(n11422) );
  OR2_X1 U11281 ( .A1(n11278), .A2(n11280), .ZN(n11423) );
  NOR2_X1 U11282 ( .A1(n8240), .A2(n8324), .ZN(n11281) );
  NAND2_X1 U11283 ( .A1(n11278), .A2(n11280), .ZN(n11421) );
  NAND2_X1 U11284 ( .A1(n11424), .A2(n11425), .ZN(n11280) );
  NAND2_X1 U11285 ( .A1(n11426), .A2(b_22_), .ZN(n11425) );
  NOR2_X1 U11286 ( .A1(n11427), .A2(n8944), .ZN(n11426) );
  NOR2_X1 U11287 ( .A1(n11275), .A2(n11276), .ZN(n11427) );
  NAND2_X1 U11288 ( .A1(n11275), .A2(n11276), .ZN(n11424) );
  NAND2_X1 U11289 ( .A1(n11428), .A2(n11429), .ZN(n11276) );
  NAND2_X1 U11290 ( .A1(n11273), .A2(n11430), .ZN(n11429) );
  OR2_X1 U11291 ( .A1(n11270), .A2(n11272), .ZN(n11430) );
  NOR2_X1 U11292 ( .A1(n8240), .A2(n8268), .ZN(n11273) );
  NAND2_X1 U11293 ( .A1(n11270), .A2(n11272), .ZN(n11428) );
  NAND2_X1 U11294 ( .A1(n11431), .A2(n11432), .ZN(n11272) );
  NAND2_X1 U11295 ( .A1(n11267), .A2(n11433), .ZN(n11432) );
  OR2_X1 U11296 ( .A1(n11268), .A2(n11269), .ZN(n11433) );
  XNOR2_X1 U11297 ( .A(n11434), .B(n11435), .ZN(n11267) );
  XNOR2_X1 U11298 ( .A(n11436), .B(n11437), .ZN(n11435) );
  NAND2_X1 U11299 ( .A1(n11269), .A2(n11268), .ZN(n11431) );
  NAND2_X1 U11300 ( .A1(n11438), .A2(n11439), .ZN(n11268) );
  NAND2_X1 U11301 ( .A1(n11265), .A2(n11440), .ZN(n11439) );
  OR2_X1 U11302 ( .A1(n11262), .A2(n11264), .ZN(n11440) );
  NOR2_X1 U11303 ( .A1(n8240), .A2(n8213), .ZN(n11265) );
  NAND2_X1 U11304 ( .A1(n11262), .A2(n11264), .ZN(n11438) );
  NAND2_X1 U11305 ( .A1(n11441), .A2(n11442), .ZN(n11264) );
  NAND2_X1 U11306 ( .A1(n11443), .A2(b_22_), .ZN(n11442) );
  NOR2_X1 U11307 ( .A1(n11444), .A2(n8939), .ZN(n11443) );
  NOR2_X1 U11308 ( .A1(n11259), .A2(n11260), .ZN(n11444) );
  NAND2_X1 U11309 ( .A1(n11259), .A2(n11260), .ZN(n11441) );
  NAND2_X1 U11310 ( .A1(n11445), .A2(n11446), .ZN(n11260) );
  NAND2_X1 U11311 ( .A1(n11257), .A2(n11447), .ZN(n11446) );
  OR2_X1 U11312 ( .A1(n11254), .A2(n11256), .ZN(n11447) );
  NOR2_X1 U11313 ( .A1(n8240), .A2(n8158), .ZN(n11257) );
  NAND2_X1 U11314 ( .A1(n11254), .A2(n11256), .ZN(n11445) );
  NAND2_X1 U11315 ( .A1(n11252), .A2(n11448), .ZN(n11256) );
  NAND2_X1 U11316 ( .A1(n11251), .A2(n11253), .ZN(n11448) );
  NAND2_X1 U11317 ( .A1(n11449), .A2(n11450), .ZN(n11253) );
  NAND2_X1 U11318 ( .A1(b_22_), .A2(a_26_), .ZN(n11450) );
  INV_X1 U11319 ( .A(n11451), .ZN(n11449) );
  XNOR2_X1 U11320 ( .A(n11452), .B(n11453), .ZN(n11251) );
  NAND2_X1 U11321 ( .A1(n11454), .A2(n11455), .ZN(n11452) );
  NAND2_X1 U11322 ( .A1(a_26_), .A2(n11451), .ZN(n11252) );
  NAND2_X1 U11323 ( .A1(n11222), .A2(n11456), .ZN(n11451) );
  NAND2_X1 U11324 ( .A1(n11221), .A2(n11223), .ZN(n11456) );
  NAND2_X1 U11325 ( .A1(n11457), .A2(n11458), .ZN(n11223) );
  NAND2_X1 U11326 ( .A1(b_22_), .A2(a_27_), .ZN(n11458) );
  INV_X1 U11327 ( .A(n11459), .ZN(n11457) );
  XOR2_X1 U11328 ( .A(n11460), .B(n11461), .Z(n11221) );
  XNOR2_X1 U11329 ( .A(n11462), .B(n11463), .ZN(n11460) );
  NAND2_X1 U11330 ( .A1(b_21_), .A2(a_28_), .ZN(n11462) );
  NAND2_X1 U11331 ( .A1(a_27_), .A2(n11459), .ZN(n11222) );
  NAND2_X1 U11332 ( .A1(n11464), .A2(n11465), .ZN(n11459) );
  NAND2_X1 U11333 ( .A1(n11466), .A2(b_22_), .ZN(n11465) );
  NOR2_X1 U11334 ( .A1(n11467), .A2(n8055), .ZN(n11466) );
  NOR2_X1 U11335 ( .A1(n11229), .A2(n11231), .ZN(n11467) );
  NAND2_X1 U11336 ( .A1(n11229), .A2(n11231), .ZN(n11464) );
  NAND2_X1 U11337 ( .A1(n11468), .A2(n11469), .ZN(n11231) );
  NAND2_X1 U11338 ( .A1(n11247), .A2(n11470), .ZN(n11469) );
  OR2_X1 U11339 ( .A1(n11248), .A2(n11249), .ZN(n11470) );
  NOR2_X1 U11340 ( .A1(n8240), .A2(n8041), .ZN(n11247) );
  NAND2_X1 U11341 ( .A1(n11249), .A2(n11248), .ZN(n11468) );
  NAND2_X1 U11342 ( .A1(n11471), .A2(n11472), .ZN(n11248) );
  NAND2_X1 U11343 ( .A1(b_20_), .A2(n11473), .ZN(n11472) );
  NAND2_X1 U11344 ( .A1(n8003), .A2(n11474), .ZN(n11473) );
  NAND2_X1 U11345 ( .A1(a_31_), .A2(n8942), .ZN(n11474) );
  NAND2_X1 U11346 ( .A1(b_21_), .A2(n11475), .ZN(n11471) );
  NAND2_X1 U11347 ( .A1(n9341), .A2(n11476), .ZN(n11475) );
  NAND2_X1 U11348 ( .A1(a_30_), .A2(n8943), .ZN(n11476) );
  AND2_X1 U11349 ( .A1(n11477), .A2(n7953), .ZN(n11249) );
  NOR2_X1 U11350 ( .A1(n8240), .A2(n8942), .ZN(n11477) );
  XOR2_X1 U11351 ( .A(n11478), .B(n11479), .Z(n11229) );
  XOR2_X1 U11352 ( .A(n11480), .B(n11481), .Z(n11478) );
  XNOR2_X1 U11353 ( .A(n11482), .B(n11483), .ZN(n11254) );
  NAND2_X1 U11354 ( .A1(n11484), .A2(n11485), .ZN(n11482) );
  XNOR2_X1 U11355 ( .A(n11486), .B(n11487), .ZN(n11259) );
  XNOR2_X1 U11356 ( .A(n11488), .B(n11489), .ZN(n11487) );
  XOR2_X1 U11357 ( .A(n11490), .B(n11491), .Z(n11262) );
  XOR2_X1 U11358 ( .A(n11492), .B(n11493), .Z(n11490) );
  NOR2_X1 U11359 ( .A1(n8939), .A2(n8942), .ZN(n11493) );
  INV_X1 U11360 ( .A(n8908), .ZN(n11269) );
  NAND2_X1 U11361 ( .A1(b_22_), .A2(a_22_), .ZN(n8908) );
  XOR2_X1 U11362 ( .A(n11494), .B(n11495), .Z(n11270) );
  XOR2_X1 U11363 ( .A(n11496), .B(n11497), .Z(n11494) );
  NOR2_X1 U11364 ( .A1(n8941), .A2(n8942), .ZN(n11497) );
  XNOR2_X1 U11365 ( .A(n11498), .B(n11499), .ZN(n11275) );
  XNOR2_X1 U11366 ( .A(n11500), .B(n8905), .ZN(n11499) );
  XOR2_X1 U11367 ( .A(n11501), .B(n11502), .Z(n11278) );
  XOR2_X1 U11368 ( .A(n11503), .B(n11504), .Z(n11501) );
  NOR2_X1 U11369 ( .A1(n8944), .A2(n8942), .ZN(n11504) );
  XNOR2_X1 U11370 ( .A(n11505), .B(n11506), .ZN(n11283) );
  XNOR2_X1 U11371 ( .A(n11507), .B(n11508), .ZN(n11506) );
  XOR2_X1 U11372 ( .A(n11509), .B(n11510), .Z(n11287) );
  XOR2_X1 U11373 ( .A(n11511), .B(n11512), .Z(n11509) );
  NOR2_X1 U11374 ( .A1(n8947), .A2(n8942), .ZN(n11512) );
  XOR2_X1 U11375 ( .A(n11513), .B(n11514), .Z(n11291) );
  XOR2_X1 U11376 ( .A(n11515), .B(n11516), .Z(n11513) );
  XOR2_X1 U11377 ( .A(n11517), .B(n11518), .Z(n11174) );
  XOR2_X1 U11378 ( .A(n11519), .B(n11520), .Z(n11517) );
  NOR2_X1 U11379 ( .A1(n8950), .A2(n8942), .ZN(n11520) );
  XOR2_X1 U11380 ( .A(n11521), .B(n11522), .Z(n11294) );
  XOR2_X1 U11381 ( .A(n11523), .B(n11524), .Z(n11521) );
  XNOR2_X1 U11382 ( .A(n11525), .B(n11526), .ZN(n11299) );
  XOR2_X1 U11383 ( .A(n11527), .B(n11528), .Z(n11526) );
  NAND2_X1 U11384 ( .A1(b_21_), .A2(a_14_), .ZN(n11528) );
  XOR2_X1 U11385 ( .A(n11529), .B(n11530), .Z(n11302) );
  XOR2_X1 U11386 ( .A(n11531), .B(n11532), .Z(n11529) );
  XOR2_X1 U11387 ( .A(n11533), .B(n11534), .Z(n11155) );
  XOR2_X1 U11388 ( .A(n11535), .B(n11536), .Z(n11533) );
  NOR2_X1 U11389 ( .A1(n8956), .A2(n8942), .ZN(n11536) );
  XOR2_X1 U11390 ( .A(n11537), .B(n11538), .Z(n11307) );
  XOR2_X1 U11391 ( .A(n11539), .B(n11540), .Z(n11537) );
  XNOR2_X1 U11392 ( .A(n11541), .B(n11542), .ZN(n11311) );
  XNOR2_X1 U11393 ( .A(n11543), .B(n11544), .ZN(n11542) );
  XOR2_X1 U11394 ( .A(n11545), .B(n11546), .Z(n11314) );
  XOR2_X1 U11395 ( .A(n11547), .B(n11548), .Z(n11545) );
  NOR2_X1 U11396 ( .A1(n8605), .A2(n8942), .ZN(n11548) );
  XOR2_X1 U11397 ( .A(n11549), .B(n11550), .Z(n11136) );
  XOR2_X1 U11398 ( .A(n11551), .B(n11552), .Z(n11549) );
  NOR2_X1 U11399 ( .A1(n8619), .A2(n8942), .ZN(n11552) );
  XOR2_X1 U11400 ( .A(n11553), .B(n11554), .Z(n11318) );
  XOR2_X1 U11401 ( .A(n11555), .B(n11556), .Z(n11553) );
  NOR2_X1 U11402 ( .A1(n8962), .A2(n8942), .ZN(n11556) );
  XOR2_X1 U11403 ( .A(n11557), .B(n11558), .Z(n11322) );
  XOR2_X1 U11404 ( .A(n11559), .B(n11560), .Z(n11557) );
  NOR2_X1 U11405 ( .A1(n8681), .A2(n8942), .ZN(n11560) );
  XOR2_X1 U11406 ( .A(n11561), .B(n11562), .Z(n11331) );
  XOR2_X1 U11407 ( .A(n11563), .B(n11564), .Z(n11561) );
  NOR2_X1 U11408 ( .A1(n8966), .A2(n8942), .ZN(n11564) );
  XNOR2_X1 U11409 ( .A(n11565), .B(n11566), .ZN(n11335) );
  XOR2_X1 U11410 ( .A(n11567), .B(n11568), .Z(n11565) );
  NOR2_X1 U11411 ( .A1(n8778), .A2(n8942), .ZN(n11568) );
  XOR2_X1 U11412 ( .A(n11569), .B(n11570), .Z(n11338) );
  XOR2_X1 U11413 ( .A(n11571), .B(n11572), .Z(n11569) );
  NOR2_X1 U11414 ( .A1(n8792), .A2(n8942), .ZN(n11572) );
  XNOR2_X1 U11415 ( .A(n11573), .B(n11574), .ZN(n11344) );
  XOR2_X1 U11416 ( .A(n11575), .B(n11576), .Z(n11573) );
  NOR2_X1 U11417 ( .A1(n8969), .A2(n8942), .ZN(n11576) );
  XNOR2_X1 U11418 ( .A(n11577), .B(n11578), .ZN(n9178) );
  XNOR2_X1 U11419 ( .A(n11579), .B(n11580), .ZN(n11577) );
  AND2_X1 U11420 ( .A1(n9171), .A2(n11348), .ZN(n11349) );
  NAND2_X1 U11421 ( .A1(n11581), .A2(n11582), .ZN(n11348) );
  XOR2_X1 U11422 ( .A(n11583), .B(n11584), .Z(n11582) );
  NOR2_X1 U11423 ( .A1(n11585), .A2(n11586), .ZN(n11581) );
  NOR2_X1 U11424 ( .A1(n11579), .A2(n11578), .ZN(n11586) );
  INV_X1 U11425 ( .A(n11587), .ZN(n11585) );
  OR2_X1 U11426 ( .A1(n9171), .A2(n9170), .ZN(n9050) );
  XNOR2_X1 U11427 ( .A(n9168), .B(n9167), .ZN(n9170) );
  NAND2_X1 U11428 ( .A1(n11588), .A2(n11589), .ZN(n9171) );
  NAND2_X1 U11429 ( .A1(n11590), .A2(n11587), .ZN(n11589) );
  NAND2_X1 U11430 ( .A1(n11580), .A2(n11591), .ZN(n11587) );
  NAND2_X1 U11431 ( .A1(n11579), .A2(n11578), .ZN(n11591) );
  NOR2_X1 U11432 ( .A1(n8942), .A2(n8974), .ZN(n11580) );
  OR2_X1 U11433 ( .A1(n11578), .A2(n11579), .ZN(n11590) );
  AND2_X1 U11434 ( .A1(n11592), .A2(n11593), .ZN(n11579) );
  NAND2_X1 U11435 ( .A1(n11594), .A2(b_21_), .ZN(n11593) );
  NOR2_X1 U11436 ( .A1(n11595), .A2(n8969), .ZN(n11594) );
  NOR2_X1 U11437 ( .A1(n11574), .A2(n11575), .ZN(n11595) );
  NAND2_X1 U11438 ( .A1(n11574), .A2(n11575), .ZN(n11592) );
  NAND2_X1 U11439 ( .A1(n11596), .A2(n11597), .ZN(n11575) );
  NAND2_X1 U11440 ( .A1(n11598), .A2(b_21_), .ZN(n11597) );
  NOR2_X1 U11441 ( .A1(n11599), .A2(n8792), .ZN(n11598) );
  NOR2_X1 U11442 ( .A1(n11570), .A2(n11571), .ZN(n11599) );
  NAND2_X1 U11443 ( .A1(n11570), .A2(n11571), .ZN(n11596) );
  NAND2_X1 U11444 ( .A1(n11600), .A2(n11601), .ZN(n11571) );
  NAND2_X1 U11445 ( .A1(n11602), .A2(b_21_), .ZN(n11601) );
  NOR2_X1 U11446 ( .A1(n11603), .A2(n8778), .ZN(n11602) );
  NOR2_X1 U11447 ( .A1(n11566), .A2(n11567), .ZN(n11603) );
  NAND2_X1 U11448 ( .A1(n11566), .A2(n11567), .ZN(n11600) );
  NAND2_X1 U11449 ( .A1(n11604), .A2(n11605), .ZN(n11567) );
  NAND2_X1 U11450 ( .A1(n11606), .A2(b_21_), .ZN(n11605) );
  NOR2_X1 U11451 ( .A1(n11607), .A2(n8966), .ZN(n11606) );
  NOR2_X1 U11452 ( .A1(n11562), .A2(n11563), .ZN(n11607) );
  NAND2_X1 U11453 ( .A1(n11562), .A2(n11563), .ZN(n11604) );
  NAND2_X1 U11454 ( .A1(n11608), .A2(n11609), .ZN(n11563) );
  NAND2_X1 U11455 ( .A1(n11610), .A2(b_21_), .ZN(n11609) );
  NOR2_X1 U11456 ( .A1(n11611), .A2(n8723), .ZN(n11610) );
  NOR2_X1 U11457 ( .A1(n11369), .A2(n11370), .ZN(n11611) );
  NAND2_X1 U11458 ( .A1(n11369), .A2(n11370), .ZN(n11608) );
  NAND2_X1 U11459 ( .A1(n11612), .A2(n11613), .ZN(n11370) );
  NAND2_X1 U11460 ( .A1(n11614), .A2(b_21_), .ZN(n11613) );
  NOR2_X1 U11461 ( .A1(n11615), .A2(n8681), .ZN(n11614) );
  NOR2_X1 U11462 ( .A1(n11558), .A2(n11559), .ZN(n11615) );
  NAND2_X1 U11463 ( .A1(n11558), .A2(n11559), .ZN(n11612) );
  NAND2_X1 U11464 ( .A1(n11616), .A2(n11617), .ZN(n11559) );
  NAND2_X1 U11465 ( .A1(n11618), .A2(b_21_), .ZN(n11617) );
  NOR2_X1 U11466 ( .A1(n11619), .A2(n8962), .ZN(n11618) );
  NOR2_X1 U11467 ( .A1(n11554), .A2(n11555), .ZN(n11619) );
  NAND2_X1 U11468 ( .A1(n11554), .A2(n11555), .ZN(n11616) );
  NAND2_X1 U11469 ( .A1(n11620), .A2(n11621), .ZN(n11555) );
  NAND2_X1 U11470 ( .A1(n11622), .A2(b_21_), .ZN(n11621) );
  NOR2_X1 U11471 ( .A1(n11623), .A2(n8619), .ZN(n11622) );
  NOR2_X1 U11472 ( .A1(n11550), .A2(n11551), .ZN(n11623) );
  NAND2_X1 U11473 ( .A1(n11550), .A2(n11551), .ZN(n11620) );
  NAND2_X1 U11474 ( .A1(n11624), .A2(n11625), .ZN(n11551) );
  NAND2_X1 U11475 ( .A1(n11626), .A2(b_21_), .ZN(n11625) );
  NOR2_X1 U11476 ( .A1(n11627), .A2(n8605), .ZN(n11626) );
  NOR2_X1 U11477 ( .A1(n11546), .A2(n11547), .ZN(n11627) );
  NAND2_X1 U11478 ( .A1(n11546), .A2(n11547), .ZN(n11624) );
  NAND2_X1 U11479 ( .A1(n11628), .A2(n11629), .ZN(n11547) );
  NAND2_X1 U11480 ( .A1(n11544), .A2(n11630), .ZN(n11629) );
  OR2_X1 U11481 ( .A1(n11543), .A2(n11541), .ZN(n11630) );
  NOR2_X1 U11482 ( .A1(n8942), .A2(n8959), .ZN(n11544) );
  NAND2_X1 U11483 ( .A1(n11541), .A2(n11543), .ZN(n11628) );
  NAND2_X1 U11484 ( .A1(n11631), .A2(n11632), .ZN(n11543) );
  NAND2_X1 U11485 ( .A1(n11540), .A2(n11633), .ZN(n11632) );
  OR2_X1 U11486 ( .A1(n11539), .A2(n11538), .ZN(n11633) );
  NOR2_X1 U11487 ( .A1(n8942), .A2(n8550), .ZN(n11540) );
  NAND2_X1 U11488 ( .A1(n11538), .A2(n11539), .ZN(n11631) );
  NAND2_X1 U11489 ( .A1(n11634), .A2(n11635), .ZN(n11539) );
  NAND2_X1 U11490 ( .A1(n11636), .A2(b_21_), .ZN(n11635) );
  NOR2_X1 U11491 ( .A1(n11637), .A2(n8956), .ZN(n11636) );
  NOR2_X1 U11492 ( .A1(n11534), .A2(n11535), .ZN(n11637) );
  NAND2_X1 U11493 ( .A1(n11534), .A2(n11535), .ZN(n11634) );
  NAND2_X1 U11494 ( .A1(n11638), .A2(n11639), .ZN(n11535) );
  NAND2_X1 U11495 ( .A1(n11532), .A2(n11640), .ZN(n11639) );
  OR2_X1 U11496 ( .A1(n11531), .A2(n11530), .ZN(n11640) );
  NOR2_X1 U11497 ( .A1(n8942), .A2(n8495), .ZN(n11532) );
  NAND2_X1 U11498 ( .A1(n11530), .A2(n11531), .ZN(n11638) );
  NAND2_X1 U11499 ( .A1(n11641), .A2(n11642), .ZN(n11531) );
  NAND2_X1 U11500 ( .A1(n11643), .A2(b_21_), .ZN(n11642) );
  NOR2_X1 U11501 ( .A1(n11644), .A2(n8953), .ZN(n11643) );
  NOR2_X1 U11502 ( .A1(n11525), .A2(n11527), .ZN(n11644) );
  NAND2_X1 U11503 ( .A1(n11525), .A2(n11527), .ZN(n11641) );
  NAND2_X1 U11504 ( .A1(n11645), .A2(n11646), .ZN(n11527) );
  NAND2_X1 U11505 ( .A1(n11524), .A2(n11647), .ZN(n11646) );
  OR2_X1 U11506 ( .A1(n11523), .A2(n11522), .ZN(n11647) );
  NOR2_X1 U11507 ( .A1(n8942), .A2(n8440), .ZN(n11524) );
  NAND2_X1 U11508 ( .A1(n11522), .A2(n11523), .ZN(n11645) );
  NAND2_X1 U11509 ( .A1(n11648), .A2(n11649), .ZN(n11523) );
  NAND2_X1 U11510 ( .A1(n11650), .A2(b_21_), .ZN(n11649) );
  NOR2_X1 U11511 ( .A1(n11651), .A2(n8950), .ZN(n11650) );
  NOR2_X1 U11512 ( .A1(n11518), .A2(n11519), .ZN(n11651) );
  NAND2_X1 U11513 ( .A1(n11518), .A2(n11519), .ZN(n11648) );
  NAND2_X1 U11514 ( .A1(n11652), .A2(n11653), .ZN(n11519) );
  NAND2_X1 U11515 ( .A1(n11516), .A2(n11654), .ZN(n11653) );
  OR2_X1 U11516 ( .A1(n11515), .A2(n11514), .ZN(n11654) );
  NOR2_X1 U11517 ( .A1(n8942), .A2(n8385), .ZN(n11516) );
  NAND2_X1 U11518 ( .A1(n11514), .A2(n11515), .ZN(n11652) );
  NAND2_X1 U11519 ( .A1(n11655), .A2(n11656), .ZN(n11515) );
  NAND2_X1 U11520 ( .A1(n11657), .A2(b_21_), .ZN(n11656) );
  NOR2_X1 U11521 ( .A1(n11658), .A2(n8947), .ZN(n11657) );
  NOR2_X1 U11522 ( .A1(n11510), .A2(n11511), .ZN(n11658) );
  NAND2_X1 U11523 ( .A1(n11510), .A2(n11511), .ZN(n11655) );
  NAND2_X1 U11524 ( .A1(n11659), .A2(n11660), .ZN(n11511) );
  NAND2_X1 U11525 ( .A1(n11508), .A2(n11661), .ZN(n11660) );
  OR2_X1 U11526 ( .A1(n11507), .A2(n11505), .ZN(n11661) );
  NOR2_X1 U11527 ( .A1(n8942), .A2(n8324), .ZN(n11508) );
  NAND2_X1 U11528 ( .A1(n11505), .A2(n11507), .ZN(n11659) );
  NAND2_X1 U11529 ( .A1(n11662), .A2(n11663), .ZN(n11507) );
  NAND2_X1 U11530 ( .A1(n11664), .A2(b_21_), .ZN(n11663) );
  NOR2_X1 U11531 ( .A1(n11665), .A2(n8944), .ZN(n11664) );
  NOR2_X1 U11532 ( .A1(n11502), .A2(n11503), .ZN(n11665) );
  NAND2_X1 U11533 ( .A1(n11502), .A2(n11503), .ZN(n11662) );
  NAND2_X1 U11534 ( .A1(n11666), .A2(n11667), .ZN(n11503) );
  NAND2_X1 U11535 ( .A1(n8905), .A2(n11668), .ZN(n11667) );
  OR2_X1 U11536 ( .A1(n11500), .A2(n11498), .ZN(n11668) );
  NOR2_X1 U11537 ( .A1(n8942), .A2(n8268), .ZN(n8905) );
  NAND2_X1 U11538 ( .A1(n11498), .A2(n11500), .ZN(n11666) );
  NAND2_X1 U11539 ( .A1(n11669), .A2(n11670), .ZN(n11500) );
  NAND2_X1 U11540 ( .A1(n11671), .A2(b_21_), .ZN(n11670) );
  NOR2_X1 U11541 ( .A1(n11672), .A2(n8941), .ZN(n11671) );
  NOR2_X1 U11542 ( .A1(n11495), .A2(n11496), .ZN(n11672) );
  NAND2_X1 U11543 ( .A1(n11495), .A2(n11496), .ZN(n11669) );
  NAND2_X1 U11544 ( .A1(n11673), .A2(n11674), .ZN(n11496) );
  NAND2_X1 U11545 ( .A1(n11437), .A2(n11675), .ZN(n11674) );
  OR2_X1 U11546 ( .A1(n11436), .A2(n11434), .ZN(n11675) );
  NOR2_X1 U11547 ( .A1(n8942), .A2(n8213), .ZN(n11437) );
  NAND2_X1 U11548 ( .A1(n11434), .A2(n11436), .ZN(n11673) );
  NAND2_X1 U11549 ( .A1(n11676), .A2(n11677), .ZN(n11436) );
  NAND2_X1 U11550 ( .A1(n11678), .A2(b_21_), .ZN(n11677) );
  NOR2_X1 U11551 ( .A1(n11679), .A2(n8939), .ZN(n11678) );
  NOR2_X1 U11552 ( .A1(n11491), .A2(n11492), .ZN(n11679) );
  NAND2_X1 U11553 ( .A1(n11491), .A2(n11492), .ZN(n11676) );
  NAND2_X1 U11554 ( .A1(n11680), .A2(n11681), .ZN(n11492) );
  NAND2_X1 U11555 ( .A1(n11489), .A2(n11682), .ZN(n11681) );
  OR2_X1 U11556 ( .A1(n11488), .A2(n11486), .ZN(n11682) );
  NOR2_X1 U11557 ( .A1(n8942), .A2(n8158), .ZN(n11489) );
  NAND2_X1 U11558 ( .A1(n11486), .A2(n11488), .ZN(n11680) );
  NAND2_X1 U11559 ( .A1(n11484), .A2(n11683), .ZN(n11488) );
  NAND2_X1 U11560 ( .A1(n11483), .A2(n11485), .ZN(n11683) );
  NAND2_X1 U11561 ( .A1(n11684), .A2(n11685), .ZN(n11485) );
  NAND2_X1 U11562 ( .A1(b_21_), .A2(a_26_), .ZN(n11685) );
  INV_X1 U11563 ( .A(n11686), .ZN(n11684) );
  XNOR2_X1 U11564 ( .A(n11687), .B(n11688), .ZN(n11483) );
  NAND2_X1 U11565 ( .A1(n11689), .A2(n11690), .ZN(n11687) );
  NAND2_X1 U11566 ( .A1(a_26_), .A2(n11686), .ZN(n11484) );
  NAND2_X1 U11567 ( .A1(n11454), .A2(n11691), .ZN(n11686) );
  NAND2_X1 U11568 ( .A1(n11453), .A2(n11455), .ZN(n11691) );
  NAND2_X1 U11569 ( .A1(n11692), .A2(n11693), .ZN(n11455) );
  NAND2_X1 U11570 ( .A1(b_21_), .A2(a_27_), .ZN(n11693) );
  INV_X1 U11571 ( .A(n11694), .ZN(n11692) );
  XOR2_X1 U11572 ( .A(n11695), .B(n11696), .Z(n11453) );
  XNOR2_X1 U11573 ( .A(n11697), .B(n11698), .ZN(n11695) );
  NAND2_X1 U11574 ( .A1(b_20_), .A2(a_28_), .ZN(n11697) );
  NAND2_X1 U11575 ( .A1(a_27_), .A2(n11694), .ZN(n11454) );
  NAND2_X1 U11576 ( .A1(n11699), .A2(n11700), .ZN(n11694) );
  NAND2_X1 U11577 ( .A1(n11701), .A2(b_21_), .ZN(n11700) );
  NOR2_X1 U11578 ( .A1(n11702), .A2(n8055), .ZN(n11701) );
  NOR2_X1 U11579 ( .A1(n11461), .A2(n11463), .ZN(n11702) );
  NAND2_X1 U11580 ( .A1(n11461), .A2(n11463), .ZN(n11699) );
  NAND2_X1 U11581 ( .A1(n11703), .A2(n11704), .ZN(n11463) );
  NAND2_X1 U11582 ( .A1(n11479), .A2(n11705), .ZN(n11704) );
  OR2_X1 U11583 ( .A1(n11480), .A2(n11481), .ZN(n11705) );
  NOR2_X1 U11584 ( .A1(n8942), .A2(n8041), .ZN(n11479) );
  NAND2_X1 U11585 ( .A1(n11481), .A2(n11480), .ZN(n11703) );
  NAND2_X1 U11586 ( .A1(n11706), .A2(n11707), .ZN(n11480) );
  NAND2_X1 U11587 ( .A1(b_19_), .A2(n11708), .ZN(n11707) );
  NAND2_X1 U11588 ( .A1(n8003), .A2(n11709), .ZN(n11708) );
  NAND2_X1 U11589 ( .A1(a_31_), .A2(n8943), .ZN(n11709) );
  NAND2_X1 U11590 ( .A1(b_20_), .A2(n11710), .ZN(n11706) );
  NAND2_X1 U11591 ( .A1(n9341), .A2(n11711), .ZN(n11710) );
  NAND2_X1 U11592 ( .A1(a_30_), .A2(n8945), .ZN(n11711) );
  AND2_X1 U11593 ( .A1(n11712), .A2(n7953), .ZN(n11481) );
  NOR2_X1 U11594 ( .A1(n8942), .A2(n8943), .ZN(n11712) );
  XOR2_X1 U11595 ( .A(n11713), .B(n11714), .Z(n11461) );
  XOR2_X1 U11596 ( .A(n11715), .B(n11716), .Z(n11713) );
  XNOR2_X1 U11597 ( .A(n11717), .B(n11718), .ZN(n11486) );
  NAND2_X1 U11598 ( .A1(n11719), .A2(n11720), .ZN(n11717) );
  XNOR2_X1 U11599 ( .A(n11721), .B(n11722), .ZN(n11491) );
  XNOR2_X1 U11600 ( .A(n11723), .B(n11724), .ZN(n11722) );
  XOR2_X1 U11601 ( .A(n11725), .B(n11726), .Z(n11434) );
  XOR2_X1 U11602 ( .A(n11727), .B(n11728), .Z(n11725) );
  NOR2_X1 U11603 ( .A1(n8939), .A2(n8943), .ZN(n11728) );
  XNOR2_X1 U11604 ( .A(n11729), .B(n11730), .ZN(n11495) );
  XNOR2_X1 U11605 ( .A(n11731), .B(n11732), .ZN(n11730) );
  XOR2_X1 U11606 ( .A(n11733), .B(n11734), .Z(n11498) );
  XOR2_X1 U11607 ( .A(n11735), .B(n11736), .Z(n11733) );
  NOR2_X1 U11608 ( .A1(n8941), .A2(n8943), .ZN(n11736) );
  XNOR2_X1 U11609 ( .A(n11737), .B(n11738), .ZN(n11502) );
  XNOR2_X1 U11610 ( .A(n11739), .B(n11740), .ZN(n11738) );
  XOR2_X1 U11611 ( .A(n11741), .B(n11742), .Z(n11505) );
  XOR2_X1 U11612 ( .A(n11743), .B(n11744), .Z(n11741) );
  XNOR2_X1 U11613 ( .A(n11745), .B(n11746), .ZN(n11510) );
  XNOR2_X1 U11614 ( .A(n11747), .B(n11748), .ZN(n11746) );
  XNOR2_X1 U11615 ( .A(n11749), .B(n11750), .ZN(n11514) );
  XOR2_X1 U11616 ( .A(n11751), .B(n11752), .Z(n11750) );
  NAND2_X1 U11617 ( .A1(b_20_), .A2(a_18_), .ZN(n11752) );
  XOR2_X1 U11618 ( .A(n11753), .B(n11754), .Z(n11518) );
  XOR2_X1 U11619 ( .A(n11755), .B(n11756), .Z(n11753) );
  XNOR2_X1 U11620 ( .A(n11757), .B(n11758), .ZN(n11522) );
  XOR2_X1 U11621 ( .A(n11759), .B(n11760), .Z(n11758) );
  NAND2_X1 U11622 ( .A1(b_20_), .A2(a_16_), .ZN(n11760) );
  XOR2_X1 U11623 ( .A(n11761), .B(n11762), .Z(n11525) );
  XOR2_X1 U11624 ( .A(n11763), .B(n11764), .Z(n11761) );
  XOR2_X1 U11625 ( .A(n11765), .B(n11766), .Z(n11530) );
  XOR2_X1 U11626 ( .A(n11767), .B(n11768), .Z(n11765) );
  NOR2_X1 U11627 ( .A1(n8953), .A2(n8943), .ZN(n11768) );
  XOR2_X1 U11628 ( .A(n11769), .B(n11770), .Z(n11534) );
  XOR2_X1 U11629 ( .A(n11771), .B(n11772), .Z(n11769) );
  XNOR2_X1 U11630 ( .A(n11773), .B(n11774), .ZN(n11538) );
  XOR2_X1 U11631 ( .A(n11775), .B(n11776), .Z(n11774) );
  NAND2_X1 U11632 ( .A1(b_20_), .A2(a_12_), .ZN(n11776) );
  XOR2_X1 U11633 ( .A(n11777), .B(n11778), .Z(n11541) );
  XOR2_X1 U11634 ( .A(n11779), .B(n11780), .Z(n11777) );
  NOR2_X1 U11635 ( .A1(n8550), .A2(n8943), .ZN(n11780) );
  XNOR2_X1 U11636 ( .A(n11781), .B(n11782), .ZN(n11546) );
  XNOR2_X1 U11637 ( .A(n11783), .B(n11784), .ZN(n11781) );
  XOR2_X1 U11638 ( .A(n11785), .B(n11786), .Z(n11550) );
  XOR2_X1 U11639 ( .A(n11787), .B(n11788), .Z(n11785) );
  XNOR2_X1 U11640 ( .A(n11789), .B(n11790), .ZN(n11554) );
  XNOR2_X1 U11641 ( .A(n11791), .B(n11792), .ZN(n11790) );
  XNOR2_X1 U11642 ( .A(n11793), .B(n11794), .ZN(n11558) );
  XOR2_X1 U11643 ( .A(n11795), .B(n11796), .Z(n11794) );
  NAND2_X1 U11644 ( .A1(b_20_), .A2(a_7_), .ZN(n11796) );
  XNOR2_X1 U11645 ( .A(n11797), .B(n11798), .ZN(n11369) );
  NAND2_X1 U11646 ( .A1(n11799), .A2(n11800), .ZN(n11797) );
  XNOR2_X1 U11647 ( .A(n11801), .B(n11802), .ZN(n11562) );
  NAND2_X1 U11648 ( .A1(n11803), .A2(n11804), .ZN(n11801) );
  XNOR2_X1 U11649 ( .A(n11805), .B(n11806), .ZN(n11566) );
  XNOR2_X1 U11650 ( .A(n11807), .B(n11808), .ZN(n11805) );
  XNOR2_X1 U11651 ( .A(n11809), .B(n11810), .ZN(n11570) );
  XOR2_X1 U11652 ( .A(n11811), .B(n11812), .Z(n11810) );
  NAND2_X1 U11653 ( .A1(b_20_), .A2(a_3_), .ZN(n11812) );
  XNOR2_X1 U11654 ( .A(n11813), .B(n11814), .ZN(n11574) );
  NAND2_X1 U11655 ( .A1(n11815), .A2(n11816), .ZN(n11813) );
  XOR2_X1 U11656 ( .A(n11817), .B(n11818), .Z(n11578) );
  XNOR2_X1 U11657 ( .A(n11819), .B(n11820), .ZN(n11817) );
  XOR2_X1 U11658 ( .A(n11821), .B(n11583), .Z(n11588) );
  XNOR2_X1 U11659 ( .A(n11822), .B(n11823), .ZN(n11583) );
  NOR2_X1 U11660 ( .A1(n8974), .A2(n8943), .ZN(n11823) );
  INV_X1 U11661 ( .A(n11584), .ZN(n11821) );
  NAND2_X1 U11662 ( .A1(n11824), .A2(n11825), .ZN(n9062) );
  XOR2_X1 U11663 ( .A(n9161), .B(n9160), .Z(n11825) );
  AND2_X1 U11664 ( .A1(n9168), .A2(n9167), .ZN(n11824) );
  XOR2_X1 U11665 ( .A(n11826), .B(n11827), .Z(n9167) );
  XOR2_X1 U11666 ( .A(n11828), .B(n11829), .Z(n11826) );
  NOR2_X1 U11667 ( .A1(n8974), .A2(n8945), .ZN(n11829) );
  NAND2_X1 U11668 ( .A1(n11830), .A2(n11831), .ZN(n9168) );
  NAND2_X1 U11669 ( .A1(n11832), .A2(b_20_), .ZN(n11831) );
  NOR2_X1 U11670 ( .A1(n11833), .A2(n8974), .ZN(n11832) );
  NOR2_X1 U11671 ( .A1(n11584), .A2(n11822), .ZN(n11833) );
  NAND2_X1 U11672 ( .A1(n11584), .A2(n11822), .ZN(n11830) );
  NAND2_X1 U11673 ( .A1(n11834), .A2(n11835), .ZN(n11822) );
  NAND2_X1 U11674 ( .A1(n11820), .A2(n11836), .ZN(n11835) );
  NAND2_X1 U11675 ( .A1(n11819), .A2(n11818), .ZN(n11836) );
  NOR2_X1 U11676 ( .A1(n8943), .A2(n8969), .ZN(n11820) );
  OR2_X1 U11677 ( .A1(n11818), .A2(n11819), .ZN(n11834) );
  AND2_X1 U11678 ( .A1(n11815), .A2(n11837), .ZN(n11819) );
  NAND2_X1 U11679 ( .A1(n11814), .A2(n11816), .ZN(n11837) );
  NAND2_X1 U11680 ( .A1(n11838), .A2(n11839), .ZN(n11816) );
  NAND2_X1 U11681 ( .A1(b_20_), .A2(a_2_), .ZN(n11839) );
  INV_X1 U11682 ( .A(n11840), .ZN(n11838) );
  XOR2_X1 U11683 ( .A(n11841), .B(n11842), .Z(n11814) );
  XOR2_X1 U11684 ( .A(n11843), .B(n11844), .Z(n11841) );
  NOR2_X1 U11685 ( .A1(n8778), .A2(n8945), .ZN(n11844) );
  NAND2_X1 U11686 ( .A1(a_2_), .A2(n11840), .ZN(n11815) );
  NAND2_X1 U11687 ( .A1(n11845), .A2(n11846), .ZN(n11840) );
  NAND2_X1 U11688 ( .A1(n11847), .A2(b_20_), .ZN(n11846) );
  NOR2_X1 U11689 ( .A1(n11848), .A2(n8778), .ZN(n11847) );
  NOR2_X1 U11690 ( .A1(n11809), .A2(n11811), .ZN(n11848) );
  NAND2_X1 U11691 ( .A1(n11809), .A2(n11811), .ZN(n11845) );
  NAND2_X1 U11692 ( .A1(n11849), .A2(n11850), .ZN(n11811) );
  NAND2_X1 U11693 ( .A1(n11808), .A2(n11851), .ZN(n11850) );
  NAND2_X1 U11694 ( .A1(n11807), .A2(n11806), .ZN(n11851) );
  NOR2_X1 U11695 ( .A1(n8943), .A2(n8966), .ZN(n11808) );
  OR2_X1 U11696 ( .A1(n11806), .A2(n11807), .ZN(n11849) );
  AND2_X1 U11697 ( .A1(n11803), .A2(n11852), .ZN(n11807) );
  NAND2_X1 U11698 ( .A1(n11802), .A2(n11804), .ZN(n11852) );
  NAND2_X1 U11699 ( .A1(n11853), .A2(n11854), .ZN(n11804) );
  NAND2_X1 U11700 ( .A1(b_20_), .A2(a_5_), .ZN(n11854) );
  INV_X1 U11701 ( .A(n11855), .ZN(n11853) );
  XOR2_X1 U11702 ( .A(n11856), .B(n11857), .Z(n11802) );
  XOR2_X1 U11703 ( .A(n11858), .B(n11859), .Z(n11856) );
  NOR2_X1 U11704 ( .A1(n8681), .A2(n8945), .ZN(n11859) );
  NAND2_X1 U11705 ( .A1(a_5_), .A2(n11855), .ZN(n11803) );
  NAND2_X1 U11706 ( .A1(n11799), .A2(n11860), .ZN(n11855) );
  NAND2_X1 U11707 ( .A1(n11798), .A2(n11800), .ZN(n11860) );
  NAND2_X1 U11708 ( .A1(n11861), .A2(n11862), .ZN(n11800) );
  NAND2_X1 U11709 ( .A1(b_20_), .A2(a_6_), .ZN(n11862) );
  INV_X1 U11710 ( .A(n11863), .ZN(n11861) );
  XOR2_X1 U11711 ( .A(n11864), .B(n11865), .Z(n11798) );
  XOR2_X1 U11712 ( .A(n11866), .B(n11867), .Z(n11864) );
  NOR2_X1 U11713 ( .A1(n8962), .A2(n8945), .ZN(n11867) );
  NAND2_X1 U11714 ( .A1(a_6_), .A2(n11863), .ZN(n11799) );
  NAND2_X1 U11715 ( .A1(n11868), .A2(n11869), .ZN(n11863) );
  NAND2_X1 U11716 ( .A1(n11870), .A2(b_20_), .ZN(n11869) );
  NOR2_X1 U11717 ( .A1(n11871), .A2(n8962), .ZN(n11870) );
  NOR2_X1 U11718 ( .A1(n11793), .A2(n11795), .ZN(n11871) );
  NAND2_X1 U11719 ( .A1(n11793), .A2(n11795), .ZN(n11868) );
  NAND2_X1 U11720 ( .A1(n11872), .A2(n11873), .ZN(n11795) );
  NAND2_X1 U11721 ( .A1(n11792), .A2(n11874), .ZN(n11873) );
  OR2_X1 U11722 ( .A1(n11791), .A2(n11789), .ZN(n11874) );
  NOR2_X1 U11723 ( .A1(n8943), .A2(n8619), .ZN(n11792) );
  NAND2_X1 U11724 ( .A1(n11789), .A2(n11791), .ZN(n11872) );
  NAND2_X1 U11725 ( .A1(n11875), .A2(n11876), .ZN(n11791) );
  NAND2_X1 U11726 ( .A1(n11788), .A2(n11877), .ZN(n11876) );
  OR2_X1 U11727 ( .A1(n11787), .A2(n11786), .ZN(n11877) );
  NOR2_X1 U11728 ( .A1(n8943), .A2(n8605), .ZN(n11788) );
  NAND2_X1 U11729 ( .A1(n11786), .A2(n11787), .ZN(n11875) );
  NAND2_X1 U11730 ( .A1(n11878), .A2(n11879), .ZN(n11787) );
  NAND2_X1 U11731 ( .A1(n11784), .A2(n11880), .ZN(n11879) );
  NAND2_X1 U11732 ( .A1(n11783), .A2(n11782), .ZN(n11880) );
  NOR2_X1 U11733 ( .A1(n8943), .A2(n8959), .ZN(n11784) );
  OR2_X1 U11734 ( .A1(n11782), .A2(n11783), .ZN(n11878) );
  AND2_X1 U11735 ( .A1(n11881), .A2(n11882), .ZN(n11783) );
  NAND2_X1 U11736 ( .A1(n11883), .A2(b_20_), .ZN(n11882) );
  NOR2_X1 U11737 ( .A1(n11884), .A2(n8550), .ZN(n11883) );
  NOR2_X1 U11738 ( .A1(n11778), .A2(n11779), .ZN(n11884) );
  NAND2_X1 U11739 ( .A1(n11778), .A2(n11779), .ZN(n11881) );
  NAND2_X1 U11740 ( .A1(n11885), .A2(n11886), .ZN(n11779) );
  NAND2_X1 U11741 ( .A1(n11887), .A2(b_20_), .ZN(n11886) );
  NOR2_X1 U11742 ( .A1(n11888), .A2(n8956), .ZN(n11887) );
  NOR2_X1 U11743 ( .A1(n11773), .A2(n11775), .ZN(n11888) );
  NAND2_X1 U11744 ( .A1(n11773), .A2(n11775), .ZN(n11885) );
  NAND2_X1 U11745 ( .A1(n11889), .A2(n11890), .ZN(n11775) );
  NAND2_X1 U11746 ( .A1(n11772), .A2(n11891), .ZN(n11890) );
  OR2_X1 U11747 ( .A1(n11771), .A2(n11770), .ZN(n11891) );
  NOR2_X1 U11748 ( .A1(n8943), .A2(n8495), .ZN(n11772) );
  NAND2_X1 U11749 ( .A1(n11770), .A2(n11771), .ZN(n11889) );
  NAND2_X1 U11750 ( .A1(n11892), .A2(n11893), .ZN(n11771) );
  NAND2_X1 U11751 ( .A1(n11894), .A2(b_20_), .ZN(n11893) );
  NOR2_X1 U11752 ( .A1(n11895), .A2(n8953), .ZN(n11894) );
  NOR2_X1 U11753 ( .A1(n11766), .A2(n11767), .ZN(n11895) );
  NAND2_X1 U11754 ( .A1(n11766), .A2(n11767), .ZN(n11892) );
  NAND2_X1 U11755 ( .A1(n11896), .A2(n11897), .ZN(n11767) );
  NAND2_X1 U11756 ( .A1(n11764), .A2(n11898), .ZN(n11897) );
  OR2_X1 U11757 ( .A1(n11763), .A2(n11762), .ZN(n11898) );
  NOR2_X1 U11758 ( .A1(n8943), .A2(n8440), .ZN(n11764) );
  NAND2_X1 U11759 ( .A1(n11762), .A2(n11763), .ZN(n11896) );
  NAND2_X1 U11760 ( .A1(n11899), .A2(n11900), .ZN(n11763) );
  NAND2_X1 U11761 ( .A1(n11901), .A2(b_20_), .ZN(n11900) );
  NOR2_X1 U11762 ( .A1(n11902), .A2(n8950), .ZN(n11901) );
  NOR2_X1 U11763 ( .A1(n11757), .A2(n11759), .ZN(n11902) );
  NAND2_X1 U11764 ( .A1(n11757), .A2(n11759), .ZN(n11899) );
  NAND2_X1 U11765 ( .A1(n11903), .A2(n11904), .ZN(n11759) );
  NAND2_X1 U11766 ( .A1(n11756), .A2(n11905), .ZN(n11904) );
  OR2_X1 U11767 ( .A1(n11755), .A2(n11754), .ZN(n11905) );
  NOR2_X1 U11768 ( .A1(n8943), .A2(n8385), .ZN(n11756) );
  NAND2_X1 U11769 ( .A1(n11754), .A2(n11755), .ZN(n11903) );
  NAND2_X1 U11770 ( .A1(n11906), .A2(n11907), .ZN(n11755) );
  NAND2_X1 U11771 ( .A1(n11908), .A2(b_20_), .ZN(n11907) );
  NOR2_X1 U11772 ( .A1(n11909), .A2(n8947), .ZN(n11908) );
  NOR2_X1 U11773 ( .A1(n11749), .A2(n11751), .ZN(n11909) );
  NAND2_X1 U11774 ( .A1(n11749), .A2(n11751), .ZN(n11906) );
  NAND2_X1 U11775 ( .A1(n11910), .A2(n11911), .ZN(n11751) );
  NAND2_X1 U11776 ( .A1(n11748), .A2(n11912), .ZN(n11911) );
  OR2_X1 U11777 ( .A1(n11747), .A2(n11745), .ZN(n11912) );
  NOR2_X1 U11778 ( .A1(n8943), .A2(n8324), .ZN(n11748) );
  NAND2_X1 U11779 ( .A1(n11745), .A2(n11747), .ZN(n11910) );
  NAND2_X1 U11780 ( .A1(n11913), .A2(n11914), .ZN(n11747) );
  NAND2_X1 U11781 ( .A1(n11742), .A2(n11915), .ZN(n11914) );
  OR2_X1 U11782 ( .A1(n11743), .A2(n11744), .ZN(n11915) );
  XNOR2_X1 U11783 ( .A(n11916), .B(n11917), .ZN(n11742) );
  XNOR2_X1 U11784 ( .A(n11918), .B(n11919), .ZN(n11917) );
  NAND2_X1 U11785 ( .A1(n11744), .A2(n11743), .ZN(n11913) );
  NAND2_X1 U11786 ( .A1(n11920), .A2(n11921), .ZN(n11743) );
  NAND2_X1 U11787 ( .A1(n11740), .A2(n11922), .ZN(n11921) );
  OR2_X1 U11788 ( .A1(n11739), .A2(n11737), .ZN(n11922) );
  NOR2_X1 U11789 ( .A1(n8943), .A2(n8268), .ZN(n11740) );
  NAND2_X1 U11790 ( .A1(n11737), .A2(n11739), .ZN(n11920) );
  NAND2_X1 U11791 ( .A1(n11923), .A2(n11924), .ZN(n11739) );
  NAND2_X1 U11792 ( .A1(n11925), .A2(b_20_), .ZN(n11924) );
  NOR2_X1 U11793 ( .A1(n11926), .A2(n8941), .ZN(n11925) );
  NOR2_X1 U11794 ( .A1(n11734), .A2(n11735), .ZN(n11926) );
  NAND2_X1 U11795 ( .A1(n11734), .A2(n11735), .ZN(n11923) );
  NAND2_X1 U11796 ( .A1(n11927), .A2(n11928), .ZN(n11735) );
  NAND2_X1 U11797 ( .A1(n11732), .A2(n11929), .ZN(n11928) );
  OR2_X1 U11798 ( .A1(n11731), .A2(n11729), .ZN(n11929) );
  NOR2_X1 U11799 ( .A1(n8943), .A2(n8213), .ZN(n11732) );
  NAND2_X1 U11800 ( .A1(n11729), .A2(n11731), .ZN(n11927) );
  NAND2_X1 U11801 ( .A1(n11930), .A2(n11931), .ZN(n11731) );
  NAND2_X1 U11802 ( .A1(n11932), .A2(b_20_), .ZN(n11931) );
  NOR2_X1 U11803 ( .A1(n11933), .A2(n8939), .ZN(n11932) );
  NOR2_X1 U11804 ( .A1(n11726), .A2(n11727), .ZN(n11933) );
  NAND2_X1 U11805 ( .A1(n11726), .A2(n11727), .ZN(n11930) );
  NAND2_X1 U11806 ( .A1(n11934), .A2(n11935), .ZN(n11727) );
  NAND2_X1 U11807 ( .A1(n11724), .A2(n11936), .ZN(n11935) );
  OR2_X1 U11808 ( .A1(n11723), .A2(n11721), .ZN(n11936) );
  NOR2_X1 U11809 ( .A1(n8943), .A2(n8158), .ZN(n11724) );
  NAND2_X1 U11810 ( .A1(n11721), .A2(n11723), .ZN(n11934) );
  NAND2_X1 U11811 ( .A1(n11719), .A2(n11937), .ZN(n11723) );
  NAND2_X1 U11812 ( .A1(n11718), .A2(n11720), .ZN(n11937) );
  NAND2_X1 U11813 ( .A1(n11938), .A2(n11939), .ZN(n11720) );
  NAND2_X1 U11814 ( .A1(b_20_), .A2(a_26_), .ZN(n11939) );
  INV_X1 U11815 ( .A(n11940), .ZN(n11938) );
  XNOR2_X1 U11816 ( .A(n11941), .B(n11942), .ZN(n11718) );
  NAND2_X1 U11817 ( .A1(n11943), .A2(n11944), .ZN(n11941) );
  NAND2_X1 U11818 ( .A1(a_26_), .A2(n11940), .ZN(n11719) );
  NAND2_X1 U11819 ( .A1(n11689), .A2(n11945), .ZN(n11940) );
  NAND2_X1 U11820 ( .A1(n11688), .A2(n11690), .ZN(n11945) );
  NAND2_X1 U11821 ( .A1(n11946), .A2(n11947), .ZN(n11690) );
  NAND2_X1 U11822 ( .A1(b_20_), .A2(a_27_), .ZN(n11947) );
  INV_X1 U11823 ( .A(n11948), .ZN(n11946) );
  XOR2_X1 U11824 ( .A(n11949), .B(n11950), .Z(n11688) );
  XNOR2_X1 U11825 ( .A(n11951), .B(n11952), .ZN(n11949) );
  NAND2_X1 U11826 ( .A1(b_19_), .A2(a_28_), .ZN(n11951) );
  NAND2_X1 U11827 ( .A1(a_27_), .A2(n11948), .ZN(n11689) );
  NAND2_X1 U11828 ( .A1(n11953), .A2(n11954), .ZN(n11948) );
  NAND2_X1 U11829 ( .A1(n11955), .A2(b_20_), .ZN(n11954) );
  NOR2_X1 U11830 ( .A1(n11956), .A2(n8055), .ZN(n11955) );
  NOR2_X1 U11831 ( .A1(n11696), .A2(n11698), .ZN(n11956) );
  NAND2_X1 U11832 ( .A1(n11696), .A2(n11698), .ZN(n11953) );
  NAND2_X1 U11833 ( .A1(n11957), .A2(n11958), .ZN(n11698) );
  NAND2_X1 U11834 ( .A1(n11714), .A2(n11959), .ZN(n11958) );
  OR2_X1 U11835 ( .A1(n11715), .A2(n11716), .ZN(n11959) );
  NOR2_X1 U11836 ( .A1(n8943), .A2(n8041), .ZN(n11714) );
  NAND2_X1 U11837 ( .A1(n11716), .A2(n11715), .ZN(n11957) );
  NAND2_X1 U11838 ( .A1(n11960), .A2(n11961), .ZN(n11715) );
  NAND2_X1 U11839 ( .A1(b_18_), .A2(n11962), .ZN(n11961) );
  NAND2_X1 U11840 ( .A1(n8003), .A2(n11963), .ZN(n11962) );
  NAND2_X1 U11841 ( .A1(a_31_), .A2(n8945), .ZN(n11963) );
  NAND2_X1 U11842 ( .A1(b_19_), .A2(n11964), .ZN(n11960) );
  NAND2_X1 U11843 ( .A1(n9341), .A2(n11965), .ZN(n11964) );
  NAND2_X1 U11844 ( .A1(a_30_), .A2(n8946), .ZN(n11965) );
  AND2_X1 U11845 ( .A1(n11966), .A2(n7953), .ZN(n11716) );
  NOR2_X1 U11846 ( .A1(n8943), .A2(n8945), .ZN(n11966) );
  XOR2_X1 U11847 ( .A(n11967), .B(n11968), .Z(n11696) );
  XOR2_X1 U11848 ( .A(n11969), .B(n11970), .Z(n11967) );
  XNOR2_X1 U11849 ( .A(n11971), .B(n11972), .ZN(n11721) );
  NAND2_X1 U11850 ( .A1(n11973), .A2(n11974), .ZN(n11971) );
  XNOR2_X1 U11851 ( .A(n11975), .B(n11976), .ZN(n11726) );
  XNOR2_X1 U11852 ( .A(n11977), .B(n11978), .ZN(n11976) );
  XOR2_X1 U11853 ( .A(n11979), .B(n11980), .Z(n11729) );
  XOR2_X1 U11854 ( .A(n11981), .B(n11982), .Z(n11979) );
  NOR2_X1 U11855 ( .A1(n8939), .A2(n8945), .ZN(n11982) );
  XNOR2_X1 U11856 ( .A(n11983), .B(n11984), .ZN(n11734) );
  XNOR2_X1 U11857 ( .A(n11985), .B(n11986), .ZN(n11984) );
  XOR2_X1 U11858 ( .A(n11987), .B(n11988), .Z(n11737) );
  XOR2_X1 U11859 ( .A(n11989), .B(n11990), .Z(n11987) );
  NOR2_X1 U11860 ( .A1(n8941), .A2(n8945), .ZN(n11990) );
  INV_X1 U11861 ( .A(n8302), .ZN(n11744) );
  NAND2_X1 U11862 ( .A1(b_20_), .A2(a_20_), .ZN(n8302) );
  XOR2_X1 U11863 ( .A(n11991), .B(n11992), .Z(n11745) );
  XOR2_X1 U11864 ( .A(n11993), .B(n11994), .Z(n11991) );
  NOR2_X1 U11865 ( .A1(n8944), .A2(n8945), .ZN(n11994) );
  XOR2_X1 U11866 ( .A(n11995), .B(n11996), .Z(n11749) );
  XOR2_X1 U11867 ( .A(n11997), .B(n11998), .Z(n11995) );
  XNOR2_X1 U11868 ( .A(n11999), .B(n12000), .ZN(n11754) );
  XOR2_X1 U11869 ( .A(n12001), .B(n12002), .Z(n12000) );
  NAND2_X1 U11870 ( .A1(b_19_), .A2(a_18_), .ZN(n12002) );
  XOR2_X1 U11871 ( .A(n12003), .B(n12004), .Z(n11757) );
  XOR2_X1 U11872 ( .A(n12005), .B(n12006), .Z(n12003) );
  XOR2_X1 U11873 ( .A(n12007), .B(n12008), .Z(n11762) );
  XOR2_X1 U11874 ( .A(n12009), .B(n12010), .Z(n12007) );
  NOR2_X1 U11875 ( .A1(n8950), .A2(n8945), .ZN(n12010) );
  XOR2_X1 U11876 ( .A(n12011), .B(n12012), .Z(n11766) );
  XOR2_X1 U11877 ( .A(n12013), .B(n12014), .Z(n12011) );
  XNOR2_X1 U11878 ( .A(n12015), .B(n12016), .ZN(n11770) );
  XOR2_X1 U11879 ( .A(n12017), .B(n12018), .Z(n12016) );
  NAND2_X1 U11880 ( .A1(b_19_), .A2(a_14_), .ZN(n12018) );
  XOR2_X1 U11881 ( .A(n12019), .B(n12020), .Z(n11773) );
  XOR2_X1 U11882 ( .A(n12021), .B(n12022), .Z(n12019) );
  XOR2_X1 U11883 ( .A(n12023), .B(n12024), .Z(n11778) );
  XOR2_X1 U11884 ( .A(n12025), .B(n12026), .Z(n12023) );
  XNOR2_X1 U11885 ( .A(n12027), .B(n12028), .ZN(n11782) );
  XOR2_X1 U11886 ( .A(n12029), .B(n12030), .Z(n12027) );
  NOR2_X1 U11887 ( .A1(n8550), .A2(n8945), .ZN(n12030) );
  XOR2_X1 U11888 ( .A(n12031), .B(n12032), .Z(n11786) );
  XOR2_X1 U11889 ( .A(n12033), .B(n12034), .Z(n12031) );
  NOR2_X1 U11890 ( .A1(n8959), .A2(n8945), .ZN(n12034) );
  XOR2_X1 U11891 ( .A(n12035), .B(n12036), .Z(n11789) );
  XOR2_X1 U11892 ( .A(n12037), .B(n12038), .Z(n12035) );
  NOR2_X1 U11893 ( .A1(n8605), .A2(n8945), .ZN(n12038) );
  XOR2_X1 U11894 ( .A(n12039), .B(n12040), .Z(n11793) );
  XOR2_X1 U11895 ( .A(n12041), .B(n12042), .Z(n12039) );
  NOR2_X1 U11896 ( .A1(n8619), .A2(n8945), .ZN(n12042) );
  XNOR2_X1 U11897 ( .A(n12043), .B(n12044), .ZN(n11806) );
  XOR2_X1 U11898 ( .A(n12045), .B(n12046), .Z(n12043) );
  NOR2_X1 U11899 ( .A1(n8723), .A2(n8945), .ZN(n12046) );
  XOR2_X1 U11900 ( .A(n12047), .B(n12048), .Z(n11809) );
  XOR2_X1 U11901 ( .A(n12049), .B(n12050), .Z(n12047) );
  NOR2_X1 U11902 ( .A1(n8966), .A2(n8945), .ZN(n12050) );
  XOR2_X1 U11903 ( .A(n12051), .B(n12052), .Z(n11818) );
  NAND2_X1 U11904 ( .A1(n12053), .A2(n12054), .ZN(n12051) );
  XOR2_X1 U11905 ( .A(n12055), .B(n12056), .Z(n11584) );
  XOR2_X1 U11906 ( .A(n12057), .B(n12058), .Z(n12055) );
  NOR2_X1 U11907 ( .A1(n8969), .A2(n8945), .ZN(n12058) );
  NAND2_X1 U11908 ( .A1(n12059), .A2(n12060), .ZN(n9067) );
  XOR2_X1 U11909 ( .A(n9163), .B(n12061), .Z(n12060) );
  AND2_X1 U11910 ( .A1(n9161), .A2(n9160), .ZN(n12059) );
  XNOR2_X1 U11911 ( .A(n12062), .B(n12063), .ZN(n9160) );
  NAND2_X1 U11912 ( .A1(n12064), .A2(n12065), .ZN(n12062) );
  NAND2_X1 U11913 ( .A1(n12066), .A2(n12067), .ZN(n9161) );
  NAND2_X1 U11914 ( .A1(n12068), .A2(b_19_), .ZN(n12067) );
  NOR2_X1 U11915 ( .A1(n12069), .A2(n8974), .ZN(n12068) );
  NOR2_X1 U11916 ( .A1(n11827), .A2(n11828), .ZN(n12069) );
  NAND2_X1 U11917 ( .A1(n11827), .A2(n11828), .ZN(n12066) );
  NAND2_X1 U11918 ( .A1(n12070), .A2(n12071), .ZN(n11828) );
  NAND2_X1 U11919 ( .A1(n12072), .A2(b_19_), .ZN(n12071) );
  NOR2_X1 U11920 ( .A1(n12073), .A2(n8969), .ZN(n12072) );
  NOR2_X1 U11921 ( .A1(n12056), .A2(n12057), .ZN(n12073) );
  NAND2_X1 U11922 ( .A1(n12056), .A2(n12057), .ZN(n12070) );
  NAND2_X1 U11923 ( .A1(n12053), .A2(n12074), .ZN(n12057) );
  NAND2_X1 U11924 ( .A1(n12052), .A2(n12054), .ZN(n12074) );
  NAND2_X1 U11925 ( .A1(n12075), .A2(n12076), .ZN(n12054) );
  NAND2_X1 U11926 ( .A1(b_19_), .A2(a_2_), .ZN(n12076) );
  INV_X1 U11927 ( .A(n12077), .ZN(n12075) );
  XNOR2_X1 U11928 ( .A(n12078), .B(n12079), .ZN(n12052) );
  NAND2_X1 U11929 ( .A1(n12080), .A2(n12081), .ZN(n12078) );
  NAND2_X1 U11930 ( .A1(a_2_), .A2(n12077), .ZN(n12053) );
  NAND2_X1 U11931 ( .A1(n12082), .A2(n12083), .ZN(n12077) );
  NAND2_X1 U11932 ( .A1(n12084), .A2(b_19_), .ZN(n12083) );
  NOR2_X1 U11933 ( .A1(n12085), .A2(n8778), .ZN(n12084) );
  NOR2_X1 U11934 ( .A1(n11842), .A2(n11843), .ZN(n12085) );
  NAND2_X1 U11935 ( .A1(n11842), .A2(n11843), .ZN(n12082) );
  NAND2_X1 U11936 ( .A1(n12086), .A2(n12087), .ZN(n11843) );
  NAND2_X1 U11937 ( .A1(n12088), .A2(b_19_), .ZN(n12087) );
  NOR2_X1 U11938 ( .A1(n12089), .A2(n8966), .ZN(n12088) );
  NOR2_X1 U11939 ( .A1(n12048), .A2(n12049), .ZN(n12089) );
  NAND2_X1 U11940 ( .A1(n12048), .A2(n12049), .ZN(n12086) );
  NAND2_X1 U11941 ( .A1(n12090), .A2(n12091), .ZN(n12049) );
  NAND2_X1 U11942 ( .A1(n12092), .A2(b_19_), .ZN(n12091) );
  NOR2_X1 U11943 ( .A1(n12093), .A2(n8723), .ZN(n12092) );
  NOR2_X1 U11944 ( .A1(n12044), .A2(n12045), .ZN(n12093) );
  NAND2_X1 U11945 ( .A1(n12044), .A2(n12045), .ZN(n12090) );
  NAND2_X1 U11946 ( .A1(n12094), .A2(n12095), .ZN(n12045) );
  NAND2_X1 U11947 ( .A1(n12096), .A2(b_19_), .ZN(n12095) );
  NOR2_X1 U11948 ( .A1(n12097), .A2(n8681), .ZN(n12096) );
  NOR2_X1 U11949 ( .A1(n11857), .A2(n11858), .ZN(n12097) );
  NAND2_X1 U11950 ( .A1(n11857), .A2(n11858), .ZN(n12094) );
  NAND2_X1 U11951 ( .A1(n12098), .A2(n12099), .ZN(n11858) );
  NAND2_X1 U11952 ( .A1(n12100), .A2(b_19_), .ZN(n12099) );
  NOR2_X1 U11953 ( .A1(n12101), .A2(n8962), .ZN(n12100) );
  NOR2_X1 U11954 ( .A1(n11865), .A2(n11866), .ZN(n12101) );
  NAND2_X1 U11955 ( .A1(n11865), .A2(n11866), .ZN(n12098) );
  NAND2_X1 U11956 ( .A1(n12102), .A2(n12103), .ZN(n11866) );
  NAND2_X1 U11957 ( .A1(n12104), .A2(b_19_), .ZN(n12103) );
  NOR2_X1 U11958 ( .A1(n12105), .A2(n8619), .ZN(n12104) );
  NOR2_X1 U11959 ( .A1(n12040), .A2(n12041), .ZN(n12105) );
  NAND2_X1 U11960 ( .A1(n12040), .A2(n12041), .ZN(n12102) );
  NAND2_X1 U11961 ( .A1(n12106), .A2(n12107), .ZN(n12041) );
  NAND2_X1 U11962 ( .A1(n12108), .A2(b_19_), .ZN(n12107) );
  NOR2_X1 U11963 ( .A1(n12109), .A2(n8605), .ZN(n12108) );
  NOR2_X1 U11964 ( .A1(n12036), .A2(n12037), .ZN(n12109) );
  NAND2_X1 U11965 ( .A1(n12036), .A2(n12037), .ZN(n12106) );
  NAND2_X1 U11966 ( .A1(n12110), .A2(n12111), .ZN(n12037) );
  NAND2_X1 U11967 ( .A1(n12112), .A2(b_19_), .ZN(n12111) );
  NOR2_X1 U11968 ( .A1(n12113), .A2(n8959), .ZN(n12112) );
  NOR2_X1 U11969 ( .A1(n12032), .A2(n12033), .ZN(n12113) );
  NAND2_X1 U11970 ( .A1(n12032), .A2(n12033), .ZN(n12110) );
  NAND2_X1 U11971 ( .A1(n12114), .A2(n12115), .ZN(n12033) );
  NAND2_X1 U11972 ( .A1(n12116), .A2(b_19_), .ZN(n12115) );
  NOR2_X1 U11973 ( .A1(n12117), .A2(n8550), .ZN(n12116) );
  NOR2_X1 U11974 ( .A1(n12028), .A2(n12029), .ZN(n12117) );
  NAND2_X1 U11975 ( .A1(n12028), .A2(n12029), .ZN(n12114) );
  NAND2_X1 U11976 ( .A1(n12118), .A2(n12119), .ZN(n12029) );
  NAND2_X1 U11977 ( .A1(n12026), .A2(n12120), .ZN(n12119) );
  OR2_X1 U11978 ( .A1(n12025), .A2(n12024), .ZN(n12120) );
  NOR2_X1 U11979 ( .A1(n8945), .A2(n8956), .ZN(n12026) );
  NAND2_X1 U11980 ( .A1(n12024), .A2(n12025), .ZN(n12118) );
  NAND2_X1 U11981 ( .A1(n12121), .A2(n12122), .ZN(n12025) );
  NAND2_X1 U11982 ( .A1(n12022), .A2(n12123), .ZN(n12122) );
  OR2_X1 U11983 ( .A1(n12021), .A2(n12020), .ZN(n12123) );
  NOR2_X1 U11984 ( .A1(n8945), .A2(n8495), .ZN(n12022) );
  NAND2_X1 U11985 ( .A1(n12020), .A2(n12021), .ZN(n12121) );
  NAND2_X1 U11986 ( .A1(n12124), .A2(n12125), .ZN(n12021) );
  NAND2_X1 U11987 ( .A1(n12126), .A2(b_19_), .ZN(n12125) );
  NOR2_X1 U11988 ( .A1(n12127), .A2(n8953), .ZN(n12126) );
  NOR2_X1 U11989 ( .A1(n12015), .A2(n12017), .ZN(n12127) );
  NAND2_X1 U11990 ( .A1(n12015), .A2(n12017), .ZN(n12124) );
  NAND2_X1 U11991 ( .A1(n12128), .A2(n12129), .ZN(n12017) );
  NAND2_X1 U11992 ( .A1(n12014), .A2(n12130), .ZN(n12129) );
  OR2_X1 U11993 ( .A1(n12013), .A2(n12012), .ZN(n12130) );
  NOR2_X1 U11994 ( .A1(n8945), .A2(n8440), .ZN(n12014) );
  NAND2_X1 U11995 ( .A1(n12012), .A2(n12013), .ZN(n12128) );
  NAND2_X1 U11996 ( .A1(n12131), .A2(n12132), .ZN(n12013) );
  NAND2_X1 U11997 ( .A1(n12133), .A2(b_19_), .ZN(n12132) );
  NOR2_X1 U11998 ( .A1(n12134), .A2(n8950), .ZN(n12133) );
  NOR2_X1 U11999 ( .A1(n12008), .A2(n12009), .ZN(n12134) );
  NAND2_X1 U12000 ( .A1(n12008), .A2(n12009), .ZN(n12131) );
  NAND2_X1 U12001 ( .A1(n12135), .A2(n12136), .ZN(n12009) );
  NAND2_X1 U12002 ( .A1(n12006), .A2(n12137), .ZN(n12136) );
  OR2_X1 U12003 ( .A1(n12005), .A2(n12004), .ZN(n12137) );
  NOR2_X1 U12004 ( .A1(n8945), .A2(n8385), .ZN(n12006) );
  NAND2_X1 U12005 ( .A1(n12004), .A2(n12005), .ZN(n12135) );
  NAND2_X1 U12006 ( .A1(n12138), .A2(n12139), .ZN(n12005) );
  NAND2_X1 U12007 ( .A1(n12140), .A2(b_19_), .ZN(n12139) );
  NOR2_X1 U12008 ( .A1(n12141), .A2(n8947), .ZN(n12140) );
  NOR2_X1 U12009 ( .A1(n11999), .A2(n12001), .ZN(n12141) );
  NAND2_X1 U12010 ( .A1(n11999), .A2(n12001), .ZN(n12138) );
  NAND2_X1 U12011 ( .A1(n12142), .A2(n12143), .ZN(n12001) );
  NAND2_X1 U12012 ( .A1(n11998), .A2(n12144), .ZN(n12143) );
  OR2_X1 U12013 ( .A1(n11997), .A2(n11996), .ZN(n12144) );
  INV_X1 U12014 ( .A(n8901), .ZN(n11998) );
  NAND2_X1 U12015 ( .A1(b_19_), .A2(a_19_), .ZN(n8901) );
  NAND2_X1 U12016 ( .A1(n11996), .A2(n11997), .ZN(n12142) );
  NAND2_X1 U12017 ( .A1(n12145), .A2(n12146), .ZN(n11997) );
  NAND2_X1 U12018 ( .A1(n12147), .A2(b_19_), .ZN(n12146) );
  NOR2_X1 U12019 ( .A1(n12148), .A2(n8944), .ZN(n12147) );
  NOR2_X1 U12020 ( .A1(n11992), .A2(n11993), .ZN(n12148) );
  NAND2_X1 U12021 ( .A1(n11992), .A2(n11993), .ZN(n12145) );
  NAND2_X1 U12022 ( .A1(n12149), .A2(n12150), .ZN(n11993) );
  NAND2_X1 U12023 ( .A1(n11919), .A2(n12151), .ZN(n12150) );
  OR2_X1 U12024 ( .A1(n11918), .A2(n11916), .ZN(n12151) );
  NOR2_X1 U12025 ( .A1(n8945), .A2(n8268), .ZN(n11919) );
  NAND2_X1 U12026 ( .A1(n11916), .A2(n11918), .ZN(n12149) );
  NAND2_X1 U12027 ( .A1(n12152), .A2(n12153), .ZN(n11918) );
  NAND2_X1 U12028 ( .A1(n12154), .A2(b_19_), .ZN(n12153) );
  NOR2_X1 U12029 ( .A1(n12155), .A2(n8941), .ZN(n12154) );
  NOR2_X1 U12030 ( .A1(n11988), .A2(n11989), .ZN(n12155) );
  NAND2_X1 U12031 ( .A1(n11988), .A2(n11989), .ZN(n12152) );
  NAND2_X1 U12032 ( .A1(n12156), .A2(n12157), .ZN(n11989) );
  NAND2_X1 U12033 ( .A1(n11986), .A2(n12158), .ZN(n12157) );
  OR2_X1 U12034 ( .A1(n11985), .A2(n11983), .ZN(n12158) );
  NOR2_X1 U12035 ( .A1(n8945), .A2(n8213), .ZN(n11986) );
  NAND2_X1 U12036 ( .A1(n11983), .A2(n11985), .ZN(n12156) );
  NAND2_X1 U12037 ( .A1(n12159), .A2(n12160), .ZN(n11985) );
  NAND2_X1 U12038 ( .A1(n12161), .A2(b_19_), .ZN(n12160) );
  NOR2_X1 U12039 ( .A1(n12162), .A2(n8939), .ZN(n12161) );
  NOR2_X1 U12040 ( .A1(n11980), .A2(n11981), .ZN(n12162) );
  NAND2_X1 U12041 ( .A1(n11980), .A2(n11981), .ZN(n12159) );
  NAND2_X1 U12042 ( .A1(n12163), .A2(n12164), .ZN(n11981) );
  NAND2_X1 U12043 ( .A1(n11978), .A2(n12165), .ZN(n12164) );
  OR2_X1 U12044 ( .A1(n11977), .A2(n11975), .ZN(n12165) );
  NOR2_X1 U12045 ( .A1(n8945), .A2(n8158), .ZN(n11978) );
  NAND2_X1 U12046 ( .A1(n11975), .A2(n11977), .ZN(n12163) );
  NAND2_X1 U12047 ( .A1(n11973), .A2(n12166), .ZN(n11977) );
  NAND2_X1 U12048 ( .A1(n11972), .A2(n11974), .ZN(n12166) );
  NAND2_X1 U12049 ( .A1(n12167), .A2(n12168), .ZN(n11974) );
  NAND2_X1 U12050 ( .A1(b_19_), .A2(a_26_), .ZN(n12168) );
  INV_X1 U12051 ( .A(n12169), .ZN(n12167) );
  XNOR2_X1 U12052 ( .A(n12170), .B(n12171), .ZN(n11972) );
  NAND2_X1 U12053 ( .A1(n12172), .A2(n12173), .ZN(n12170) );
  NAND2_X1 U12054 ( .A1(a_26_), .A2(n12169), .ZN(n11973) );
  NAND2_X1 U12055 ( .A1(n11943), .A2(n12174), .ZN(n12169) );
  NAND2_X1 U12056 ( .A1(n11942), .A2(n11944), .ZN(n12174) );
  NAND2_X1 U12057 ( .A1(n12175), .A2(n12176), .ZN(n11944) );
  NAND2_X1 U12058 ( .A1(b_19_), .A2(a_27_), .ZN(n12176) );
  INV_X1 U12059 ( .A(n12177), .ZN(n12175) );
  XOR2_X1 U12060 ( .A(n12178), .B(n12179), .Z(n11942) );
  XNOR2_X1 U12061 ( .A(n12180), .B(n12181), .ZN(n12178) );
  NAND2_X1 U12062 ( .A1(b_18_), .A2(a_28_), .ZN(n12180) );
  NAND2_X1 U12063 ( .A1(a_27_), .A2(n12177), .ZN(n11943) );
  NAND2_X1 U12064 ( .A1(n12182), .A2(n12183), .ZN(n12177) );
  NAND2_X1 U12065 ( .A1(n12184), .A2(b_19_), .ZN(n12183) );
  NOR2_X1 U12066 ( .A1(n12185), .A2(n8055), .ZN(n12184) );
  NOR2_X1 U12067 ( .A1(n11950), .A2(n11952), .ZN(n12185) );
  NAND2_X1 U12068 ( .A1(n11950), .A2(n11952), .ZN(n12182) );
  NAND2_X1 U12069 ( .A1(n12186), .A2(n12187), .ZN(n11952) );
  NAND2_X1 U12070 ( .A1(n11968), .A2(n12188), .ZN(n12187) );
  OR2_X1 U12071 ( .A1(n11969), .A2(n11970), .ZN(n12188) );
  NOR2_X1 U12072 ( .A1(n8945), .A2(n8041), .ZN(n11968) );
  NAND2_X1 U12073 ( .A1(n11970), .A2(n11969), .ZN(n12186) );
  NAND2_X1 U12074 ( .A1(n12189), .A2(n12190), .ZN(n11969) );
  NAND2_X1 U12075 ( .A1(b_17_), .A2(n12191), .ZN(n12190) );
  NAND2_X1 U12076 ( .A1(n8003), .A2(n12192), .ZN(n12191) );
  NAND2_X1 U12077 ( .A1(a_31_), .A2(n8946), .ZN(n12192) );
  NAND2_X1 U12078 ( .A1(b_18_), .A2(n12193), .ZN(n12189) );
  NAND2_X1 U12079 ( .A1(n9341), .A2(n12194), .ZN(n12193) );
  NAND2_X1 U12080 ( .A1(a_30_), .A2(n8948), .ZN(n12194) );
  AND2_X1 U12081 ( .A1(n12195), .A2(n7953), .ZN(n11970) );
  NOR2_X1 U12082 ( .A1(n8945), .A2(n8946), .ZN(n12195) );
  XOR2_X1 U12083 ( .A(n12196), .B(n12197), .Z(n11950) );
  XOR2_X1 U12084 ( .A(n12198), .B(n12199), .Z(n12196) );
  XNOR2_X1 U12085 ( .A(n12200), .B(n12201), .ZN(n11975) );
  NAND2_X1 U12086 ( .A1(n12202), .A2(n12203), .ZN(n12200) );
  XNOR2_X1 U12087 ( .A(n12204), .B(n12205), .ZN(n11980) );
  XNOR2_X1 U12088 ( .A(n12206), .B(n12207), .ZN(n12205) );
  XOR2_X1 U12089 ( .A(n12208), .B(n12209), .Z(n11983) );
  XOR2_X1 U12090 ( .A(n12210), .B(n12211), .Z(n12208) );
  NOR2_X1 U12091 ( .A1(n8939), .A2(n8946), .ZN(n12211) );
  XNOR2_X1 U12092 ( .A(n12212), .B(n12213), .ZN(n11988) );
  XOR2_X1 U12093 ( .A(n12214), .B(n12215), .Z(n12213) );
  NAND2_X1 U12094 ( .A1(b_18_), .A2(a_23_), .ZN(n12215) );
  XNOR2_X1 U12095 ( .A(n12216), .B(n12217), .ZN(n11916) );
  NAND2_X1 U12096 ( .A1(n12218), .A2(n12219), .ZN(n12216) );
  XOR2_X1 U12097 ( .A(n12220), .B(n12221), .Z(n11992) );
  XOR2_X1 U12098 ( .A(n12222), .B(n12223), .Z(n12220) );
  XOR2_X1 U12099 ( .A(n12224), .B(n12225), .Z(n11996) );
  XOR2_X1 U12100 ( .A(n12226), .B(n12227), .Z(n12224) );
  NOR2_X1 U12101 ( .A1(n8944), .A2(n8946), .ZN(n12227) );
  XNOR2_X1 U12102 ( .A(n12228), .B(n12229), .ZN(n11999) );
  XNOR2_X1 U12103 ( .A(n12230), .B(n12231), .ZN(n12229) );
  XOR2_X1 U12104 ( .A(n12232), .B(n12233), .Z(n12004) );
  XOR2_X1 U12105 ( .A(n12234), .B(n12235), .Z(n12232) );
  XNOR2_X1 U12106 ( .A(n12236), .B(n12237), .ZN(n12008) );
  XNOR2_X1 U12107 ( .A(n12238), .B(n12239), .ZN(n12237) );
  XNOR2_X1 U12108 ( .A(n12240), .B(n12241), .ZN(n12012) );
  XOR2_X1 U12109 ( .A(n12242), .B(n12243), .Z(n12241) );
  NAND2_X1 U12110 ( .A1(b_18_), .A2(a_16_), .ZN(n12243) );
  XOR2_X1 U12111 ( .A(n12244), .B(n12245), .Z(n12015) );
  XOR2_X1 U12112 ( .A(n12246), .B(n12247), .Z(n12244) );
  XOR2_X1 U12113 ( .A(n12248), .B(n12249), .Z(n12020) );
  XOR2_X1 U12114 ( .A(n12250), .B(n12251), .Z(n12248) );
  NOR2_X1 U12115 ( .A1(n8953), .A2(n8946), .ZN(n12251) );
  XOR2_X1 U12116 ( .A(n12252), .B(n12253), .Z(n12024) );
  XOR2_X1 U12117 ( .A(n12254), .B(n12255), .Z(n12252) );
  NOR2_X1 U12118 ( .A1(n8495), .A2(n8946), .ZN(n12255) );
  XNOR2_X1 U12119 ( .A(n12256), .B(n12257), .ZN(n12028) );
  XNOR2_X1 U12120 ( .A(n12258), .B(n12259), .ZN(n12256) );
  XOR2_X1 U12121 ( .A(n12260), .B(n12261), .Z(n12032) );
  XOR2_X1 U12122 ( .A(n12262), .B(n12263), .Z(n12260) );
  XNOR2_X1 U12123 ( .A(n12264), .B(n12265), .ZN(n12036) );
  XNOR2_X1 U12124 ( .A(n12266), .B(n12267), .ZN(n12265) );
  XNOR2_X1 U12125 ( .A(n12268), .B(n12269), .ZN(n12040) );
  XOR2_X1 U12126 ( .A(n12270), .B(n12271), .Z(n12269) );
  NAND2_X1 U12127 ( .A1(b_18_), .A2(a_9_), .ZN(n12271) );
  XNOR2_X1 U12128 ( .A(n12272), .B(n12273), .ZN(n11865) );
  NAND2_X1 U12129 ( .A1(n12274), .A2(n12275), .ZN(n12272) );
  XNOR2_X1 U12130 ( .A(n12276), .B(n12277), .ZN(n11857) );
  NAND2_X1 U12131 ( .A1(n12278), .A2(n12279), .ZN(n12276) );
  XNOR2_X1 U12132 ( .A(n12280), .B(n12281), .ZN(n12044) );
  XNOR2_X1 U12133 ( .A(n12282), .B(n12283), .ZN(n12280) );
  XOR2_X1 U12134 ( .A(n12284), .B(n12285), .Z(n12048) );
  XOR2_X1 U12135 ( .A(n12286), .B(n12287), .Z(n12284) );
  NOR2_X1 U12136 ( .A1(n8723), .A2(n8946), .ZN(n12287) );
  XNOR2_X1 U12137 ( .A(n12288), .B(n12289), .ZN(n11842) );
  NAND2_X1 U12138 ( .A1(n12290), .A2(n12291), .ZN(n12288) );
  XNOR2_X1 U12139 ( .A(n12292), .B(n12293), .ZN(n12056) );
  NAND2_X1 U12140 ( .A1(n12294), .A2(n12295), .ZN(n12292) );
  XOR2_X1 U12141 ( .A(n12296), .B(n12297), .Z(n11827) );
  NOR2_X1 U12142 ( .A1(n12298), .A2(n12299), .ZN(n12297) );
  NOR2_X1 U12143 ( .A1(n12300), .A2(n12301), .ZN(n12298) );
  NOR2_X1 U12144 ( .A1(n8969), .A2(n8946), .ZN(n12300) );
  NAND2_X1 U12145 ( .A1(n12302), .A2(n12303), .ZN(n9073) );
  NAND2_X1 U12146 ( .A1(n12304), .A2(n9162), .ZN(n12303) );
  INV_X1 U12147 ( .A(n9163), .ZN(n12304) );
  XOR2_X1 U12148 ( .A(n9153), .B(n12305), .Z(n12302) );
  NAND2_X1 U12149 ( .A1(n12306), .A2(n12307), .ZN(n9074) );
  XOR2_X1 U12150 ( .A(n9153), .B(n9152), .Z(n12307) );
  NOR2_X1 U12151 ( .A1(n12061), .A2(n9163), .ZN(n12306) );
  XNOR2_X1 U12152 ( .A(n12308), .B(n12309), .ZN(n9163) );
  XOR2_X1 U12153 ( .A(n12310), .B(n12311), .Z(n12308) );
  NOR2_X1 U12154 ( .A1(n8974), .A2(n8948), .ZN(n12311) );
  INV_X1 U12155 ( .A(n9162), .ZN(n12061) );
  NAND2_X1 U12156 ( .A1(n12064), .A2(n12312), .ZN(n9162) );
  NAND2_X1 U12157 ( .A1(n12063), .A2(n12065), .ZN(n12312) );
  NAND2_X1 U12158 ( .A1(n12313), .A2(n12314), .ZN(n12065) );
  NAND2_X1 U12159 ( .A1(b_18_), .A2(a_0_), .ZN(n12314) );
  XOR2_X1 U12160 ( .A(n12315), .B(n12316), .Z(n12063) );
  XOR2_X1 U12161 ( .A(n12317), .B(n12318), .Z(n12315) );
  NOR2_X1 U12162 ( .A1(n8969), .A2(n8948), .ZN(n12318) );
  OR2_X1 U12163 ( .A1(n8974), .A2(n12313), .ZN(n12064) );
  NOR2_X1 U12164 ( .A1(n12299), .A2(n12319), .ZN(n12313) );
  AND2_X1 U12165 ( .A1(n12296), .A2(n12320), .ZN(n12319) );
  NAND2_X1 U12166 ( .A1(n12321), .A2(n12322), .ZN(n12320) );
  NAND2_X1 U12167 ( .A1(b_18_), .A2(a_1_), .ZN(n12322) );
  XOR2_X1 U12168 ( .A(n12323), .B(n12324), .Z(n12296) );
  XOR2_X1 U12169 ( .A(n12325), .B(n12326), .Z(n12323) );
  NOR2_X1 U12170 ( .A1(n8792), .A2(n8948), .ZN(n12326) );
  NOR2_X1 U12171 ( .A1(n8969), .A2(n12321), .ZN(n12299) );
  INV_X1 U12172 ( .A(n12301), .ZN(n12321) );
  NAND2_X1 U12173 ( .A1(n12294), .A2(n12327), .ZN(n12301) );
  NAND2_X1 U12174 ( .A1(n12293), .A2(n12295), .ZN(n12327) );
  NAND2_X1 U12175 ( .A1(n12328), .A2(n12329), .ZN(n12295) );
  NAND2_X1 U12176 ( .A1(b_18_), .A2(a_2_), .ZN(n12329) );
  INV_X1 U12177 ( .A(n12330), .ZN(n12328) );
  XOR2_X1 U12178 ( .A(n12331), .B(n12332), .Z(n12293) );
  XOR2_X1 U12179 ( .A(n12333), .B(n12334), .Z(n12331) );
  NOR2_X1 U12180 ( .A1(n8778), .A2(n8948), .ZN(n12334) );
  NAND2_X1 U12181 ( .A1(a_2_), .A2(n12330), .ZN(n12294) );
  NAND2_X1 U12182 ( .A1(n12080), .A2(n12335), .ZN(n12330) );
  NAND2_X1 U12183 ( .A1(n12079), .A2(n12081), .ZN(n12335) );
  NAND2_X1 U12184 ( .A1(n12336), .A2(n12337), .ZN(n12081) );
  NAND2_X1 U12185 ( .A1(b_18_), .A2(a_3_), .ZN(n12337) );
  INV_X1 U12186 ( .A(n12338), .ZN(n12336) );
  XOR2_X1 U12187 ( .A(n12339), .B(n12340), .Z(n12079) );
  XOR2_X1 U12188 ( .A(n12341), .B(n12342), .Z(n12339) );
  NOR2_X1 U12189 ( .A1(n8966), .A2(n8948), .ZN(n12342) );
  NAND2_X1 U12190 ( .A1(a_3_), .A2(n12338), .ZN(n12080) );
  NAND2_X1 U12191 ( .A1(n12290), .A2(n12343), .ZN(n12338) );
  NAND2_X1 U12192 ( .A1(n12289), .A2(n12291), .ZN(n12343) );
  NAND2_X1 U12193 ( .A1(n12344), .A2(n12345), .ZN(n12291) );
  NAND2_X1 U12194 ( .A1(b_18_), .A2(a_4_), .ZN(n12345) );
  INV_X1 U12195 ( .A(n12346), .ZN(n12344) );
  XOR2_X1 U12196 ( .A(n12347), .B(n12348), .Z(n12289) );
  XOR2_X1 U12197 ( .A(n12349), .B(n12350), .Z(n12347) );
  NOR2_X1 U12198 ( .A1(n8723), .A2(n8948), .ZN(n12350) );
  NAND2_X1 U12199 ( .A1(a_4_), .A2(n12346), .ZN(n12290) );
  NAND2_X1 U12200 ( .A1(n12351), .A2(n12352), .ZN(n12346) );
  NAND2_X1 U12201 ( .A1(n12353), .A2(b_18_), .ZN(n12352) );
  NOR2_X1 U12202 ( .A1(n12354), .A2(n8723), .ZN(n12353) );
  NOR2_X1 U12203 ( .A1(n12285), .A2(n12286), .ZN(n12354) );
  NAND2_X1 U12204 ( .A1(n12285), .A2(n12286), .ZN(n12351) );
  NAND2_X1 U12205 ( .A1(n12355), .A2(n12356), .ZN(n12286) );
  NAND2_X1 U12206 ( .A1(n12283), .A2(n12357), .ZN(n12356) );
  NAND2_X1 U12207 ( .A1(n12282), .A2(n12281), .ZN(n12357) );
  NOR2_X1 U12208 ( .A1(n8946), .A2(n8681), .ZN(n12283) );
  OR2_X1 U12209 ( .A1(n12281), .A2(n12282), .ZN(n12355) );
  AND2_X1 U12210 ( .A1(n12278), .A2(n12358), .ZN(n12282) );
  NAND2_X1 U12211 ( .A1(n12277), .A2(n12279), .ZN(n12358) );
  NAND2_X1 U12212 ( .A1(n12359), .A2(n12360), .ZN(n12279) );
  NAND2_X1 U12213 ( .A1(b_18_), .A2(a_7_), .ZN(n12360) );
  INV_X1 U12214 ( .A(n12361), .ZN(n12359) );
  XOR2_X1 U12215 ( .A(n12362), .B(n12363), .Z(n12277) );
  XOR2_X1 U12216 ( .A(n12364), .B(n12365), .Z(n12362) );
  NOR2_X1 U12217 ( .A1(n8619), .A2(n8948), .ZN(n12365) );
  NAND2_X1 U12218 ( .A1(a_7_), .A2(n12361), .ZN(n12278) );
  NAND2_X1 U12219 ( .A1(n12274), .A2(n12366), .ZN(n12361) );
  NAND2_X1 U12220 ( .A1(n12273), .A2(n12275), .ZN(n12366) );
  NAND2_X1 U12221 ( .A1(n12367), .A2(n12368), .ZN(n12275) );
  NAND2_X1 U12222 ( .A1(b_18_), .A2(a_8_), .ZN(n12368) );
  INV_X1 U12223 ( .A(n12369), .ZN(n12367) );
  XNOR2_X1 U12224 ( .A(n12370), .B(n12371), .ZN(n12273) );
  XOR2_X1 U12225 ( .A(n12372), .B(n12373), .Z(n12371) );
  NAND2_X1 U12226 ( .A1(b_17_), .A2(a_9_), .ZN(n12373) );
  NAND2_X1 U12227 ( .A1(a_8_), .A2(n12369), .ZN(n12274) );
  NAND2_X1 U12228 ( .A1(n12374), .A2(n12375), .ZN(n12369) );
  NAND2_X1 U12229 ( .A1(n12376), .A2(b_18_), .ZN(n12375) );
  NOR2_X1 U12230 ( .A1(n12377), .A2(n8605), .ZN(n12376) );
  NOR2_X1 U12231 ( .A1(n12270), .A2(n12268), .ZN(n12377) );
  NAND2_X1 U12232 ( .A1(n12268), .A2(n12270), .ZN(n12374) );
  NAND2_X1 U12233 ( .A1(n12378), .A2(n12379), .ZN(n12270) );
  NAND2_X1 U12234 ( .A1(n12267), .A2(n12380), .ZN(n12379) );
  OR2_X1 U12235 ( .A1(n12266), .A2(n12264), .ZN(n12380) );
  NOR2_X1 U12236 ( .A1(n8946), .A2(n8959), .ZN(n12267) );
  NAND2_X1 U12237 ( .A1(n12264), .A2(n12266), .ZN(n12378) );
  NAND2_X1 U12238 ( .A1(n12381), .A2(n12382), .ZN(n12266) );
  NAND2_X1 U12239 ( .A1(n12263), .A2(n12383), .ZN(n12382) );
  OR2_X1 U12240 ( .A1(n12261), .A2(n12262), .ZN(n12383) );
  NOR2_X1 U12241 ( .A1(n8946), .A2(n8550), .ZN(n12263) );
  NAND2_X1 U12242 ( .A1(n12261), .A2(n12262), .ZN(n12381) );
  NAND2_X1 U12243 ( .A1(n12384), .A2(n12385), .ZN(n12262) );
  NAND2_X1 U12244 ( .A1(n12259), .A2(n12386), .ZN(n12385) );
  NAND2_X1 U12245 ( .A1(n12258), .A2(n12257), .ZN(n12386) );
  NOR2_X1 U12246 ( .A1(n8946), .A2(n8956), .ZN(n12259) );
  OR2_X1 U12247 ( .A1(n12257), .A2(n12258), .ZN(n12384) );
  AND2_X1 U12248 ( .A1(n12387), .A2(n12388), .ZN(n12258) );
  NAND2_X1 U12249 ( .A1(n12389), .A2(b_18_), .ZN(n12388) );
  NOR2_X1 U12250 ( .A1(n12390), .A2(n8495), .ZN(n12389) );
  NOR2_X1 U12251 ( .A1(n12253), .A2(n12254), .ZN(n12390) );
  NAND2_X1 U12252 ( .A1(n12253), .A2(n12254), .ZN(n12387) );
  NAND2_X1 U12253 ( .A1(n12391), .A2(n12392), .ZN(n12254) );
  NAND2_X1 U12254 ( .A1(n12393), .A2(b_18_), .ZN(n12392) );
  NOR2_X1 U12255 ( .A1(n12394), .A2(n8953), .ZN(n12393) );
  NOR2_X1 U12256 ( .A1(n12249), .A2(n12250), .ZN(n12394) );
  NAND2_X1 U12257 ( .A1(n12249), .A2(n12250), .ZN(n12391) );
  NAND2_X1 U12258 ( .A1(n12395), .A2(n12396), .ZN(n12250) );
  NAND2_X1 U12259 ( .A1(n12247), .A2(n12397), .ZN(n12396) );
  OR2_X1 U12260 ( .A1(n12245), .A2(n12246), .ZN(n12397) );
  NOR2_X1 U12261 ( .A1(n8946), .A2(n8440), .ZN(n12247) );
  NAND2_X1 U12262 ( .A1(n12245), .A2(n12246), .ZN(n12395) );
  NAND2_X1 U12263 ( .A1(n12398), .A2(n12399), .ZN(n12246) );
  NAND2_X1 U12264 ( .A1(n12400), .A2(b_18_), .ZN(n12399) );
  NOR2_X1 U12265 ( .A1(n12401), .A2(n8950), .ZN(n12400) );
  NOR2_X1 U12266 ( .A1(n12240), .A2(n12242), .ZN(n12401) );
  NAND2_X1 U12267 ( .A1(n12240), .A2(n12242), .ZN(n12398) );
  NAND2_X1 U12268 ( .A1(n12402), .A2(n12403), .ZN(n12242) );
  NAND2_X1 U12269 ( .A1(n12239), .A2(n12404), .ZN(n12403) );
  OR2_X1 U12270 ( .A1(n12236), .A2(n12238), .ZN(n12404) );
  NOR2_X1 U12271 ( .A1(n8946), .A2(n8385), .ZN(n12239) );
  NAND2_X1 U12272 ( .A1(n12236), .A2(n12238), .ZN(n12402) );
  NAND2_X1 U12273 ( .A1(n12405), .A2(n12406), .ZN(n12238) );
  NAND2_X1 U12274 ( .A1(n12233), .A2(n12407), .ZN(n12406) );
  OR2_X1 U12275 ( .A1(n12234), .A2(n12235), .ZN(n12407) );
  XNOR2_X1 U12276 ( .A(n12408), .B(n12409), .ZN(n12233) );
  XNOR2_X1 U12277 ( .A(n12410), .B(n12411), .ZN(n12409) );
  NAND2_X1 U12278 ( .A1(n12235), .A2(n12234), .ZN(n12405) );
  NAND2_X1 U12279 ( .A1(n12412), .A2(n12413), .ZN(n12234) );
  NAND2_X1 U12280 ( .A1(n12231), .A2(n12414), .ZN(n12413) );
  OR2_X1 U12281 ( .A1(n12228), .A2(n12230), .ZN(n12414) );
  NOR2_X1 U12282 ( .A1(n8946), .A2(n8324), .ZN(n12231) );
  NAND2_X1 U12283 ( .A1(n12228), .A2(n12230), .ZN(n12412) );
  NAND2_X1 U12284 ( .A1(n12415), .A2(n12416), .ZN(n12230) );
  NAND2_X1 U12285 ( .A1(n12417), .A2(b_18_), .ZN(n12416) );
  NOR2_X1 U12286 ( .A1(n12418), .A2(n8944), .ZN(n12417) );
  NOR2_X1 U12287 ( .A1(n12225), .A2(n12226), .ZN(n12418) );
  NAND2_X1 U12288 ( .A1(n12225), .A2(n12226), .ZN(n12415) );
  NAND2_X1 U12289 ( .A1(n12419), .A2(n12420), .ZN(n12226) );
  NAND2_X1 U12290 ( .A1(n12223), .A2(n12421), .ZN(n12420) );
  OR2_X1 U12291 ( .A1(n12221), .A2(n12222), .ZN(n12421) );
  NOR2_X1 U12292 ( .A1(n8946), .A2(n8268), .ZN(n12223) );
  NAND2_X1 U12293 ( .A1(n12221), .A2(n12222), .ZN(n12419) );
  NAND2_X1 U12294 ( .A1(n12218), .A2(n12422), .ZN(n12222) );
  NAND2_X1 U12295 ( .A1(n12217), .A2(n12219), .ZN(n12422) );
  NAND2_X1 U12296 ( .A1(n12423), .A2(n12424), .ZN(n12219) );
  NAND2_X1 U12297 ( .A1(b_18_), .A2(a_22_), .ZN(n12424) );
  INV_X1 U12298 ( .A(n12425), .ZN(n12423) );
  XNOR2_X1 U12299 ( .A(n12426), .B(n12427), .ZN(n12217) );
  XNOR2_X1 U12300 ( .A(n12428), .B(n12429), .ZN(n12427) );
  NAND2_X1 U12301 ( .A1(a_22_), .A2(n12425), .ZN(n12218) );
  NAND2_X1 U12302 ( .A1(n12430), .A2(n12431), .ZN(n12425) );
  NAND2_X1 U12303 ( .A1(n12432), .A2(b_18_), .ZN(n12431) );
  NOR2_X1 U12304 ( .A1(n12433), .A2(n8213), .ZN(n12432) );
  NOR2_X1 U12305 ( .A1(n12214), .A2(n12212), .ZN(n12433) );
  NAND2_X1 U12306 ( .A1(n12212), .A2(n12214), .ZN(n12430) );
  NAND2_X1 U12307 ( .A1(n12434), .A2(n12435), .ZN(n12214) );
  NAND2_X1 U12308 ( .A1(n12436), .A2(b_18_), .ZN(n12435) );
  NOR2_X1 U12309 ( .A1(n12437), .A2(n8939), .ZN(n12436) );
  NOR2_X1 U12310 ( .A1(n12209), .A2(n12210), .ZN(n12437) );
  NAND2_X1 U12311 ( .A1(n12209), .A2(n12210), .ZN(n12434) );
  NAND2_X1 U12312 ( .A1(n12438), .A2(n12439), .ZN(n12210) );
  NAND2_X1 U12313 ( .A1(n12207), .A2(n12440), .ZN(n12439) );
  OR2_X1 U12314 ( .A1(n12204), .A2(n12206), .ZN(n12440) );
  NOR2_X1 U12315 ( .A1(n8946), .A2(n8158), .ZN(n12207) );
  NAND2_X1 U12316 ( .A1(n12204), .A2(n12206), .ZN(n12438) );
  NAND2_X1 U12317 ( .A1(n12202), .A2(n12441), .ZN(n12206) );
  NAND2_X1 U12318 ( .A1(n12201), .A2(n12203), .ZN(n12441) );
  NAND2_X1 U12319 ( .A1(n12442), .A2(n12443), .ZN(n12203) );
  NAND2_X1 U12320 ( .A1(b_18_), .A2(a_26_), .ZN(n12443) );
  INV_X1 U12321 ( .A(n12444), .ZN(n12442) );
  XNOR2_X1 U12322 ( .A(n12445), .B(n12446), .ZN(n12201) );
  NAND2_X1 U12323 ( .A1(n12447), .A2(n12448), .ZN(n12445) );
  NAND2_X1 U12324 ( .A1(a_26_), .A2(n12444), .ZN(n12202) );
  NAND2_X1 U12325 ( .A1(n12172), .A2(n12449), .ZN(n12444) );
  NAND2_X1 U12326 ( .A1(n12171), .A2(n12173), .ZN(n12449) );
  NAND2_X1 U12327 ( .A1(n12450), .A2(n12451), .ZN(n12173) );
  NAND2_X1 U12328 ( .A1(b_18_), .A2(a_27_), .ZN(n12451) );
  INV_X1 U12329 ( .A(n12452), .ZN(n12450) );
  XOR2_X1 U12330 ( .A(n12453), .B(n12454), .Z(n12171) );
  XNOR2_X1 U12331 ( .A(n12455), .B(n12456), .ZN(n12453) );
  NAND2_X1 U12332 ( .A1(b_17_), .A2(a_28_), .ZN(n12455) );
  NAND2_X1 U12333 ( .A1(a_27_), .A2(n12452), .ZN(n12172) );
  NAND2_X1 U12334 ( .A1(n12457), .A2(n12458), .ZN(n12452) );
  NAND2_X1 U12335 ( .A1(n12459), .A2(b_18_), .ZN(n12458) );
  NOR2_X1 U12336 ( .A1(n12460), .A2(n8055), .ZN(n12459) );
  NOR2_X1 U12337 ( .A1(n12179), .A2(n12181), .ZN(n12460) );
  NAND2_X1 U12338 ( .A1(n12179), .A2(n12181), .ZN(n12457) );
  NAND2_X1 U12339 ( .A1(n12461), .A2(n12462), .ZN(n12181) );
  NAND2_X1 U12340 ( .A1(n12197), .A2(n12463), .ZN(n12462) );
  OR2_X1 U12341 ( .A1(n12198), .A2(n12199), .ZN(n12463) );
  NOR2_X1 U12342 ( .A1(n8946), .A2(n8041), .ZN(n12197) );
  NAND2_X1 U12343 ( .A1(n12199), .A2(n12198), .ZN(n12461) );
  NAND2_X1 U12344 ( .A1(n12464), .A2(n12465), .ZN(n12198) );
  NAND2_X1 U12345 ( .A1(b_16_), .A2(n12466), .ZN(n12465) );
  NAND2_X1 U12346 ( .A1(n8003), .A2(n12467), .ZN(n12466) );
  NAND2_X1 U12347 ( .A1(a_31_), .A2(n8948), .ZN(n12467) );
  NAND2_X1 U12348 ( .A1(b_17_), .A2(n12468), .ZN(n12464) );
  NAND2_X1 U12349 ( .A1(n9341), .A2(n12469), .ZN(n12468) );
  NAND2_X1 U12350 ( .A1(a_30_), .A2(n8949), .ZN(n12469) );
  AND2_X1 U12351 ( .A1(n12470), .A2(n7953), .ZN(n12199) );
  NOR2_X1 U12352 ( .A1(n8946), .A2(n8948), .ZN(n12470) );
  XOR2_X1 U12353 ( .A(n12471), .B(n12472), .Z(n12179) );
  XOR2_X1 U12354 ( .A(n12473), .B(n12474), .Z(n12471) );
  XNOR2_X1 U12355 ( .A(n12475), .B(n12476), .ZN(n12204) );
  NAND2_X1 U12356 ( .A1(n12477), .A2(n12478), .ZN(n12475) );
  XNOR2_X1 U12357 ( .A(n12479), .B(n12480), .ZN(n12209) );
  XNOR2_X1 U12358 ( .A(n12481), .B(n12482), .ZN(n12480) );
  XOR2_X1 U12359 ( .A(n12483), .B(n12484), .Z(n12212) );
  XOR2_X1 U12360 ( .A(n12485), .B(n12486), .Z(n12483) );
  NOR2_X1 U12361 ( .A1(n8939), .A2(n8948), .ZN(n12486) );
  XOR2_X1 U12362 ( .A(n12487), .B(n12488), .Z(n12221) );
  XOR2_X1 U12363 ( .A(n12489), .B(n12490), .Z(n12487) );
  NOR2_X1 U12364 ( .A1(n8941), .A2(n8948), .ZN(n12490) );
  XNOR2_X1 U12365 ( .A(n12491), .B(n12492), .ZN(n12225) );
  XNOR2_X1 U12366 ( .A(n12493), .B(n12494), .ZN(n12492) );
  XOR2_X1 U12367 ( .A(n12495), .B(n12496), .Z(n12228) );
  XOR2_X1 U12368 ( .A(n12497), .B(n12498), .Z(n12495) );
  NOR2_X1 U12369 ( .A1(n8944), .A2(n8948), .ZN(n12498) );
  INV_X1 U12370 ( .A(n8357), .ZN(n12235) );
  NAND2_X1 U12371 ( .A1(b_18_), .A2(a_18_), .ZN(n8357) );
  XOR2_X1 U12372 ( .A(n12499), .B(n12500), .Z(n12236) );
  XOR2_X1 U12373 ( .A(n12501), .B(n12502), .Z(n12499) );
  NOR2_X1 U12374 ( .A1(n8947), .A2(n8948), .ZN(n12502) );
  XOR2_X1 U12375 ( .A(n12503), .B(n12504), .Z(n12240) );
  XOR2_X1 U12376 ( .A(n12505), .B(n12506), .Z(n12503) );
  XOR2_X1 U12377 ( .A(n12507), .B(n12508), .Z(n12245) );
  XOR2_X1 U12378 ( .A(n12509), .B(n12510), .Z(n12507) );
  NOR2_X1 U12379 ( .A1(n8950), .A2(n8948), .ZN(n12510) );
  XOR2_X1 U12380 ( .A(n12511), .B(n12512), .Z(n12249) );
  XOR2_X1 U12381 ( .A(n12513), .B(n12514), .Z(n12511) );
  XOR2_X1 U12382 ( .A(n12515), .B(n12516), .Z(n12253) );
  XOR2_X1 U12383 ( .A(n12517), .B(n12518), .Z(n12515) );
  XNOR2_X1 U12384 ( .A(n12519), .B(n12520), .ZN(n12257) );
  XOR2_X1 U12385 ( .A(n12521), .B(n12522), .Z(n12519) );
  NOR2_X1 U12386 ( .A1(n8495), .A2(n8948), .ZN(n12522) );
  XNOR2_X1 U12387 ( .A(n12523), .B(n12524), .ZN(n12261) );
  XOR2_X1 U12388 ( .A(n12525), .B(n12526), .Z(n12524) );
  NAND2_X1 U12389 ( .A1(b_17_), .A2(a_12_), .ZN(n12526) );
  XOR2_X1 U12390 ( .A(n12527), .B(n12528), .Z(n12264) );
  XOR2_X1 U12391 ( .A(n12529), .B(n12530), .Z(n12527) );
  NOR2_X1 U12392 ( .A1(n8550), .A2(n8948), .ZN(n12530) );
  XOR2_X1 U12393 ( .A(n12531), .B(n12532), .Z(n12268) );
  XOR2_X1 U12394 ( .A(n12533), .B(n12534), .Z(n12531) );
  NOR2_X1 U12395 ( .A1(n8959), .A2(n8948), .ZN(n12534) );
  XOR2_X1 U12396 ( .A(n12535), .B(n12536), .Z(n12281) );
  XOR2_X1 U12397 ( .A(n12537), .B(n12538), .Z(n12536) );
  NAND2_X1 U12398 ( .A1(b_17_), .A2(a_7_), .ZN(n12538) );
  XNOR2_X1 U12399 ( .A(n12539), .B(n12540), .ZN(n12285) );
  XOR2_X1 U12400 ( .A(n12541), .B(n12542), .Z(n12540) );
  NAND2_X1 U12401 ( .A1(b_17_), .A2(a_6_), .ZN(n12542) );
  NAND2_X1 U12402 ( .A1(n12543), .A2(n12544), .ZN(n9080) );
  XOR2_X1 U12403 ( .A(n12545), .B(n9154), .Z(n12544) );
  AND2_X1 U12404 ( .A1(n9153), .A2(n9152), .ZN(n12543) );
  INV_X1 U12405 ( .A(n12305), .ZN(n9152) );
  XOR2_X1 U12406 ( .A(n12546), .B(n12547), .Z(n12305) );
  NAND2_X1 U12407 ( .A1(n12548), .A2(n12549), .ZN(n12546) );
  NAND2_X1 U12408 ( .A1(n12550), .A2(n12551), .ZN(n9153) );
  NAND2_X1 U12409 ( .A1(n12552), .A2(b_17_), .ZN(n12551) );
  NOR2_X1 U12410 ( .A1(n12553), .A2(n8974), .ZN(n12552) );
  NOR2_X1 U12411 ( .A1(n12309), .A2(n12310), .ZN(n12553) );
  NAND2_X1 U12412 ( .A1(n12309), .A2(n12310), .ZN(n12550) );
  NAND2_X1 U12413 ( .A1(n12554), .A2(n12555), .ZN(n12310) );
  NAND2_X1 U12414 ( .A1(n12556), .A2(b_17_), .ZN(n12555) );
  NOR2_X1 U12415 ( .A1(n12557), .A2(n8969), .ZN(n12556) );
  NOR2_X1 U12416 ( .A1(n12316), .A2(n12317), .ZN(n12557) );
  NAND2_X1 U12417 ( .A1(n12316), .A2(n12317), .ZN(n12554) );
  NAND2_X1 U12418 ( .A1(n12558), .A2(n12559), .ZN(n12317) );
  NAND2_X1 U12419 ( .A1(n12560), .A2(b_17_), .ZN(n12559) );
  NOR2_X1 U12420 ( .A1(n12561), .A2(n8792), .ZN(n12560) );
  NOR2_X1 U12421 ( .A1(n12324), .A2(n12325), .ZN(n12561) );
  NAND2_X1 U12422 ( .A1(n12324), .A2(n12325), .ZN(n12558) );
  NAND2_X1 U12423 ( .A1(n12562), .A2(n12563), .ZN(n12325) );
  NAND2_X1 U12424 ( .A1(n12564), .A2(b_17_), .ZN(n12563) );
  NOR2_X1 U12425 ( .A1(n12565), .A2(n8778), .ZN(n12564) );
  NOR2_X1 U12426 ( .A1(n12332), .A2(n12333), .ZN(n12565) );
  NAND2_X1 U12427 ( .A1(n12332), .A2(n12333), .ZN(n12562) );
  NAND2_X1 U12428 ( .A1(n12566), .A2(n12567), .ZN(n12333) );
  NAND2_X1 U12429 ( .A1(n12568), .A2(b_17_), .ZN(n12567) );
  NOR2_X1 U12430 ( .A1(n12569), .A2(n8966), .ZN(n12568) );
  NOR2_X1 U12431 ( .A1(n12340), .A2(n12341), .ZN(n12569) );
  NAND2_X1 U12432 ( .A1(n12340), .A2(n12341), .ZN(n12566) );
  NAND2_X1 U12433 ( .A1(n12570), .A2(n12571), .ZN(n12341) );
  NAND2_X1 U12434 ( .A1(n12572), .A2(b_17_), .ZN(n12571) );
  NOR2_X1 U12435 ( .A1(n12573), .A2(n8723), .ZN(n12572) );
  NOR2_X1 U12436 ( .A1(n12348), .A2(n12349), .ZN(n12573) );
  NAND2_X1 U12437 ( .A1(n12348), .A2(n12349), .ZN(n12570) );
  NAND2_X1 U12438 ( .A1(n12574), .A2(n12575), .ZN(n12349) );
  NAND2_X1 U12439 ( .A1(n12576), .A2(b_17_), .ZN(n12575) );
  NOR2_X1 U12440 ( .A1(n12577), .A2(n8681), .ZN(n12576) );
  NOR2_X1 U12441 ( .A1(n12539), .A2(n12541), .ZN(n12577) );
  NAND2_X1 U12442 ( .A1(n12539), .A2(n12541), .ZN(n12574) );
  NAND2_X1 U12443 ( .A1(n12578), .A2(n12579), .ZN(n12541) );
  NAND2_X1 U12444 ( .A1(n12580), .A2(b_17_), .ZN(n12579) );
  NOR2_X1 U12445 ( .A1(n12581), .A2(n8962), .ZN(n12580) );
  NOR2_X1 U12446 ( .A1(n12535), .A2(n12537), .ZN(n12581) );
  NAND2_X1 U12447 ( .A1(n12535), .A2(n12537), .ZN(n12578) );
  NAND2_X1 U12448 ( .A1(n12582), .A2(n12583), .ZN(n12537) );
  NAND2_X1 U12449 ( .A1(n12584), .A2(b_17_), .ZN(n12583) );
  NOR2_X1 U12450 ( .A1(n12585), .A2(n8619), .ZN(n12584) );
  NOR2_X1 U12451 ( .A1(n12363), .A2(n12364), .ZN(n12585) );
  NAND2_X1 U12452 ( .A1(n12363), .A2(n12364), .ZN(n12582) );
  NAND2_X1 U12453 ( .A1(n12586), .A2(n12587), .ZN(n12364) );
  NAND2_X1 U12454 ( .A1(n12588), .A2(b_17_), .ZN(n12587) );
  NOR2_X1 U12455 ( .A1(n12589), .A2(n8605), .ZN(n12588) );
  NOR2_X1 U12456 ( .A1(n12370), .A2(n12372), .ZN(n12589) );
  NAND2_X1 U12457 ( .A1(n12370), .A2(n12372), .ZN(n12586) );
  NAND2_X1 U12458 ( .A1(n12590), .A2(n12591), .ZN(n12372) );
  NAND2_X1 U12459 ( .A1(n12592), .A2(b_17_), .ZN(n12591) );
  NOR2_X1 U12460 ( .A1(n12593), .A2(n8959), .ZN(n12592) );
  NOR2_X1 U12461 ( .A1(n12532), .A2(n12533), .ZN(n12593) );
  NAND2_X1 U12462 ( .A1(n12532), .A2(n12533), .ZN(n12590) );
  NAND2_X1 U12463 ( .A1(n12594), .A2(n12595), .ZN(n12533) );
  NAND2_X1 U12464 ( .A1(n12596), .A2(b_17_), .ZN(n12595) );
  NOR2_X1 U12465 ( .A1(n12597), .A2(n8550), .ZN(n12596) );
  NOR2_X1 U12466 ( .A1(n12528), .A2(n12529), .ZN(n12597) );
  NAND2_X1 U12467 ( .A1(n12528), .A2(n12529), .ZN(n12594) );
  NAND2_X1 U12468 ( .A1(n12598), .A2(n12599), .ZN(n12529) );
  NAND2_X1 U12469 ( .A1(n12600), .A2(b_17_), .ZN(n12599) );
  NOR2_X1 U12470 ( .A1(n12601), .A2(n8956), .ZN(n12600) );
  NOR2_X1 U12471 ( .A1(n12523), .A2(n12525), .ZN(n12601) );
  NAND2_X1 U12472 ( .A1(n12523), .A2(n12525), .ZN(n12598) );
  NAND2_X1 U12473 ( .A1(n12602), .A2(n12603), .ZN(n12525) );
  NAND2_X1 U12474 ( .A1(n12604), .A2(b_17_), .ZN(n12603) );
  NOR2_X1 U12475 ( .A1(n12605), .A2(n8495), .ZN(n12604) );
  NOR2_X1 U12476 ( .A1(n12520), .A2(n12521), .ZN(n12605) );
  NAND2_X1 U12477 ( .A1(n12520), .A2(n12521), .ZN(n12602) );
  NAND2_X1 U12478 ( .A1(n12606), .A2(n12607), .ZN(n12521) );
  NAND2_X1 U12479 ( .A1(n12518), .A2(n12608), .ZN(n12607) );
  OR2_X1 U12480 ( .A1(n12517), .A2(n12516), .ZN(n12608) );
  NOR2_X1 U12481 ( .A1(n8948), .A2(n8953), .ZN(n12518) );
  NAND2_X1 U12482 ( .A1(n12516), .A2(n12517), .ZN(n12606) );
  NAND2_X1 U12483 ( .A1(n12609), .A2(n12610), .ZN(n12517) );
  NAND2_X1 U12484 ( .A1(n12514), .A2(n12611), .ZN(n12610) );
  OR2_X1 U12485 ( .A1(n12513), .A2(n12512), .ZN(n12611) );
  NOR2_X1 U12486 ( .A1(n8948), .A2(n8440), .ZN(n12514) );
  NAND2_X1 U12487 ( .A1(n12512), .A2(n12513), .ZN(n12609) );
  NAND2_X1 U12488 ( .A1(n12612), .A2(n12613), .ZN(n12513) );
  NAND2_X1 U12489 ( .A1(n12614), .A2(b_17_), .ZN(n12613) );
  NOR2_X1 U12490 ( .A1(n12615), .A2(n8950), .ZN(n12614) );
  NOR2_X1 U12491 ( .A1(n12508), .A2(n12509), .ZN(n12615) );
  NAND2_X1 U12492 ( .A1(n12508), .A2(n12509), .ZN(n12612) );
  NAND2_X1 U12493 ( .A1(n12616), .A2(n12617), .ZN(n12509) );
  NAND2_X1 U12494 ( .A1(n12506), .A2(n12618), .ZN(n12617) );
  OR2_X1 U12495 ( .A1(n12505), .A2(n12504), .ZN(n12618) );
  INV_X1 U12496 ( .A(n8897), .ZN(n12506) );
  NAND2_X1 U12497 ( .A1(b_17_), .A2(a_17_), .ZN(n8897) );
  NAND2_X1 U12498 ( .A1(n12504), .A2(n12505), .ZN(n12616) );
  NAND2_X1 U12499 ( .A1(n12619), .A2(n12620), .ZN(n12505) );
  NAND2_X1 U12500 ( .A1(n12621), .A2(b_17_), .ZN(n12620) );
  NOR2_X1 U12501 ( .A1(n12622), .A2(n8947), .ZN(n12621) );
  NOR2_X1 U12502 ( .A1(n12500), .A2(n12501), .ZN(n12622) );
  NAND2_X1 U12503 ( .A1(n12500), .A2(n12501), .ZN(n12619) );
  NAND2_X1 U12504 ( .A1(n12623), .A2(n12624), .ZN(n12501) );
  NAND2_X1 U12505 ( .A1(n12411), .A2(n12625), .ZN(n12624) );
  OR2_X1 U12506 ( .A1(n12410), .A2(n12408), .ZN(n12625) );
  NOR2_X1 U12507 ( .A1(n8948), .A2(n8324), .ZN(n12411) );
  NAND2_X1 U12508 ( .A1(n12408), .A2(n12410), .ZN(n12623) );
  NAND2_X1 U12509 ( .A1(n12626), .A2(n12627), .ZN(n12410) );
  NAND2_X1 U12510 ( .A1(n12628), .A2(b_17_), .ZN(n12627) );
  NOR2_X1 U12511 ( .A1(n12629), .A2(n8944), .ZN(n12628) );
  NOR2_X1 U12512 ( .A1(n12496), .A2(n12497), .ZN(n12629) );
  NAND2_X1 U12513 ( .A1(n12496), .A2(n12497), .ZN(n12626) );
  NAND2_X1 U12514 ( .A1(n12630), .A2(n12631), .ZN(n12497) );
  NAND2_X1 U12515 ( .A1(n12494), .A2(n12632), .ZN(n12631) );
  OR2_X1 U12516 ( .A1(n12493), .A2(n12491), .ZN(n12632) );
  NOR2_X1 U12517 ( .A1(n8948), .A2(n8268), .ZN(n12494) );
  NAND2_X1 U12518 ( .A1(n12491), .A2(n12493), .ZN(n12630) );
  NAND2_X1 U12519 ( .A1(n12633), .A2(n12634), .ZN(n12493) );
  NAND2_X1 U12520 ( .A1(n12635), .A2(b_17_), .ZN(n12634) );
  NOR2_X1 U12521 ( .A1(n12636), .A2(n8941), .ZN(n12635) );
  NOR2_X1 U12522 ( .A1(n12488), .A2(n12489), .ZN(n12636) );
  NAND2_X1 U12523 ( .A1(n12488), .A2(n12489), .ZN(n12633) );
  NAND2_X1 U12524 ( .A1(n12637), .A2(n12638), .ZN(n12489) );
  NAND2_X1 U12525 ( .A1(n12429), .A2(n12639), .ZN(n12638) );
  OR2_X1 U12526 ( .A1(n12428), .A2(n12426), .ZN(n12639) );
  NOR2_X1 U12527 ( .A1(n8948), .A2(n8213), .ZN(n12429) );
  NAND2_X1 U12528 ( .A1(n12426), .A2(n12428), .ZN(n12637) );
  NAND2_X1 U12529 ( .A1(n12640), .A2(n12641), .ZN(n12428) );
  NAND2_X1 U12530 ( .A1(n12642), .A2(b_17_), .ZN(n12641) );
  NOR2_X1 U12531 ( .A1(n12643), .A2(n8939), .ZN(n12642) );
  NOR2_X1 U12532 ( .A1(n12484), .A2(n12485), .ZN(n12643) );
  NAND2_X1 U12533 ( .A1(n12484), .A2(n12485), .ZN(n12640) );
  NAND2_X1 U12534 ( .A1(n12644), .A2(n12645), .ZN(n12485) );
  NAND2_X1 U12535 ( .A1(n12482), .A2(n12646), .ZN(n12645) );
  OR2_X1 U12536 ( .A1(n12481), .A2(n12479), .ZN(n12646) );
  NOR2_X1 U12537 ( .A1(n8948), .A2(n8158), .ZN(n12482) );
  NAND2_X1 U12538 ( .A1(n12479), .A2(n12481), .ZN(n12644) );
  NAND2_X1 U12539 ( .A1(n12477), .A2(n12647), .ZN(n12481) );
  NAND2_X1 U12540 ( .A1(n12476), .A2(n12478), .ZN(n12647) );
  NAND2_X1 U12541 ( .A1(n12648), .A2(n12649), .ZN(n12478) );
  NAND2_X1 U12542 ( .A1(b_17_), .A2(a_26_), .ZN(n12649) );
  INV_X1 U12543 ( .A(n12650), .ZN(n12648) );
  XNOR2_X1 U12544 ( .A(n12651), .B(n12652), .ZN(n12476) );
  NAND2_X1 U12545 ( .A1(n12653), .A2(n12654), .ZN(n12651) );
  NAND2_X1 U12546 ( .A1(a_26_), .A2(n12650), .ZN(n12477) );
  NAND2_X1 U12547 ( .A1(n12447), .A2(n12655), .ZN(n12650) );
  NAND2_X1 U12548 ( .A1(n12446), .A2(n12448), .ZN(n12655) );
  NAND2_X1 U12549 ( .A1(n12656), .A2(n12657), .ZN(n12448) );
  NAND2_X1 U12550 ( .A1(b_17_), .A2(a_27_), .ZN(n12657) );
  INV_X1 U12551 ( .A(n12658), .ZN(n12656) );
  XOR2_X1 U12552 ( .A(n12659), .B(n12660), .Z(n12446) );
  XNOR2_X1 U12553 ( .A(n12661), .B(n12662), .ZN(n12659) );
  NAND2_X1 U12554 ( .A1(b_16_), .A2(a_28_), .ZN(n12661) );
  NAND2_X1 U12555 ( .A1(a_27_), .A2(n12658), .ZN(n12447) );
  NAND2_X1 U12556 ( .A1(n12663), .A2(n12664), .ZN(n12658) );
  NAND2_X1 U12557 ( .A1(n12665), .A2(b_17_), .ZN(n12664) );
  NOR2_X1 U12558 ( .A1(n12666), .A2(n8055), .ZN(n12665) );
  NOR2_X1 U12559 ( .A1(n12454), .A2(n12456), .ZN(n12666) );
  NAND2_X1 U12560 ( .A1(n12454), .A2(n12456), .ZN(n12663) );
  NAND2_X1 U12561 ( .A1(n12667), .A2(n12668), .ZN(n12456) );
  NAND2_X1 U12562 ( .A1(n12472), .A2(n12669), .ZN(n12668) );
  OR2_X1 U12563 ( .A1(n12473), .A2(n12474), .ZN(n12669) );
  NOR2_X1 U12564 ( .A1(n8948), .A2(n8041), .ZN(n12472) );
  NAND2_X1 U12565 ( .A1(n12474), .A2(n12473), .ZN(n12667) );
  NAND2_X1 U12566 ( .A1(n12670), .A2(n12671), .ZN(n12473) );
  NAND2_X1 U12567 ( .A1(b_15_), .A2(n12672), .ZN(n12671) );
  NAND2_X1 U12568 ( .A1(n8003), .A2(n12673), .ZN(n12672) );
  NAND2_X1 U12569 ( .A1(a_31_), .A2(n8949), .ZN(n12673) );
  NAND2_X1 U12570 ( .A1(b_16_), .A2(n12674), .ZN(n12670) );
  NAND2_X1 U12571 ( .A1(n9341), .A2(n12675), .ZN(n12674) );
  NAND2_X1 U12572 ( .A1(a_30_), .A2(n8951), .ZN(n12675) );
  AND2_X1 U12573 ( .A1(n12676), .A2(n7953), .ZN(n12474) );
  NOR2_X1 U12574 ( .A1(n8948), .A2(n8949), .ZN(n12676) );
  XOR2_X1 U12575 ( .A(n12677), .B(n12678), .Z(n12454) );
  XOR2_X1 U12576 ( .A(n12679), .B(n12680), .Z(n12677) );
  XNOR2_X1 U12577 ( .A(n12681), .B(n12682), .ZN(n12479) );
  NAND2_X1 U12578 ( .A1(n12683), .A2(n12684), .ZN(n12681) );
  XNOR2_X1 U12579 ( .A(n12685), .B(n12686), .ZN(n12484) );
  XNOR2_X1 U12580 ( .A(n12687), .B(n12688), .ZN(n12686) );
  XOR2_X1 U12581 ( .A(n12689), .B(n12690), .Z(n12426) );
  XOR2_X1 U12582 ( .A(n12691), .B(n12692), .Z(n12689) );
  NOR2_X1 U12583 ( .A1(n8939), .A2(n8949), .ZN(n12692) );
  XNOR2_X1 U12584 ( .A(n12693), .B(n12694), .ZN(n12488) );
  XNOR2_X1 U12585 ( .A(n12695), .B(n12696), .ZN(n12694) );
  XOR2_X1 U12586 ( .A(n12697), .B(n12698), .Z(n12491) );
  XOR2_X1 U12587 ( .A(n12699), .B(n12700), .Z(n12697) );
  NOR2_X1 U12588 ( .A1(n8941), .A2(n8949), .ZN(n12700) );
  XNOR2_X1 U12589 ( .A(n12701), .B(n12702), .ZN(n12496) );
  XNOR2_X1 U12590 ( .A(n12703), .B(n12704), .ZN(n12702) );
  XOR2_X1 U12591 ( .A(n12705), .B(n12706), .Z(n12408) );
  XOR2_X1 U12592 ( .A(n12707), .B(n12708), .Z(n12705) );
  NOR2_X1 U12593 ( .A1(n8944), .A2(n8949), .ZN(n12708) );
  XOR2_X1 U12594 ( .A(n12709), .B(n12710), .Z(n12500) );
  XOR2_X1 U12595 ( .A(n12711), .B(n12712), .Z(n12709) );
  XOR2_X1 U12596 ( .A(n12713), .B(n12714), .Z(n12504) );
  XOR2_X1 U12597 ( .A(n12715), .B(n12716), .Z(n12713) );
  NOR2_X1 U12598 ( .A1(n8947), .A2(n8949), .ZN(n12716) );
  XOR2_X1 U12599 ( .A(n12717), .B(n12718), .Z(n12508) );
  XOR2_X1 U12600 ( .A(n12719), .B(n12720), .Z(n12717) );
  XOR2_X1 U12601 ( .A(n12721), .B(n12722), .Z(n12512) );
  XOR2_X1 U12602 ( .A(n12723), .B(n12724), .Z(n12721) );
  XNOR2_X1 U12603 ( .A(n12725), .B(n12726), .ZN(n12516) );
  XOR2_X1 U12604 ( .A(n12727), .B(n12728), .Z(n12726) );
  NAND2_X1 U12605 ( .A1(b_16_), .A2(a_15_), .ZN(n12728) );
  XNOR2_X1 U12606 ( .A(n12729), .B(n12730), .ZN(n12520) );
  XNOR2_X1 U12607 ( .A(n12731), .B(n12732), .ZN(n12729) );
  XNOR2_X1 U12608 ( .A(n12733), .B(n12734), .ZN(n12523) );
  XNOR2_X1 U12609 ( .A(n12735), .B(n12736), .ZN(n12734) );
  XNOR2_X1 U12610 ( .A(n12737), .B(n12738), .ZN(n12528) );
  XNOR2_X1 U12611 ( .A(n12739), .B(n12740), .ZN(n12737) );
  XNOR2_X1 U12612 ( .A(n12741), .B(n12742), .ZN(n12532) );
  XNOR2_X1 U12613 ( .A(n12743), .B(n12744), .ZN(n12742) );
  XNOR2_X1 U12614 ( .A(n12745), .B(n12746), .ZN(n12370) );
  XOR2_X1 U12615 ( .A(n12747), .B(n12748), .Z(n12746) );
  NAND2_X1 U12616 ( .A1(b_16_), .A2(a_10_), .ZN(n12748) );
  XNOR2_X1 U12617 ( .A(n12749), .B(n12750), .ZN(n12363) );
  NAND2_X1 U12618 ( .A1(n12751), .A2(n12752), .ZN(n12749) );
  XNOR2_X1 U12619 ( .A(n12753), .B(n12754), .ZN(n12535) );
  XNOR2_X1 U12620 ( .A(n12755), .B(n12756), .ZN(n12753) );
  XNOR2_X1 U12621 ( .A(n12757), .B(n12758), .ZN(n12539) );
  XNOR2_X1 U12622 ( .A(n12759), .B(n12760), .ZN(n12758) );
  XNOR2_X1 U12623 ( .A(n12761), .B(n12762), .ZN(n12348) );
  XNOR2_X1 U12624 ( .A(n12763), .B(n12764), .ZN(n12762) );
  XNOR2_X1 U12625 ( .A(n12765), .B(n12766), .ZN(n12340) );
  XOR2_X1 U12626 ( .A(n12767), .B(n12768), .Z(n12766) );
  NAND2_X1 U12627 ( .A1(b_16_), .A2(a_5_), .ZN(n12768) );
  XOR2_X1 U12628 ( .A(n12769), .B(n12770), .Z(n12332) );
  XOR2_X1 U12629 ( .A(n12771), .B(n12772), .Z(n12769) );
  XNOR2_X1 U12630 ( .A(n12773), .B(n12774), .ZN(n12324) );
  XNOR2_X1 U12631 ( .A(n12775), .B(n12776), .ZN(n12774) );
  XNOR2_X1 U12632 ( .A(n12777), .B(n12778), .ZN(n12316) );
  XOR2_X1 U12633 ( .A(n12779), .B(n12780), .Z(n12778) );
  NAND2_X1 U12634 ( .A1(b_16_), .A2(a_2_), .ZN(n12780) );
  XNOR2_X1 U12635 ( .A(n12781), .B(n12782), .ZN(n12309) );
  NAND2_X1 U12636 ( .A1(n12783), .A2(n12784), .ZN(n12781) );
  NAND2_X1 U12637 ( .A1(n12785), .A2(n12786), .ZN(n9085) );
  NAND2_X1 U12638 ( .A1(n9154), .A2(n12545), .ZN(n12786) );
  NAND2_X1 U12639 ( .A1(n12787), .A2(n9154), .ZN(n9086) );
  XOR2_X1 U12640 ( .A(n12788), .B(n12789), .Z(n9154) );
  XOR2_X1 U12641 ( .A(n12790), .B(n12791), .Z(n12788) );
  NOR2_X1 U12642 ( .A1(n8974), .A2(n8951), .ZN(n12791) );
  NOR2_X1 U12643 ( .A1(n9155), .A2(n12785), .ZN(n12787) );
  XOR2_X1 U12644 ( .A(n12792), .B(n12793), .Z(n12785) );
  INV_X1 U12645 ( .A(n12545), .ZN(n9155) );
  NAND2_X1 U12646 ( .A1(n12548), .A2(n12794), .ZN(n12545) );
  NAND2_X1 U12647 ( .A1(n12547), .A2(n12549), .ZN(n12794) );
  NAND2_X1 U12648 ( .A1(n12795), .A2(n12796), .ZN(n12549) );
  NAND2_X1 U12649 ( .A1(b_16_), .A2(a_0_), .ZN(n12796) );
  INV_X1 U12650 ( .A(n12797), .ZN(n12795) );
  XNOR2_X1 U12651 ( .A(n12798), .B(n12799), .ZN(n12547) );
  NAND2_X1 U12652 ( .A1(n12800), .A2(n12801), .ZN(n12798) );
  NAND2_X1 U12653 ( .A1(a_0_), .A2(n12797), .ZN(n12548) );
  NAND2_X1 U12654 ( .A1(n12783), .A2(n12802), .ZN(n12797) );
  NAND2_X1 U12655 ( .A1(n12782), .A2(n12784), .ZN(n12802) );
  NAND2_X1 U12656 ( .A1(n12803), .A2(n12804), .ZN(n12784) );
  NAND2_X1 U12657 ( .A1(b_16_), .A2(a_1_), .ZN(n12804) );
  INV_X1 U12658 ( .A(n12805), .ZN(n12803) );
  XOR2_X1 U12659 ( .A(n12806), .B(n12807), .Z(n12782) );
  XOR2_X1 U12660 ( .A(n12808), .B(n12809), .Z(n12806) );
  NOR2_X1 U12661 ( .A1(n8792), .A2(n8951), .ZN(n12809) );
  NAND2_X1 U12662 ( .A1(a_1_), .A2(n12805), .ZN(n12783) );
  NAND2_X1 U12663 ( .A1(n12810), .A2(n12811), .ZN(n12805) );
  NAND2_X1 U12664 ( .A1(n12812), .A2(b_16_), .ZN(n12811) );
  NOR2_X1 U12665 ( .A1(n12813), .A2(n8792), .ZN(n12812) );
  NOR2_X1 U12666 ( .A1(n12777), .A2(n12779), .ZN(n12813) );
  NAND2_X1 U12667 ( .A1(n12777), .A2(n12779), .ZN(n12810) );
  NAND2_X1 U12668 ( .A1(n12814), .A2(n12815), .ZN(n12779) );
  NAND2_X1 U12669 ( .A1(n12776), .A2(n12816), .ZN(n12815) );
  OR2_X1 U12670 ( .A1(n12775), .A2(n12773), .ZN(n12816) );
  NOR2_X1 U12671 ( .A1(n8949), .A2(n8778), .ZN(n12776) );
  NAND2_X1 U12672 ( .A1(n12773), .A2(n12775), .ZN(n12814) );
  NAND2_X1 U12673 ( .A1(n12817), .A2(n12818), .ZN(n12775) );
  NAND2_X1 U12674 ( .A1(n12772), .A2(n12819), .ZN(n12818) );
  OR2_X1 U12675 ( .A1(n12770), .A2(n12771), .ZN(n12819) );
  NOR2_X1 U12676 ( .A1(n8949), .A2(n8966), .ZN(n12772) );
  NAND2_X1 U12677 ( .A1(n12770), .A2(n12771), .ZN(n12817) );
  NAND2_X1 U12678 ( .A1(n12820), .A2(n12821), .ZN(n12771) );
  NAND2_X1 U12679 ( .A1(n12822), .A2(b_16_), .ZN(n12821) );
  NOR2_X1 U12680 ( .A1(n12823), .A2(n8723), .ZN(n12822) );
  NOR2_X1 U12681 ( .A1(n12765), .A2(n12767), .ZN(n12823) );
  NAND2_X1 U12682 ( .A1(n12765), .A2(n12767), .ZN(n12820) );
  NAND2_X1 U12683 ( .A1(n12824), .A2(n12825), .ZN(n12767) );
  NAND2_X1 U12684 ( .A1(n12764), .A2(n12826), .ZN(n12825) );
  OR2_X1 U12685 ( .A1(n12763), .A2(n12761), .ZN(n12826) );
  NOR2_X1 U12686 ( .A1(n8949), .A2(n8681), .ZN(n12764) );
  NAND2_X1 U12687 ( .A1(n12761), .A2(n12763), .ZN(n12824) );
  NAND2_X1 U12688 ( .A1(n12827), .A2(n12828), .ZN(n12763) );
  NAND2_X1 U12689 ( .A1(n12760), .A2(n12829), .ZN(n12828) );
  OR2_X1 U12690 ( .A1(n12759), .A2(n12757), .ZN(n12829) );
  NOR2_X1 U12691 ( .A1(n8949), .A2(n8962), .ZN(n12760) );
  NAND2_X1 U12692 ( .A1(n12757), .A2(n12759), .ZN(n12827) );
  NAND2_X1 U12693 ( .A1(n12830), .A2(n12831), .ZN(n12759) );
  NAND2_X1 U12694 ( .A1(n12756), .A2(n12832), .ZN(n12831) );
  NAND2_X1 U12695 ( .A1(n12755), .A2(n12754), .ZN(n12832) );
  NOR2_X1 U12696 ( .A1(n8949), .A2(n8619), .ZN(n12756) );
  OR2_X1 U12697 ( .A1(n12754), .A2(n12755), .ZN(n12830) );
  AND2_X1 U12698 ( .A1(n12751), .A2(n12833), .ZN(n12755) );
  NAND2_X1 U12699 ( .A1(n12750), .A2(n12752), .ZN(n12833) );
  NAND2_X1 U12700 ( .A1(n12834), .A2(n12835), .ZN(n12752) );
  NAND2_X1 U12701 ( .A1(b_16_), .A2(a_9_), .ZN(n12835) );
  INV_X1 U12702 ( .A(n12836), .ZN(n12834) );
  XOR2_X1 U12703 ( .A(n12837), .B(n12838), .Z(n12750) );
  XOR2_X1 U12704 ( .A(n12839), .B(n12840), .Z(n12837) );
  NOR2_X1 U12705 ( .A1(n8959), .A2(n8951), .ZN(n12840) );
  NAND2_X1 U12706 ( .A1(a_9_), .A2(n12836), .ZN(n12751) );
  NAND2_X1 U12707 ( .A1(n12841), .A2(n12842), .ZN(n12836) );
  NAND2_X1 U12708 ( .A1(n12843), .A2(b_16_), .ZN(n12842) );
  NOR2_X1 U12709 ( .A1(n12844), .A2(n8959), .ZN(n12843) );
  NOR2_X1 U12710 ( .A1(n12745), .A2(n12747), .ZN(n12844) );
  NAND2_X1 U12711 ( .A1(n12745), .A2(n12747), .ZN(n12841) );
  NAND2_X1 U12712 ( .A1(n12845), .A2(n12846), .ZN(n12747) );
  NAND2_X1 U12713 ( .A1(n12744), .A2(n12847), .ZN(n12846) );
  OR2_X1 U12714 ( .A1(n12741), .A2(n12743), .ZN(n12847) );
  NOR2_X1 U12715 ( .A1(n8949), .A2(n8550), .ZN(n12744) );
  NAND2_X1 U12716 ( .A1(n12741), .A2(n12743), .ZN(n12845) );
  NAND2_X1 U12717 ( .A1(n12848), .A2(n12849), .ZN(n12743) );
  NAND2_X1 U12718 ( .A1(n12740), .A2(n12850), .ZN(n12849) );
  NAND2_X1 U12719 ( .A1(n12739), .A2(n12738), .ZN(n12850) );
  NOR2_X1 U12720 ( .A1(n8949), .A2(n8956), .ZN(n12740) );
  OR2_X1 U12721 ( .A1(n12738), .A2(n12739), .ZN(n12848) );
  AND2_X1 U12722 ( .A1(n12851), .A2(n12852), .ZN(n12739) );
  NAND2_X1 U12723 ( .A1(n12736), .A2(n12853), .ZN(n12852) );
  OR2_X1 U12724 ( .A1(n12733), .A2(n12735), .ZN(n12853) );
  NOR2_X1 U12725 ( .A1(n8949), .A2(n8495), .ZN(n12736) );
  NAND2_X1 U12726 ( .A1(n12733), .A2(n12735), .ZN(n12851) );
  NAND2_X1 U12727 ( .A1(n12854), .A2(n12855), .ZN(n12735) );
  NAND2_X1 U12728 ( .A1(n12732), .A2(n12856), .ZN(n12855) );
  NAND2_X1 U12729 ( .A1(n12731), .A2(n12730), .ZN(n12856) );
  NOR2_X1 U12730 ( .A1(n8949), .A2(n8953), .ZN(n12732) );
  OR2_X1 U12731 ( .A1(n12730), .A2(n12731), .ZN(n12854) );
  AND2_X1 U12732 ( .A1(n12857), .A2(n12858), .ZN(n12731) );
  NAND2_X1 U12733 ( .A1(n12859), .A2(b_16_), .ZN(n12858) );
  NOR2_X1 U12734 ( .A1(n12860), .A2(n8440), .ZN(n12859) );
  NOR2_X1 U12735 ( .A1(n12725), .A2(n12727), .ZN(n12860) );
  NAND2_X1 U12736 ( .A1(n12725), .A2(n12727), .ZN(n12857) );
  NAND2_X1 U12737 ( .A1(n12861), .A2(n12862), .ZN(n12727) );
  NAND2_X1 U12738 ( .A1(n12722), .A2(n12863), .ZN(n12862) );
  OR2_X1 U12739 ( .A1(n12723), .A2(n12724), .ZN(n12863) );
  XOR2_X1 U12740 ( .A(n12864), .B(n12865), .Z(n12722) );
  XOR2_X1 U12741 ( .A(n12866), .B(n12867), .Z(n12864) );
  NAND2_X1 U12742 ( .A1(n12724), .A2(n12723), .ZN(n12861) );
  NAND2_X1 U12743 ( .A1(n12868), .A2(n12869), .ZN(n12723) );
  NAND2_X1 U12744 ( .A1(n12720), .A2(n12870), .ZN(n12869) );
  OR2_X1 U12745 ( .A1(n12718), .A2(n12719), .ZN(n12870) );
  NOR2_X1 U12746 ( .A1(n8949), .A2(n8385), .ZN(n12720) );
  NAND2_X1 U12747 ( .A1(n12718), .A2(n12719), .ZN(n12868) );
  NAND2_X1 U12748 ( .A1(n12871), .A2(n12872), .ZN(n12719) );
  NAND2_X1 U12749 ( .A1(n12873), .A2(b_16_), .ZN(n12872) );
  NOR2_X1 U12750 ( .A1(n12874), .A2(n8947), .ZN(n12873) );
  NOR2_X1 U12751 ( .A1(n12714), .A2(n12715), .ZN(n12874) );
  NAND2_X1 U12752 ( .A1(n12714), .A2(n12715), .ZN(n12871) );
  NAND2_X1 U12753 ( .A1(n12875), .A2(n12876), .ZN(n12715) );
  NAND2_X1 U12754 ( .A1(n12712), .A2(n12877), .ZN(n12876) );
  OR2_X1 U12755 ( .A1(n12710), .A2(n12711), .ZN(n12877) );
  NOR2_X1 U12756 ( .A1(n8949), .A2(n8324), .ZN(n12712) );
  NAND2_X1 U12757 ( .A1(n12710), .A2(n12711), .ZN(n12875) );
  NAND2_X1 U12758 ( .A1(n12878), .A2(n12879), .ZN(n12711) );
  NAND2_X1 U12759 ( .A1(n12880), .A2(b_16_), .ZN(n12879) );
  NOR2_X1 U12760 ( .A1(n12881), .A2(n8944), .ZN(n12880) );
  NOR2_X1 U12761 ( .A1(n12706), .A2(n12707), .ZN(n12881) );
  NAND2_X1 U12762 ( .A1(n12706), .A2(n12707), .ZN(n12878) );
  NAND2_X1 U12763 ( .A1(n12882), .A2(n12883), .ZN(n12707) );
  NAND2_X1 U12764 ( .A1(n12704), .A2(n12884), .ZN(n12883) );
  OR2_X1 U12765 ( .A1(n12701), .A2(n12703), .ZN(n12884) );
  NOR2_X1 U12766 ( .A1(n8949), .A2(n8268), .ZN(n12704) );
  NAND2_X1 U12767 ( .A1(n12701), .A2(n12703), .ZN(n12882) );
  NAND2_X1 U12768 ( .A1(n12885), .A2(n12886), .ZN(n12703) );
  NAND2_X1 U12769 ( .A1(n12887), .A2(b_16_), .ZN(n12886) );
  NOR2_X1 U12770 ( .A1(n12888), .A2(n8941), .ZN(n12887) );
  NOR2_X1 U12771 ( .A1(n12698), .A2(n12699), .ZN(n12888) );
  NAND2_X1 U12772 ( .A1(n12698), .A2(n12699), .ZN(n12885) );
  NAND2_X1 U12773 ( .A1(n12889), .A2(n12890), .ZN(n12699) );
  NAND2_X1 U12774 ( .A1(n12696), .A2(n12891), .ZN(n12890) );
  OR2_X1 U12775 ( .A1(n12693), .A2(n12695), .ZN(n12891) );
  NOR2_X1 U12776 ( .A1(n8949), .A2(n8213), .ZN(n12696) );
  NAND2_X1 U12777 ( .A1(n12693), .A2(n12695), .ZN(n12889) );
  NAND2_X1 U12778 ( .A1(n12892), .A2(n12893), .ZN(n12695) );
  NAND2_X1 U12779 ( .A1(n12894), .A2(b_16_), .ZN(n12893) );
  NOR2_X1 U12780 ( .A1(n12895), .A2(n8939), .ZN(n12894) );
  NOR2_X1 U12781 ( .A1(n12690), .A2(n12691), .ZN(n12895) );
  NAND2_X1 U12782 ( .A1(n12690), .A2(n12691), .ZN(n12892) );
  NAND2_X1 U12783 ( .A1(n12896), .A2(n12897), .ZN(n12691) );
  NAND2_X1 U12784 ( .A1(n12688), .A2(n12898), .ZN(n12897) );
  OR2_X1 U12785 ( .A1(n12685), .A2(n12687), .ZN(n12898) );
  NOR2_X1 U12786 ( .A1(n8949), .A2(n8158), .ZN(n12688) );
  NAND2_X1 U12787 ( .A1(n12685), .A2(n12687), .ZN(n12896) );
  NAND2_X1 U12788 ( .A1(n12683), .A2(n12899), .ZN(n12687) );
  NAND2_X1 U12789 ( .A1(n12682), .A2(n12684), .ZN(n12899) );
  NAND2_X1 U12790 ( .A1(n12900), .A2(n12901), .ZN(n12684) );
  NAND2_X1 U12791 ( .A1(b_16_), .A2(a_26_), .ZN(n12901) );
  INV_X1 U12792 ( .A(n12902), .ZN(n12900) );
  XNOR2_X1 U12793 ( .A(n12903), .B(n12904), .ZN(n12682) );
  NAND2_X1 U12794 ( .A1(n12905), .A2(n12906), .ZN(n12903) );
  NAND2_X1 U12795 ( .A1(a_26_), .A2(n12902), .ZN(n12683) );
  NAND2_X1 U12796 ( .A1(n12653), .A2(n12907), .ZN(n12902) );
  NAND2_X1 U12797 ( .A1(n12652), .A2(n12654), .ZN(n12907) );
  NAND2_X1 U12798 ( .A1(n12908), .A2(n12909), .ZN(n12654) );
  NAND2_X1 U12799 ( .A1(b_16_), .A2(a_27_), .ZN(n12909) );
  INV_X1 U12800 ( .A(n12910), .ZN(n12908) );
  XOR2_X1 U12801 ( .A(n12911), .B(n12912), .Z(n12652) );
  XNOR2_X1 U12802 ( .A(n12913), .B(n12914), .ZN(n12911) );
  NAND2_X1 U12803 ( .A1(b_15_), .A2(a_28_), .ZN(n12913) );
  NAND2_X1 U12804 ( .A1(a_27_), .A2(n12910), .ZN(n12653) );
  NAND2_X1 U12805 ( .A1(n12915), .A2(n12916), .ZN(n12910) );
  NAND2_X1 U12806 ( .A1(n12917), .A2(b_16_), .ZN(n12916) );
  NOR2_X1 U12807 ( .A1(n12918), .A2(n8055), .ZN(n12917) );
  NOR2_X1 U12808 ( .A1(n12660), .A2(n12662), .ZN(n12918) );
  NAND2_X1 U12809 ( .A1(n12660), .A2(n12662), .ZN(n12915) );
  NAND2_X1 U12810 ( .A1(n12919), .A2(n12920), .ZN(n12662) );
  NAND2_X1 U12811 ( .A1(n12678), .A2(n12921), .ZN(n12920) );
  OR2_X1 U12812 ( .A1(n12679), .A2(n12680), .ZN(n12921) );
  NOR2_X1 U12813 ( .A1(n8949), .A2(n8041), .ZN(n12678) );
  NAND2_X1 U12814 ( .A1(n12680), .A2(n12679), .ZN(n12919) );
  NAND2_X1 U12815 ( .A1(n12922), .A2(n12923), .ZN(n12679) );
  NAND2_X1 U12816 ( .A1(b_14_), .A2(n12924), .ZN(n12923) );
  NAND2_X1 U12817 ( .A1(n8003), .A2(n12925), .ZN(n12924) );
  NAND2_X1 U12818 ( .A1(a_31_), .A2(n8951), .ZN(n12925) );
  NAND2_X1 U12819 ( .A1(b_15_), .A2(n12926), .ZN(n12922) );
  NAND2_X1 U12820 ( .A1(n9341), .A2(n12927), .ZN(n12926) );
  NAND2_X1 U12821 ( .A1(a_30_), .A2(n8952), .ZN(n12927) );
  AND2_X1 U12822 ( .A1(n12928), .A2(n7953), .ZN(n12680) );
  NOR2_X1 U12823 ( .A1(n8949), .A2(n8951), .ZN(n12928) );
  XOR2_X1 U12824 ( .A(n12929), .B(n12930), .Z(n12660) );
  XOR2_X1 U12825 ( .A(n12931), .B(n12932), .Z(n12929) );
  XNOR2_X1 U12826 ( .A(n12933), .B(n12934), .ZN(n12685) );
  NAND2_X1 U12827 ( .A1(n12935), .A2(n12936), .ZN(n12933) );
  XNOR2_X1 U12828 ( .A(n12937), .B(n12938), .ZN(n12690) );
  XNOR2_X1 U12829 ( .A(n12939), .B(n12940), .ZN(n12938) );
  XOR2_X1 U12830 ( .A(n12941), .B(n12942), .Z(n12693) );
  XOR2_X1 U12831 ( .A(n12943), .B(n12944), .Z(n12941) );
  NOR2_X1 U12832 ( .A1(n8939), .A2(n8951), .ZN(n12944) );
  XNOR2_X1 U12833 ( .A(n12945), .B(n12946), .ZN(n12698) );
  XNOR2_X1 U12834 ( .A(n12947), .B(n12948), .ZN(n12946) );
  XOR2_X1 U12835 ( .A(n12949), .B(n12950), .Z(n12701) );
  XOR2_X1 U12836 ( .A(n12951), .B(n12952), .Z(n12949) );
  NOR2_X1 U12837 ( .A1(n8941), .A2(n8951), .ZN(n12952) );
  XNOR2_X1 U12838 ( .A(n12953), .B(n12954), .ZN(n12706) );
  XNOR2_X1 U12839 ( .A(n12955), .B(n12956), .ZN(n12954) );
  XOR2_X1 U12840 ( .A(n12957), .B(n12958), .Z(n12710) );
  XOR2_X1 U12841 ( .A(n12959), .B(n12960), .Z(n12957) );
  NOR2_X1 U12842 ( .A1(n8944), .A2(n8951), .ZN(n12960) );
  XNOR2_X1 U12843 ( .A(n12961), .B(n12962), .ZN(n12714) );
  XNOR2_X1 U12844 ( .A(n12963), .B(n12964), .ZN(n12962) );
  XOR2_X1 U12845 ( .A(n12965), .B(n12966), .Z(n12718) );
  XOR2_X1 U12846 ( .A(n12967), .B(n12968), .Z(n12965) );
  NOR2_X1 U12847 ( .A1(n8947), .A2(n8951), .ZN(n12968) );
  INV_X1 U12848 ( .A(n8418), .ZN(n12724) );
  NAND2_X1 U12849 ( .A1(b_16_), .A2(a_16_), .ZN(n8418) );
  XOR2_X1 U12850 ( .A(n12969), .B(n12970), .Z(n12725) );
  XOR2_X1 U12851 ( .A(n12971), .B(n12972), .Z(n12969) );
  XNOR2_X1 U12852 ( .A(n12973), .B(n12974), .ZN(n12730) );
  XOR2_X1 U12853 ( .A(n12975), .B(n12976), .Z(n12973) );
  XOR2_X1 U12854 ( .A(n12977), .B(n12978), .Z(n12733) );
  XNOR2_X1 U12855 ( .A(n12979), .B(n12980), .ZN(n12977) );
  NAND2_X1 U12856 ( .A1(b_15_), .A2(a_14_), .ZN(n12979) );
  XNOR2_X1 U12857 ( .A(n12981), .B(n12982), .ZN(n12738) );
  XOR2_X1 U12858 ( .A(n12983), .B(n12984), .Z(n12981) );
  NOR2_X1 U12859 ( .A1(n8495), .A2(n8951), .ZN(n12984) );
  XNOR2_X1 U12860 ( .A(n12985), .B(n12986), .ZN(n12741) );
  XOR2_X1 U12861 ( .A(n12987), .B(n12988), .Z(n12986) );
  NAND2_X1 U12862 ( .A1(b_15_), .A2(a_12_), .ZN(n12988) );
  XNOR2_X1 U12863 ( .A(n12989), .B(n12990), .ZN(n12745) );
  XOR2_X1 U12864 ( .A(n12991), .B(n12992), .Z(n12990) );
  NAND2_X1 U12865 ( .A1(b_15_), .A2(a_11_), .ZN(n12992) );
  XNOR2_X1 U12866 ( .A(n12993), .B(n12994), .ZN(n12754) );
  XOR2_X1 U12867 ( .A(n12995), .B(n12996), .Z(n12993) );
  NOR2_X1 U12868 ( .A1(n8605), .A2(n8951), .ZN(n12996) );
  XOR2_X1 U12869 ( .A(n12997), .B(n12998), .Z(n12757) );
  XOR2_X1 U12870 ( .A(n12999), .B(n13000), .Z(n12997) );
  NOR2_X1 U12871 ( .A1(n8619), .A2(n8951), .ZN(n13000) );
  XOR2_X1 U12872 ( .A(n13001), .B(n13002), .Z(n12761) );
  XOR2_X1 U12873 ( .A(n13003), .B(n13004), .Z(n13001) );
  NOR2_X1 U12874 ( .A1(n8962), .A2(n8951), .ZN(n13004) );
  XNOR2_X1 U12875 ( .A(n13005), .B(n13006), .ZN(n12765) );
  XOR2_X1 U12876 ( .A(n13007), .B(n13008), .Z(n13006) );
  NAND2_X1 U12877 ( .A1(b_15_), .A2(a_6_), .ZN(n13008) );
  XNOR2_X1 U12878 ( .A(n13009), .B(n13010), .ZN(n12770) );
  XOR2_X1 U12879 ( .A(n13011), .B(n13012), .Z(n13010) );
  NAND2_X1 U12880 ( .A1(b_15_), .A2(a_5_), .ZN(n13012) );
  XOR2_X1 U12881 ( .A(n13013), .B(n13014), .Z(n12773) );
  XOR2_X1 U12882 ( .A(n13015), .B(n13016), .Z(n13013) );
  NOR2_X1 U12883 ( .A1(n8966), .A2(n8951), .ZN(n13016) );
  XOR2_X1 U12884 ( .A(n13017), .B(n13018), .Z(n12777) );
  XOR2_X1 U12885 ( .A(n13019), .B(n13020), .Z(n13017) );
  NOR2_X1 U12886 ( .A1(n8778), .A2(n8951), .ZN(n13020) );
  NAND2_X1 U12887 ( .A1(n13021), .A2(n13022), .ZN(n9091) );
  NAND2_X1 U12888 ( .A1(n13023), .A2(n12792), .ZN(n13022) );
  XNOR2_X1 U12889 ( .A(n13024), .B(n13025), .ZN(n13021) );
  NAND2_X1 U12890 ( .A1(n13026), .A2(n13027), .ZN(n9092) );
  AND2_X1 U12891 ( .A1(n9146), .A2(n12792), .ZN(n13027) );
  NAND2_X1 U12892 ( .A1(n13028), .A2(n13029), .ZN(n12792) );
  NAND2_X1 U12893 ( .A1(n13030), .A2(b_15_), .ZN(n13029) );
  NOR2_X1 U12894 ( .A1(n13031), .A2(n8974), .ZN(n13030) );
  NOR2_X1 U12895 ( .A1(n12790), .A2(n12789), .ZN(n13031) );
  NAND2_X1 U12896 ( .A1(n12789), .A2(n12790), .ZN(n13028) );
  NAND2_X1 U12897 ( .A1(n12800), .A2(n13032), .ZN(n12790) );
  NAND2_X1 U12898 ( .A1(n12799), .A2(n12801), .ZN(n13032) );
  NAND2_X1 U12899 ( .A1(n13033), .A2(n13034), .ZN(n12801) );
  NAND2_X1 U12900 ( .A1(b_15_), .A2(a_1_), .ZN(n13034) );
  INV_X1 U12901 ( .A(n13035), .ZN(n13033) );
  XNOR2_X1 U12902 ( .A(n13036), .B(n13037), .ZN(n12799) );
  NAND2_X1 U12903 ( .A1(n13038), .A2(n13039), .ZN(n13036) );
  NAND2_X1 U12904 ( .A1(a_1_), .A2(n13035), .ZN(n12800) );
  NAND2_X1 U12905 ( .A1(n13040), .A2(n13041), .ZN(n13035) );
  NAND2_X1 U12906 ( .A1(n13042), .A2(b_15_), .ZN(n13041) );
  NOR2_X1 U12907 ( .A1(n13043), .A2(n8792), .ZN(n13042) );
  NOR2_X1 U12908 ( .A1(n12808), .A2(n12807), .ZN(n13043) );
  NAND2_X1 U12909 ( .A1(n12807), .A2(n12808), .ZN(n13040) );
  NAND2_X1 U12910 ( .A1(n13044), .A2(n13045), .ZN(n12808) );
  NAND2_X1 U12911 ( .A1(n13046), .A2(b_15_), .ZN(n13045) );
  NOR2_X1 U12912 ( .A1(n13047), .A2(n8778), .ZN(n13046) );
  NOR2_X1 U12913 ( .A1(n13019), .A2(n13018), .ZN(n13047) );
  NAND2_X1 U12914 ( .A1(n13018), .A2(n13019), .ZN(n13044) );
  NAND2_X1 U12915 ( .A1(n13048), .A2(n13049), .ZN(n13019) );
  NAND2_X1 U12916 ( .A1(n13050), .A2(b_15_), .ZN(n13049) );
  NOR2_X1 U12917 ( .A1(n13051), .A2(n8966), .ZN(n13050) );
  NOR2_X1 U12918 ( .A1(n13015), .A2(n13014), .ZN(n13051) );
  NAND2_X1 U12919 ( .A1(n13014), .A2(n13015), .ZN(n13048) );
  NAND2_X1 U12920 ( .A1(n13052), .A2(n13053), .ZN(n13015) );
  NAND2_X1 U12921 ( .A1(n13054), .A2(b_15_), .ZN(n13053) );
  NOR2_X1 U12922 ( .A1(n13055), .A2(n8723), .ZN(n13054) );
  NOR2_X1 U12923 ( .A1(n13009), .A2(n13011), .ZN(n13055) );
  NAND2_X1 U12924 ( .A1(n13009), .A2(n13011), .ZN(n13052) );
  NAND2_X1 U12925 ( .A1(n13056), .A2(n13057), .ZN(n13011) );
  NAND2_X1 U12926 ( .A1(n13058), .A2(b_15_), .ZN(n13057) );
  NOR2_X1 U12927 ( .A1(n13059), .A2(n8681), .ZN(n13058) );
  NOR2_X1 U12928 ( .A1(n13007), .A2(n13005), .ZN(n13059) );
  NAND2_X1 U12929 ( .A1(n13005), .A2(n13007), .ZN(n13056) );
  NAND2_X1 U12930 ( .A1(n13060), .A2(n13061), .ZN(n13007) );
  NAND2_X1 U12931 ( .A1(n13062), .A2(b_15_), .ZN(n13061) );
  NOR2_X1 U12932 ( .A1(n13063), .A2(n8962), .ZN(n13062) );
  NOR2_X1 U12933 ( .A1(n13003), .A2(n13002), .ZN(n13063) );
  NAND2_X1 U12934 ( .A1(n13002), .A2(n13003), .ZN(n13060) );
  NAND2_X1 U12935 ( .A1(n13064), .A2(n13065), .ZN(n13003) );
  NAND2_X1 U12936 ( .A1(n13066), .A2(b_15_), .ZN(n13065) );
  NOR2_X1 U12937 ( .A1(n13067), .A2(n8619), .ZN(n13066) );
  NOR2_X1 U12938 ( .A1(n12999), .A2(n12998), .ZN(n13067) );
  NAND2_X1 U12939 ( .A1(n12998), .A2(n12999), .ZN(n13064) );
  NAND2_X1 U12940 ( .A1(n13068), .A2(n13069), .ZN(n12999) );
  NAND2_X1 U12941 ( .A1(n13070), .A2(b_15_), .ZN(n13069) );
  NOR2_X1 U12942 ( .A1(n13071), .A2(n8605), .ZN(n13070) );
  NOR2_X1 U12943 ( .A1(n12995), .A2(n12994), .ZN(n13071) );
  NAND2_X1 U12944 ( .A1(n12994), .A2(n12995), .ZN(n13068) );
  NAND2_X1 U12945 ( .A1(n13072), .A2(n13073), .ZN(n12995) );
  NAND2_X1 U12946 ( .A1(n13074), .A2(b_15_), .ZN(n13073) );
  NOR2_X1 U12947 ( .A1(n13075), .A2(n8959), .ZN(n13074) );
  NOR2_X1 U12948 ( .A1(n12839), .A2(n12838), .ZN(n13075) );
  NAND2_X1 U12949 ( .A1(n12838), .A2(n12839), .ZN(n13072) );
  NAND2_X1 U12950 ( .A1(n13076), .A2(n13077), .ZN(n12839) );
  NAND2_X1 U12951 ( .A1(n13078), .A2(b_15_), .ZN(n13077) );
  NOR2_X1 U12952 ( .A1(n13079), .A2(n8550), .ZN(n13078) );
  NOR2_X1 U12953 ( .A1(n12991), .A2(n12989), .ZN(n13079) );
  NAND2_X1 U12954 ( .A1(n12989), .A2(n12991), .ZN(n13076) );
  NAND2_X1 U12955 ( .A1(n13080), .A2(n13081), .ZN(n12991) );
  NAND2_X1 U12956 ( .A1(n13082), .A2(b_15_), .ZN(n13081) );
  NOR2_X1 U12957 ( .A1(n13083), .A2(n8956), .ZN(n13082) );
  NOR2_X1 U12958 ( .A1(n12985), .A2(n12987), .ZN(n13083) );
  NAND2_X1 U12959 ( .A1(n12985), .A2(n12987), .ZN(n13080) );
  NAND2_X1 U12960 ( .A1(n13084), .A2(n13085), .ZN(n12987) );
  NAND2_X1 U12961 ( .A1(n13086), .A2(b_15_), .ZN(n13085) );
  NOR2_X1 U12962 ( .A1(n13087), .A2(n8495), .ZN(n13086) );
  NOR2_X1 U12963 ( .A1(n12983), .A2(n12982), .ZN(n13087) );
  NAND2_X1 U12964 ( .A1(n12982), .A2(n12983), .ZN(n13084) );
  NAND2_X1 U12965 ( .A1(n13088), .A2(n13089), .ZN(n12983) );
  NAND2_X1 U12966 ( .A1(n13090), .A2(b_15_), .ZN(n13089) );
  NOR2_X1 U12967 ( .A1(n13091), .A2(n8953), .ZN(n13090) );
  NOR2_X1 U12968 ( .A1(n12978), .A2(n12980), .ZN(n13091) );
  NAND2_X1 U12969 ( .A1(n12978), .A2(n12980), .ZN(n13088) );
  NAND2_X1 U12970 ( .A1(n13092), .A2(n13093), .ZN(n12980) );
  NAND2_X1 U12971 ( .A1(n12974), .A2(n13094), .ZN(n13093) );
  OR2_X1 U12972 ( .A1(n12975), .A2(n12976), .ZN(n13094) );
  XNOR2_X1 U12973 ( .A(n13095), .B(n13096), .ZN(n12974) );
  XNOR2_X1 U12974 ( .A(n13097), .B(n13098), .ZN(n13095) );
  NAND2_X1 U12975 ( .A1(n12976), .A2(n12975), .ZN(n13092) );
  NAND2_X1 U12976 ( .A1(n13099), .A2(n13100), .ZN(n12975) );
  NAND2_X1 U12977 ( .A1(n12972), .A2(n13101), .ZN(n13100) );
  OR2_X1 U12978 ( .A1(n12970), .A2(n12971), .ZN(n13101) );
  NOR2_X1 U12979 ( .A1(n8951), .A2(n8950), .ZN(n12972) );
  NAND2_X1 U12980 ( .A1(n12970), .A2(n12971), .ZN(n13099) );
  NAND2_X1 U12981 ( .A1(n13102), .A2(n13103), .ZN(n12971) );
  NAND2_X1 U12982 ( .A1(n12867), .A2(n13104), .ZN(n13103) );
  OR2_X1 U12983 ( .A1(n12865), .A2(n12866), .ZN(n13104) );
  NOR2_X1 U12984 ( .A1(n8951), .A2(n8385), .ZN(n12867) );
  NAND2_X1 U12985 ( .A1(n12865), .A2(n12866), .ZN(n13102) );
  NAND2_X1 U12986 ( .A1(n13105), .A2(n13106), .ZN(n12866) );
  NAND2_X1 U12987 ( .A1(n13107), .A2(b_15_), .ZN(n13106) );
  NOR2_X1 U12988 ( .A1(n13108), .A2(n8947), .ZN(n13107) );
  NOR2_X1 U12989 ( .A1(n12966), .A2(n12967), .ZN(n13108) );
  NAND2_X1 U12990 ( .A1(n12966), .A2(n12967), .ZN(n13105) );
  NAND2_X1 U12991 ( .A1(n13109), .A2(n13110), .ZN(n12967) );
  NAND2_X1 U12992 ( .A1(n12964), .A2(n13111), .ZN(n13110) );
  OR2_X1 U12993 ( .A1(n12961), .A2(n12963), .ZN(n13111) );
  NOR2_X1 U12994 ( .A1(n8951), .A2(n8324), .ZN(n12964) );
  NAND2_X1 U12995 ( .A1(n12961), .A2(n12963), .ZN(n13109) );
  NAND2_X1 U12996 ( .A1(n13112), .A2(n13113), .ZN(n12963) );
  NAND2_X1 U12997 ( .A1(n13114), .A2(b_15_), .ZN(n13113) );
  NOR2_X1 U12998 ( .A1(n13115), .A2(n8944), .ZN(n13114) );
  NOR2_X1 U12999 ( .A1(n12958), .A2(n12959), .ZN(n13115) );
  NAND2_X1 U13000 ( .A1(n12958), .A2(n12959), .ZN(n13112) );
  NAND2_X1 U13001 ( .A1(n13116), .A2(n13117), .ZN(n12959) );
  NAND2_X1 U13002 ( .A1(n12956), .A2(n13118), .ZN(n13117) );
  OR2_X1 U13003 ( .A1(n12953), .A2(n12955), .ZN(n13118) );
  NOR2_X1 U13004 ( .A1(n8951), .A2(n8268), .ZN(n12956) );
  NAND2_X1 U13005 ( .A1(n12953), .A2(n12955), .ZN(n13116) );
  NAND2_X1 U13006 ( .A1(n13119), .A2(n13120), .ZN(n12955) );
  NAND2_X1 U13007 ( .A1(n13121), .A2(b_15_), .ZN(n13120) );
  NOR2_X1 U13008 ( .A1(n13122), .A2(n8941), .ZN(n13121) );
  NOR2_X1 U13009 ( .A1(n12950), .A2(n12951), .ZN(n13122) );
  NAND2_X1 U13010 ( .A1(n12950), .A2(n12951), .ZN(n13119) );
  NAND2_X1 U13011 ( .A1(n13123), .A2(n13124), .ZN(n12951) );
  NAND2_X1 U13012 ( .A1(n12948), .A2(n13125), .ZN(n13124) );
  OR2_X1 U13013 ( .A1(n12945), .A2(n12947), .ZN(n13125) );
  NOR2_X1 U13014 ( .A1(n8951), .A2(n8213), .ZN(n12948) );
  NAND2_X1 U13015 ( .A1(n12945), .A2(n12947), .ZN(n13123) );
  NAND2_X1 U13016 ( .A1(n13126), .A2(n13127), .ZN(n12947) );
  NAND2_X1 U13017 ( .A1(n13128), .A2(b_15_), .ZN(n13127) );
  NOR2_X1 U13018 ( .A1(n13129), .A2(n8939), .ZN(n13128) );
  NOR2_X1 U13019 ( .A1(n12942), .A2(n12943), .ZN(n13129) );
  NAND2_X1 U13020 ( .A1(n12942), .A2(n12943), .ZN(n13126) );
  NAND2_X1 U13021 ( .A1(n13130), .A2(n13131), .ZN(n12943) );
  NAND2_X1 U13022 ( .A1(n12940), .A2(n13132), .ZN(n13131) );
  OR2_X1 U13023 ( .A1(n12937), .A2(n12939), .ZN(n13132) );
  NOR2_X1 U13024 ( .A1(n8951), .A2(n8158), .ZN(n12940) );
  NAND2_X1 U13025 ( .A1(n12937), .A2(n12939), .ZN(n13130) );
  NAND2_X1 U13026 ( .A1(n12935), .A2(n13133), .ZN(n12939) );
  NAND2_X1 U13027 ( .A1(n12934), .A2(n12936), .ZN(n13133) );
  NAND2_X1 U13028 ( .A1(n13134), .A2(n13135), .ZN(n12936) );
  NAND2_X1 U13029 ( .A1(b_15_), .A2(a_26_), .ZN(n13135) );
  INV_X1 U13030 ( .A(n13136), .ZN(n13134) );
  XNOR2_X1 U13031 ( .A(n13137), .B(n13138), .ZN(n12934) );
  NAND2_X1 U13032 ( .A1(n13139), .A2(n13140), .ZN(n13137) );
  NAND2_X1 U13033 ( .A1(a_26_), .A2(n13136), .ZN(n12935) );
  NAND2_X1 U13034 ( .A1(n12905), .A2(n13141), .ZN(n13136) );
  NAND2_X1 U13035 ( .A1(n12904), .A2(n12906), .ZN(n13141) );
  NAND2_X1 U13036 ( .A1(n13142), .A2(n13143), .ZN(n12906) );
  NAND2_X1 U13037 ( .A1(b_15_), .A2(a_27_), .ZN(n13143) );
  INV_X1 U13038 ( .A(n13144), .ZN(n13142) );
  XOR2_X1 U13039 ( .A(n13145), .B(n13146), .Z(n12904) );
  XNOR2_X1 U13040 ( .A(n13147), .B(n13148), .ZN(n13145) );
  NAND2_X1 U13041 ( .A1(b_14_), .A2(a_28_), .ZN(n13147) );
  NAND2_X1 U13042 ( .A1(a_27_), .A2(n13144), .ZN(n12905) );
  NAND2_X1 U13043 ( .A1(n13149), .A2(n13150), .ZN(n13144) );
  NAND2_X1 U13044 ( .A1(n13151), .A2(b_15_), .ZN(n13150) );
  NOR2_X1 U13045 ( .A1(n13152), .A2(n8055), .ZN(n13151) );
  NOR2_X1 U13046 ( .A1(n12912), .A2(n12914), .ZN(n13152) );
  NAND2_X1 U13047 ( .A1(n12912), .A2(n12914), .ZN(n13149) );
  NAND2_X1 U13048 ( .A1(n13153), .A2(n13154), .ZN(n12914) );
  NAND2_X1 U13049 ( .A1(n12930), .A2(n13155), .ZN(n13154) );
  OR2_X1 U13050 ( .A1(n12931), .A2(n12932), .ZN(n13155) );
  NOR2_X1 U13051 ( .A1(n8951), .A2(n8041), .ZN(n12930) );
  NAND2_X1 U13052 ( .A1(n12932), .A2(n12931), .ZN(n13153) );
  NAND2_X1 U13053 ( .A1(n13156), .A2(n13157), .ZN(n12931) );
  NAND2_X1 U13054 ( .A1(b_13_), .A2(n13158), .ZN(n13157) );
  NAND2_X1 U13055 ( .A1(n8003), .A2(n13159), .ZN(n13158) );
  NAND2_X1 U13056 ( .A1(a_31_), .A2(n8952), .ZN(n13159) );
  NAND2_X1 U13057 ( .A1(b_14_), .A2(n13160), .ZN(n13156) );
  NAND2_X1 U13058 ( .A1(n9341), .A2(n13161), .ZN(n13160) );
  NAND2_X1 U13059 ( .A1(a_30_), .A2(n8954), .ZN(n13161) );
  AND2_X1 U13060 ( .A1(n13162), .A2(n7953), .ZN(n12932) );
  NOR2_X1 U13061 ( .A1(n8951), .A2(n8952), .ZN(n13162) );
  XOR2_X1 U13062 ( .A(n13163), .B(n13164), .Z(n12912) );
  XOR2_X1 U13063 ( .A(n13165), .B(n13166), .Z(n13163) );
  XNOR2_X1 U13064 ( .A(n13167), .B(n13168), .ZN(n12937) );
  NAND2_X1 U13065 ( .A1(n13169), .A2(n13170), .ZN(n13167) );
  XNOR2_X1 U13066 ( .A(n13171), .B(n13172), .ZN(n12942) );
  XNOR2_X1 U13067 ( .A(n13173), .B(n13174), .ZN(n13172) );
  XOR2_X1 U13068 ( .A(n13175), .B(n13176), .Z(n12945) );
  XOR2_X1 U13069 ( .A(n13177), .B(n13178), .Z(n13175) );
  NOR2_X1 U13070 ( .A1(n8939), .A2(n8952), .ZN(n13178) );
  XNOR2_X1 U13071 ( .A(n13179), .B(n13180), .ZN(n12950) );
  XNOR2_X1 U13072 ( .A(n13181), .B(n13182), .ZN(n13180) );
  XOR2_X1 U13073 ( .A(n13183), .B(n13184), .Z(n12953) );
  XOR2_X1 U13074 ( .A(n13185), .B(n13186), .Z(n13183) );
  NOR2_X1 U13075 ( .A1(n8941), .A2(n8952), .ZN(n13186) );
  XNOR2_X1 U13076 ( .A(n13187), .B(n13188), .ZN(n12958) );
  XNOR2_X1 U13077 ( .A(n13189), .B(n13190), .ZN(n13188) );
  XOR2_X1 U13078 ( .A(n13191), .B(n13192), .Z(n12961) );
  XOR2_X1 U13079 ( .A(n13193), .B(n13194), .Z(n13191) );
  NOR2_X1 U13080 ( .A1(n8944), .A2(n8952), .ZN(n13194) );
  XNOR2_X1 U13081 ( .A(n13195), .B(n13196), .ZN(n12966) );
  XNOR2_X1 U13082 ( .A(n13197), .B(n13198), .ZN(n13196) );
  XOR2_X1 U13083 ( .A(n13199), .B(n13200), .Z(n12865) );
  XOR2_X1 U13084 ( .A(n13201), .B(n13202), .Z(n13199) );
  NOR2_X1 U13085 ( .A1(n8947), .A2(n8952), .ZN(n13202) );
  XOR2_X1 U13086 ( .A(n13203), .B(n13204), .Z(n12970) );
  XOR2_X1 U13087 ( .A(n13205), .B(n13206), .Z(n13203) );
  NOR2_X1 U13088 ( .A1(n8385), .A2(n8952), .ZN(n13206) );
  INV_X1 U13089 ( .A(n8893), .ZN(n12976) );
  NAND2_X1 U13090 ( .A1(b_15_), .A2(a_15_), .ZN(n8893) );
  XOR2_X1 U13091 ( .A(n13207), .B(n13208), .Z(n12978) );
  XOR2_X1 U13092 ( .A(n13209), .B(n13210), .Z(n13207) );
  XNOR2_X1 U13093 ( .A(n13211), .B(n13212), .ZN(n12982) );
  XOR2_X1 U13094 ( .A(n13213), .B(n8473), .Z(n13212) );
  XNOR2_X1 U13095 ( .A(n13214), .B(n13215), .ZN(n12985) );
  XOR2_X1 U13096 ( .A(n13216), .B(n13217), .Z(n13215) );
  NAND2_X1 U13097 ( .A1(b_14_), .A2(a_13_), .ZN(n13217) );
  XNOR2_X1 U13098 ( .A(n13218), .B(n13219), .ZN(n12989) );
  NAND2_X1 U13099 ( .A1(n13220), .A2(n13221), .ZN(n13218) );
  XNOR2_X1 U13100 ( .A(n13222), .B(n13223), .ZN(n12838) );
  NAND2_X1 U13101 ( .A1(n13224), .A2(n13225), .ZN(n13222) );
  XNOR2_X1 U13102 ( .A(n13226), .B(n13227), .ZN(n12994) );
  NAND2_X1 U13103 ( .A1(n13228), .A2(n13229), .ZN(n13226) );
  XNOR2_X1 U13104 ( .A(n13230), .B(n13231), .ZN(n12998) );
  XNOR2_X1 U13105 ( .A(n13232), .B(n13233), .ZN(n13230) );
  XNOR2_X1 U13106 ( .A(n13234), .B(n13235), .ZN(n13002) );
  XOR2_X1 U13107 ( .A(n13236), .B(n13237), .Z(n13235) );
  NAND2_X1 U13108 ( .A1(b_14_), .A2(a_8_), .ZN(n13237) );
  XNOR2_X1 U13109 ( .A(n13238), .B(n13239), .ZN(n13005) );
  NAND2_X1 U13110 ( .A1(n13240), .A2(n13241), .ZN(n13238) );
  XNOR2_X1 U13111 ( .A(n13242), .B(n13243), .ZN(n13009) );
  NAND2_X1 U13112 ( .A1(n13244), .A2(n13245), .ZN(n13242) );
  XNOR2_X1 U13113 ( .A(n13246), .B(n13247), .ZN(n13014) );
  XNOR2_X1 U13114 ( .A(n13248), .B(n13249), .ZN(n13246) );
  XOR2_X1 U13115 ( .A(n13250), .B(n13251), .Z(n13018) );
  XNOR2_X1 U13116 ( .A(n13252), .B(n13253), .ZN(n13250) );
  NAND2_X1 U13117 ( .A1(b_14_), .A2(a_4_), .ZN(n13252) );
  XNOR2_X1 U13118 ( .A(n13254), .B(n13255), .ZN(n12807) );
  NAND2_X1 U13119 ( .A1(n13256), .A2(n13257), .ZN(n13254) );
  XNOR2_X1 U13120 ( .A(n13258), .B(n13259), .ZN(n12789) );
  NAND2_X1 U13121 ( .A1(n13260), .A2(n13261), .ZN(n13258) );
  NOR2_X1 U13122 ( .A1(n13262), .A2(n12793), .ZN(n13026) );
  INV_X1 U13123 ( .A(n13023), .ZN(n12793) );
  XNOR2_X1 U13124 ( .A(n13263), .B(n13264), .ZN(n13023) );
  NAND2_X1 U13125 ( .A1(n13265), .A2(n13266), .ZN(n13263) );
  NOR2_X1 U13126 ( .A1(n13024), .A2(n13025), .ZN(n13262) );
  OR2_X1 U13127 ( .A1(n9146), .A2(n9145), .ZN(n9097) );
  NAND2_X1 U13128 ( .A1(n9141), .A2(n13267), .ZN(n9145) );
  NAND2_X1 U13129 ( .A1(n13268), .A2(n13269), .ZN(n13267) );
  INV_X1 U13130 ( .A(n13270), .ZN(n13269) );
  XOR2_X1 U13131 ( .A(n13271), .B(n13272), .Z(n13268) );
  NAND2_X1 U13132 ( .A1(n13024), .A2(n13025), .ZN(n9146) );
  NAND2_X1 U13133 ( .A1(n13265), .A2(n13273), .ZN(n13025) );
  NAND2_X1 U13134 ( .A1(n13264), .A2(n13266), .ZN(n13273) );
  NAND2_X1 U13135 ( .A1(n13274), .A2(n13275), .ZN(n13266) );
  NAND2_X1 U13136 ( .A1(b_14_), .A2(a_0_), .ZN(n13275) );
  INV_X1 U13137 ( .A(n13276), .ZN(n13274) );
  XOR2_X1 U13138 ( .A(n13277), .B(n13278), .Z(n13264) );
  XOR2_X1 U13139 ( .A(n13279), .B(n13280), .Z(n13277) );
  NOR2_X1 U13140 ( .A1(n8969), .A2(n8954), .ZN(n13280) );
  NAND2_X1 U13141 ( .A1(a_0_), .A2(n13276), .ZN(n13265) );
  NAND2_X1 U13142 ( .A1(n13260), .A2(n13281), .ZN(n13276) );
  NAND2_X1 U13143 ( .A1(n13259), .A2(n13261), .ZN(n13281) );
  NAND2_X1 U13144 ( .A1(n13282), .A2(n13283), .ZN(n13261) );
  NAND2_X1 U13145 ( .A1(b_14_), .A2(a_1_), .ZN(n13283) );
  INV_X1 U13146 ( .A(n13284), .ZN(n13282) );
  XOR2_X1 U13147 ( .A(n13285), .B(n13286), .Z(n13259) );
  XOR2_X1 U13148 ( .A(n13287), .B(n13288), .Z(n13285) );
  NOR2_X1 U13149 ( .A1(n8792), .A2(n8954), .ZN(n13288) );
  NAND2_X1 U13150 ( .A1(a_1_), .A2(n13284), .ZN(n13260) );
  NAND2_X1 U13151 ( .A1(n13038), .A2(n13289), .ZN(n13284) );
  NAND2_X1 U13152 ( .A1(n13037), .A2(n13039), .ZN(n13289) );
  NAND2_X1 U13153 ( .A1(n13290), .A2(n13291), .ZN(n13039) );
  NAND2_X1 U13154 ( .A1(b_14_), .A2(a_2_), .ZN(n13291) );
  INV_X1 U13155 ( .A(n13292), .ZN(n13290) );
  XOR2_X1 U13156 ( .A(n13293), .B(n13294), .Z(n13037) );
  XOR2_X1 U13157 ( .A(n13295), .B(n13296), .Z(n13293) );
  NOR2_X1 U13158 ( .A1(n8778), .A2(n8954), .ZN(n13296) );
  NAND2_X1 U13159 ( .A1(a_2_), .A2(n13292), .ZN(n13038) );
  NAND2_X1 U13160 ( .A1(n13256), .A2(n13297), .ZN(n13292) );
  NAND2_X1 U13161 ( .A1(n13255), .A2(n13257), .ZN(n13297) );
  NAND2_X1 U13162 ( .A1(n13298), .A2(n13299), .ZN(n13257) );
  NAND2_X1 U13163 ( .A1(b_14_), .A2(a_3_), .ZN(n13299) );
  INV_X1 U13164 ( .A(n13300), .ZN(n13298) );
  XNOR2_X1 U13165 ( .A(n13301), .B(n13302), .ZN(n13255) );
  XOR2_X1 U13166 ( .A(n13303), .B(n13304), .Z(n13302) );
  NAND2_X1 U13167 ( .A1(b_13_), .A2(a_4_), .ZN(n13304) );
  NAND2_X1 U13168 ( .A1(a_3_), .A2(n13300), .ZN(n13256) );
  NAND2_X1 U13169 ( .A1(n13305), .A2(n13306), .ZN(n13300) );
  NAND2_X1 U13170 ( .A1(n13307), .A2(b_14_), .ZN(n13306) );
  NOR2_X1 U13171 ( .A1(n13308), .A2(n8966), .ZN(n13307) );
  NOR2_X1 U13172 ( .A1(n13251), .A2(n13253), .ZN(n13308) );
  NAND2_X1 U13173 ( .A1(n13251), .A2(n13253), .ZN(n13305) );
  NAND2_X1 U13174 ( .A1(n13309), .A2(n13310), .ZN(n13253) );
  NAND2_X1 U13175 ( .A1(n13249), .A2(n13311), .ZN(n13310) );
  NAND2_X1 U13176 ( .A1(n13248), .A2(n13247), .ZN(n13311) );
  NOR2_X1 U13177 ( .A1(n8952), .A2(n8723), .ZN(n13249) );
  OR2_X1 U13178 ( .A1(n13247), .A2(n13248), .ZN(n13309) );
  AND2_X1 U13179 ( .A1(n13244), .A2(n13312), .ZN(n13248) );
  NAND2_X1 U13180 ( .A1(n13243), .A2(n13245), .ZN(n13312) );
  NAND2_X1 U13181 ( .A1(n13313), .A2(n13314), .ZN(n13245) );
  NAND2_X1 U13182 ( .A1(b_14_), .A2(a_6_), .ZN(n13314) );
  INV_X1 U13183 ( .A(n13315), .ZN(n13313) );
  XOR2_X1 U13184 ( .A(n13316), .B(n13317), .Z(n13243) );
  XOR2_X1 U13185 ( .A(n13318), .B(n13319), .Z(n13316) );
  NOR2_X1 U13186 ( .A1(n8962), .A2(n8954), .ZN(n13319) );
  NAND2_X1 U13187 ( .A1(a_6_), .A2(n13315), .ZN(n13244) );
  NAND2_X1 U13188 ( .A1(n13240), .A2(n13320), .ZN(n13315) );
  NAND2_X1 U13189 ( .A1(n13239), .A2(n13241), .ZN(n13320) );
  NAND2_X1 U13190 ( .A1(n13321), .A2(n13322), .ZN(n13241) );
  NAND2_X1 U13191 ( .A1(b_14_), .A2(a_7_), .ZN(n13322) );
  INV_X1 U13192 ( .A(n13323), .ZN(n13321) );
  XOR2_X1 U13193 ( .A(n13324), .B(n13325), .Z(n13239) );
  XOR2_X1 U13194 ( .A(n13326), .B(n13327), .Z(n13324) );
  NOR2_X1 U13195 ( .A1(n8619), .A2(n8954), .ZN(n13327) );
  NAND2_X1 U13196 ( .A1(a_7_), .A2(n13323), .ZN(n13240) );
  NAND2_X1 U13197 ( .A1(n13328), .A2(n13329), .ZN(n13323) );
  NAND2_X1 U13198 ( .A1(n13330), .A2(b_14_), .ZN(n13329) );
  NOR2_X1 U13199 ( .A1(n13331), .A2(n8619), .ZN(n13330) );
  NOR2_X1 U13200 ( .A1(n13234), .A2(n13236), .ZN(n13331) );
  NAND2_X1 U13201 ( .A1(n13234), .A2(n13236), .ZN(n13328) );
  NAND2_X1 U13202 ( .A1(n13332), .A2(n13333), .ZN(n13236) );
  NAND2_X1 U13203 ( .A1(n13233), .A2(n13334), .ZN(n13333) );
  NAND2_X1 U13204 ( .A1(n13232), .A2(n13231), .ZN(n13334) );
  NOR2_X1 U13205 ( .A1(n8952), .A2(n8605), .ZN(n13233) );
  OR2_X1 U13206 ( .A1(n13231), .A2(n13232), .ZN(n13332) );
  AND2_X1 U13207 ( .A1(n13228), .A2(n13335), .ZN(n13232) );
  NAND2_X1 U13208 ( .A1(n13227), .A2(n13229), .ZN(n13335) );
  NAND2_X1 U13209 ( .A1(n13336), .A2(n13337), .ZN(n13229) );
  NAND2_X1 U13210 ( .A1(b_14_), .A2(a_10_), .ZN(n13337) );
  INV_X1 U13211 ( .A(n13338), .ZN(n13336) );
  XOR2_X1 U13212 ( .A(n13339), .B(n13340), .Z(n13227) );
  XOR2_X1 U13213 ( .A(n13341), .B(n13342), .Z(n13339) );
  NOR2_X1 U13214 ( .A1(n8550), .A2(n8954), .ZN(n13342) );
  NAND2_X1 U13215 ( .A1(a_10_), .A2(n13338), .ZN(n13228) );
  NAND2_X1 U13216 ( .A1(n13224), .A2(n13343), .ZN(n13338) );
  NAND2_X1 U13217 ( .A1(n13223), .A2(n13225), .ZN(n13343) );
  NAND2_X1 U13218 ( .A1(n13344), .A2(n13345), .ZN(n13225) );
  NAND2_X1 U13219 ( .A1(b_14_), .A2(a_11_), .ZN(n13345) );
  INV_X1 U13220 ( .A(n13346), .ZN(n13344) );
  XOR2_X1 U13221 ( .A(n13347), .B(n13348), .Z(n13223) );
  XNOR2_X1 U13222 ( .A(n13349), .B(n13350), .ZN(n13347) );
  NAND2_X1 U13223 ( .A1(b_13_), .A2(a_12_), .ZN(n13349) );
  NAND2_X1 U13224 ( .A1(a_11_), .A2(n13346), .ZN(n13224) );
  NAND2_X1 U13225 ( .A1(n13220), .A2(n13351), .ZN(n13346) );
  NAND2_X1 U13226 ( .A1(n13219), .A2(n13221), .ZN(n13351) );
  NAND2_X1 U13227 ( .A1(n13352), .A2(n13353), .ZN(n13221) );
  NAND2_X1 U13228 ( .A1(b_14_), .A2(a_12_), .ZN(n13353) );
  INV_X1 U13229 ( .A(n13354), .ZN(n13352) );
  XOR2_X1 U13230 ( .A(n13355), .B(n13356), .Z(n13219) );
  XOR2_X1 U13231 ( .A(n13357), .B(n13358), .Z(n13355) );
  NAND2_X1 U13232 ( .A1(a_12_), .A2(n13354), .ZN(n13220) );
  NAND2_X1 U13233 ( .A1(n13359), .A2(n13360), .ZN(n13354) );
  NAND2_X1 U13234 ( .A1(n13361), .A2(b_14_), .ZN(n13360) );
  NOR2_X1 U13235 ( .A1(n13362), .A2(n8495), .ZN(n13361) );
  NOR2_X1 U13236 ( .A1(n13214), .A2(n13216), .ZN(n13362) );
  NAND2_X1 U13237 ( .A1(n13214), .A2(n13216), .ZN(n13359) );
  NAND2_X1 U13238 ( .A1(n13363), .A2(n13364), .ZN(n13216) );
  NAND2_X1 U13239 ( .A1(n13365), .A2(n13366), .ZN(n13364) );
  OR2_X1 U13240 ( .A1(n13213), .A2(n13211), .ZN(n13366) );
  INV_X1 U13241 ( .A(n8473), .ZN(n13365) );
  NAND2_X1 U13242 ( .A1(b_14_), .A2(a_14_), .ZN(n8473) );
  NAND2_X1 U13243 ( .A1(n13211), .A2(n13213), .ZN(n13363) );
  NAND2_X1 U13244 ( .A1(n13367), .A2(n13368), .ZN(n13213) );
  NAND2_X1 U13245 ( .A1(n13210), .A2(n13369), .ZN(n13368) );
  OR2_X1 U13246 ( .A1(n13209), .A2(n13208), .ZN(n13369) );
  NOR2_X1 U13247 ( .A1(n8952), .A2(n8440), .ZN(n13210) );
  NAND2_X1 U13248 ( .A1(n13208), .A2(n13209), .ZN(n13367) );
  NAND2_X1 U13249 ( .A1(n13370), .A2(n13371), .ZN(n13209) );
  NAND2_X1 U13250 ( .A1(n13098), .A2(n13372), .ZN(n13371) );
  NAND2_X1 U13251 ( .A1(n13097), .A2(n13096), .ZN(n13372) );
  NOR2_X1 U13252 ( .A1(n8952), .A2(n8950), .ZN(n13098) );
  OR2_X1 U13253 ( .A1(n13096), .A2(n13097), .ZN(n13370) );
  AND2_X1 U13254 ( .A1(n13373), .A2(n13374), .ZN(n13097) );
  NAND2_X1 U13255 ( .A1(n13375), .A2(b_14_), .ZN(n13374) );
  NOR2_X1 U13256 ( .A1(n13376), .A2(n8385), .ZN(n13375) );
  NOR2_X1 U13257 ( .A1(n13204), .A2(n13205), .ZN(n13376) );
  NAND2_X1 U13258 ( .A1(n13204), .A2(n13205), .ZN(n13373) );
  NAND2_X1 U13259 ( .A1(n13377), .A2(n13378), .ZN(n13205) );
  NAND2_X1 U13260 ( .A1(n13379), .A2(b_14_), .ZN(n13378) );
  NOR2_X1 U13261 ( .A1(n13380), .A2(n8947), .ZN(n13379) );
  NOR2_X1 U13262 ( .A1(n13200), .A2(n13201), .ZN(n13380) );
  NAND2_X1 U13263 ( .A1(n13200), .A2(n13201), .ZN(n13377) );
  NAND2_X1 U13264 ( .A1(n13381), .A2(n13382), .ZN(n13201) );
  NAND2_X1 U13265 ( .A1(n13198), .A2(n13383), .ZN(n13382) );
  OR2_X1 U13266 ( .A1(n13197), .A2(n13195), .ZN(n13383) );
  NOR2_X1 U13267 ( .A1(n8952), .A2(n8324), .ZN(n13198) );
  NAND2_X1 U13268 ( .A1(n13195), .A2(n13197), .ZN(n13381) );
  NAND2_X1 U13269 ( .A1(n13384), .A2(n13385), .ZN(n13197) );
  NAND2_X1 U13270 ( .A1(n13386), .A2(b_14_), .ZN(n13385) );
  NOR2_X1 U13271 ( .A1(n13387), .A2(n8944), .ZN(n13386) );
  NOR2_X1 U13272 ( .A1(n13192), .A2(n13193), .ZN(n13387) );
  NAND2_X1 U13273 ( .A1(n13192), .A2(n13193), .ZN(n13384) );
  NAND2_X1 U13274 ( .A1(n13388), .A2(n13389), .ZN(n13193) );
  NAND2_X1 U13275 ( .A1(n13190), .A2(n13390), .ZN(n13389) );
  OR2_X1 U13276 ( .A1(n13189), .A2(n13187), .ZN(n13390) );
  NOR2_X1 U13277 ( .A1(n8952), .A2(n8268), .ZN(n13190) );
  NAND2_X1 U13278 ( .A1(n13187), .A2(n13189), .ZN(n13388) );
  NAND2_X1 U13279 ( .A1(n13391), .A2(n13392), .ZN(n13189) );
  NAND2_X1 U13280 ( .A1(n13393), .A2(b_14_), .ZN(n13392) );
  NOR2_X1 U13281 ( .A1(n13394), .A2(n8941), .ZN(n13393) );
  NOR2_X1 U13282 ( .A1(n13184), .A2(n13185), .ZN(n13394) );
  NAND2_X1 U13283 ( .A1(n13184), .A2(n13185), .ZN(n13391) );
  NAND2_X1 U13284 ( .A1(n13395), .A2(n13396), .ZN(n13185) );
  NAND2_X1 U13285 ( .A1(n13182), .A2(n13397), .ZN(n13396) );
  OR2_X1 U13286 ( .A1(n13181), .A2(n13179), .ZN(n13397) );
  NOR2_X1 U13287 ( .A1(n8952), .A2(n8213), .ZN(n13182) );
  NAND2_X1 U13288 ( .A1(n13179), .A2(n13181), .ZN(n13395) );
  NAND2_X1 U13289 ( .A1(n13398), .A2(n13399), .ZN(n13181) );
  NAND2_X1 U13290 ( .A1(n13400), .A2(b_14_), .ZN(n13399) );
  NOR2_X1 U13291 ( .A1(n13401), .A2(n8939), .ZN(n13400) );
  NOR2_X1 U13292 ( .A1(n13176), .A2(n13177), .ZN(n13401) );
  NAND2_X1 U13293 ( .A1(n13176), .A2(n13177), .ZN(n13398) );
  NAND2_X1 U13294 ( .A1(n13402), .A2(n13403), .ZN(n13177) );
  NAND2_X1 U13295 ( .A1(n13174), .A2(n13404), .ZN(n13403) );
  OR2_X1 U13296 ( .A1(n13173), .A2(n13171), .ZN(n13404) );
  NOR2_X1 U13297 ( .A1(n8952), .A2(n8158), .ZN(n13174) );
  NAND2_X1 U13298 ( .A1(n13171), .A2(n13173), .ZN(n13402) );
  NAND2_X1 U13299 ( .A1(n13169), .A2(n13405), .ZN(n13173) );
  NAND2_X1 U13300 ( .A1(n13168), .A2(n13170), .ZN(n13405) );
  NAND2_X1 U13301 ( .A1(n13406), .A2(n13407), .ZN(n13170) );
  NAND2_X1 U13302 ( .A1(b_14_), .A2(a_26_), .ZN(n13407) );
  INV_X1 U13303 ( .A(n13408), .ZN(n13406) );
  XNOR2_X1 U13304 ( .A(n13409), .B(n13410), .ZN(n13168) );
  NAND2_X1 U13305 ( .A1(n13411), .A2(n13412), .ZN(n13409) );
  NAND2_X1 U13306 ( .A1(a_26_), .A2(n13408), .ZN(n13169) );
  NAND2_X1 U13307 ( .A1(n13139), .A2(n13413), .ZN(n13408) );
  NAND2_X1 U13308 ( .A1(n13138), .A2(n13140), .ZN(n13413) );
  NAND2_X1 U13309 ( .A1(n13414), .A2(n13415), .ZN(n13140) );
  NAND2_X1 U13310 ( .A1(b_14_), .A2(a_27_), .ZN(n13415) );
  INV_X1 U13311 ( .A(n13416), .ZN(n13414) );
  XOR2_X1 U13312 ( .A(n13417), .B(n13418), .Z(n13138) );
  XNOR2_X1 U13313 ( .A(n13419), .B(n13420), .ZN(n13417) );
  NAND2_X1 U13314 ( .A1(b_13_), .A2(a_28_), .ZN(n13419) );
  NAND2_X1 U13315 ( .A1(a_27_), .A2(n13416), .ZN(n13139) );
  NAND2_X1 U13316 ( .A1(n13421), .A2(n13422), .ZN(n13416) );
  NAND2_X1 U13317 ( .A1(n13423), .A2(b_14_), .ZN(n13422) );
  NOR2_X1 U13318 ( .A1(n13424), .A2(n8055), .ZN(n13423) );
  NOR2_X1 U13319 ( .A1(n13146), .A2(n13148), .ZN(n13424) );
  NAND2_X1 U13320 ( .A1(n13146), .A2(n13148), .ZN(n13421) );
  NAND2_X1 U13321 ( .A1(n13425), .A2(n13426), .ZN(n13148) );
  NAND2_X1 U13322 ( .A1(n13164), .A2(n13427), .ZN(n13426) );
  OR2_X1 U13323 ( .A1(n13165), .A2(n13166), .ZN(n13427) );
  NOR2_X1 U13324 ( .A1(n8952), .A2(n8041), .ZN(n13164) );
  NAND2_X1 U13325 ( .A1(n13166), .A2(n13165), .ZN(n13425) );
  NAND2_X1 U13326 ( .A1(n13428), .A2(n13429), .ZN(n13165) );
  NAND2_X1 U13327 ( .A1(b_12_), .A2(n13430), .ZN(n13429) );
  NAND2_X1 U13328 ( .A1(n8003), .A2(n13431), .ZN(n13430) );
  NAND2_X1 U13329 ( .A1(a_31_), .A2(n8954), .ZN(n13431) );
  NAND2_X1 U13330 ( .A1(b_13_), .A2(n13432), .ZN(n13428) );
  NAND2_X1 U13331 ( .A1(n9341), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U13332 ( .A1(a_30_), .A2(n8955), .ZN(n13433) );
  AND2_X1 U13333 ( .A1(n13434), .A2(n7953), .ZN(n13166) );
  NOR2_X1 U13334 ( .A1(n8952), .A2(n8954), .ZN(n13434) );
  XOR2_X1 U13335 ( .A(n13435), .B(n13436), .Z(n13146) );
  XOR2_X1 U13336 ( .A(n13437), .B(n13438), .Z(n13435) );
  XNOR2_X1 U13337 ( .A(n13439), .B(n13440), .ZN(n13171) );
  NAND2_X1 U13338 ( .A1(n13441), .A2(n13442), .ZN(n13439) );
  XNOR2_X1 U13339 ( .A(n13443), .B(n13444), .ZN(n13176) );
  XNOR2_X1 U13340 ( .A(n13445), .B(n13446), .ZN(n13444) );
  XOR2_X1 U13341 ( .A(n13447), .B(n13448), .Z(n13179) );
  XOR2_X1 U13342 ( .A(n13449), .B(n13450), .Z(n13447) );
  NOR2_X1 U13343 ( .A1(n8939), .A2(n8954), .ZN(n13450) );
  XNOR2_X1 U13344 ( .A(n13451), .B(n13452), .ZN(n13184) );
  XNOR2_X1 U13345 ( .A(n13453), .B(n13454), .ZN(n13452) );
  XOR2_X1 U13346 ( .A(n13455), .B(n13456), .Z(n13187) );
  XOR2_X1 U13347 ( .A(n13457), .B(n13458), .Z(n13455) );
  NOR2_X1 U13348 ( .A1(n8941), .A2(n8954), .ZN(n13458) );
  XNOR2_X1 U13349 ( .A(n13459), .B(n13460), .ZN(n13192) );
  XNOR2_X1 U13350 ( .A(n13461), .B(n13462), .ZN(n13460) );
  XOR2_X1 U13351 ( .A(n13463), .B(n13464), .Z(n13195) );
  XOR2_X1 U13352 ( .A(n13465), .B(n13466), .Z(n13463) );
  NOR2_X1 U13353 ( .A1(n8944), .A2(n8954), .ZN(n13466) );
  XNOR2_X1 U13354 ( .A(n13467), .B(n13468), .ZN(n13200) );
  XNOR2_X1 U13355 ( .A(n13469), .B(n13470), .ZN(n13468) );
  XOR2_X1 U13356 ( .A(n13471), .B(n13472), .Z(n13204) );
  XOR2_X1 U13357 ( .A(n13473), .B(n13474), .Z(n13471) );
  XNOR2_X1 U13358 ( .A(n13475), .B(n13476), .ZN(n13096) );
  XOR2_X1 U13359 ( .A(n13477), .B(n13478), .Z(n13475) );
  NOR2_X1 U13360 ( .A1(n8385), .A2(n8954), .ZN(n13478) );
  XOR2_X1 U13361 ( .A(n13479), .B(n13480), .Z(n13208) );
  XOR2_X1 U13362 ( .A(n13481), .B(n13482), .Z(n13479) );
  NOR2_X1 U13363 ( .A1(n8950), .A2(n8954), .ZN(n13482) );
  XOR2_X1 U13364 ( .A(n13483), .B(n13484), .Z(n13211) );
  XOR2_X1 U13365 ( .A(n13485), .B(n13486), .Z(n13483) );
  NOR2_X1 U13366 ( .A1(n8440), .A2(n8954), .ZN(n13486) );
  XOR2_X1 U13367 ( .A(n13487), .B(n13488), .Z(n13214) );
  XOR2_X1 U13368 ( .A(n13489), .B(n13490), .Z(n13487) );
  NOR2_X1 U13369 ( .A1(n8953), .A2(n8954), .ZN(n13490) );
  XNOR2_X1 U13370 ( .A(n13491), .B(n13492), .ZN(n13231) );
  XOR2_X1 U13371 ( .A(n13493), .B(n13494), .Z(n13491) );
  NOR2_X1 U13372 ( .A1(n8959), .A2(n8954), .ZN(n13494) );
  XOR2_X1 U13373 ( .A(n13495), .B(n13496), .Z(n13234) );
  XOR2_X1 U13374 ( .A(n13497), .B(n13498), .Z(n13495) );
  NOR2_X1 U13375 ( .A1(n8605), .A2(n8954), .ZN(n13498) );
  XOR2_X1 U13376 ( .A(n13499), .B(n13500), .Z(n13247) );
  XOR2_X1 U13377 ( .A(n13501), .B(n13502), .Z(n13500) );
  NAND2_X1 U13378 ( .A1(b_13_), .A2(a_6_), .ZN(n13502) );
  XNOR2_X1 U13379 ( .A(n13503), .B(n13504), .ZN(n13251) );
  XOR2_X1 U13380 ( .A(n13505), .B(n13506), .Z(n13504) );
  NAND2_X1 U13381 ( .A1(b_13_), .A2(a_5_), .ZN(n13506) );
  XNOR2_X1 U13382 ( .A(n13507), .B(n13508), .ZN(n13024) );
  XNOR2_X1 U13383 ( .A(n13509), .B(n13510), .ZN(n13508) );
  OR2_X1 U13384 ( .A1(n13511), .A2(n9141), .ZN(n9104) );
  NAND2_X1 U13385 ( .A1(n13512), .A2(n13270), .ZN(n9141) );
  NAND2_X1 U13386 ( .A1(n13513), .A2(n13514), .ZN(n13270) );
  NAND2_X1 U13387 ( .A1(n13510), .A2(n13515), .ZN(n13514) );
  OR2_X1 U13388 ( .A1(n13509), .A2(n13507), .ZN(n13515) );
  NOR2_X1 U13389 ( .A1(n8954), .A2(n8974), .ZN(n13510) );
  NAND2_X1 U13390 ( .A1(n13507), .A2(n13509), .ZN(n13513) );
  NAND2_X1 U13391 ( .A1(n13516), .A2(n13517), .ZN(n13509) );
  NAND2_X1 U13392 ( .A1(n13518), .A2(b_13_), .ZN(n13517) );
  NOR2_X1 U13393 ( .A1(n13519), .A2(n8969), .ZN(n13518) );
  NOR2_X1 U13394 ( .A1(n13278), .A2(n13279), .ZN(n13519) );
  NAND2_X1 U13395 ( .A1(n13278), .A2(n13279), .ZN(n13516) );
  NAND2_X1 U13396 ( .A1(n13520), .A2(n13521), .ZN(n13279) );
  NAND2_X1 U13397 ( .A1(n13522), .A2(b_13_), .ZN(n13521) );
  NOR2_X1 U13398 ( .A1(n13523), .A2(n8792), .ZN(n13522) );
  NOR2_X1 U13399 ( .A1(n13286), .A2(n13287), .ZN(n13523) );
  NAND2_X1 U13400 ( .A1(n13286), .A2(n13287), .ZN(n13520) );
  NAND2_X1 U13401 ( .A1(n13524), .A2(n13525), .ZN(n13287) );
  NAND2_X1 U13402 ( .A1(n13526), .A2(b_13_), .ZN(n13525) );
  NOR2_X1 U13403 ( .A1(n13527), .A2(n8778), .ZN(n13526) );
  NOR2_X1 U13404 ( .A1(n13294), .A2(n13295), .ZN(n13527) );
  NAND2_X1 U13405 ( .A1(n13294), .A2(n13295), .ZN(n13524) );
  NAND2_X1 U13406 ( .A1(n13528), .A2(n13529), .ZN(n13295) );
  NAND2_X1 U13407 ( .A1(n13530), .A2(b_13_), .ZN(n13529) );
  NOR2_X1 U13408 ( .A1(n13531), .A2(n8966), .ZN(n13530) );
  NOR2_X1 U13409 ( .A1(n13301), .A2(n13303), .ZN(n13531) );
  NAND2_X1 U13410 ( .A1(n13301), .A2(n13303), .ZN(n13528) );
  NAND2_X1 U13411 ( .A1(n13532), .A2(n13533), .ZN(n13303) );
  NAND2_X1 U13412 ( .A1(n13534), .A2(b_13_), .ZN(n13533) );
  NOR2_X1 U13413 ( .A1(n13535), .A2(n8723), .ZN(n13534) );
  NOR2_X1 U13414 ( .A1(n13503), .A2(n13505), .ZN(n13535) );
  NAND2_X1 U13415 ( .A1(n13503), .A2(n13505), .ZN(n13532) );
  NAND2_X1 U13416 ( .A1(n13536), .A2(n13537), .ZN(n13505) );
  NAND2_X1 U13417 ( .A1(n13538), .A2(b_13_), .ZN(n13537) );
  NOR2_X1 U13418 ( .A1(n13539), .A2(n8681), .ZN(n13538) );
  NOR2_X1 U13419 ( .A1(n13499), .A2(n13501), .ZN(n13539) );
  NAND2_X1 U13420 ( .A1(n13499), .A2(n13501), .ZN(n13536) );
  NAND2_X1 U13421 ( .A1(n13540), .A2(n13541), .ZN(n13501) );
  NAND2_X1 U13422 ( .A1(n13542), .A2(b_13_), .ZN(n13541) );
  NOR2_X1 U13423 ( .A1(n13543), .A2(n8962), .ZN(n13542) );
  NOR2_X1 U13424 ( .A1(n13317), .A2(n13318), .ZN(n13543) );
  NAND2_X1 U13425 ( .A1(n13317), .A2(n13318), .ZN(n13540) );
  NAND2_X1 U13426 ( .A1(n13544), .A2(n13545), .ZN(n13318) );
  NAND2_X1 U13427 ( .A1(n13546), .A2(b_13_), .ZN(n13545) );
  NOR2_X1 U13428 ( .A1(n13547), .A2(n8619), .ZN(n13546) );
  NOR2_X1 U13429 ( .A1(n13325), .A2(n13326), .ZN(n13547) );
  NAND2_X1 U13430 ( .A1(n13325), .A2(n13326), .ZN(n13544) );
  NAND2_X1 U13431 ( .A1(n13548), .A2(n13549), .ZN(n13326) );
  NAND2_X1 U13432 ( .A1(n13550), .A2(b_13_), .ZN(n13549) );
  NOR2_X1 U13433 ( .A1(n13551), .A2(n8605), .ZN(n13550) );
  NOR2_X1 U13434 ( .A1(n13496), .A2(n13497), .ZN(n13551) );
  NAND2_X1 U13435 ( .A1(n13496), .A2(n13497), .ZN(n13548) );
  NAND2_X1 U13436 ( .A1(n13552), .A2(n13553), .ZN(n13497) );
  NAND2_X1 U13437 ( .A1(n13554), .A2(b_13_), .ZN(n13553) );
  NOR2_X1 U13438 ( .A1(n13555), .A2(n8959), .ZN(n13554) );
  NOR2_X1 U13439 ( .A1(n13492), .A2(n13493), .ZN(n13555) );
  NAND2_X1 U13440 ( .A1(n13492), .A2(n13493), .ZN(n13552) );
  NAND2_X1 U13441 ( .A1(n13556), .A2(n13557), .ZN(n13493) );
  NAND2_X1 U13442 ( .A1(n13558), .A2(b_13_), .ZN(n13557) );
  NOR2_X1 U13443 ( .A1(n13559), .A2(n8550), .ZN(n13558) );
  NOR2_X1 U13444 ( .A1(n13340), .A2(n13341), .ZN(n13559) );
  NAND2_X1 U13445 ( .A1(n13340), .A2(n13341), .ZN(n13556) );
  NAND2_X1 U13446 ( .A1(n13560), .A2(n13561), .ZN(n13341) );
  NAND2_X1 U13447 ( .A1(n13562), .A2(b_13_), .ZN(n13561) );
  NOR2_X1 U13448 ( .A1(n13563), .A2(n8956), .ZN(n13562) );
  NOR2_X1 U13449 ( .A1(n13348), .A2(n13350), .ZN(n13563) );
  NAND2_X1 U13450 ( .A1(n13348), .A2(n13350), .ZN(n13560) );
  NAND2_X1 U13451 ( .A1(n13564), .A2(n13565), .ZN(n13350) );
  NAND2_X1 U13452 ( .A1(n13356), .A2(n13566), .ZN(n13565) );
  OR2_X1 U13453 ( .A1(n13357), .A2(n13358), .ZN(n13566) );
  XNOR2_X1 U13454 ( .A(n13567), .B(n13568), .ZN(n13356) );
  NAND2_X1 U13455 ( .A1(n13569), .A2(n13570), .ZN(n13567) );
  NAND2_X1 U13456 ( .A1(n13358), .A2(n13357), .ZN(n13564) );
  NAND2_X1 U13457 ( .A1(n13571), .A2(n13572), .ZN(n13357) );
  NAND2_X1 U13458 ( .A1(n13573), .A2(b_13_), .ZN(n13572) );
  NOR2_X1 U13459 ( .A1(n13574), .A2(n8953), .ZN(n13573) );
  NOR2_X1 U13460 ( .A1(n13488), .A2(n13489), .ZN(n13574) );
  NAND2_X1 U13461 ( .A1(n13488), .A2(n13489), .ZN(n13571) );
  NAND2_X1 U13462 ( .A1(n13575), .A2(n13576), .ZN(n13489) );
  NAND2_X1 U13463 ( .A1(n13577), .A2(b_13_), .ZN(n13576) );
  NOR2_X1 U13464 ( .A1(n13578), .A2(n8440), .ZN(n13577) );
  NOR2_X1 U13465 ( .A1(n13484), .A2(n13485), .ZN(n13578) );
  NAND2_X1 U13466 ( .A1(n13484), .A2(n13485), .ZN(n13575) );
  NAND2_X1 U13467 ( .A1(n13579), .A2(n13580), .ZN(n13485) );
  NAND2_X1 U13468 ( .A1(n13581), .A2(b_13_), .ZN(n13580) );
  NOR2_X1 U13469 ( .A1(n13582), .A2(n8950), .ZN(n13581) );
  NOR2_X1 U13470 ( .A1(n13480), .A2(n13481), .ZN(n13582) );
  NAND2_X1 U13471 ( .A1(n13480), .A2(n13481), .ZN(n13579) );
  NAND2_X1 U13472 ( .A1(n13583), .A2(n13584), .ZN(n13481) );
  NAND2_X1 U13473 ( .A1(n13585), .A2(b_13_), .ZN(n13584) );
  NOR2_X1 U13474 ( .A1(n13586), .A2(n8385), .ZN(n13585) );
  NOR2_X1 U13475 ( .A1(n13476), .A2(n13477), .ZN(n13586) );
  NAND2_X1 U13476 ( .A1(n13476), .A2(n13477), .ZN(n13583) );
  NAND2_X1 U13477 ( .A1(n13587), .A2(n13588), .ZN(n13477) );
  NAND2_X1 U13478 ( .A1(n13474), .A2(n13589), .ZN(n13588) );
  OR2_X1 U13479 ( .A1(n13473), .A2(n13472), .ZN(n13589) );
  NOR2_X1 U13480 ( .A1(n8954), .A2(n8947), .ZN(n13474) );
  NAND2_X1 U13481 ( .A1(n13472), .A2(n13473), .ZN(n13587) );
  NAND2_X1 U13482 ( .A1(n13590), .A2(n13591), .ZN(n13473) );
  NAND2_X1 U13483 ( .A1(n13470), .A2(n13592), .ZN(n13591) );
  OR2_X1 U13484 ( .A1(n13469), .A2(n13467), .ZN(n13592) );
  NOR2_X1 U13485 ( .A1(n8954), .A2(n8324), .ZN(n13470) );
  NAND2_X1 U13486 ( .A1(n13467), .A2(n13469), .ZN(n13590) );
  NAND2_X1 U13487 ( .A1(n13593), .A2(n13594), .ZN(n13469) );
  NAND2_X1 U13488 ( .A1(n13595), .A2(b_13_), .ZN(n13594) );
  NOR2_X1 U13489 ( .A1(n13596), .A2(n8944), .ZN(n13595) );
  NOR2_X1 U13490 ( .A1(n13464), .A2(n13465), .ZN(n13596) );
  NAND2_X1 U13491 ( .A1(n13464), .A2(n13465), .ZN(n13593) );
  NAND2_X1 U13492 ( .A1(n13597), .A2(n13598), .ZN(n13465) );
  NAND2_X1 U13493 ( .A1(n13462), .A2(n13599), .ZN(n13598) );
  OR2_X1 U13494 ( .A1(n13461), .A2(n13459), .ZN(n13599) );
  NOR2_X1 U13495 ( .A1(n8954), .A2(n8268), .ZN(n13462) );
  NAND2_X1 U13496 ( .A1(n13459), .A2(n13461), .ZN(n13597) );
  NAND2_X1 U13497 ( .A1(n13600), .A2(n13601), .ZN(n13461) );
  NAND2_X1 U13498 ( .A1(n13602), .A2(b_13_), .ZN(n13601) );
  NOR2_X1 U13499 ( .A1(n13603), .A2(n8941), .ZN(n13602) );
  NOR2_X1 U13500 ( .A1(n13456), .A2(n13457), .ZN(n13603) );
  NAND2_X1 U13501 ( .A1(n13456), .A2(n13457), .ZN(n13600) );
  NAND2_X1 U13502 ( .A1(n13604), .A2(n13605), .ZN(n13457) );
  NAND2_X1 U13503 ( .A1(n13454), .A2(n13606), .ZN(n13605) );
  OR2_X1 U13504 ( .A1(n13453), .A2(n13451), .ZN(n13606) );
  NOR2_X1 U13505 ( .A1(n8954), .A2(n8213), .ZN(n13454) );
  NAND2_X1 U13506 ( .A1(n13451), .A2(n13453), .ZN(n13604) );
  NAND2_X1 U13507 ( .A1(n13607), .A2(n13608), .ZN(n13453) );
  NAND2_X1 U13508 ( .A1(n13609), .A2(b_13_), .ZN(n13608) );
  NOR2_X1 U13509 ( .A1(n13610), .A2(n8939), .ZN(n13609) );
  NOR2_X1 U13510 ( .A1(n13448), .A2(n13449), .ZN(n13610) );
  NAND2_X1 U13511 ( .A1(n13448), .A2(n13449), .ZN(n13607) );
  NAND2_X1 U13512 ( .A1(n13611), .A2(n13612), .ZN(n13449) );
  NAND2_X1 U13513 ( .A1(n13446), .A2(n13613), .ZN(n13612) );
  OR2_X1 U13514 ( .A1(n13445), .A2(n13443), .ZN(n13613) );
  NOR2_X1 U13515 ( .A1(n8954), .A2(n8158), .ZN(n13446) );
  NAND2_X1 U13516 ( .A1(n13443), .A2(n13445), .ZN(n13611) );
  NAND2_X1 U13517 ( .A1(n13441), .A2(n13614), .ZN(n13445) );
  NAND2_X1 U13518 ( .A1(n13440), .A2(n13442), .ZN(n13614) );
  NAND2_X1 U13519 ( .A1(n13615), .A2(n13616), .ZN(n13442) );
  NAND2_X1 U13520 ( .A1(b_13_), .A2(a_26_), .ZN(n13616) );
  INV_X1 U13521 ( .A(n13617), .ZN(n13615) );
  XNOR2_X1 U13522 ( .A(n13618), .B(n13619), .ZN(n13440) );
  NAND2_X1 U13523 ( .A1(n13620), .A2(n13621), .ZN(n13618) );
  NAND2_X1 U13524 ( .A1(a_26_), .A2(n13617), .ZN(n13441) );
  NAND2_X1 U13525 ( .A1(n13411), .A2(n13622), .ZN(n13617) );
  NAND2_X1 U13526 ( .A1(n13410), .A2(n13412), .ZN(n13622) );
  NAND2_X1 U13527 ( .A1(n13623), .A2(n13624), .ZN(n13412) );
  NAND2_X1 U13528 ( .A1(b_13_), .A2(a_27_), .ZN(n13624) );
  INV_X1 U13529 ( .A(n13625), .ZN(n13623) );
  XOR2_X1 U13530 ( .A(n13626), .B(n13627), .Z(n13410) );
  XNOR2_X1 U13531 ( .A(n13628), .B(n13629), .ZN(n13626) );
  NAND2_X1 U13532 ( .A1(b_12_), .A2(a_28_), .ZN(n13628) );
  NAND2_X1 U13533 ( .A1(a_27_), .A2(n13625), .ZN(n13411) );
  NAND2_X1 U13534 ( .A1(n13630), .A2(n13631), .ZN(n13625) );
  NAND2_X1 U13535 ( .A1(n13632), .A2(b_13_), .ZN(n13631) );
  NOR2_X1 U13536 ( .A1(n13633), .A2(n8055), .ZN(n13632) );
  NOR2_X1 U13537 ( .A1(n13418), .A2(n13420), .ZN(n13633) );
  NAND2_X1 U13538 ( .A1(n13418), .A2(n13420), .ZN(n13630) );
  NAND2_X1 U13539 ( .A1(n13634), .A2(n13635), .ZN(n13420) );
  NAND2_X1 U13540 ( .A1(n13436), .A2(n13636), .ZN(n13635) );
  OR2_X1 U13541 ( .A1(n13437), .A2(n13438), .ZN(n13636) );
  NOR2_X1 U13542 ( .A1(n8954), .A2(n8041), .ZN(n13436) );
  NAND2_X1 U13543 ( .A1(n13438), .A2(n13437), .ZN(n13634) );
  NAND2_X1 U13544 ( .A1(n13637), .A2(n13638), .ZN(n13437) );
  NAND2_X1 U13545 ( .A1(b_11_), .A2(n13639), .ZN(n13638) );
  NAND2_X1 U13546 ( .A1(n8003), .A2(n13640), .ZN(n13639) );
  NAND2_X1 U13547 ( .A1(a_31_), .A2(n8955), .ZN(n13640) );
  NAND2_X1 U13548 ( .A1(b_12_), .A2(n13641), .ZN(n13637) );
  NAND2_X1 U13549 ( .A1(n9341), .A2(n13642), .ZN(n13641) );
  NAND2_X1 U13550 ( .A1(a_30_), .A2(n8957), .ZN(n13642) );
  AND2_X1 U13551 ( .A1(n13643), .A2(n7953), .ZN(n13438) );
  NOR2_X1 U13552 ( .A1(n8954), .A2(n8955), .ZN(n13643) );
  XOR2_X1 U13553 ( .A(n13644), .B(n13645), .Z(n13418) );
  XOR2_X1 U13554 ( .A(n13646), .B(n13647), .Z(n13644) );
  XNOR2_X1 U13555 ( .A(n13648), .B(n13649), .ZN(n13443) );
  NAND2_X1 U13556 ( .A1(n13650), .A2(n13651), .ZN(n13648) );
  XNOR2_X1 U13557 ( .A(n13652), .B(n13653), .ZN(n13448) );
  XNOR2_X1 U13558 ( .A(n13654), .B(n13655), .ZN(n13653) );
  XOR2_X1 U13559 ( .A(n13656), .B(n13657), .Z(n13451) );
  XOR2_X1 U13560 ( .A(n13658), .B(n13659), .Z(n13656) );
  NOR2_X1 U13561 ( .A1(n8939), .A2(n8955), .ZN(n13659) );
  XNOR2_X1 U13562 ( .A(n13660), .B(n13661), .ZN(n13456) );
  XNOR2_X1 U13563 ( .A(n13662), .B(n13663), .ZN(n13661) );
  XOR2_X1 U13564 ( .A(n13664), .B(n13665), .Z(n13459) );
  XOR2_X1 U13565 ( .A(n13666), .B(n13667), .Z(n13664) );
  NOR2_X1 U13566 ( .A1(n8941), .A2(n8955), .ZN(n13667) );
  XNOR2_X1 U13567 ( .A(n13668), .B(n13669), .ZN(n13464) );
  XNOR2_X1 U13568 ( .A(n13670), .B(n13671), .ZN(n13669) );
  XOR2_X1 U13569 ( .A(n13672), .B(n13673), .Z(n13467) );
  XOR2_X1 U13570 ( .A(n13674), .B(n13675), .Z(n13672) );
  NOR2_X1 U13571 ( .A1(n8944), .A2(n8955), .ZN(n13675) );
  XOR2_X1 U13572 ( .A(n13676), .B(n13677), .Z(n13472) );
  XOR2_X1 U13573 ( .A(n13678), .B(n13679), .Z(n13676) );
  NOR2_X1 U13574 ( .A1(n8324), .A2(n8955), .ZN(n13679) );
  XNOR2_X1 U13575 ( .A(n13680), .B(n13681), .ZN(n13476) );
  XNOR2_X1 U13576 ( .A(n13682), .B(n13683), .ZN(n13680) );
  XOR2_X1 U13577 ( .A(n13684), .B(n13685), .Z(n13480) );
  XOR2_X1 U13578 ( .A(n13686), .B(n13687), .Z(n13684) );
  XNOR2_X1 U13579 ( .A(n13688), .B(n13689), .ZN(n13484) );
  XNOR2_X1 U13580 ( .A(n13690), .B(n13691), .ZN(n13688) );
  XNOR2_X1 U13581 ( .A(n13692), .B(n13693), .ZN(n13488) );
  XOR2_X1 U13582 ( .A(n13694), .B(n13695), .Z(n13693) );
  NAND2_X1 U13583 ( .A1(b_12_), .A2(a_15_), .ZN(n13695) );
  INV_X1 U13584 ( .A(n8889), .ZN(n13358) );
  NAND2_X1 U13585 ( .A1(b_13_), .A2(a_13_), .ZN(n8889) );
  XNOR2_X1 U13586 ( .A(n13696), .B(n13697), .ZN(n13348) );
  NAND2_X1 U13587 ( .A1(n13698), .A2(n13699), .ZN(n13696) );
  XOR2_X1 U13588 ( .A(n13700), .B(n13701), .Z(n13340) );
  XOR2_X1 U13589 ( .A(n13702), .B(n13703), .Z(n13700) );
  XNOR2_X1 U13590 ( .A(n13704), .B(n13705), .ZN(n13492) );
  NAND2_X1 U13591 ( .A1(n13706), .A2(n13707), .ZN(n13704) );
  XNOR2_X1 U13592 ( .A(n13708), .B(n13709), .ZN(n13496) );
  XNOR2_X1 U13593 ( .A(n13710), .B(n13711), .ZN(n13708) );
  XNOR2_X1 U13594 ( .A(n13712), .B(n13713), .ZN(n13325) );
  XOR2_X1 U13595 ( .A(n13714), .B(n13715), .Z(n13713) );
  NAND2_X1 U13596 ( .A1(b_12_), .A2(a_9_), .ZN(n13715) );
  XNOR2_X1 U13597 ( .A(n13716), .B(n13717), .ZN(n13317) );
  NAND2_X1 U13598 ( .A1(n13718), .A2(n13719), .ZN(n13716) );
  XNOR2_X1 U13599 ( .A(n13720), .B(n13721), .ZN(n13499) );
  NAND2_X1 U13600 ( .A1(n13722), .A2(n13723), .ZN(n13720) );
  XNOR2_X1 U13601 ( .A(n13724), .B(n13725), .ZN(n13503) );
  NAND2_X1 U13602 ( .A1(n13726), .A2(n13727), .ZN(n13724) );
  XNOR2_X1 U13603 ( .A(n13728), .B(n13729), .ZN(n13301) );
  NAND2_X1 U13604 ( .A1(n13730), .A2(n13731), .ZN(n13728) );
  XNOR2_X1 U13605 ( .A(n13732), .B(n13733), .ZN(n13294) );
  NAND2_X1 U13606 ( .A1(n13734), .A2(n13735), .ZN(n13732) );
  XNOR2_X1 U13607 ( .A(n13736), .B(n13737), .ZN(n13286) );
  NAND2_X1 U13608 ( .A1(n13738), .A2(n13739), .ZN(n13736) );
  XNOR2_X1 U13609 ( .A(n13740), .B(n13741), .ZN(n13278) );
  XNOR2_X1 U13610 ( .A(n13742), .B(n13743), .ZN(n13740) );
  XNOR2_X1 U13611 ( .A(n13744), .B(n13745), .ZN(n13507) );
  XNOR2_X1 U13612 ( .A(n13746), .B(n13747), .ZN(n13744) );
  XOR2_X1 U13613 ( .A(n13748), .B(n13272), .Z(n13512) );
  XNOR2_X1 U13614 ( .A(n13749), .B(n13750), .ZN(n13272) );
  NOR2_X1 U13615 ( .A1(n8974), .A2(n8955), .ZN(n13750) );
  INV_X1 U13616 ( .A(n13271), .ZN(n13748) );
  NAND2_X1 U13617 ( .A1(n9138), .A2(n13751), .ZN(n13511) );
  OR2_X1 U13618 ( .A1(n9143), .A2(n9142), .ZN(n13751) );
  OR2_X1 U13619 ( .A1(n9138), .A2(n9137), .ZN(n9109) );
  NAND2_X1 U13620 ( .A1(n9135), .A2(n13752), .ZN(n9137) );
  NAND2_X1 U13621 ( .A1(n13753), .A2(n13754), .ZN(n13752) );
  INV_X1 U13622 ( .A(n13755), .ZN(n13754) );
  XOR2_X1 U13623 ( .A(n13756), .B(n13757), .Z(n13753) );
  NAND2_X1 U13624 ( .A1(n9143), .A2(n9142), .ZN(n9138) );
  NAND2_X1 U13625 ( .A1(n13758), .A2(n13759), .ZN(n9142) );
  NAND2_X1 U13626 ( .A1(n13760), .A2(b_12_), .ZN(n13759) );
  NOR2_X1 U13627 ( .A1(n13761), .A2(n8974), .ZN(n13760) );
  NOR2_X1 U13628 ( .A1(n13271), .A2(n13749), .ZN(n13761) );
  NAND2_X1 U13629 ( .A1(n13271), .A2(n13749), .ZN(n13758) );
  NAND2_X1 U13630 ( .A1(n13762), .A2(n13763), .ZN(n13749) );
  NAND2_X1 U13631 ( .A1(n13747), .A2(n13764), .ZN(n13763) );
  NAND2_X1 U13632 ( .A1(n13746), .A2(n13745), .ZN(n13764) );
  NOR2_X1 U13633 ( .A1(n8955), .A2(n8969), .ZN(n13747) );
  OR2_X1 U13634 ( .A1(n13745), .A2(n13746), .ZN(n13762) );
  AND2_X1 U13635 ( .A1(n13765), .A2(n13766), .ZN(n13746) );
  NAND2_X1 U13636 ( .A1(n13743), .A2(n13767), .ZN(n13766) );
  NAND2_X1 U13637 ( .A1(n13742), .A2(n13741), .ZN(n13767) );
  NOR2_X1 U13638 ( .A1(n8955), .A2(n8792), .ZN(n13743) );
  OR2_X1 U13639 ( .A1(n13741), .A2(n13742), .ZN(n13765) );
  AND2_X1 U13640 ( .A1(n13738), .A2(n13768), .ZN(n13742) );
  NAND2_X1 U13641 ( .A1(n13737), .A2(n13739), .ZN(n13768) );
  NAND2_X1 U13642 ( .A1(n13769), .A2(n13770), .ZN(n13739) );
  NAND2_X1 U13643 ( .A1(b_12_), .A2(a_3_), .ZN(n13770) );
  INV_X1 U13644 ( .A(n13771), .ZN(n13769) );
  XOR2_X1 U13645 ( .A(n13772), .B(n13773), .Z(n13737) );
  XOR2_X1 U13646 ( .A(n13774), .B(n13775), .Z(n13772) );
  NOR2_X1 U13647 ( .A1(n8966), .A2(n8957), .ZN(n13775) );
  NAND2_X1 U13648 ( .A1(a_3_), .A2(n13771), .ZN(n13738) );
  NAND2_X1 U13649 ( .A1(n13734), .A2(n13776), .ZN(n13771) );
  NAND2_X1 U13650 ( .A1(n13733), .A2(n13735), .ZN(n13776) );
  NAND2_X1 U13651 ( .A1(n13777), .A2(n13778), .ZN(n13735) );
  NAND2_X1 U13652 ( .A1(b_12_), .A2(a_4_), .ZN(n13778) );
  INV_X1 U13653 ( .A(n13779), .ZN(n13777) );
  XOR2_X1 U13654 ( .A(n13780), .B(n13781), .Z(n13733) );
  XOR2_X1 U13655 ( .A(n13782), .B(n13783), .Z(n13780) );
  NOR2_X1 U13656 ( .A1(n8723), .A2(n8957), .ZN(n13783) );
  NAND2_X1 U13657 ( .A1(a_4_), .A2(n13779), .ZN(n13734) );
  NAND2_X1 U13658 ( .A1(n13730), .A2(n13784), .ZN(n13779) );
  NAND2_X1 U13659 ( .A1(n13729), .A2(n13731), .ZN(n13784) );
  NAND2_X1 U13660 ( .A1(n13785), .A2(n13786), .ZN(n13731) );
  NAND2_X1 U13661 ( .A1(b_12_), .A2(a_5_), .ZN(n13786) );
  INV_X1 U13662 ( .A(n13787), .ZN(n13785) );
  XOR2_X1 U13663 ( .A(n13788), .B(n13789), .Z(n13729) );
  XOR2_X1 U13664 ( .A(n13790), .B(n13791), .Z(n13788) );
  NOR2_X1 U13665 ( .A1(n8681), .A2(n8957), .ZN(n13791) );
  NAND2_X1 U13666 ( .A1(a_5_), .A2(n13787), .ZN(n13730) );
  NAND2_X1 U13667 ( .A1(n13726), .A2(n13792), .ZN(n13787) );
  NAND2_X1 U13668 ( .A1(n13725), .A2(n13727), .ZN(n13792) );
  NAND2_X1 U13669 ( .A1(n13793), .A2(n13794), .ZN(n13727) );
  NAND2_X1 U13670 ( .A1(b_12_), .A2(a_6_), .ZN(n13794) );
  INV_X1 U13671 ( .A(n13795), .ZN(n13793) );
  XOR2_X1 U13672 ( .A(n13796), .B(n13797), .Z(n13725) );
  XOR2_X1 U13673 ( .A(n13798), .B(n13799), .Z(n13796) );
  NOR2_X1 U13674 ( .A1(n8962), .A2(n8957), .ZN(n13799) );
  NAND2_X1 U13675 ( .A1(a_6_), .A2(n13795), .ZN(n13726) );
  NAND2_X1 U13676 ( .A1(n13722), .A2(n13800), .ZN(n13795) );
  NAND2_X1 U13677 ( .A1(n13721), .A2(n13723), .ZN(n13800) );
  NAND2_X1 U13678 ( .A1(n13801), .A2(n13802), .ZN(n13723) );
  NAND2_X1 U13679 ( .A1(b_12_), .A2(a_7_), .ZN(n13802) );
  INV_X1 U13680 ( .A(n13803), .ZN(n13801) );
  XNOR2_X1 U13681 ( .A(n13804), .B(n13805), .ZN(n13721) );
  XOR2_X1 U13682 ( .A(n13806), .B(n13807), .Z(n13805) );
  NAND2_X1 U13683 ( .A1(b_11_), .A2(a_8_), .ZN(n13807) );
  NAND2_X1 U13684 ( .A1(a_7_), .A2(n13803), .ZN(n13722) );
  NAND2_X1 U13685 ( .A1(n13718), .A2(n13808), .ZN(n13803) );
  NAND2_X1 U13686 ( .A1(n13717), .A2(n13719), .ZN(n13808) );
  NAND2_X1 U13687 ( .A1(n13809), .A2(n13810), .ZN(n13719) );
  NAND2_X1 U13688 ( .A1(b_12_), .A2(a_8_), .ZN(n13810) );
  INV_X1 U13689 ( .A(n13811), .ZN(n13809) );
  XOR2_X1 U13690 ( .A(n13812), .B(n13813), .Z(n13717) );
  XOR2_X1 U13691 ( .A(n13814), .B(n13815), .Z(n13812) );
  NOR2_X1 U13692 ( .A1(n8605), .A2(n8957), .ZN(n13815) );
  NAND2_X1 U13693 ( .A1(a_8_), .A2(n13811), .ZN(n13718) );
  NAND2_X1 U13694 ( .A1(n13816), .A2(n13817), .ZN(n13811) );
  NAND2_X1 U13695 ( .A1(n13818), .A2(b_12_), .ZN(n13817) );
  NOR2_X1 U13696 ( .A1(n13819), .A2(n8605), .ZN(n13818) );
  NOR2_X1 U13697 ( .A1(n13712), .A2(n13714), .ZN(n13819) );
  NAND2_X1 U13698 ( .A1(n13712), .A2(n13714), .ZN(n13816) );
  NAND2_X1 U13699 ( .A1(n13820), .A2(n13821), .ZN(n13714) );
  NAND2_X1 U13700 ( .A1(n13711), .A2(n13822), .ZN(n13821) );
  NAND2_X1 U13701 ( .A1(n13710), .A2(n13709), .ZN(n13822) );
  NOR2_X1 U13702 ( .A1(n8955), .A2(n8959), .ZN(n13711) );
  OR2_X1 U13703 ( .A1(n13709), .A2(n13710), .ZN(n13820) );
  AND2_X1 U13704 ( .A1(n13706), .A2(n13823), .ZN(n13710) );
  NAND2_X1 U13705 ( .A1(n13705), .A2(n13707), .ZN(n13823) );
  NAND2_X1 U13706 ( .A1(n13824), .A2(n13825), .ZN(n13707) );
  NAND2_X1 U13707 ( .A1(b_12_), .A2(a_11_), .ZN(n13825) );
  INV_X1 U13708 ( .A(n13826), .ZN(n13824) );
  XOR2_X1 U13709 ( .A(n13827), .B(n13828), .Z(n13705) );
  XOR2_X1 U13710 ( .A(n13829), .B(n13830), .Z(n13827) );
  NOR2_X1 U13711 ( .A1(n8956), .A2(n8957), .ZN(n13830) );
  NAND2_X1 U13712 ( .A1(a_11_), .A2(n13826), .ZN(n13706) );
  NAND2_X1 U13713 ( .A1(n13831), .A2(n13832), .ZN(n13826) );
  NAND2_X1 U13714 ( .A1(n13701), .A2(n13833), .ZN(n13832) );
  OR2_X1 U13715 ( .A1(n13702), .A2(n13703), .ZN(n13833) );
  XOR2_X1 U13716 ( .A(n13834), .B(n13835), .Z(n13701) );
  XOR2_X1 U13717 ( .A(n13836), .B(n13837), .Z(n13834) );
  NOR2_X1 U13718 ( .A1(n8495), .A2(n8957), .ZN(n13837) );
  NAND2_X1 U13719 ( .A1(n13703), .A2(n13702), .ZN(n13831) );
  NAND2_X1 U13720 ( .A1(n13698), .A2(n13838), .ZN(n13702) );
  NAND2_X1 U13721 ( .A1(n13697), .A2(n13699), .ZN(n13838) );
  NAND2_X1 U13722 ( .A1(n13839), .A2(n13840), .ZN(n13699) );
  NAND2_X1 U13723 ( .A1(b_12_), .A2(a_13_), .ZN(n13840) );
  INV_X1 U13724 ( .A(n13841), .ZN(n13839) );
  XNOR2_X1 U13725 ( .A(n13842), .B(n13843), .ZN(n13697) );
  XOR2_X1 U13726 ( .A(n13844), .B(n13845), .Z(n13843) );
  NAND2_X1 U13727 ( .A1(b_11_), .A2(a_14_), .ZN(n13845) );
  NAND2_X1 U13728 ( .A1(a_13_), .A2(n13841), .ZN(n13698) );
  NAND2_X1 U13729 ( .A1(n13569), .A2(n13846), .ZN(n13841) );
  NAND2_X1 U13730 ( .A1(n13568), .A2(n13570), .ZN(n13846) );
  NAND2_X1 U13731 ( .A1(n13847), .A2(n13848), .ZN(n13570) );
  NAND2_X1 U13732 ( .A1(b_12_), .A2(a_14_), .ZN(n13848) );
  INV_X1 U13733 ( .A(n13849), .ZN(n13847) );
  XOR2_X1 U13734 ( .A(n13850), .B(n13851), .Z(n13568) );
  XOR2_X1 U13735 ( .A(n13852), .B(n13853), .Z(n13850) );
  NOR2_X1 U13736 ( .A1(n8440), .A2(n8957), .ZN(n13853) );
  NAND2_X1 U13737 ( .A1(a_14_), .A2(n13849), .ZN(n13569) );
  NAND2_X1 U13738 ( .A1(n13854), .A2(n13855), .ZN(n13849) );
  NAND2_X1 U13739 ( .A1(n13856), .A2(b_12_), .ZN(n13855) );
  NOR2_X1 U13740 ( .A1(n13857), .A2(n8440), .ZN(n13856) );
  NOR2_X1 U13741 ( .A1(n13692), .A2(n13694), .ZN(n13857) );
  NAND2_X1 U13742 ( .A1(n13692), .A2(n13694), .ZN(n13854) );
  NAND2_X1 U13743 ( .A1(n13858), .A2(n13859), .ZN(n13694) );
  NAND2_X1 U13744 ( .A1(n13691), .A2(n13860), .ZN(n13859) );
  NAND2_X1 U13745 ( .A1(n13690), .A2(n13689), .ZN(n13860) );
  NOR2_X1 U13746 ( .A1(n8955), .A2(n8950), .ZN(n13691) );
  OR2_X1 U13747 ( .A1(n13689), .A2(n13690), .ZN(n13858) );
  AND2_X1 U13748 ( .A1(n13861), .A2(n13862), .ZN(n13690) );
  NAND2_X1 U13749 ( .A1(n13687), .A2(n13863), .ZN(n13862) );
  OR2_X1 U13750 ( .A1(n13686), .A2(n13685), .ZN(n13863) );
  NOR2_X1 U13751 ( .A1(n8955), .A2(n8385), .ZN(n13687) );
  NAND2_X1 U13752 ( .A1(n13685), .A2(n13686), .ZN(n13861) );
  NAND2_X1 U13753 ( .A1(n13864), .A2(n13865), .ZN(n13686) );
  NAND2_X1 U13754 ( .A1(n13683), .A2(n13866), .ZN(n13865) );
  NAND2_X1 U13755 ( .A1(n13682), .A2(n13681), .ZN(n13866) );
  NOR2_X1 U13756 ( .A1(n8955), .A2(n8947), .ZN(n13683) );
  OR2_X1 U13757 ( .A1(n13681), .A2(n13682), .ZN(n13864) );
  AND2_X1 U13758 ( .A1(n13867), .A2(n13868), .ZN(n13682) );
  NAND2_X1 U13759 ( .A1(n13869), .A2(b_12_), .ZN(n13868) );
  NOR2_X1 U13760 ( .A1(n13870), .A2(n8324), .ZN(n13869) );
  NOR2_X1 U13761 ( .A1(n13677), .A2(n13678), .ZN(n13870) );
  NAND2_X1 U13762 ( .A1(n13677), .A2(n13678), .ZN(n13867) );
  NAND2_X1 U13763 ( .A1(n13871), .A2(n13872), .ZN(n13678) );
  NAND2_X1 U13764 ( .A1(n13873), .A2(b_12_), .ZN(n13872) );
  NOR2_X1 U13765 ( .A1(n13874), .A2(n8944), .ZN(n13873) );
  NOR2_X1 U13766 ( .A1(n13673), .A2(n13674), .ZN(n13874) );
  NAND2_X1 U13767 ( .A1(n13673), .A2(n13674), .ZN(n13871) );
  NAND2_X1 U13768 ( .A1(n13875), .A2(n13876), .ZN(n13674) );
  NAND2_X1 U13769 ( .A1(n13671), .A2(n13877), .ZN(n13876) );
  OR2_X1 U13770 ( .A1(n13670), .A2(n13668), .ZN(n13877) );
  NOR2_X1 U13771 ( .A1(n8955), .A2(n8268), .ZN(n13671) );
  NAND2_X1 U13772 ( .A1(n13668), .A2(n13670), .ZN(n13875) );
  NAND2_X1 U13773 ( .A1(n13878), .A2(n13879), .ZN(n13670) );
  NAND2_X1 U13774 ( .A1(n13880), .A2(b_12_), .ZN(n13879) );
  NOR2_X1 U13775 ( .A1(n13881), .A2(n8941), .ZN(n13880) );
  NOR2_X1 U13776 ( .A1(n13665), .A2(n13666), .ZN(n13881) );
  NAND2_X1 U13777 ( .A1(n13665), .A2(n13666), .ZN(n13878) );
  NAND2_X1 U13778 ( .A1(n13882), .A2(n13883), .ZN(n13666) );
  NAND2_X1 U13779 ( .A1(n13663), .A2(n13884), .ZN(n13883) );
  OR2_X1 U13780 ( .A1(n13662), .A2(n13660), .ZN(n13884) );
  NOR2_X1 U13781 ( .A1(n8955), .A2(n8213), .ZN(n13663) );
  NAND2_X1 U13782 ( .A1(n13660), .A2(n13662), .ZN(n13882) );
  NAND2_X1 U13783 ( .A1(n13885), .A2(n13886), .ZN(n13662) );
  NAND2_X1 U13784 ( .A1(n13887), .A2(b_12_), .ZN(n13886) );
  NOR2_X1 U13785 ( .A1(n13888), .A2(n8939), .ZN(n13887) );
  NOR2_X1 U13786 ( .A1(n13657), .A2(n13658), .ZN(n13888) );
  NAND2_X1 U13787 ( .A1(n13657), .A2(n13658), .ZN(n13885) );
  NAND2_X1 U13788 ( .A1(n13889), .A2(n13890), .ZN(n13658) );
  NAND2_X1 U13789 ( .A1(n13655), .A2(n13891), .ZN(n13890) );
  OR2_X1 U13790 ( .A1(n13654), .A2(n13652), .ZN(n13891) );
  NOR2_X1 U13791 ( .A1(n8955), .A2(n8158), .ZN(n13655) );
  NAND2_X1 U13792 ( .A1(n13652), .A2(n13654), .ZN(n13889) );
  NAND2_X1 U13793 ( .A1(n13650), .A2(n13892), .ZN(n13654) );
  NAND2_X1 U13794 ( .A1(n13649), .A2(n13651), .ZN(n13892) );
  NAND2_X1 U13795 ( .A1(n13893), .A2(n13894), .ZN(n13651) );
  NAND2_X1 U13796 ( .A1(b_12_), .A2(a_26_), .ZN(n13894) );
  INV_X1 U13797 ( .A(n13895), .ZN(n13893) );
  XNOR2_X1 U13798 ( .A(n13896), .B(n13897), .ZN(n13649) );
  NAND2_X1 U13799 ( .A1(n13898), .A2(n13899), .ZN(n13896) );
  NAND2_X1 U13800 ( .A1(a_26_), .A2(n13895), .ZN(n13650) );
  NAND2_X1 U13801 ( .A1(n13620), .A2(n13900), .ZN(n13895) );
  NAND2_X1 U13802 ( .A1(n13619), .A2(n13621), .ZN(n13900) );
  NAND2_X1 U13803 ( .A1(n13901), .A2(n13902), .ZN(n13621) );
  NAND2_X1 U13804 ( .A1(b_12_), .A2(a_27_), .ZN(n13902) );
  INV_X1 U13805 ( .A(n13903), .ZN(n13901) );
  XOR2_X1 U13806 ( .A(n13904), .B(n13905), .Z(n13619) );
  XNOR2_X1 U13807 ( .A(n13906), .B(n13907), .ZN(n13904) );
  NAND2_X1 U13808 ( .A1(b_11_), .A2(a_28_), .ZN(n13906) );
  NAND2_X1 U13809 ( .A1(a_27_), .A2(n13903), .ZN(n13620) );
  NAND2_X1 U13810 ( .A1(n13908), .A2(n13909), .ZN(n13903) );
  NAND2_X1 U13811 ( .A1(n13910), .A2(b_12_), .ZN(n13909) );
  NOR2_X1 U13812 ( .A1(n13911), .A2(n8055), .ZN(n13910) );
  NOR2_X1 U13813 ( .A1(n13627), .A2(n13629), .ZN(n13911) );
  NAND2_X1 U13814 ( .A1(n13627), .A2(n13629), .ZN(n13908) );
  NAND2_X1 U13815 ( .A1(n13912), .A2(n13913), .ZN(n13629) );
  NAND2_X1 U13816 ( .A1(n13645), .A2(n13914), .ZN(n13913) );
  OR2_X1 U13817 ( .A1(n13646), .A2(n13647), .ZN(n13914) );
  NOR2_X1 U13818 ( .A1(n8955), .A2(n8041), .ZN(n13645) );
  NAND2_X1 U13819 ( .A1(n13647), .A2(n13646), .ZN(n13912) );
  NAND2_X1 U13820 ( .A1(n13915), .A2(n13916), .ZN(n13646) );
  NAND2_X1 U13821 ( .A1(b_10_), .A2(n13917), .ZN(n13916) );
  NAND2_X1 U13822 ( .A1(n8003), .A2(n13918), .ZN(n13917) );
  NAND2_X1 U13823 ( .A1(a_31_), .A2(n8957), .ZN(n13918) );
  NAND2_X1 U13824 ( .A1(b_11_), .A2(n13919), .ZN(n13915) );
  NAND2_X1 U13825 ( .A1(n9341), .A2(n13920), .ZN(n13919) );
  NAND2_X1 U13826 ( .A1(a_30_), .A2(n8958), .ZN(n13920) );
  AND2_X1 U13827 ( .A1(n13921), .A2(n7953), .ZN(n13647) );
  NOR2_X1 U13828 ( .A1(n8955), .A2(n8957), .ZN(n13921) );
  XOR2_X1 U13829 ( .A(n13922), .B(n13923), .Z(n13627) );
  XOR2_X1 U13830 ( .A(n13924), .B(n13925), .Z(n13922) );
  XNOR2_X1 U13831 ( .A(n13926), .B(n13927), .ZN(n13652) );
  NAND2_X1 U13832 ( .A1(n13928), .A2(n13929), .ZN(n13926) );
  XNOR2_X1 U13833 ( .A(n13930), .B(n13931), .ZN(n13657) );
  XNOR2_X1 U13834 ( .A(n13932), .B(n13933), .ZN(n13931) );
  XOR2_X1 U13835 ( .A(n13934), .B(n13935), .Z(n13660) );
  XOR2_X1 U13836 ( .A(n13936), .B(n13937), .Z(n13934) );
  NOR2_X1 U13837 ( .A1(n8939), .A2(n8957), .ZN(n13937) );
  XNOR2_X1 U13838 ( .A(n13938), .B(n13939), .ZN(n13665) );
  XNOR2_X1 U13839 ( .A(n13940), .B(n13941), .ZN(n13939) );
  XOR2_X1 U13840 ( .A(n13942), .B(n13943), .Z(n13668) );
  XOR2_X1 U13841 ( .A(n13944), .B(n13945), .Z(n13942) );
  NOR2_X1 U13842 ( .A1(n8941), .A2(n8957), .ZN(n13945) );
  XNOR2_X1 U13843 ( .A(n13946), .B(n13947), .ZN(n13673) );
  XNOR2_X1 U13844 ( .A(n13948), .B(n13949), .ZN(n13947) );
  XOR2_X1 U13845 ( .A(n13950), .B(n13951), .Z(n13677) );
  XOR2_X1 U13846 ( .A(n13952), .B(n13953), .Z(n13950) );
  XNOR2_X1 U13847 ( .A(n13954), .B(n13955), .ZN(n13681) );
  XOR2_X1 U13848 ( .A(n13956), .B(n13957), .Z(n13954) );
  NOR2_X1 U13849 ( .A1(n8324), .A2(n8957), .ZN(n13957) );
  XNOR2_X1 U13850 ( .A(n13958), .B(n13959), .ZN(n13685) );
  NAND2_X1 U13851 ( .A1(n13960), .A2(n13961), .ZN(n13958) );
  XNOR2_X1 U13852 ( .A(n13962), .B(n13963), .ZN(n13689) );
  XOR2_X1 U13853 ( .A(n13964), .B(n13965), .Z(n13962) );
  NOR2_X1 U13854 ( .A1(n8385), .A2(n8957), .ZN(n13965) );
  XNOR2_X1 U13855 ( .A(n13966), .B(n13967), .ZN(n13692) );
  XOR2_X1 U13856 ( .A(n13968), .B(n13969), .Z(n13967) );
  NAND2_X1 U13857 ( .A1(b_11_), .A2(a_16_), .ZN(n13969) );
  INV_X1 U13858 ( .A(n8528), .ZN(n13703) );
  NAND2_X1 U13859 ( .A1(b_12_), .A2(a_12_), .ZN(n8528) );
  XNOR2_X1 U13860 ( .A(n13970), .B(n13971), .ZN(n13709) );
  XOR2_X1 U13861 ( .A(n13972), .B(n13973), .Z(n13970) );
  XOR2_X1 U13862 ( .A(n13974), .B(n13975), .Z(n13712) );
  XNOR2_X1 U13863 ( .A(n13976), .B(n13977), .ZN(n13974) );
  NAND2_X1 U13864 ( .A1(b_11_), .A2(a_10_), .ZN(n13976) );
  XOR2_X1 U13865 ( .A(n13978), .B(n13979), .Z(n13741) );
  XOR2_X1 U13866 ( .A(n13980), .B(n13981), .Z(n13979) );
  NAND2_X1 U13867 ( .A1(b_11_), .A2(a_3_), .ZN(n13981) );
  XOR2_X1 U13868 ( .A(n13982), .B(n13983), .Z(n13745) );
  XOR2_X1 U13869 ( .A(n13984), .B(n13985), .Z(n13983) );
  NAND2_X1 U13870 ( .A1(b_11_), .A2(a_2_), .ZN(n13985) );
  XNOR2_X1 U13871 ( .A(n13986), .B(n13987), .ZN(n13271) );
  XOR2_X1 U13872 ( .A(n13988), .B(n13989), .Z(n13987) );
  NAND2_X1 U13873 ( .A1(b_11_), .A2(a_1_), .ZN(n13989) );
  XOR2_X1 U13874 ( .A(n13990), .B(n13991), .Z(n9143) );
  XOR2_X1 U13875 ( .A(n13992), .B(n13993), .Z(n13990) );
  OR2_X1 U13876 ( .A1(n9135), .A2(n9134), .ZN(n9116) );
  XNOR2_X1 U13877 ( .A(n13994), .B(n13995), .ZN(n9134) );
  NAND2_X1 U13878 ( .A1(n13996), .A2(n13755), .ZN(n9135) );
  NAND2_X1 U13879 ( .A1(n13997), .A2(n13998), .ZN(n13755) );
  NAND2_X1 U13880 ( .A1(n13993), .A2(n13999), .ZN(n13998) );
  OR2_X1 U13881 ( .A1(n13992), .A2(n13991), .ZN(n13999) );
  NOR2_X1 U13882 ( .A1(n8957), .A2(n8974), .ZN(n13993) );
  NAND2_X1 U13883 ( .A1(n13991), .A2(n13992), .ZN(n13997) );
  NAND2_X1 U13884 ( .A1(n14000), .A2(n14001), .ZN(n13992) );
  NAND2_X1 U13885 ( .A1(n14002), .A2(b_11_), .ZN(n14001) );
  NOR2_X1 U13886 ( .A1(n14003), .A2(n8969), .ZN(n14002) );
  NOR2_X1 U13887 ( .A1(n13986), .A2(n13988), .ZN(n14003) );
  NAND2_X1 U13888 ( .A1(n13986), .A2(n13988), .ZN(n14000) );
  NAND2_X1 U13889 ( .A1(n14004), .A2(n14005), .ZN(n13988) );
  NAND2_X1 U13890 ( .A1(n14006), .A2(b_11_), .ZN(n14005) );
  NOR2_X1 U13891 ( .A1(n14007), .A2(n8792), .ZN(n14006) );
  NOR2_X1 U13892 ( .A1(n13982), .A2(n13984), .ZN(n14007) );
  NAND2_X1 U13893 ( .A1(n13982), .A2(n13984), .ZN(n14004) );
  NAND2_X1 U13894 ( .A1(n14008), .A2(n14009), .ZN(n13984) );
  NAND2_X1 U13895 ( .A1(n14010), .A2(b_11_), .ZN(n14009) );
  NOR2_X1 U13896 ( .A1(n14011), .A2(n8778), .ZN(n14010) );
  NOR2_X1 U13897 ( .A1(n13978), .A2(n13980), .ZN(n14011) );
  NAND2_X1 U13898 ( .A1(n13978), .A2(n13980), .ZN(n14008) );
  NAND2_X1 U13899 ( .A1(n14012), .A2(n14013), .ZN(n13980) );
  NAND2_X1 U13900 ( .A1(n14014), .A2(b_11_), .ZN(n14013) );
  NOR2_X1 U13901 ( .A1(n14015), .A2(n8966), .ZN(n14014) );
  NOR2_X1 U13902 ( .A1(n13773), .A2(n13774), .ZN(n14015) );
  NAND2_X1 U13903 ( .A1(n13773), .A2(n13774), .ZN(n14012) );
  NAND2_X1 U13904 ( .A1(n14016), .A2(n14017), .ZN(n13774) );
  NAND2_X1 U13905 ( .A1(n14018), .A2(b_11_), .ZN(n14017) );
  NOR2_X1 U13906 ( .A1(n14019), .A2(n8723), .ZN(n14018) );
  NOR2_X1 U13907 ( .A1(n13781), .A2(n13782), .ZN(n14019) );
  NAND2_X1 U13908 ( .A1(n13781), .A2(n13782), .ZN(n14016) );
  NAND2_X1 U13909 ( .A1(n14020), .A2(n14021), .ZN(n13782) );
  NAND2_X1 U13910 ( .A1(n14022), .A2(b_11_), .ZN(n14021) );
  NOR2_X1 U13911 ( .A1(n14023), .A2(n8681), .ZN(n14022) );
  NOR2_X1 U13912 ( .A1(n13789), .A2(n13790), .ZN(n14023) );
  NAND2_X1 U13913 ( .A1(n13789), .A2(n13790), .ZN(n14020) );
  NAND2_X1 U13914 ( .A1(n14024), .A2(n14025), .ZN(n13790) );
  NAND2_X1 U13915 ( .A1(n14026), .A2(b_11_), .ZN(n14025) );
  NOR2_X1 U13916 ( .A1(n14027), .A2(n8962), .ZN(n14026) );
  NOR2_X1 U13917 ( .A1(n13797), .A2(n13798), .ZN(n14027) );
  NAND2_X1 U13918 ( .A1(n13797), .A2(n13798), .ZN(n14024) );
  NAND2_X1 U13919 ( .A1(n14028), .A2(n14029), .ZN(n13798) );
  NAND2_X1 U13920 ( .A1(n14030), .A2(b_11_), .ZN(n14029) );
  NOR2_X1 U13921 ( .A1(n14031), .A2(n8619), .ZN(n14030) );
  NOR2_X1 U13922 ( .A1(n13804), .A2(n13806), .ZN(n14031) );
  NAND2_X1 U13923 ( .A1(n13804), .A2(n13806), .ZN(n14028) );
  NAND2_X1 U13924 ( .A1(n14032), .A2(n14033), .ZN(n13806) );
  NAND2_X1 U13925 ( .A1(n14034), .A2(b_11_), .ZN(n14033) );
  NOR2_X1 U13926 ( .A1(n14035), .A2(n8605), .ZN(n14034) );
  NOR2_X1 U13927 ( .A1(n13813), .A2(n13814), .ZN(n14035) );
  NAND2_X1 U13928 ( .A1(n13813), .A2(n13814), .ZN(n14032) );
  NAND2_X1 U13929 ( .A1(n14036), .A2(n14037), .ZN(n13814) );
  NAND2_X1 U13930 ( .A1(n14038), .A2(b_11_), .ZN(n14037) );
  NOR2_X1 U13931 ( .A1(n14039), .A2(n8959), .ZN(n14038) );
  NOR2_X1 U13932 ( .A1(n13975), .A2(n13977), .ZN(n14039) );
  NAND2_X1 U13933 ( .A1(n13975), .A2(n13977), .ZN(n14036) );
  NAND2_X1 U13934 ( .A1(n14040), .A2(n14041), .ZN(n13977) );
  NAND2_X1 U13935 ( .A1(n13971), .A2(n14042), .ZN(n14041) );
  OR2_X1 U13936 ( .A1(n13972), .A2(n13973), .ZN(n14042) );
  XNOR2_X1 U13937 ( .A(n14043), .B(n14044), .ZN(n13971) );
  NAND2_X1 U13938 ( .A1(n14045), .A2(n14046), .ZN(n14043) );
  NAND2_X1 U13939 ( .A1(n13973), .A2(n13972), .ZN(n14040) );
  NAND2_X1 U13940 ( .A1(n14047), .A2(n14048), .ZN(n13972) );
  NAND2_X1 U13941 ( .A1(n14049), .A2(b_11_), .ZN(n14048) );
  NOR2_X1 U13942 ( .A1(n14050), .A2(n8956), .ZN(n14049) );
  NOR2_X1 U13943 ( .A1(n13828), .A2(n13829), .ZN(n14050) );
  NAND2_X1 U13944 ( .A1(n13828), .A2(n13829), .ZN(n14047) );
  NAND2_X1 U13945 ( .A1(n14051), .A2(n14052), .ZN(n13829) );
  NAND2_X1 U13946 ( .A1(n14053), .A2(b_11_), .ZN(n14052) );
  NOR2_X1 U13947 ( .A1(n14054), .A2(n8495), .ZN(n14053) );
  NOR2_X1 U13948 ( .A1(n13835), .A2(n13836), .ZN(n14054) );
  NAND2_X1 U13949 ( .A1(n13835), .A2(n13836), .ZN(n14051) );
  NAND2_X1 U13950 ( .A1(n14055), .A2(n14056), .ZN(n13836) );
  NAND2_X1 U13951 ( .A1(n14057), .A2(b_11_), .ZN(n14056) );
  NOR2_X1 U13952 ( .A1(n14058), .A2(n8953), .ZN(n14057) );
  NOR2_X1 U13953 ( .A1(n13842), .A2(n13844), .ZN(n14058) );
  NAND2_X1 U13954 ( .A1(n13842), .A2(n13844), .ZN(n14055) );
  NAND2_X1 U13955 ( .A1(n14059), .A2(n14060), .ZN(n13844) );
  NAND2_X1 U13956 ( .A1(n14061), .A2(b_11_), .ZN(n14060) );
  NOR2_X1 U13957 ( .A1(n14062), .A2(n8440), .ZN(n14061) );
  NOR2_X1 U13958 ( .A1(n13851), .A2(n13852), .ZN(n14062) );
  NAND2_X1 U13959 ( .A1(n13851), .A2(n13852), .ZN(n14059) );
  NAND2_X1 U13960 ( .A1(n14063), .A2(n14064), .ZN(n13852) );
  NAND2_X1 U13961 ( .A1(n14065), .A2(b_11_), .ZN(n14064) );
  NOR2_X1 U13962 ( .A1(n14066), .A2(n8950), .ZN(n14065) );
  NOR2_X1 U13963 ( .A1(n13966), .A2(n13968), .ZN(n14066) );
  NAND2_X1 U13964 ( .A1(n13966), .A2(n13968), .ZN(n14063) );
  NAND2_X1 U13965 ( .A1(n14067), .A2(n14068), .ZN(n13968) );
  NAND2_X1 U13966 ( .A1(n14069), .A2(b_11_), .ZN(n14068) );
  NOR2_X1 U13967 ( .A1(n14070), .A2(n8385), .ZN(n14069) );
  NOR2_X1 U13968 ( .A1(n13963), .A2(n13964), .ZN(n14070) );
  NAND2_X1 U13969 ( .A1(n13963), .A2(n13964), .ZN(n14067) );
  NAND2_X1 U13970 ( .A1(n13960), .A2(n14071), .ZN(n13964) );
  NAND2_X1 U13971 ( .A1(n13959), .A2(n13961), .ZN(n14071) );
  NAND2_X1 U13972 ( .A1(n14072), .A2(n14073), .ZN(n13961) );
  NAND2_X1 U13973 ( .A1(b_11_), .A2(a_18_), .ZN(n14073) );
  INV_X1 U13974 ( .A(n14074), .ZN(n14072) );
  XNOR2_X1 U13975 ( .A(n14075), .B(n14076), .ZN(n13959) );
  XNOR2_X1 U13976 ( .A(n14077), .B(n14078), .ZN(n14075) );
  NAND2_X1 U13977 ( .A1(a_18_), .A2(n14074), .ZN(n13960) );
  NAND2_X1 U13978 ( .A1(n14079), .A2(n14080), .ZN(n14074) );
  NAND2_X1 U13979 ( .A1(n14081), .A2(b_11_), .ZN(n14080) );
  NOR2_X1 U13980 ( .A1(n14082), .A2(n8324), .ZN(n14081) );
  NOR2_X1 U13981 ( .A1(n13955), .A2(n13956), .ZN(n14082) );
  NAND2_X1 U13982 ( .A1(n13955), .A2(n13956), .ZN(n14079) );
  NAND2_X1 U13983 ( .A1(n14083), .A2(n14084), .ZN(n13956) );
  NAND2_X1 U13984 ( .A1(n13953), .A2(n14085), .ZN(n14084) );
  OR2_X1 U13985 ( .A1(n13952), .A2(n13951), .ZN(n14085) );
  NOR2_X1 U13986 ( .A1(n8957), .A2(n8944), .ZN(n13953) );
  NAND2_X1 U13987 ( .A1(n13951), .A2(n13952), .ZN(n14083) );
  NAND2_X1 U13988 ( .A1(n14086), .A2(n14087), .ZN(n13952) );
  NAND2_X1 U13989 ( .A1(n13949), .A2(n14088), .ZN(n14087) );
  OR2_X1 U13990 ( .A1(n13948), .A2(n13946), .ZN(n14088) );
  NOR2_X1 U13991 ( .A1(n8957), .A2(n8268), .ZN(n13949) );
  NAND2_X1 U13992 ( .A1(n13946), .A2(n13948), .ZN(n14086) );
  NAND2_X1 U13993 ( .A1(n14089), .A2(n14090), .ZN(n13948) );
  NAND2_X1 U13994 ( .A1(n14091), .A2(b_11_), .ZN(n14090) );
  NOR2_X1 U13995 ( .A1(n14092), .A2(n8941), .ZN(n14091) );
  NOR2_X1 U13996 ( .A1(n13943), .A2(n13944), .ZN(n14092) );
  NAND2_X1 U13997 ( .A1(n13943), .A2(n13944), .ZN(n14089) );
  NAND2_X1 U13998 ( .A1(n14093), .A2(n14094), .ZN(n13944) );
  NAND2_X1 U13999 ( .A1(n13941), .A2(n14095), .ZN(n14094) );
  OR2_X1 U14000 ( .A1(n13940), .A2(n13938), .ZN(n14095) );
  NOR2_X1 U14001 ( .A1(n8957), .A2(n8213), .ZN(n13941) );
  NAND2_X1 U14002 ( .A1(n13938), .A2(n13940), .ZN(n14093) );
  NAND2_X1 U14003 ( .A1(n14096), .A2(n14097), .ZN(n13940) );
  NAND2_X1 U14004 ( .A1(n14098), .A2(b_11_), .ZN(n14097) );
  NOR2_X1 U14005 ( .A1(n14099), .A2(n8939), .ZN(n14098) );
  NOR2_X1 U14006 ( .A1(n13935), .A2(n13936), .ZN(n14099) );
  NAND2_X1 U14007 ( .A1(n13935), .A2(n13936), .ZN(n14096) );
  NAND2_X1 U14008 ( .A1(n14100), .A2(n14101), .ZN(n13936) );
  NAND2_X1 U14009 ( .A1(n13933), .A2(n14102), .ZN(n14101) );
  OR2_X1 U14010 ( .A1(n13932), .A2(n13930), .ZN(n14102) );
  NOR2_X1 U14011 ( .A1(n8957), .A2(n8158), .ZN(n13933) );
  NAND2_X1 U14012 ( .A1(n13930), .A2(n13932), .ZN(n14100) );
  NAND2_X1 U14013 ( .A1(n13928), .A2(n14103), .ZN(n13932) );
  NAND2_X1 U14014 ( .A1(n13927), .A2(n13929), .ZN(n14103) );
  NAND2_X1 U14015 ( .A1(n14104), .A2(n14105), .ZN(n13929) );
  NAND2_X1 U14016 ( .A1(b_11_), .A2(a_26_), .ZN(n14105) );
  INV_X1 U14017 ( .A(n14106), .ZN(n14104) );
  XNOR2_X1 U14018 ( .A(n14107), .B(n14108), .ZN(n13927) );
  NAND2_X1 U14019 ( .A1(n14109), .A2(n14110), .ZN(n14107) );
  NAND2_X1 U14020 ( .A1(a_26_), .A2(n14106), .ZN(n13928) );
  NAND2_X1 U14021 ( .A1(n13898), .A2(n14111), .ZN(n14106) );
  NAND2_X1 U14022 ( .A1(n13897), .A2(n13899), .ZN(n14111) );
  NAND2_X1 U14023 ( .A1(n14112), .A2(n14113), .ZN(n13899) );
  NAND2_X1 U14024 ( .A1(b_11_), .A2(a_27_), .ZN(n14113) );
  INV_X1 U14025 ( .A(n14114), .ZN(n14112) );
  XOR2_X1 U14026 ( .A(n14115), .B(n14116), .Z(n13897) );
  XNOR2_X1 U14027 ( .A(n14117), .B(n14118), .ZN(n14115) );
  NAND2_X1 U14028 ( .A1(b_10_), .A2(a_28_), .ZN(n14117) );
  NAND2_X1 U14029 ( .A1(a_27_), .A2(n14114), .ZN(n13898) );
  NAND2_X1 U14030 ( .A1(n14119), .A2(n14120), .ZN(n14114) );
  NAND2_X1 U14031 ( .A1(n14121), .A2(b_11_), .ZN(n14120) );
  NOR2_X1 U14032 ( .A1(n14122), .A2(n8055), .ZN(n14121) );
  NOR2_X1 U14033 ( .A1(n13905), .A2(n13907), .ZN(n14122) );
  NAND2_X1 U14034 ( .A1(n13905), .A2(n13907), .ZN(n14119) );
  NAND2_X1 U14035 ( .A1(n14123), .A2(n14124), .ZN(n13907) );
  NAND2_X1 U14036 ( .A1(n13923), .A2(n14125), .ZN(n14124) );
  OR2_X1 U14037 ( .A1(n13924), .A2(n13925), .ZN(n14125) );
  NOR2_X1 U14038 ( .A1(n8957), .A2(n8041), .ZN(n13923) );
  NAND2_X1 U14039 ( .A1(n13925), .A2(n13924), .ZN(n14123) );
  NAND2_X1 U14040 ( .A1(n14126), .A2(n14127), .ZN(n13924) );
  NAND2_X1 U14041 ( .A1(b_10_), .A2(n14128), .ZN(n14127) );
  NAND2_X1 U14042 ( .A1(n9341), .A2(n14129), .ZN(n14128) );
  NAND2_X1 U14043 ( .A1(a_30_), .A2(n8960), .ZN(n14129) );
  NAND2_X1 U14044 ( .A1(b_9_), .A2(n14130), .ZN(n14126) );
  NAND2_X1 U14045 ( .A1(n8003), .A2(n14131), .ZN(n14130) );
  NAND2_X1 U14046 ( .A1(a_31_), .A2(n8958), .ZN(n14131) );
  AND2_X1 U14047 ( .A1(n14132), .A2(n7953), .ZN(n13925) );
  NOR2_X1 U14048 ( .A1(n8957), .A2(n8958), .ZN(n14132) );
  XOR2_X1 U14049 ( .A(n14133), .B(n14134), .Z(n13905) );
  XOR2_X1 U14050 ( .A(n14135), .B(n14136), .Z(n14133) );
  XNOR2_X1 U14051 ( .A(n14137), .B(n14138), .ZN(n13930) );
  NAND2_X1 U14052 ( .A1(n14139), .A2(n14140), .ZN(n14137) );
  XNOR2_X1 U14053 ( .A(n14141), .B(n14142), .ZN(n13935) );
  XNOR2_X1 U14054 ( .A(n14143), .B(n14144), .ZN(n14142) );
  XOR2_X1 U14055 ( .A(n14145), .B(n14146), .Z(n13938) );
  XOR2_X1 U14056 ( .A(n14147), .B(n14148), .Z(n14145) );
  NOR2_X1 U14057 ( .A1(n8939), .A2(n8958), .ZN(n14148) );
  XNOR2_X1 U14058 ( .A(n14149), .B(n14150), .ZN(n13943) );
  XNOR2_X1 U14059 ( .A(n14151), .B(n14152), .ZN(n14150) );
  XOR2_X1 U14060 ( .A(n14153), .B(n14154), .Z(n13946) );
  XOR2_X1 U14061 ( .A(n14155), .B(n14156), .Z(n14153) );
  NOR2_X1 U14062 ( .A1(n8941), .A2(n8958), .ZN(n14156) );
  XNOR2_X1 U14063 ( .A(n14157), .B(n14158), .ZN(n13951) );
  XOR2_X1 U14064 ( .A(n14159), .B(n14160), .Z(n14158) );
  NAND2_X1 U14065 ( .A1(b_10_), .A2(a_21_), .ZN(n14160) );
  XNOR2_X1 U14066 ( .A(n14161), .B(n14162), .ZN(n13955) );
  XNOR2_X1 U14067 ( .A(n14163), .B(n14164), .ZN(n14162) );
  XNOR2_X1 U14068 ( .A(n14165), .B(n14166), .ZN(n13963) );
  XNOR2_X1 U14069 ( .A(n14167), .B(n14168), .ZN(n14166) );
  XNOR2_X1 U14070 ( .A(n14169), .B(n14170), .ZN(n13966) );
  XOR2_X1 U14071 ( .A(n14171), .B(n14172), .Z(n14170) );
  NAND2_X1 U14072 ( .A1(b_10_), .A2(a_17_), .ZN(n14172) );
  XNOR2_X1 U14073 ( .A(n14173), .B(n14174), .ZN(n13851) );
  NAND2_X1 U14074 ( .A1(n14175), .A2(n14176), .ZN(n14173) );
  XNOR2_X1 U14075 ( .A(n14177), .B(n14178), .ZN(n13842) );
  NAND2_X1 U14076 ( .A1(n14179), .A2(n14180), .ZN(n14177) );
  XNOR2_X1 U14077 ( .A(n14181), .B(n14182), .ZN(n13835) );
  NAND2_X1 U14078 ( .A1(n14183), .A2(n14184), .ZN(n14181) );
  XNOR2_X1 U14079 ( .A(n14185), .B(n14186), .ZN(n13828) );
  NAND2_X1 U14080 ( .A1(n14187), .A2(n14188), .ZN(n14185) );
  INV_X1 U14081 ( .A(n8885), .ZN(n13973) );
  NAND2_X1 U14082 ( .A1(b_11_), .A2(a_11_), .ZN(n8885) );
  XNOR2_X1 U14083 ( .A(n14189), .B(n14190), .ZN(n13975) );
  NAND2_X1 U14084 ( .A1(n14191), .A2(n14192), .ZN(n14189) );
  XNOR2_X1 U14085 ( .A(n14193), .B(n14194), .ZN(n13813) );
  XOR2_X1 U14086 ( .A(n8583), .B(n14195), .Z(n14194) );
  XNOR2_X1 U14087 ( .A(n14196), .B(n14197), .ZN(n13804) );
  NAND2_X1 U14088 ( .A1(n14198), .A2(n14199), .ZN(n14196) );
  XNOR2_X1 U14089 ( .A(n14200), .B(n14201), .ZN(n13797) );
  NAND2_X1 U14090 ( .A1(n14202), .A2(n14203), .ZN(n14200) );
  XNOR2_X1 U14091 ( .A(n14204), .B(n14205), .ZN(n13789) );
  XNOR2_X1 U14092 ( .A(n14206), .B(n14207), .ZN(n14204) );
  XNOR2_X1 U14093 ( .A(n14208), .B(n14209), .ZN(n13781) );
  XNOR2_X1 U14094 ( .A(n14210), .B(n14211), .ZN(n14208) );
  XNOR2_X1 U14095 ( .A(n14212), .B(n14213), .ZN(n13773) );
  XNOR2_X1 U14096 ( .A(n14214), .B(n14215), .ZN(n14213) );
  XNOR2_X1 U14097 ( .A(n14216), .B(n14217), .ZN(n13978) );
  XNOR2_X1 U14098 ( .A(n14218), .B(n14219), .ZN(n14217) );
  XNOR2_X1 U14099 ( .A(n14220), .B(n14221), .ZN(n13982) );
  XNOR2_X1 U14100 ( .A(n14222), .B(n14223), .ZN(n14221) );
  XNOR2_X1 U14101 ( .A(n14224), .B(n14225), .ZN(n13986) );
  XNOR2_X1 U14102 ( .A(n14226), .B(n14227), .ZN(n14225) );
  XOR2_X1 U14103 ( .A(n14228), .B(n14229), .Z(n13991) );
  XOR2_X1 U14104 ( .A(n14230), .B(n14231), .Z(n14228) );
  NOR2_X1 U14105 ( .A1(n8969), .A2(n8958), .ZN(n14231) );
  XOR2_X1 U14106 ( .A(n14232), .B(n13757), .Z(n13996) );
  XNOR2_X1 U14107 ( .A(n14233), .B(n14234), .ZN(n13757) );
  NOR2_X1 U14108 ( .A1(n8974), .A2(n8958), .ZN(n14234) );
  INV_X1 U14109 ( .A(n13756), .ZN(n14232) );
  NAND2_X1 U14110 ( .A1(n14235), .A2(n14236), .ZN(n7963) );
  OR2_X1 U14111 ( .A1(n14236), .A2(n14235), .ZN(n7962) );
  NAND2_X1 U14112 ( .A1(n14237), .A2(n14238), .ZN(n14235) );
  NAND2_X1 U14113 ( .A1(n14239), .A2(n14240), .ZN(n14238) );
  INV_X1 U14114 ( .A(n14241), .ZN(n14240) );
  XOR2_X1 U14115 ( .A(n14242), .B(n14243), .Z(n14239) );
  NAND2_X1 U14116 ( .A1(n13995), .A2(n13994), .ZN(n14236) );
  NAND2_X1 U14117 ( .A1(n14244), .A2(n14245), .ZN(n13994) );
  NAND2_X1 U14118 ( .A1(n14246), .A2(b_10_), .ZN(n14245) );
  NOR2_X1 U14119 ( .A1(n14247), .A2(n8974), .ZN(n14246) );
  NOR2_X1 U14120 ( .A1(n13756), .A2(n14233), .ZN(n14247) );
  NAND2_X1 U14121 ( .A1(n13756), .A2(n14233), .ZN(n14244) );
  NAND2_X1 U14122 ( .A1(n14248), .A2(n14249), .ZN(n14233) );
  NAND2_X1 U14123 ( .A1(n14250), .A2(b_10_), .ZN(n14249) );
  NOR2_X1 U14124 ( .A1(n14251), .A2(n8969), .ZN(n14250) );
  NOR2_X1 U14125 ( .A1(n14229), .A2(n14230), .ZN(n14251) );
  NAND2_X1 U14126 ( .A1(n14229), .A2(n14230), .ZN(n14248) );
  NAND2_X1 U14127 ( .A1(n14252), .A2(n14253), .ZN(n14230) );
  NAND2_X1 U14128 ( .A1(n14227), .A2(n14254), .ZN(n14253) );
  OR2_X1 U14129 ( .A1(n14226), .A2(n14224), .ZN(n14254) );
  NOR2_X1 U14130 ( .A1(n8958), .A2(n8792), .ZN(n14227) );
  NAND2_X1 U14131 ( .A1(n14224), .A2(n14226), .ZN(n14252) );
  NAND2_X1 U14132 ( .A1(n14255), .A2(n14256), .ZN(n14226) );
  NAND2_X1 U14133 ( .A1(n14223), .A2(n14257), .ZN(n14256) );
  OR2_X1 U14134 ( .A1(n14222), .A2(n14220), .ZN(n14257) );
  NOR2_X1 U14135 ( .A1(n8958), .A2(n8778), .ZN(n14223) );
  NAND2_X1 U14136 ( .A1(n14220), .A2(n14222), .ZN(n14255) );
  NAND2_X1 U14137 ( .A1(n14258), .A2(n14259), .ZN(n14222) );
  NAND2_X1 U14138 ( .A1(n14219), .A2(n14260), .ZN(n14259) );
  OR2_X1 U14139 ( .A1(n14218), .A2(n14216), .ZN(n14260) );
  NOR2_X1 U14140 ( .A1(n8958), .A2(n8966), .ZN(n14219) );
  NAND2_X1 U14141 ( .A1(n14216), .A2(n14218), .ZN(n14258) );
  NAND2_X1 U14142 ( .A1(n14261), .A2(n14262), .ZN(n14218) );
  NAND2_X1 U14143 ( .A1(n14215), .A2(n14263), .ZN(n14262) );
  OR2_X1 U14144 ( .A1(n14214), .A2(n14212), .ZN(n14263) );
  NOR2_X1 U14145 ( .A1(n8958), .A2(n8723), .ZN(n14215) );
  NAND2_X1 U14146 ( .A1(n14212), .A2(n14214), .ZN(n14261) );
  NAND2_X1 U14147 ( .A1(n14264), .A2(n14265), .ZN(n14214) );
  NAND2_X1 U14148 ( .A1(n14210), .A2(n14266), .ZN(n14265) );
  NAND2_X1 U14149 ( .A1(n14211), .A2(n14209), .ZN(n14266) );
  NOR2_X1 U14150 ( .A1(n8958), .A2(n8681), .ZN(n14210) );
  OR2_X1 U14151 ( .A1(n14209), .A2(n14211), .ZN(n14264) );
  AND2_X1 U14152 ( .A1(n14267), .A2(n14268), .ZN(n14211) );
  NAND2_X1 U14153 ( .A1(n14207), .A2(n14269), .ZN(n14268) );
  NAND2_X1 U14154 ( .A1(n14206), .A2(n14205), .ZN(n14269) );
  NOR2_X1 U14155 ( .A1(n8958), .A2(n8962), .ZN(n14207) );
  OR2_X1 U14156 ( .A1(n14205), .A2(n14206), .ZN(n14267) );
  AND2_X1 U14157 ( .A1(n14202), .A2(n14270), .ZN(n14206) );
  NAND2_X1 U14158 ( .A1(n14201), .A2(n14203), .ZN(n14270) );
  NAND2_X1 U14159 ( .A1(n14271), .A2(n14272), .ZN(n14203) );
  NAND2_X1 U14160 ( .A1(b_10_), .A2(a_8_), .ZN(n14272) );
  INV_X1 U14161 ( .A(n14273), .ZN(n14271) );
  XOR2_X1 U14162 ( .A(n14274), .B(n14275), .Z(n14201) );
  XOR2_X1 U14163 ( .A(n14276), .B(n14277), .Z(n14274) );
  NAND2_X1 U14164 ( .A1(a_8_), .A2(n14273), .ZN(n14202) );
  NAND2_X1 U14165 ( .A1(n14198), .A2(n14278), .ZN(n14273) );
  NAND2_X1 U14166 ( .A1(n14197), .A2(n14199), .ZN(n14278) );
  NAND2_X1 U14167 ( .A1(n14279), .A2(n14280), .ZN(n14199) );
  NAND2_X1 U14168 ( .A1(b_10_), .A2(a_9_), .ZN(n14280) );
  INV_X1 U14169 ( .A(n14281), .ZN(n14279) );
  XOR2_X1 U14170 ( .A(n14282), .B(n14283), .Z(n14197) );
  XOR2_X1 U14171 ( .A(n14284), .B(n14285), .Z(n14282) );
  NOR2_X1 U14172 ( .A1(n8959), .A2(n8960), .ZN(n14285) );
  NAND2_X1 U14173 ( .A1(a_9_), .A2(n14281), .ZN(n14198) );
  NAND2_X1 U14174 ( .A1(n14286), .A2(n14287), .ZN(n14281) );
  NAND2_X1 U14175 ( .A1(n14193), .A2(n14288), .ZN(n14287) );
  OR2_X1 U14176 ( .A1(n14195), .A2(n14289), .ZN(n14288) );
  XOR2_X1 U14177 ( .A(n14290), .B(n14291), .Z(n14193) );
  XOR2_X1 U14178 ( .A(n14292), .B(n14293), .Z(n14290) );
  NOR2_X1 U14179 ( .A1(n8550), .A2(n8960), .ZN(n14293) );
  NAND2_X1 U14180 ( .A1(n14289), .A2(n14195), .ZN(n14286) );
  NAND2_X1 U14181 ( .A1(n14191), .A2(n14294), .ZN(n14195) );
  NAND2_X1 U14182 ( .A1(n14190), .A2(n14192), .ZN(n14294) );
  NAND2_X1 U14183 ( .A1(n14295), .A2(n14296), .ZN(n14192) );
  NAND2_X1 U14184 ( .A1(b_10_), .A2(a_11_), .ZN(n14296) );
  INV_X1 U14185 ( .A(n14297), .ZN(n14295) );
  XNOR2_X1 U14186 ( .A(n14298), .B(n14299), .ZN(n14190) );
  XOR2_X1 U14187 ( .A(n14300), .B(n14301), .Z(n14299) );
  NAND2_X1 U14188 ( .A1(b_9_), .A2(a_12_), .ZN(n14301) );
  NAND2_X1 U14189 ( .A1(a_11_), .A2(n14297), .ZN(n14191) );
  NAND2_X1 U14190 ( .A1(n14045), .A2(n14302), .ZN(n14297) );
  NAND2_X1 U14191 ( .A1(n14044), .A2(n14046), .ZN(n14302) );
  NAND2_X1 U14192 ( .A1(n14303), .A2(n14304), .ZN(n14046) );
  NAND2_X1 U14193 ( .A1(b_10_), .A2(a_12_), .ZN(n14304) );
  INV_X1 U14194 ( .A(n14305), .ZN(n14303) );
  XNOR2_X1 U14195 ( .A(n14306), .B(n14307), .ZN(n14044) );
  XOR2_X1 U14196 ( .A(n14308), .B(n14309), .Z(n14307) );
  NAND2_X1 U14197 ( .A1(b_9_), .A2(a_13_), .ZN(n14309) );
  NAND2_X1 U14198 ( .A1(a_12_), .A2(n14305), .ZN(n14045) );
  NAND2_X1 U14199 ( .A1(n14187), .A2(n14310), .ZN(n14305) );
  NAND2_X1 U14200 ( .A1(n14186), .A2(n14188), .ZN(n14310) );
  NAND2_X1 U14201 ( .A1(n14311), .A2(n14312), .ZN(n14188) );
  NAND2_X1 U14202 ( .A1(b_10_), .A2(a_13_), .ZN(n14312) );
  INV_X1 U14203 ( .A(n14313), .ZN(n14311) );
  XNOR2_X1 U14204 ( .A(n14314), .B(n14315), .ZN(n14186) );
  XOR2_X1 U14205 ( .A(n14316), .B(n14317), .Z(n14315) );
  NAND2_X1 U14206 ( .A1(b_9_), .A2(a_14_), .ZN(n14317) );
  NAND2_X1 U14207 ( .A1(a_13_), .A2(n14313), .ZN(n14187) );
  NAND2_X1 U14208 ( .A1(n14183), .A2(n14318), .ZN(n14313) );
  NAND2_X1 U14209 ( .A1(n14182), .A2(n14184), .ZN(n14318) );
  NAND2_X1 U14210 ( .A1(n14319), .A2(n14320), .ZN(n14184) );
  NAND2_X1 U14211 ( .A1(b_10_), .A2(a_14_), .ZN(n14320) );
  INV_X1 U14212 ( .A(n14321), .ZN(n14319) );
  XNOR2_X1 U14213 ( .A(n14322), .B(n14323), .ZN(n14182) );
  XOR2_X1 U14214 ( .A(n14324), .B(n14325), .Z(n14323) );
  NAND2_X1 U14215 ( .A1(b_9_), .A2(a_15_), .ZN(n14325) );
  NAND2_X1 U14216 ( .A1(a_14_), .A2(n14321), .ZN(n14183) );
  NAND2_X1 U14217 ( .A1(n14179), .A2(n14326), .ZN(n14321) );
  NAND2_X1 U14218 ( .A1(n14178), .A2(n14180), .ZN(n14326) );
  NAND2_X1 U14219 ( .A1(n14327), .A2(n14328), .ZN(n14180) );
  NAND2_X1 U14220 ( .A1(b_10_), .A2(a_15_), .ZN(n14328) );
  INV_X1 U14221 ( .A(n14329), .ZN(n14327) );
  XOR2_X1 U14222 ( .A(n14330), .B(n14331), .Z(n14178) );
  XOR2_X1 U14223 ( .A(n14332), .B(n14333), .Z(n14330) );
  NOR2_X1 U14224 ( .A1(n8950), .A2(n8960), .ZN(n14333) );
  NAND2_X1 U14225 ( .A1(a_15_), .A2(n14329), .ZN(n14179) );
  NAND2_X1 U14226 ( .A1(n14175), .A2(n14334), .ZN(n14329) );
  NAND2_X1 U14227 ( .A1(n14174), .A2(n14176), .ZN(n14334) );
  NAND2_X1 U14228 ( .A1(n14335), .A2(n14336), .ZN(n14176) );
  NAND2_X1 U14229 ( .A1(b_10_), .A2(a_16_), .ZN(n14336) );
  INV_X1 U14230 ( .A(n14337), .ZN(n14335) );
  XOR2_X1 U14231 ( .A(n14338), .B(n14339), .Z(n14174) );
  XOR2_X1 U14232 ( .A(n14340), .B(n14341), .Z(n14338) );
  NOR2_X1 U14233 ( .A1(n8385), .A2(n8960), .ZN(n14341) );
  NAND2_X1 U14234 ( .A1(a_16_), .A2(n14337), .ZN(n14175) );
  NAND2_X1 U14235 ( .A1(n14342), .A2(n14343), .ZN(n14337) );
  NAND2_X1 U14236 ( .A1(n14344), .A2(b_10_), .ZN(n14343) );
  NOR2_X1 U14237 ( .A1(n14345), .A2(n8385), .ZN(n14344) );
  NOR2_X1 U14238 ( .A1(n14171), .A2(n14169), .ZN(n14345) );
  NAND2_X1 U14239 ( .A1(n14169), .A2(n14171), .ZN(n14342) );
  NAND2_X1 U14240 ( .A1(n14346), .A2(n14347), .ZN(n14171) );
  NAND2_X1 U14241 ( .A1(n14168), .A2(n14348), .ZN(n14347) );
  OR2_X1 U14242 ( .A1(n14167), .A2(n14165), .ZN(n14348) );
  NOR2_X1 U14243 ( .A1(n8958), .A2(n8947), .ZN(n14168) );
  NAND2_X1 U14244 ( .A1(n14165), .A2(n14167), .ZN(n14346) );
  NAND2_X1 U14245 ( .A1(n14349), .A2(n14350), .ZN(n14167) );
  NAND2_X1 U14246 ( .A1(n14077), .A2(n14351), .ZN(n14350) );
  NAND2_X1 U14247 ( .A1(n14078), .A2(n14076), .ZN(n14351) );
  NOR2_X1 U14248 ( .A1(n8958), .A2(n8324), .ZN(n14077) );
  OR2_X1 U14249 ( .A1(n14076), .A2(n14078), .ZN(n14349) );
  AND2_X1 U14250 ( .A1(n14352), .A2(n14353), .ZN(n14078) );
  NAND2_X1 U14251 ( .A1(n14164), .A2(n14354), .ZN(n14353) );
  OR2_X1 U14252 ( .A1(n14163), .A2(n14161), .ZN(n14354) );
  NOR2_X1 U14253 ( .A1(n8958), .A2(n8944), .ZN(n14164) );
  NAND2_X1 U14254 ( .A1(n14161), .A2(n14163), .ZN(n14352) );
  NAND2_X1 U14255 ( .A1(n14355), .A2(n14356), .ZN(n14163) );
  NAND2_X1 U14256 ( .A1(n14357), .A2(b_10_), .ZN(n14356) );
  NOR2_X1 U14257 ( .A1(n14358), .A2(n8268), .ZN(n14357) );
  NOR2_X1 U14258 ( .A1(n14157), .A2(n14159), .ZN(n14358) );
  NAND2_X1 U14259 ( .A1(n14157), .A2(n14159), .ZN(n14355) );
  NAND2_X1 U14260 ( .A1(n14359), .A2(n14360), .ZN(n14159) );
  NAND2_X1 U14261 ( .A1(n14361), .A2(b_10_), .ZN(n14360) );
  NOR2_X1 U14262 ( .A1(n14362), .A2(n8941), .ZN(n14361) );
  NOR2_X1 U14263 ( .A1(n14154), .A2(n14155), .ZN(n14362) );
  NAND2_X1 U14264 ( .A1(n14154), .A2(n14155), .ZN(n14359) );
  NAND2_X1 U14265 ( .A1(n14363), .A2(n14364), .ZN(n14155) );
  NAND2_X1 U14266 ( .A1(n14152), .A2(n14365), .ZN(n14364) );
  OR2_X1 U14267 ( .A1(n14149), .A2(n14151), .ZN(n14365) );
  NOR2_X1 U14268 ( .A1(n8958), .A2(n8213), .ZN(n14152) );
  NAND2_X1 U14269 ( .A1(n14149), .A2(n14151), .ZN(n14363) );
  NAND2_X1 U14270 ( .A1(n14366), .A2(n14367), .ZN(n14151) );
  NAND2_X1 U14271 ( .A1(n14368), .A2(b_10_), .ZN(n14367) );
  NOR2_X1 U14272 ( .A1(n14369), .A2(n8939), .ZN(n14368) );
  NOR2_X1 U14273 ( .A1(n14146), .A2(n14147), .ZN(n14369) );
  NAND2_X1 U14274 ( .A1(n14146), .A2(n14147), .ZN(n14366) );
  NAND2_X1 U14275 ( .A1(n14370), .A2(n14371), .ZN(n14147) );
  NAND2_X1 U14276 ( .A1(n14144), .A2(n14372), .ZN(n14371) );
  OR2_X1 U14277 ( .A1(n14141), .A2(n14143), .ZN(n14372) );
  NOR2_X1 U14278 ( .A1(n8958), .A2(n8158), .ZN(n14144) );
  NAND2_X1 U14279 ( .A1(n14141), .A2(n14143), .ZN(n14370) );
  NAND2_X1 U14280 ( .A1(n14139), .A2(n14373), .ZN(n14143) );
  NAND2_X1 U14281 ( .A1(n14138), .A2(n14140), .ZN(n14373) );
  NAND2_X1 U14282 ( .A1(n14374), .A2(n14375), .ZN(n14140) );
  NAND2_X1 U14283 ( .A1(b_10_), .A2(a_26_), .ZN(n14375) );
  INV_X1 U14284 ( .A(n14376), .ZN(n14374) );
  XNOR2_X1 U14285 ( .A(n14377), .B(n14378), .ZN(n14138) );
  NAND2_X1 U14286 ( .A1(n14379), .A2(n14380), .ZN(n14377) );
  NAND2_X1 U14287 ( .A1(a_26_), .A2(n14376), .ZN(n14139) );
  NAND2_X1 U14288 ( .A1(n14109), .A2(n14381), .ZN(n14376) );
  NAND2_X1 U14289 ( .A1(n14108), .A2(n14110), .ZN(n14381) );
  NAND2_X1 U14290 ( .A1(n14382), .A2(n14383), .ZN(n14110) );
  NAND2_X1 U14291 ( .A1(b_10_), .A2(a_27_), .ZN(n14383) );
  INV_X1 U14292 ( .A(n14384), .ZN(n14382) );
  XOR2_X1 U14293 ( .A(n14385), .B(n14386), .Z(n14108) );
  XNOR2_X1 U14294 ( .A(n14387), .B(n14388), .ZN(n14385) );
  NAND2_X1 U14295 ( .A1(b_9_), .A2(a_28_), .ZN(n14387) );
  NAND2_X1 U14296 ( .A1(a_27_), .A2(n14384), .ZN(n14109) );
  NAND2_X1 U14297 ( .A1(n14389), .A2(n14390), .ZN(n14384) );
  NAND2_X1 U14298 ( .A1(n14391), .A2(b_10_), .ZN(n14390) );
  NOR2_X1 U14299 ( .A1(n14392), .A2(n8055), .ZN(n14391) );
  NOR2_X1 U14300 ( .A1(n14116), .A2(n14118), .ZN(n14392) );
  NAND2_X1 U14301 ( .A1(n14116), .A2(n14118), .ZN(n14389) );
  NAND2_X1 U14302 ( .A1(n14393), .A2(n14394), .ZN(n14118) );
  NAND2_X1 U14303 ( .A1(n14134), .A2(n14395), .ZN(n14394) );
  OR2_X1 U14304 ( .A1(n14135), .A2(n14136), .ZN(n14395) );
  NOR2_X1 U14305 ( .A1(n8958), .A2(n8041), .ZN(n14134) );
  NAND2_X1 U14306 ( .A1(n14136), .A2(n14135), .ZN(n14393) );
  NAND2_X1 U14307 ( .A1(n14396), .A2(n14397), .ZN(n14135) );
  NAND2_X1 U14308 ( .A1(b_8_), .A2(n14398), .ZN(n14397) );
  NAND2_X1 U14309 ( .A1(n8003), .A2(n14399), .ZN(n14398) );
  NAND2_X1 U14310 ( .A1(a_31_), .A2(n8960), .ZN(n14399) );
  NAND2_X1 U14311 ( .A1(b_9_), .A2(n14400), .ZN(n14396) );
  NAND2_X1 U14312 ( .A1(n9341), .A2(n14401), .ZN(n14400) );
  NAND2_X1 U14313 ( .A1(a_30_), .A2(n8961), .ZN(n14401) );
  AND2_X1 U14314 ( .A1(n14402), .A2(n7953), .ZN(n14136) );
  NOR2_X1 U14315 ( .A1(n8958), .A2(n8960), .ZN(n14402) );
  XOR2_X1 U14316 ( .A(n14403), .B(n14404), .Z(n14116) );
  XOR2_X1 U14317 ( .A(n14405), .B(n14406), .Z(n14403) );
  XNOR2_X1 U14318 ( .A(n14407), .B(n14408), .ZN(n14141) );
  NAND2_X1 U14319 ( .A1(n14409), .A2(n14410), .ZN(n14407) );
  XNOR2_X1 U14320 ( .A(n14411), .B(n14412), .ZN(n14146) );
  XNOR2_X1 U14321 ( .A(n14413), .B(n14414), .ZN(n14412) );
  XOR2_X1 U14322 ( .A(n14415), .B(n14416), .Z(n14149) );
  XOR2_X1 U14323 ( .A(n14417), .B(n14418), .Z(n14415) );
  NOR2_X1 U14324 ( .A1(n8939), .A2(n8960), .ZN(n14418) );
  XNOR2_X1 U14325 ( .A(n14419), .B(n14420), .ZN(n14154) );
  XNOR2_X1 U14326 ( .A(n14421), .B(n14422), .ZN(n14420) );
  XOR2_X1 U14327 ( .A(n14423), .B(n14424), .Z(n14157) );
  XOR2_X1 U14328 ( .A(n14425), .B(n14426), .Z(n14423) );
  XOR2_X1 U14329 ( .A(n14427), .B(n14428), .Z(n14161) );
  XOR2_X1 U14330 ( .A(n14429), .B(n14430), .Z(n14427) );
  NOR2_X1 U14331 ( .A1(n8268), .A2(n8960), .ZN(n14430) );
  XNOR2_X1 U14332 ( .A(n14431), .B(n14432), .ZN(n14076) );
  XOR2_X1 U14333 ( .A(n14433), .B(n14434), .Z(n14431) );
  NOR2_X1 U14334 ( .A1(n8944), .A2(n8960), .ZN(n14434) );
  XOR2_X1 U14335 ( .A(n14435), .B(n14436), .Z(n14165) );
  XOR2_X1 U14336 ( .A(n14437), .B(n14438), .Z(n14435) );
  NOR2_X1 U14337 ( .A1(n8324), .A2(n8960), .ZN(n14438) );
  XOR2_X1 U14338 ( .A(n14439), .B(n14440), .Z(n14169) );
  XOR2_X1 U14339 ( .A(n14441), .B(n14442), .Z(n14439) );
  NOR2_X1 U14340 ( .A1(n8947), .A2(n8960), .ZN(n14442) );
  INV_X1 U14341 ( .A(n8583), .ZN(n14289) );
  NAND2_X1 U14342 ( .A1(b_10_), .A2(a_10_), .ZN(n8583) );
  XNOR2_X1 U14343 ( .A(n14443), .B(n14444), .ZN(n14205) );
  XNOR2_X1 U14344 ( .A(n14445), .B(n14446), .ZN(n14443) );
  NAND2_X1 U14345 ( .A1(b_9_), .A2(a_8_), .ZN(n14445) );
  XNOR2_X1 U14346 ( .A(n14447), .B(n14448), .ZN(n14209) );
  XOR2_X1 U14347 ( .A(n14449), .B(n14450), .Z(n14447) );
  NOR2_X1 U14348 ( .A1(n8962), .A2(n8960), .ZN(n14450) );
  XOR2_X1 U14349 ( .A(n14451), .B(n14452), .Z(n14212) );
  XOR2_X1 U14350 ( .A(n14453), .B(n14454), .Z(n14451) );
  NOR2_X1 U14351 ( .A1(n8681), .A2(n8960), .ZN(n14454) );
  XOR2_X1 U14352 ( .A(n14455), .B(n14456), .Z(n14216) );
  XOR2_X1 U14353 ( .A(n14457), .B(n14458), .Z(n14455) );
  NOR2_X1 U14354 ( .A1(n8723), .A2(n8960), .ZN(n14458) );
  XOR2_X1 U14355 ( .A(n14459), .B(n14460), .Z(n14220) );
  XOR2_X1 U14356 ( .A(n14461), .B(n14462), .Z(n14459) );
  NOR2_X1 U14357 ( .A1(n8966), .A2(n8960), .ZN(n14462) );
  XNOR2_X1 U14358 ( .A(n14463), .B(n14464), .ZN(n14224) );
  XOR2_X1 U14359 ( .A(n14465), .B(n14466), .Z(n14464) );
  NAND2_X1 U14360 ( .A1(b_9_), .A2(a_3_), .ZN(n14466) );
  XNOR2_X1 U14361 ( .A(n14467), .B(n14468), .ZN(n14229) );
  XOR2_X1 U14362 ( .A(n14469), .B(n14470), .Z(n14468) );
  NAND2_X1 U14363 ( .A1(b_9_), .A2(a_2_), .ZN(n14470) );
  XOR2_X1 U14364 ( .A(n14471), .B(n14472), .Z(n13756) );
  XOR2_X1 U14365 ( .A(n14473), .B(n14474), .Z(n14471) );
  NOR2_X1 U14366 ( .A1(n8969), .A2(n8960), .ZN(n14474) );
  XOR2_X1 U14367 ( .A(n14475), .B(n14476), .Z(n13995) );
  XOR2_X1 U14368 ( .A(n14477), .B(n14478), .Z(n14475) );
  NAND2_X1 U14369 ( .A1(n14479), .A2(n14237), .ZN(n7968) );
  OR2_X1 U14370 ( .A1(n14237), .A2(n14479), .ZN(n7969) );
  XNOR2_X1 U14371 ( .A(n14480), .B(n14481), .ZN(n14479) );
  NAND2_X1 U14372 ( .A1(n14482), .A2(n14241), .ZN(n14237) );
  NAND2_X1 U14373 ( .A1(n14483), .A2(n14484), .ZN(n14241) );
  NAND2_X1 U14374 ( .A1(n14478), .A2(n14485), .ZN(n14484) );
  OR2_X1 U14375 ( .A1(n14476), .A2(n14477), .ZN(n14485) );
  NOR2_X1 U14376 ( .A1(n8960), .A2(n8974), .ZN(n14478) );
  NAND2_X1 U14377 ( .A1(n14476), .A2(n14477), .ZN(n14483) );
  NAND2_X1 U14378 ( .A1(n14486), .A2(n14487), .ZN(n14477) );
  NAND2_X1 U14379 ( .A1(n14488), .A2(b_9_), .ZN(n14487) );
  NOR2_X1 U14380 ( .A1(n14489), .A2(n8969), .ZN(n14488) );
  NOR2_X1 U14381 ( .A1(n14473), .A2(n14472), .ZN(n14489) );
  NAND2_X1 U14382 ( .A1(n14472), .A2(n14473), .ZN(n14486) );
  NAND2_X1 U14383 ( .A1(n14490), .A2(n14491), .ZN(n14473) );
  NAND2_X1 U14384 ( .A1(n14492), .A2(b_9_), .ZN(n14491) );
  NOR2_X1 U14385 ( .A1(n14493), .A2(n8792), .ZN(n14492) );
  NOR2_X1 U14386 ( .A1(n14469), .A2(n14467), .ZN(n14493) );
  NAND2_X1 U14387 ( .A1(n14467), .A2(n14469), .ZN(n14490) );
  NAND2_X1 U14388 ( .A1(n14494), .A2(n14495), .ZN(n14469) );
  NAND2_X1 U14389 ( .A1(n14496), .A2(b_9_), .ZN(n14495) );
  NOR2_X1 U14390 ( .A1(n14497), .A2(n8778), .ZN(n14496) );
  NOR2_X1 U14391 ( .A1(n14465), .A2(n14463), .ZN(n14497) );
  NAND2_X1 U14392 ( .A1(n14463), .A2(n14465), .ZN(n14494) );
  NAND2_X1 U14393 ( .A1(n14498), .A2(n14499), .ZN(n14465) );
  NAND2_X1 U14394 ( .A1(n14500), .A2(b_9_), .ZN(n14499) );
  NOR2_X1 U14395 ( .A1(n14501), .A2(n8966), .ZN(n14500) );
  NOR2_X1 U14396 ( .A1(n14461), .A2(n14460), .ZN(n14501) );
  NAND2_X1 U14397 ( .A1(n14460), .A2(n14461), .ZN(n14498) );
  NAND2_X1 U14398 ( .A1(n14502), .A2(n14503), .ZN(n14461) );
  NAND2_X1 U14399 ( .A1(n14504), .A2(b_9_), .ZN(n14503) );
  NOR2_X1 U14400 ( .A1(n14505), .A2(n8723), .ZN(n14504) );
  NOR2_X1 U14401 ( .A1(n14457), .A2(n14456), .ZN(n14505) );
  NAND2_X1 U14402 ( .A1(n14456), .A2(n14457), .ZN(n14502) );
  NAND2_X1 U14403 ( .A1(n14506), .A2(n14507), .ZN(n14457) );
  NAND2_X1 U14404 ( .A1(n14508), .A2(b_9_), .ZN(n14507) );
  NOR2_X1 U14405 ( .A1(n14509), .A2(n8681), .ZN(n14508) );
  NOR2_X1 U14406 ( .A1(n14453), .A2(n14452), .ZN(n14509) );
  NAND2_X1 U14407 ( .A1(n14452), .A2(n14453), .ZN(n14506) );
  NAND2_X1 U14408 ( .A1(n14510), .A2(n14511), .ZN(n14453) );
  NAND2_X1 U14409 ( .A1(n14512), .A2(b_9_), .ZN(n14511) );
  NOR2_X1 U14410 ( .A1(n14513), .A2(n8962), .ZN(n14512) );
  NOR2_X1 U14411 ( .A1(n14449), .A2(n14448), .ZN(n14513) );
  NAND2_X1 U14412 ( .A1(n14448), .A2(n14449), .ZN(n14510) );
  NAND2_X1 U14413 ( .A1(n14514), .A2(n14515), .ZN(n14449) );
  NAND2_X1 U14414 ( .A1(n14516), .A2(b_9_), .ZN(n14515) );
  NOR2_X1 U14415 ( .A1(n14517), .A2(n8619), .ZN(n14516) );
  NOR2_X1 U14416 ( .A1(n14446), .A2(n14444), .ZN(n14517) );
  NAND2_X1 U14417 ( .A1(n14444), .A2(n14446), .ZN(n14514) );
  NAND2_X1 U14418 ( .A1(n14518), .A2(n14519), .ZN(n14446) );
  NAND2_X1 U14419 ( .A1(n14275), .A2(n14520), .ZN(n14519) );
  OR2_X1 U14420 ( .A1(n14276), .A2(n14277), .ZN(n14520) );
  XNOR2_X1 U14421 ( .A(n14521), .B(n14522), .ZN(n14275) );
  XNOR2_X1 U14422 ( .A(n14523), .B(n14524), .ZN(n14522) );
  NAND2_X1 U14423 ( .A1(n14277), .A2(n14276), .ZN(n14518) );
  NAND2_X1 U14424 ( .A1(n14525), .A2(n14526), .ZN(n14276) );
  NAND2_X1 U14425 ( .A1(n14527), .A2(b_9_), .ZN(n14526) );
  NOR2_X1 U14426 ( .A1(n14528), .A2(n8959), .ZN(n14527) );
  NOR2_X1 U14427 ( .A1(n14284), .A2(n14283), .ZN(n14528) );
  NAND2_X1 U14428 ( .A1(n14283), .A2(n14284), .ZN(n14525) );
  NAND2_X1 U14429 ( .A1(n14529), .A2(n14530), .ZN(n14284) );
  NAND2_X1 U14430 ( .A1(n14531), .A2(b_9_), .ZN(n14530) );
  NOR2_X1 U14431 ( .A1(n14532), .A2(n8550), .ZN(n14531) );
  NOR2_X1 U14432 ( .A1(n14291), .A2(n14292), .ZN(n14532) );
  NAND2_X1 U14433 ( .A1(n14291), .A2(n14292), .ZN(n14529) );
  NAND2_X1 U14434 ( .A1(n14533), .A2(n14534), .ZN(n14292) );
  NAND2_X1 U14435 ( .A1(n14535), .A2(b_9_), .ZN(n14534) );
  NOR2_X1 U14436 ( .A1(n14536), .A2(n8956), .ZN(n14535) );
  NOR2_X1 U14437 ( .A1(n14300), .A2(n14298), .ZN(n14536) );
  NAND2_X1 U14438 ( .A1(n14298), .A2(n14300), .ZN(n14533) );
  NAND2_X1 U14439 ( .A1(n14537), .A2(n14538), .ZN(n14300) );
  NAND2_X1 U14440 ( .A1(n14539), .A2(b_9_), .ZN(n14538) );
  NOR2_X1 U14441 ( .A1(n14540), .A2(n8495), .ZN(n14539) );
  NOR2_X1 U14442 ( .A1(n14306), .A2(n14308), .ZN(n14540) );
  NAND2_X1 U14443 ( .A1(n14306), .A2(n14308), .ZN(n14537) );
  NAND2_X1 U14444 ( .A1(n14541), .A2(n14542), .ZN(n14308) );
  NAND2_X1 U14445 ( .A1(n14543), .A2(b_9_), .ZN(n14542) );
  NOR2_X1 U14446 ( .A1(n14544), .A2(n8953), .ZN(n14543) );
  NOR2_X1 U14447 ( .A1(n14316), .A2(n14314), .ZN(n14544) );
  NAND2_X1 U14448 ( .A1(n14314), .A2(n14316), .ZN(n14541) );
  NAND2_X1 U14449 ( .A1(n14545), .A2(n14546), .ZN(n14316) );
  NAND2_X1 U14450 ( .A1(n14547), .A2(b_9_), .ZN(n14546) );
  NOR2_X1 U14451 ( .A1(n14548), .A2(n8440), .ZN(n14547) );
  NOR2_X1 U14452 ( .A1(n14324), .A2(n14322), .ZN(n14548) );
  NAND2_X1 U14453 ( .A1(n14322), .A2(n14324), .ZN(n14545) );
  NAND2_X1 U14454 ( .A1(n14549), .A2(n14550), .ZN(n14324) );
  NAND2_X1 U14455 ( .A1(n14551), .A2(b_9_), .ZN(n14550) );
  NOR2_X1 U14456 ( .A1(n14552), .A2(n8950), .ZN(n14551) );
  NOR2_X1 U14457 ( .A1(n14331), .A2(n14332), .ZN(n14552) );
  NAND2_X1 U14458 ( .A1(n14331), .A2(n14332), .ZN(n14549) );
  NAND2_X1 U14459 ( .A1(n14553), .A2(n14554), .ZN(n14332) );
  NAND2_X1 U14460 ( .A1(n14555), .A2(b_9_), .ZN(n14554) );
  NOR2_X1 U14461 ( .A1(n14556), .A2(n8385), .ZN(n14555) );
  NOR2_X1 U14462 ( .A1(n14339), .A2(n14340), .ZN(n14556) );
  NAND2_X1 U14463 ( .A1(n14339), .A2(n14340), .ZN(n14553) );
  NAND2_X1 U14464 ( .A1(n14557), .A2(n14558), .ZN(n14340) );
  NAND2_X1 U14465 ( .A1(n14559), .A2(b_9_), .ZN(n14558) );
  NOR2_X1 U14466 ( .A1(n14560), .A2(n8947), .ZN(n14559) );
  NOR2_X1 U14467 ( .A1(n14440), .A2(n14441), .ZN(n14560) );
  NAND2_X1 U14468 ( .A1(n14440), .A2(n14441), .ZN(n14557) );
  NAND2_X1 U14469 ( .A1(n14561), .A2(n14562), .ZN(n14441) );
  NAND2_X1 U14470 ( .A1(n14563), .A2(b_9_), .ZN(n14562) );
  NOR2_X1 U14471 ( .A1(n14564), .A2(n8324), .ZN(n14563) );
  NOR2_X1 U14472 ( .A1(n14437), .A2(n14436), .ZN(n14564) );
  NAND2_X1 U14473 ( .A1(n14436), .A2(n14437), .ZN(n14561) );
  NAND2_X1 U14474 ( .A1(n14565), .A2(n14566), .ZN(n14437) );
  NAND2_X1 U14475 ( .A1(n14567), .A2(b_9_), .ZN(n14566) );
  NOR2_X1 U14476 ( .A1(n14568), .A2(n8944), .ZN(n14567) );
  NOR2_X1 U14477 ( .A1(n14433), .A2(n14432), .ZN(n14568) );
  NAND2_X1 U14478 ( .A1(n14432), .A2(n14433), .ZN(n14565) );
  NAND2_X1 U14479 ( .A1(n14569), .A2(n14570), .ZN(n14433) );
  NAND2_X1 U14480 ( .A1(n14571), .A2(b_9_), .ZN(n14570) );
  NOR2_X1 U14481 ( .A1(n14572), .A2(n8268), .ZN(n14571) );
  NOR2_X1 U14482 ( .A1(n14429), .A2(n14428), .ZN(n14572) );
  NAND2_X1 U14483 ( .A1(n14428), .A2(n14429), .ZN(n14569) );
  NAND2_X1 U14484 ( .A1(n14573), .A2(n14574), .ZN(n14429) );
  NAND2_X1 U14485 ( .A1(n14426), .A2(n14575), .ZN(n14574) );
  OR2_X1 U14486 ( .A1(n14424), .A2(n14425), .ZN(n14575) );
  NOR2_X1 U14487 ( .A1(n8960), .A2(n8941), .ZN(n14426) );
  NAND2_X1 U14488 ( .A1(n14424), .A2(n14425), .ZN(n14573) );
  NAND2_X1 U14489 ( .A1(n14576), .A2(n14577), .ZN(n14425) );
  NAND2_X1 U14490 ( .A1(n14422), .A2(n14578), .ZN(n14577) );
  OR2_X1 U14491 ( .A1(n14419), .A2(n14421), .ZN(n14578) );
  NOR2_X1 U14492 ( .A1(n8960), .A2(n8213), .ZN(n14422) );
  NAND2_X1 U14493 ( .A1(n14419), .A2(n14421), .ZN(n14576) );
  NAND2_X1 U14494 ( .A1(n14579), .A2(n14580), .ZN(n14421) );
  NAND2_X1 U14495 ( .A1(n14581), .A2(b_9_), .ZN(n14580) );
  NOR2_X1 U14496 ( .A1(n14582), .A2(n8939), .ZN(n14581) );
  NOR2_X1 U14497 ( .A1(n14416), .A2(n14417), .ZN(n14582) );
  NAND2_X1 U14498 ( .A1(n14416), .A2(n14417), .ZN(n14579) );
  NAND2_X1 U14499 ( .A1(n14583), .A2(n14584), .ZN(n14417) );
  NAND2_X1 U14500 ( .A1(n14414), .A2(n14585), .ZN(n14584) );
  OR2_X1 U14501 ( .A1(n14411), .A2(n14413), .ZN(n14585) );
  NOR2_X1 U14502 ( .A1(n8960), .A2(n8158), .ZN(n14414) );
  NAND2_X1 U14503 ( .A1(n14411), .A2(n14413), .ZN(n14583) );
  NAND2_X1 U14504 ( .A1(n14409), .A2(n14586), .ZN(n14413) );
  NAND2_X1 U14505 ( .A1(n14408), .A2(n14410), .ZN(n14586) );
  NAND2_X1 U14506 ( .A1(n14587), .A2(n14588), .ZN(n14410) );
  NAND2_X1 U14507 ( .A1(b_9_), .A2(a_26_), .ZN(n14588) );
  INV_X1 U14508 ( .A(n14589), .ZN(n14587) );
  XNOR2_X1 U14509 ( .A(n14590), .B(n14591), .ZN(n14408) );
  NAND2_X1 U14510 ( .A1(n14592), .A2(n14593), .ZN(n14590) );
  NAND2_X1 U14511 ( .A1(a_26_), .A2(n14589), .ZN(n14409) );
  NAND2_X1 U14512 ( .A1(n14379), .A2(n14594), .ZN(n14589) );
  NAND2_X1 U14513 ( .A1(n14378), .A2(n14380), .ZN(n14594) );
  NAND2_X1 U14514 ( .A1(n14595), .A2(n14596), .ZN(n14380) );
  NAND2_X1 U14515 ( .A1(b_9_), .A2(a_27_), .ZN(n14596) );
  INV_X1 U14516 ( .A(n14597), .ZN(n14595) );
  XOR2_X1 U14517 ( .A(n14598), .B(n14599), .Z(n14378) );
  XNOR2_X1 U14518 ( .A(n14600), .B(n14601), .ZN(n14598) );
  NAND2_X1 U14519 ( .A1(b_8_), .A2(a_28_), .ZN(n14600) );
  NAND2_X1 U14520 ( .A1(a_27_), .A2(n14597), .ZN(n14379) );
  NAND2_X1 U14521 ( .A1(n14602), .A2(n14603), .ZN(n14597) );
  NAND2_X1 U14522 ( .A1(n14604), .A2(b_9_), .ZN(n14603) );
  NOR2_X1 U14523 ( .A1(n14605), .A2(n8055), .ZN(n14604) );
  NOR2_X1 U14524 ( .A1(n14386), .A2(n14388), .ZN(n14605) );
  NAND2_X1 U14525 ( .A1(n14386), .A2(n14388), .ZN(n14602) );
  NAND2_X1 U14526 ( .A1(n14606), .A2(n14607), .ZN(n14388) );
  NAND2_X1 U14527 ( .A1(n14404), .A2(n14608), .ZN(n14607) );
  OR2_X1 U14528 ( .A1(n14405), .A2(n14406), .ZN(n14608) );
  NOR2_X1 U14529 ( .A1(n8960), .A2(n8041), .ZN(n14404) );
  NAND2_X1 U14530 ( .A1(n14406), .A2(n14405), .ZN(n14606) );
  NAND2_X1 U14531 ( .A1(n14609), .A2(n14610), .ZN(n14405) );
  NAND2_X1 U14532 ( .A1(b_7_), .A2(n14611), .ZN(n14610) );
  NAND2_X1 U14533 ( .A1(n8003), .A2(n14612), .ZN(n14611) );
  NAND2_X1 U14534 ( .A1(a_31_), .A2(n8961), .ZN(n14612) );
  NAND2_X1 U14535 ( .A1(b_8_), .A2(n14613), .ZN(n14609) );
  NAND2_X1 U14536 ( .A1(n9341), .A2(n14614), .ZN(n14613) );
  NAND2_X1 U14537 ( .A1(a_30_), .A2(n8667), .ZN(n14614) );
  AND2_X1 U14538 ( .A1(n14615), .A2(n7953), .ZN(n14406) );
  NOR2_X1 U14539 ( .A1(n8960), .A2(n8961), .ZN(n14615) );
  XOR2_X1 U14540 ( .A(n14616), .B(n14617), .Z(n14386) );
  XOR2_X1 U14541 ( .A(n14618), .B(n14619), .Z(n14616) );
  XNOR2_X1 U14542 ( .A(n14620), .B(n14621), .ZN(n14411) );
  NAND2_X1 U14543 ( .A1(n14622), .A2(n14623), .ZN(n14620) );
  XNOR2_X1 U14544 ( .A(n14624), .B(n14625), .ZN(n14416) );
  XNOR2_X1 U14545 ( .A(n14626), .B(n14627), .ZN(n14625) );
  XOR2_X1 U14546 ( .A(n14628), .B(n14629), .Z(n14419) );
  XOR2_X1 U14547 ( .A(n14630), .B(n14631), .Z(n14628) );
  NOR2_X1 U14548 ( .A1(n8939), .A2(n8961), .ZN(n14631) );
  XNOR2_X1 U14549 ( .A(n14632), .B(n14633), .ZN(n14424) );
  XOR2_X1 U14550 ( .A(n14634), .B(n14635), .Z(n14633) );
  NAND2_X1 U14551 ( .A1(b_8_), .A2(a_23_), .ZN(n14635) );
  XNOR2_X1 U14552 ( .A(n14636), .B(n14637), .ZN(n14428) );
  XNOR2_X1 U14553 ( .A(n14638), .B(n14639), .ZN(n14637) );
  XNOR2_X1 U14554 ( .A(n14640), .B(n14641), .ZN(n14432) );
  XNOR2_X1 U14555 ( .A(n14642), .B(n14643), .ZN(n14640) );
  XNOR2_X1 U14556 ( .A(n14644), .B(n14645), .ZN(n14436) );
  XNOR2_X1 U14557 ( .A(n14646), .B(n14647), .ZN(n14644) );
  XOR2_X1 U14558 ( .A(n14648), .B(n14649), .Z(n14440) );
  XOR2_X1 U14559 ( .A(n14650), .B(n14651), .Z(n14648) );
  XOR2_X1 U14560 ( .A(n14652), .B(n14653), .Z(n14339) );
  XOR2_X1 U14561 ( .A(n14654), .B(n14655), .Z(n14652) );
  NOR2_X1 U14562 ( .A1(n8947), .A2(n8961), .ZN(n14655) );
  XNOR2_X1 U14563 ( .A(n14656), .B(n14657), .ZN(n14331) );
  NAND2_X1 U14564 ( .A1(n14658), .A2(n14659), .ZN(n14656) );
  XNOR2_X1 U14565 ( .A(n14660), .B(n14661), .ZN(n14322) );
  NAND2_X1 U14566 ( .A1(n14662), .A2(n14663), .ZN(n14660) );
  XNOR2_X1 U14567 ( .A(n14664), .B(n14665), .ZN(n14314) );
  XNOR2_X1 U14568 ( .A(n14666), .B(n14667), .ZN(n14665) );
  XNOR2_X1 U14569 ( .A(n14668), .B(n14669), .ZN(n14306) );
  XOR2_X1 U14570 ( .A(n14670), .B(n14671), .Z(n14669) );
  NAND2_X1 U14571 ( .A1(b_8_), .A2(a_14_), .ZN(n14671) );
  XNOR2_X1 U14572 ( .A(n14672), .B(n14673), .ZN(n14298) );
  XNOR2_X1 U14573 ( .A(n14674), .B(n14675), .ZN(n14672) );
  XNOR2_X1 U14574 ( .A(n14676), .B(n14677), .ZN(n14291) );
  XNOR2_X1 U14575 ( .A(n14678), .B(n14679), .ZN(n14677) );
  XNOR2_X1 U14576 ( .A(n14680), .B(n14681), .ZN(n14283) );
  XNOR2_X1 U14577 ( .A(n14682), .B(n14683), .ZN(n14680) );
  INV_X1 U14578 ( .A(n8881), .ZN(n14277) );
  NAND2_X1 U14579 ( .A1(b_9_), .A2(a_9_), .ZN(n8881) );
  XNOR2_X1 U14580 ( .A(n14684), .B(n14685), .ZN(n14444) );
  XNOR2_X1 U14581 ( .A(n14686), .B(n14687), .ZN(n14685) );
  XNOR2_X1 U14582 ( .A(n14688), .B(n14689), .ZN(n14448) );
  XOR2_X1 U14583 ( .A(n14690), .B(n8639), .Z(n14689) );
  XNOR2_X1 U14584 ( .A(n14691), .B(n14692), .ZN(n14452) );
  XNOR2_X1 U14585 ( .A(n14693), .B(n14694), .ZN(n14692) );
  XNOR2_X1 U14586 ( .A(n14695), .B(n14696), .ZN(n14456) );
  XNOR2_X1 U14587 ( .A(n14697), .B(n14698), .ZN(n14696) );
  XOR2_X1 U14588 ( .A(n14699), .B(n14700), .Z(n14460) );
  XOR2_X1 U14589 ( .A(n14701), .B(n14702), .Z(n14699) );
  NOR2_X1 U14590 ( .A1(n8723), .A2(n8961), .ZN(n14702) );
  XNOR2_X1 U14591 ( .A(n14703), .B(n14704), .ZN(n14463) );
  XOR2_X1 U14592 ( .A(n14705), .B(n14706), .Z(n14704) );
  NAND2_X1 U14593 ( .A1(b_8_), .A2(a_4_), .ZN(n14706) );
  XOR2_X1 U14594 ( .A(n14707), .B(n14708), .Z(n14467) );
  XOR2_X1 U14595 ( .A(n14709), .B(n14710), .Z(n14707) );
  NOR2_X1 U14596 ( .A1(n8778), .A2(n8961), .ZN(n14710) );
  XOR2_X1 U14597 ( .A(n14711), .B(n14712), .Z(n14472) );
  XOR2_X1 U14598 ( .A(n14713), .B(n14714), .Z(n14711) );
  NOR2_X1 U14599 ( .A1(n8792), .A2(n8961), .ZN(n14714) );
  XOR2_X1 U14600 ( .A(n14715), .B(n14716), .Z(n14476) );
  XOR2_X1 U14601 ( .A(n14717), .B(n14718), .Z(n14715) );
  NOR2_X1 U14602 ( .A1(n8969), .A2(n8961), .ZN(n14718) );
  XOR2_X1 U14603 ( .A(n14719), .B(n14242), .Z(n14482) );
  XNOR2_X1 U14604 ( .A(n14720), .B(n14721), .ZN(n14242) );
  NOR2_X1 U14605 ( .A1(n8974), .A2(n8961), .ZN(n14721) );
  INV_X1 U14606 ( .A(n14243), .ZN(n14719) );
  NAND2_X1 U14607 ( .A1(n14722), .A2(n14723), .ZN(n7975) );
  OR2_X1 U14608 ( .A1(n14723), .A2(n14722), .ZN(n7974) );
  NAND2_X1 U14609 ( .A1(n14724), .A2(n14725), .ZN(n14722) );
  NAND2_X1 U14610 ( .A1(n14726), .A2(n14727), .ZN(n14725) );
  XOR2_X1 U14611 ( .A(n14728), .B(n14729), .Z(n14727) );
  INV_X1 U14612 ( .A(n14730), .ZN(n14726) );
  OR2_X1 U14613 ( .A1(n14481), .A2(n14480), .ZN(n14723) );
  AND2_X1 U14614 ( .A1(n14731), .A2(n14732), .ZN(n14480) );
  NAND2_X1 U14615 ( .A1(n14733), .A2(b_8_), .ZN(n14732) );
  NOR2_X1 U14616 ( .A1(n14734), .A2(n8974), .ZN(n14733) );
  NOR2_X1 U14617 ( .A1(n14243), .A2(n14720), .ZN(n14734) );
  NAND2_X1 U14618 ( .A1(n14243), .A2(n14720), .ZN(n14731) );
  NAND2_X1 U14619 ( .A1(n14735), .A2(n14736), .ZN(n14720) );
  NAND2_X1 U14620 ( .A1(n14737), .A2(b_8_), .ZN(n14736) );
  NOR2_X1 U14621 ( .A1(n14738), .A2(n8969), .ZN(n14737) );
  NOR2_X1 U14622 ( .A1(n14716), .A2(n14717), .ZN(n14738) );
  NAND2_X1 U14623 ( .A1(n14716), .A2(n14717), .ZN(n14735) );
  NAND2_X1 U14624 ( .A1(n14739), .A2(n14740), .ZN(n14717) );
  NAND2_X1 U14625 ( .A1(n14741), .A2(b_8_), .ZN(n14740) );
  NOR2_X1 U14626 ( .A1(n14742), .A2(n8792), .ZN(n14741) );
  NOR2_X1 U14627 ( .A1(n14712), .A2(n14713), .ZN(n14742) );
  NAND2_X1 U14628 ( .A1(n14712), .A2(n14713), .ZN(n14739) );
  NAND2_X1 U14629 ( .A1(n14743), .A2(n14744), .ZN(n14713) );
  NAND2_X1 U14630 ( .A1(n14745), .A2(b_8_), .ZN(n14744) );
  NOR2_X1 U14631 ( .A1(n14746), .A2(n8778), .ZN(n14745) );
  NOR2_X1 U14632 ( .A1(n14708), .A2(n14709), .ZN(n14746) );
  NAND2_X1 U14633 ( .A1(n14708), .A2(n14709), .ZN(n14743) );
  NAND2_X1 U14634 ( .A1(n14747), .A2(n14748), .ZN(n14709) );
  NAND2_X1 U14635 ( .A1(n14749), .A2(b_8_), .ZN(n14748) );
  NOR2_X1 U14636 ( .A1(n14750), .A2(n8966), .ZN(n14749) );
  NOR2_X1 U14637 ( .A1(n14703), .A2(n14705), .ZN(n14750) );
  NAND2_X1 U14638 ( .A1(n14703), .A2(n14705), .ZN(n14747) );
  NAND2_X1 U14639 ( .A1(n14751), .A2(n14752), .ZN(n14705) );
  NAND2_X1 U14640 ( .A1(n14753), .A2(b_8_), .ZN(n14752) );
  NOR2_X1 U14641 ( .A1(n14754), .A2(n8723), .ZN(n14753) );
  NOR2_X1 U14642 ( .A1(n14700), .A2(n14701), .ZN(n14754) );
  NAND2_X1 U14643 ( .A1(n14700), .A2(n14701), .ZN(n14751) );
  NAND2_X1 U14644 ( .A1(n14755), .A2(n14756), .ZN(n14701) );
  NAND2_X1 U14645 ( .A1(n14698), .A2(n14757), .ZN(n14756) );
  OR2_X1 U14646 ( .A1(n14697), .A2(n14695), .ZN(n14757) );
  NOR2_X1 U14647 ( .A1(n8961), .A2(n8681), .ZN(n14698) );
  NAND2_X1 U14648 ( .A1(n14695), .A2(n14697), .ZN(n14755) );
  NAND2_X1 U14649 ( .A1(n14758), .A2(n14759), .ZN(n14697) );
  NAND2_X1 U14650 ( .A1(n14694), .A2(n14760), .ZN(n14759) );
  OR2_X1 U14651 ( .A1(n14693), .A2(n14691), .ZN(n14760) );
  NOR2_X1 U14652 ( .A1(n8961), .A2(n8962), .ZN(n14694) );
  NAND2_X1 U14653 ( .A1(n14691), .A2(n14693), .ZN(n14758) );
  NAND2_X1 U14654 ( .A1(n14761), .A2(n14762), .ZN(n14693) );
  NAND2_X1 U14655 ( .A1(n14763), .A2(n14764), .ZN(n14762) );
  OR2_X1 U14656 ( .A1(n14690), .A2(n14688), .ZN(n14764) );
  INV_X1 U14657 ( .A(n8639), .ZN(n14763) );
  NAND2_X1 U14658 ( .A1(b_8_), .A2(a_8_), .ZN(n8639) );
  NAND2_X1 U14659 ( .A1(n14688), .A2(n14690), .ZN(n14761) );
  NAND2_X1 U14660 ( .A1(n14765), .A2(n14766), .ZN(n14690) );
  NAND2_X1 U14661 ( .A1(n14687), .A2(n14767), .ZN(n14766) );
  OR2_X1 U14662 ( .A1(n14686), .A2(n14684), .ZN(n14767) );
  NOR2_X1 U14663 ( .A1(n8961), .A2(n8605), .ZN(n14687) );
  NAND2_X1 U14664 ( .A1(n14684), .A2(n14686), .ZN(n14765) );
  NAND2_X1 U14665 ( .A1(n14768), .A2(n14769), .ZN(n14686) );
  NAND2_X1 U14666 ( .A1(n14524), .A2(n14770), .ZN(n14769) );
  OR2_X1 U14667 ( .A1(n14523), .A2(n14521), .ZN(n14770) );
  NOR2_X1 U14668 ( .A1(n8961), .A2(n8959), .ZN(n14524) );
  NAND2_X1 U14669 ( .A1(n14521), .A2(n14523), .ZN(n14768) );
  NAND2_X1 U14670 ( .A1(n14771), .A2(n14772), .ZN(n14523) );
  NAND2_X1 U14671 ( .A1(n14683), .A2(n14773), .ZN(n14772) );
  NAND2_X1 U14672 ( .A1(n14682), .A2(n14681), .ZN(n14773) );
  NOR2_X1 U14673 ( .A1(n8961), .A2(n8550), .ZN(n14683) );
  OR2_X1 U14674 ( .A1(n14681), .A2(n14682), .ZN(n14771) );
  AND2_X1 U14675 ( .A1(n14774), .A2(n14775), .ZN(n14682) );
  NAND2_X1 U14676 ( .A1(n14679), .A2(n14776), .ZN(n14775) );
  OR2_X1 U14677 ( .A1(n14676), .A2(n14678), .ZN(n14776) );
  NOR2_X1 U14678 ( .A1(n8961), .A2(n8956), .ZN(n14679) );
  NAND2_X1 U14679 ( .A1(n14676), .A2(n14678), .ZN(n14774) );
  NAND2_X1 U14680 ( .A1(n14777), .A2(n14778), .ZN(n14678) );
  NAND2_X1 U14681 ( .A1(n14674), .A2(n14779), .ZN(n14778) );
  NAND2_X1 U14682 ( .A1(n14675), .A2(n14673), .ZN(n14779) );
  NOR2_X1 U14683 ( .A1(n8961), .A2(n8495), .ZN(n14674) );
  OR2_X1 U14684 ( .A1(n14673), .A2(n14675), .ZN(n14777) );
  AND2_X1 U14685 ( .A1(n14780), .A2(n14781), .ZN(n14675) );
  NAND2_X1 U14686 ( .A1(n14782), .A2(b_8_), .ZN(n14781) );
  NOR2_X1 U14687 ( .A1(n14783), .A2(n8953), .ZN(n14782) );
  NOR2_X1 U14688 ( .A1(n14670), .A2(n14668), .ZN(n14783) );
  NAND2_X1 U14689 ( .A1(n14668), .A2(n14670), .ZN(n14780) );
  NAND2_X1 U14690 ( .A1(n14784), .A2(n14785), .ZN(n14670) );
  NAND2_X1 U14691 ( .A1(n14667), .A2(n14786), .ZN(n14785) );
  OR2_X1 U14692 ( .A1(n14666), .A2(n14664), .ZN(n14786) );
  NOR2_X1 U14693 ( .A1(n8961), .A2(n8440), .ZN(n14667) );
  NAND2_X1 U14694 ( .A1(n14664), .A2(n14666), .ZN(n14784) );
  NAND2_X1 U14695 ( .A1(n14662), .A2(n14787), .ZN(n14666) );
  NAND2_X1 U14696 ( .A1(n14661), .A2(n14663), .ZN(n14787) );
  NAND2_X1 U14697 ( .A1(n14788), .A2(n14789), .ZN(n14663) );
  NAND2_X1 U14698 ( .A1(b_8_), .A2(a_16_), .ZN(n14789) );
  INV_X1 U14699 ( .A(n14790), .ZN(n14788) );
  XOR2_X1 U14700 ( .A(n14791), .B(n14792), .Z(n14661) );
  XNOR2_X1 U14701 ( .A(n14793), .B(n14794), .ZN(n14791) );
  NAND2_X1 U14702 ( .A1(b_7_), .A2(a_17_), .ZN(n14793) );
  NAND2_X1 U14703 ( .A1(a_16_), .A2(n14790), .ZN(n14662) );
  NAND2_X1 U14704 ( .A1(n14658), .A2(n14795), .ZN(n14790) );
  NAND2_X1 U14705 ( .A1(n14657), .A2(n14659), .ZN(n14795) );
  NAND2_X1 U14706 ( .A1(n14796), .A2(n14797), .ZN(n14659) );
  NAND2_X1 U14707 ( .A1(b_8_), .A2(a_17_), .ZN(n14797) );
  INV_X1 U14708 ( .A(n14798), .ZN(n14796) );
  XNOR2_X1 U14709 ( .A(n14799), .B(n14800), .ZN(n14657) );
  XOR2_X1 U14710 ( .A(n14801), .B(n14802), .Z(n14800) );
  NAND2_X1 U14711 ( .A1(b_7_), .A2(a_18_), .ZN(n14802) );
  NAND2_X1 U14712 ( .A1(a_17_), .A2(n14798), .ZN(n14658) );
  NAND2_X1 U14713 ( .A1(n14803), .A2(n14804), .ZN(n14798) );
  NAND2_X1 U14714 ( .A1(n14805), .A2(b_8_), .ZN(n14804) );
  NOR2_X1 U14715 ( .A1(n14806), .A2(n8947), .ZN(n14805) );
  NOR2_X1 U14716 ( .A1(n14654), .A2(n14653), .ZN(n14806) );
  NAND2_X1 U14717 ( .A1(n14653), .A2(n14654), .ZN(n14803) );
  NAND2_X1 U14718 ( .A1(n14807), .A2(n14808), .ZN(n14654) );
  NAND2_X1 U14719 ( .A1(n14651), .A2(n14809), .ZN(n14808) );
  OR2_X1 U14720 ( .A1(n14649), .A2(n14650), .ZN(n14809) );
  NOR2_X1 U14721 ( .A1(n8961), .A2(n8324), .ZN(n14651) );
  NAND2_X1 U14722 ( .A1(n14649), .A2(n14650), .ZN(n14807) );
  NAND2_X1 U14723 ( .A1(n14810), .A2(n14811), .ZN(n14650) );
  NAND2_X1 U14724 ( .A1(n14647), .A2(n14812), .ZN(n14811) );
  NAND2_X1 U14725 ( .A1(n14646), .A2(n14645), .ZN(n14812) );
  NOR2_X1 U14726 ( .A1(n8961), .A2(n8944), .ZN(n14647) );
  OR2_X1 U14727 ( .A1(n14645), .A2(n14646), .ZN(n14810) );
  AND2_X1 U14728 ( .A1(n14813), .A2(n14814), .ZN(n14646) );
  NAND2_X1 U14729 ( .A1(n14642), .A2(n14815), .ZN(n14814) );
  NAND2_X1 U14730 ( .A1(n14643), .A2(n14641), .ZN(n14815) );
  NOR2_X1 U14731 ( .A1(n8961), .A2(n8268), .ZN(n14642) );
  OR2_X1 U14732 ( .A1(n14641), .A2(n14643), .ZN(n14813) );
  AND2_X1 U14733 ( .A1(n14816), .A2(n14817), .ZN(n14643) );
  NAND2_X1 U14734 ( .A1(n14639), .A2(n14818), .ZN(n14817) );
  OR2_X1 U14735 ( .A1(n14638), .A2(n14636), .ZN(n14818) );
  NOR2_X1 U14736 ( .A1(n8961), .A2(n8941), .ZN(n14639) );
  NAND2_X1 U14737 ( .A1(n14636), .A2(n14638), .ZN(n14816) );
  NAND2_X1 U14738 ( .A1(n14819), .A2(n14820), .ZN(n14638) );
  NAND2_X1 U14739 ( .A1(n14821), .A2(b_8_), .ZN(n14820) );
  NOR2_X1 U14740 ( .A1(n14822), .A2(n8213), .ZN(n14821) );
  NOR2_X1 U14741 ( .A1(n14632), .A2(n14634), .ZN(n14822) );
  NAND2_X1 U14742 ( .A1(n14632), .A2(n14634), .ZN(n14819) );
  NAND2_X1 U14743 ( .A1(n14823), .A2(n14824), .ZN(n14634) );
  NAND2_X1 U14744 ( .A1(n14825), .A2(b_8_), .ZN(n14824) );
  NOR2_X1 U14745 ( .A1(n14826), .A2(n8939), .ZN(n14825) );
  NOR2_X1 U14746 ( .A1(n14629), .A2(n14630), .ZN(n14826) );
  NAND2_X1 U14747 ( .A1(n14629), .A2(n14630), .ZN(n14823) );
  NAND2_X1 U14748 ( .A1(n14827), .A2(n14828), .ZN(n14630) );
  NAND2_X1 U14749 ( .A1(n14627), .A2(n14829), .ZN(n14828) );
  OR2_X1 U14750 ( .A1(n14624), .A2(n14626), .ZN(n14829) );
  NOR2_X1 U14751 ( .A1(n8961), .A2(n8158), .ZN(n14627) );
  NAND2_X1 U14752 ( .A1(n14624), .A2(n14626), .ZN(n14827) );
  NAND2_X1 U14753 ( .A1(n14622), .A2(n14830), .ZN(n14626) );
  NAND2_X1 U14754 ( .A1(n14621), .A2(n14623), .ZN(n14830) );
  NAND2_X1 U14755 ( .A1(n14831), .A2(n14832), .ZN(n14623) );
  NAND2_X1 U14756 ( .A1(b_8_), .A2(a_26_), .ZN(n14832) );
  INV_X1 U14757 ( .A(n14833), .ZN(n14831) );
  XNOR2_X1 U14758 ( .A(n14834), .B(n14835), .ZN(n14621) );
  NAND2_X1 U14759 ( .A1(n14836), .A2(n14837), .ZN(n14834) );
  NAND2_X1 U14760 ( .A1(a_26_), .A2(n14833), .ZN(n14622) );
  NAND2_X1 U14761 ( .A1(n14592), .A2(n14838), .ZN(n14833) );
  NAND2_X1 U14762 ( .A1(n14591), .A2(n14593), .ZN(n14838) );
  NAND2_X1 U14763 ( .A1(n14839), .A2(n14840), .ZN(n14593) );
  NAND2_X1 U14764 ( .A1(b_8_), .A2(a_27_), .ZN(n14840) );
  INV_X1 U14765 ( .A(n14841), .ZN(n14839) );
  XOR2_X1 U14766 ( .A(n14842), .B(n14843), .Z(n14591) );
  XNOR2_X1 U14767 ( .A(n14844), .B(n14845), .ZN(n14842) );
  NAND2_X1 U14768 ( .A1(b_7_), .A2(a_28_), .ZN(n14844) );
  NAND2_X1 U14769 ( .A1(a_27_), .A2(n14841), .ZN(n14592) );
  NAND2_X1 U14770 ( .A1(n14846), .A2(n14847), .ZN(n14841) );
  NAND2_X1 U14771 ( .A1(n14848), .A2(b_8_), .ZN(n14847) );
  NOR2_X1 U14772 ( .A1(n14849), .A2(n8055), .ZN(n14848) );
  NOR2_X1 U14773 ( .A1(n14599), .A2(n14601), .ZN(n14849) );
  NAND2_X1 U14774 ( .A1(n14599), .A2(n14601), .ZN(n14846) );
  NAND2_X1 U14775 ( .A1(n14850), .A2(n14851), .ZN(n14601) );
  NAND2_X1 U14776 ( .A1(n14617), .A2(n14852), .ZN(n14851) );
  OR2_X1 U14777 ( .A1(n14618), .A2(n14619), .ZN(n14852) );
  NOR2_X1 U14778 ( .A1(n8961), .A2(n8041), .ZN(n14617) );
  NAND2_X1 U14779 ( .A1(n14619), .A2(n14618), .ZN(n14850) );
  NAND2_X1 U14780 ( .A1(n14853), .A2(n14854), .ZN(n14618) );
  NAND2_X1 U14781 ( .A1(b_6_), .A2(n14855), .ZN(n14854) );
  NAND2_X1 U14782 ( .A1(n8003), .A2(n14856), .ZN(n14855) );
  NAND2_X1 U14783 ( .A1(a_31_), .A2(n8667), .ZN(n14856) );
  NAND2_X1 U14784 ( .A1(b_7_), .A2(n14857), .ZN(n14853) );
  NAND2_X1 U14785 ( .A1(n9341), .A2(n14858), .ZN(n14857) );
  NAND2_X1 U14786 ( .A1(a_30_), .A2(n8963), .ZN(n14858) );
  AND2_X1 U14787 ( .A1(n14859), .A2(n7953), .ZN(n14619) );
  NOR2_X1 U14788 ( .A1(n8961), .A2(n8667), .ZN(n14859) );
  XOR2_X1 U14789 ( .A(n14860), .B(n14861), .Z(n14599) );
  XOR2_X1 U14790 ( .A(n14862), .B(n14863), .Z(n14860) );
  XNOR2_X1 U14791 ( .A(n14864), .B(n14865), .ZN(n14624) );
  NAND2_X1 U14792 ( .A1(n14866), .A2(n14867), .ZN(n14864) );
  XNOR2_X1 U14793 ( .A(n14868), .B(n14869), .ZN(n14629) );
  XNOR2_X1 U14794 ( .A(n14870), .B(n14871), .ZN(n14869) );
  XOR2_X1 U14795 ( .A(n14872), .B(n14873), .Z(n14632) );
  XOR2_X1 U14796 ( .A(n14874), .B(n14875), .Z(n14872) );
  XOR2_X1 U14797 ( .A(n14876), .B(n14877), .Z(n14636) );
  XOR2_X1 U14798 ( .A(n14878), .B(n14879), .Z(n14876) );
  NOR2_X1 U14799 ( .A1(n8213), .A2(n8667), .ZN(n14879) );
  XOR2_X1 U14800 ( .A(n14880), .B(n14881), .Z(n14641) );
  NAND2_X1 U14801 ( .A1(n14882), .A2(n14883), .ZN(n14880) );
  XNOR2_X1 U14802 ( .A(n14884), .B(n14885), .ZN(n14645) );
  XOR2_X1 U14803 ( .A(n14886), .B(n14887), .Z(n14884) );
  NOR2_X1 U14804 ( .A1(n8268), .A2(n8667), .ZN(n14887) );
  XNOR2_X1 U14805 ( .A(n14888), .B(n14889), .ZN(n14649) );
  XOR2_X1 U14806 ( .A(n14890), .B(n14891), .Z(n14889) );
  NAND2_X1 U14807 ( .A1(b_7_), .A2(a_20_), .ZN(n14891) );
  XNOR2_X1 U14808 ( .A(n14892), .B(n14893), .ZN(n14653) );
  XOR2_X1 U14809 ( .A(n14894), .B(n14895), .Z(n14893) );
  NAND2_X1 U14810 ( .A1(b_7_), .A2(a_19_), .ZN(n14895) );
  XOR2_X1 U14811 ( .A(n14896), .B(n14897), .Z(n14664) );
  XOR2_X1 U14812 ( .A(n14898), .B(n14899), .Z(n14896) );
  NOR2_X1 U14813 ( .A1(n8950), .A2(n8667), .ZN(n14899) );
  XOR2_X1 U14814 ( .A(n14900), .B(n14901), .Z(n14668) );
  XOR2_X1 U14815 ( .A(n14902), .B(n14903), .Z(n14900) );
  NOR2_X1 U14816 ( .A1(n8440), .A2(n8667), .ZN(n14903) );
  XNOR2_X1 U14817 ( .A(n14904), .B(n14905), .ZN(n14673) );
  XOR2_X1 U14818 ( .A(n14906), .B(n14907), .Z(n14904) );
  NOR2_X1 U14819 ( .A1(n8953), .A2(n8667), .ZN(n14907) );
  XOR2_X1 U14820 ( .A(n14908), .B(n14909), .Z(n14676) );
  XOR2_X1 U14821 ( .A(n14910), .B(n14911), .Z(n14908) );
  NOR2_X1 U14822 ( .A1(n8495), .A2(n8667), .ZN(n14911) );
  XNOR2_X1 U14823 ( .A(n14912), .B(n14913), .ZN(n14681) );
  XOR2_X1 U14824 ( .A(n14914), .B(n14915), .Z(n14912) );
  NOR2_X1 U14825 ( .A1(n8956), .A2(n8667), .ZN(n14915) );
  XOR2_X1 U14826 ( .A(n14916), .B(n14917), .Z(n14521) );
  XOR2_X1 U14827 ( .A(n14918), .B(n14919), .Z(n14916) );
  NOR2_X1 U14828 ( .A1(n8550), .A2(n8667), .ZN(n14919) );
  XOR2_X1 U14829 ( .A(n14920), .B(n14921), .Z(n14684) );
  XOR2_X1 U14830 ( .A(n14922), .B(n14923), .Z(n14920) );
  NOR2_X1 U14831 ( .A1(n8959), .A2(n8667), .ZN(n14923) );
  XOR2_X1 U14832 ( .A(n14924), .B(n14925), .Z(n14688) );
  XOR2_X1 U14833 ( .A(n14926), .B(n14927), .Z(n14924) );
  NOR2_X1 U14834 ( .A1(n8605), .A2(n8667), .ZN(n14927) );
  XOR2_X1 U14835 ( .A(n14928), .B(n14929), .Z(n14691) );
  XOR2_X1 U14836 ( .A(n14930), .B(n14931), .Z(n14928) );
  NOR2_X1 U14837 ( .A1(n8619), .A2(n8667), .ZN(n14931) );
  XOR2_X1 U14838 ( .A(n14932), .B(n14933), .Z(n14695) );
  XOR2_X1 U14839 ( .A(n14934), .B(n14935), .Z(n14932) );
  XOR2_X1 U14840 ( .A(n14936), .B(n14937), .Z(n14700) );
  XNOR2_X1 U14841 ( .A(n14938), .B(n14939), .ZN(n14936) );
  NAND2_X1 U14842 ( .A1(b_7_), .A2(a_6_), .ZN(n14938) );
  XOR2_X1 U14843 ( .A(n14940), .B(n14941), .Z(n14703) );
  XOR2_X1 U14844 ( .A(n14942), .B(n14943), .Z(n14940) );
  NOR2_X1 U14845 ( .A1(n8723), .A2(n8667), .ZN(n14943) );
  XOR2_X1 U14846 ( .A(n14944), .B(n14945), .Z(n14708) );
  XOR2_X1 U14847 ( .A(n14946), .B(n14947), .Z(n14944) );
  NOR2_X1 U14848 ( .A1(n8966), .A2(n8667), .ZN(n14947) );
  XOR2_X1 U14849 ( .A(n14948), .B(n14949), .Z(n14712) );
  XOR2_X1 U14850 ( .A(n14950), .B(n14951), .Z(n14948) );
  NOR2_X1 U14851 ( .A1(n8778), .A2(n8667), .ZN(n14951) );
  XOR2_X1 U14852 ( .A(n14952), .B(n14953), .Z(n14716) );
  XOR2_X1 U14853 ( .A(n14954), .B(n14955), .Z(n14952) );
  NOR2_X1 U14854 ( .A1(n8792), .A2(n8667), .ZN(n14955) );
  XNOR2_X1 U14855 ( .A(n14956), .B(n14957), .ZN(n14243) );
  XOR2_X1 U14856 ( .A(n14958), .B(n14959), .Z(n14957) );
  NAND2_X1 U14857 ( .A1(b_7_), .A2(a_1_), .ZN(n14959) );
  XOR2_X1 U14858 ( .A(n14960), .B(n14961), .Z(n14481) );
  XNOR2_X1 U14859 ( .A(n14962), .B(n14963), .ZN(n14961) );
  NAND2_X1 U14860 ( .A1(n14964), .A2(n14724), .ZN(n7980) );
  OR2_X1 U14861 ( .A1(n14724), .A2(n14964), .ZN(n7981) );
  XNOR2_X1 U14862 ( .A(n14965), .B(n14966), .ZN(n14964) );
  NAND2_X1 U14863 ( .A1(n14967), .A2(n14730), .ZN(n14724) );
  NAND2_X1 U14864 ( .A1(n14968), .A2(n14969), .ZN(n14730) );
  NAND2_X1 U14865 ( .A1(n14963), .A2(n14970), .ZN(n14969) );
  OR2_X1 U14866 ( .A1(n14960), .A2(n14962), .ZN(n14970) );
  NOR2_X1 U14867 ( .A1(n8667), .A2(n8974), .ZN(n14963) );
  NAND2_X1 U14868 ( .A1(n14960), .A2(n14962), .ZN(n14968) );
  NAND2_X1 U14869 ( .A1(n14971), .A2(n14972), .ZN(n14962) );
  NAND2_X1 U14870 ( .A1(n14973), .A2(b_7_), .ZN(n14972) );
  NOR2_X1 U14871 ( .A1(n14974), .A2(n8969), .ZN(n14973) );
  NOR2_X1 U14872 ( .A1(n14958), .A2(n14956), .ZN(n14974) );
  NAND2_X1 U14873 ( .A1(n14956), .A2(n14958), .ZN(n14971) );
  NAND2_X1 U14874 ( .A1(n14975), .A2(n14976), .ZN(n14958) );
  NAND2_X1 U14875 ( .A1(n14977), .A2(b_7_), .ZN(n14976) );
  NOR2_X1 U14876 ( .A1(n14978), .A2(n8792), .ZN(n14977) );
  NOR2_X1 U14877 ( .A1(n14954), .A2(n14953), .ZN(n14978) );
  NAND2_X1 U14878 ( .A1(n14953), .A2(n14954), .ZN(n14975) );
  NAND2_X1 U14879 ( .A1(n14979), .A2(n14980), .ZN(n14954) );
  NAND2_X1 U14880 ( .A1(n14981), .A2(b_7_), .ZN(n14980) );
  NOR2_X1 U14881 ( .A1(n14982), .A2(n8778), .ZN(n14981) );
  NOR2_X1 U14882 ( .A1(n14950), .A2(n14949), .ZN(n14982) );
  NAND2_X1 U14883 ( .A1(n14949), .A2(n14950), .ZN(n14979) );
  NAND2_X1 U14884 ( .A1(n14983), .A2(n14984), .ZN(n14950) );
  NAND2_X1 U14885 ( .A1(n14985), .A2(b_7_), .ZN(n14984) );
  NOR2_X1 U14886 ( .A1(n14986), .A2(n8966), .ZN(n14985) );
  NOR2_X1 U14887 ( .A1(n14946), .A2(n14945), .ZN(n14986) );
  NAND2_X1 U14888 ( .A1(n14945), .A2(n14946), .ZN(n14983) );
  NAND2_X1 U14889 ( .A1(n14987), .A2(n14988), .ZN(n14946) );
  NAND2_X1 U14890 ( .A1(n14989), .A2(b_7_), .ZN(n14988) );
  NOR2_X1 U14891 ( .A1(n14990), .A2(n8723), .ZN(n14989) );
  NOR2_X1 U14892 ( .A1(n14942), .A2(n14941), .ZN(n14990) );
  NAND2_X1 U14893 ( .A1(n14941), .A2(n14942), .ZN(n14987) );
  NAND2_X1 U14894 ( .A1(n14991), .A2(n14992), .ZN(n14942) );
  NAND2_X1 U14895 ( .A1(n14993), .A2(b_7_), .ZN(n14992) );
  NOR2_X1 U14896 ( .A1(n14994), .A2(n8681), .ZN(n14993) );
  NOR2_X1 U14897 ( .A1(n14939), .A2(n14937), .ZN(n14994) );
  NAND2_X1 U14898 ( .A1(n14937), .A2(n14939), .ZN(n14991) );
  NAND2_X1 U14899 ( .A1(n14995), .A2(n14996), .ZN(n14939) );
  NAND2_X1 U14900 ( .A1(n14933), .A2(n14997), .ZN(n14996) );
  OR2_X1 U14901 ( .A1(n14934), .A2(n14935), .ZN(n14997) );
  XOR2_X1 U14902 ( .A(n14998), .B(n14999), .Z(n14933) );
  XOR2_X1 U14903 ( .A(n15000), .B(n15001), .Z(n14998) );
  NOR2_X1 U14904 ( .A1(n8619), .A2(n8963), .ZN(n15001) );
  NAND2_X1 U14905 ( .A1(n14935), .A2(n14934), .ZN(n14995) );
  NAND2_X1 U14906 ( .A1(n15002), .A2(n15003), .ZN(n14934) );
  NAND2_X1 U14907 ( .A1(n15004), .A2(b_7_), .ZN(n15003) );
  NOR2_X1 U14908 ( .A1(n15005), .A2(n8619), .ZN(n15004) );
  NOR2_X1 U14909 ( .A1(n14930), .A2(n14929), .ZN(n15005) );
  NAND2_X1 U14910 ( .A1(n14929), .A2(n14930), .ZN(n15002) );
  NAND2_X1 U14911 ( .A1(n15006), .A2(n15007), .ZN(n14930) );
  NAND2_X1 U14912 ( .A1(n15008), .A2(b_7_), .ZN(n15007) );
  NOR2_X1 U14913 ( .A1(n15009), .A2(n8605), .ZN(n15008) );
  NOR2_X1 U14914 ( .A1(n14926), .A2(n14925), .ZN(n15009) );
  NAND2_X1 U14915 ( .A1(n14925), .A2(n14926), .ZN(n15006) );
  NAND2_X1 U14916 ( .A1(n15010), .A2(n15011), .ZN(n14926) );
  NAND2_X1 U14917 ( .A1(n15012), .A2(b_7_), .ZN(n15011) );
  NOR2_X1 U14918 ( .A1(n15013), .A2(n8959), .ZN(n15012) );
  NOR2_X1 U14919 ( .A1(n14922), .A2(n14921), .ZN(n15013) );
  NAND2_X1 U14920 ( .A1(n14921), .A2(n14922), .ZN(n15010) );
  NAND2_X1 U14921 ( .A1(n15014), .A2(n15015), .ZN(n14922) );
  NAND2_X1 U14922 ( .A1(n15016), .A2(b_7_), .ZN(n15015) );
  NOR2_X1 U14923 ( .A1(n15017), .A2(n8550), .ZN(n15016) );
  NOR2_X1 U14924 ( .A1(n14918), .A2(n14917), .ZN(n15017) );
  NAND2_X1 U14925 ( .A1(n14917), .A2(n14918), .ZN(n15014) );
  NAND2_X1 U14926 ( .A1(n15018), .A2(n15019), .ZN(n14918) );
  NAND2_X1 U14927 ( .A1(n15020), .A2(b_7_), .ZN(n15019) );
  NOR2_X1 U14928 ( .A1(n15021), .A2(n8956), .ZN(n15020) );
  NOR2_X1 U14929 ( .A1(n14914), .A2(n14913), .ZN(n15021) );
  NAND2_X1 U14930 ( .A1(n14913), .A2(n14914), .ZN(n15018) );
  NAND2_X1 U14931 ( .A1(n15022), .A2(n15023), .ZN(n14914) );
  NAND2_X1 U14932 ( .A1(n15024), .A2(b_7_), .ZN(n15023) );
  NOR2_X1 U14933 ( .A1(n15025), .A2(n8495), .ZN(n15024) );
  NOR2_X1 U14934 ( .A1(n14909), .A2(n14910), .ZN(n15025) );
  NAND2_X1 U14935 ( .A1(n14909), .A2(n14910), .ZN(n15022) );
  NAND2_X1 U14936 ( .A1(n15026), .A2(n15027), .ZN(n14910) );
  NAND2_X1 U14937 ( .A1(n15028), .A2(b_7_), .ZN(n15027) );
  NOR2_X1 U14938 ( .A1(n15029), .A2(n8953), .ZN(n15028) );
  NOR2_X1 U14939 ( .A1(n14906), .A2(n14905), .ZN(n15029) );
  NAND2_X1 U14940 ( .A1(n14905), .A2(n14906), .ZN(n15026) );
  NAND2_X1 U14941 ( .A1(n15030), .A2(n15031), .ZN(n14906) );
  NAND2_X1 U14942 ( .A1(n15032), .A2(b_7_), .ZN(n15031) );
  NOR2_X1 U14943 ( .A1(n15033), .A2(n8440), .ZN(n15032) );
  NOR2_X1 U14944 ( .A1(n14901), .A2(n14902), .ZN(n15033) );
  NAND2_X1 U14945 ( .A1(n14901), .A2(n14902), .ZN(n15030) );
  NAND2_X1 U14946 ( .A1(n15034), .A2(n15035), .ZN(n14902) );
  NAND2_X1 U14947 ( .A1(n15036), .A2(b_7_), .ZN(n15035) );
  NOR2_X1 U14948 ( .A1(n15037), .A2(n8950), .ZN(n15036) );
  NOR2_X1 U14949 ( .A1(n14898), .A2(n14897), .ZN(n15037) );
  NAND2_X1 U14950 ( .A1(n14897), .A2(n14898), .ZN(n15034) );
  NAND2_X1 U14951 ( .A1(n15038), .A2(n15039), .ZN(n14898) );
  NAND2_X1 U14952 ( .A1(n15040), .A2(b_7_), .ZN(n15039) );
  NOR2_X1 U14953 ( .A1(n15041), .A2(n8385), .ZN(n15040) );
  NOR2_X1 U14954 ( .A1(n14792), .A2(n14794), .ZN(n15041) );
  NAND2_X1 U14955 ( .A1(n14792), .A2(n14794), .ZN(n15038) );
  NAND2_X1 U14956 ( .A1(n15042), .A2(n15043), .ZN(n14794) );
  NAND2_X1 U14957 ( .A1(n15044), .A2(b_7_), .ZN(n15043) );
  NOR2_X1 U14958 ( .A1(n15045), .A2(n8947), .ZN(n15044) );
  NOR2_X1 U14959 ( .A1(n14801), .A2(n14799), .ZN(n15045) );
  NAND2_X1 U14960 ( .A1(n14799), .A2(n14801), .ZN(n15042) );
  NAND2_X1 U14961 ( .A1(n15046), .A2(n15047), .ZN(n14801) );
  NAND2_X1 U14962 ( .A1(n15048), .A2(b_7_), .ZN(n15047) );
  NOR2_X1 U14963 ( .A1(n15049), .A2(n8324), .ZN(n15048) );
  NOR2_X1 U14964 ( .A1(n14892), .A2(n14894), .ZN(n15049) );
  NAND2_X1 U14965 ( .A1(n14892), .A2(n14894), .ZN(n15046) );
  NAND2_X1 U14966 ( .A1(n15050), .A2(n15051), .ZN(n14894) );
  NAND2_X1 U14967 ( .A1(n15052), .A2(b_7_), .ZN(n15051) );
  NOR2_X1 U14968 ( .A1(n15053), .A2(n8944), .ZN(n15052) );
  NOR2_X1 U14969 ( .A1(n14888), .A2(n14890), .ZN(n15053) );
  NAND2_X1 U14970 ( .A1(n14888), .A2(n14890), .ZN(n15050) );
  NAND2_X1 U14971 ( .A1(n15054), .A2(n15055), .ZN(n14890) );
  NAND2_X1 U14972 ( .A1(n15056), .A2(b_7_), .ZN(n15055) );
  NOR2_X1 U14973 ( .A1(n15057), .A2(n8268), .ZN(n15056) );
  NOR2_X1 U14974 ( .A1(n14886), .A2(n14885), .ZN(n15057) );
  NAND2_X1 U14975 ( .A1(n14885), .A2(n14886), .ZN(n15054) );
  NAND2_X1 U14976 ( .A1(n14882), .A2(n15058), .ZN(n14886) );
  NAND2_X1 U14977 ( .A1(n14881), .A2(n14883), .ZN(n15058) );
  NAND2_X1 U14978 ( .A1(n15059), .A2(n15060), .ZN(n14883) );
  NAND2_X1 U14979 ( .A1(b_7_), .A2(a_22_), .ZN(n15060) );
  INV_X1 U14980 ( .A(n15061), .ZN(n15059) );
  XOR2_X1 U14981 ( .A(n15062), .B(n15063), .Z(n14881) );
  XNOR2_X1 U14982 ( .A(n15064), .B(n15065), .ZN(n15062) );
  NAND2_X1 U14983 ( .A1(b_6_), .A2(a_23_), .ZN(n15064) );
  NAND2_X1 U14984 ( .A1(a_22_), .A2(n15061), .ZN(n14882) );
  NAND2_X1 U14985 ( .A1(n15066), .A2(n15067), .ZN(n15061) );
  NAND2_X1 U14986 ( .A1(n15068), .A2(b_7_), .ZN(n15067) );
  NOR2_X1 U14987 ( .A1(n15069), .A2(n8213), .ZN(n15068) );
  NOR2_X1 U14988 ( .A1(n14878), .A2(n14877), .ZN(n15069) );
  NAND2_X1 U14989 ( .A1(n14877), .A2(n14878), .ZN(n15066) );
  NAND2_X1 U14990 ( .A1(n15070), .A2(n15071), .ZN(n14878) );
  NAND2_X1 U14991 ( .A1(n14875), .A2(n15072), .ZN(n15071) );
  OR2_X1 U14992 ( .A1(n14873), .A2(n14874), .ZN(n15072) );
  NOR2_X1 U14993 ( .A1(n8667), .A2(n8939), .ZN(n14875) );
  NAND2_X1 U14994 ( .A1(n14873), .A2(n14874), .ZN(n15070) );
  NAND2_X1 U14995 ( .A1(n15073), .A2(n15074), .ZN(n14874) );
  NAND2_X1 U14996 ( .A1(n14871), .A2(n15075), .ZN(n15074) );
  OR2_X1 U14997 ( .A1(n14868), .A2(n14870), .ZN(n15075) );
  NOR2_X1 U14998 ( .A1(n8667), .A2(n8158), .ZN(n14871) );
  NAND2_X1 U14999 ( .A1(n14868), .A2(n14870), .ZN(n15073) );
  NAND2_X1 U15000 ( .A1(n14866), .A2(n15076), .ZN(n14870) );
  NAND2_X1 U15001 ( .A1(n14865), .A2(n14867), .ZN(n15076) );
  NAND2_X1 U15002 ( .A1(n15077), .A2(n15078), .ZN(n14867) );
  NAND2_X1 U15003 ( .A1(b_7_), .A2(a_26_), .ZN(n15078) );
  INV_X1 U15004 ( .A(n15079), .ZN(n15077) );
  XNOR2_X1 U15005 ( .A(n15080), .B(n15081), .ZN(n14865) );
  NAND2_X1 U15006 ( .A1(n15082), .A2(n15083), .ZN(n15080) );
  NAND2_X1 U15007 ( .A1(a_26_), .A2(n15079), .ZN(n14866) );
  NAND2_X1 U15008 ( .A1(n14836), .A2(n15084), .ZN(n15079) );
  NAND2_X1 U15009 ( .A1(n14835), .A2(n14837), .ZN(n15084) );
  NAND2_X1 U15010 ( .A1(n15085), .A2(n15086), .ZN(n14837) );
  NAND2_X1 U15011 ( .A1(b_7_), .A2(a_27_), .ZN(n15086) );
  INV_X1 U15012 ( .A(n15087), .ZN(n15085) );
  XOR2_X1 U15013 ( .A(n15088), .B(n15089), .Z(n14835) );
  XNOR2_X1 U15014 ( .A(n15090), .B(n15091), .ZN(n15088) );
  NAND2_X1 U15015 ( .A1(b_6_), .A2(a_28_), .ZN(n15090) );
  NAND2_X1 U15016 ( .A1(a_27_), .A2(n15087), .ZN(n14836) );
  NAND2_X1 U15017 ( .A1(n15092), .A2(n15093), .ZN(n15087) );
  NAND2_X1 U15018 ( .A1(n15094), .A2(b_7_), .ZN(n15093) );
  NOR2_X1 U15019 ( .A1(n15095), .A2(n8055), .ZN(n15094) );
  NOR2_X1 U15020 ( .A1(n14843), .A2(n14845), .ZN(n15095) );
  NAND2_X1 U15021 ( .A1(n14843), .A2(n14845), .ZN(n15092) );
  NAND2_X1 U15022 ( .A1(n15096), .A2(n15097), .ZN(n14845) );
  NAND2_X1 U15023 ( .A1(n14861), .A2(n15098), .ZN(n15097) );
  OR2_X1 U15024 ( .A1(n14862), .A2(n14863), .ZN(n15098) );
  NOR2_X1 U15025 ( .A1(n8667), .A2(n8041), .ZN(n14861) );
  NAND2_X1 U15026 ( .A1(n14863), .A2(n14862), .ZN(n15096) );
  NAND2_X1 U15027 ( .A1(n15099), .A2(n15100), .ZN(n14862) );
  NAND2_X1 U15028 ( .A1(b_5_), .A2(n15101), .ZN(n15100) );
  NAND2_X1 U15029 ( .A1(n8003), .A2(n15102), .ZN(n15101) );
  NAND2_X1 U15030 ( .A1(a_31_), .A2(n8963), .ZN(n15102) );
  NAND2_X1 U15031 ( .A1(b_6_), .A2(n15103), .ZN(n15099) );
  NAND2_X1 U15032 ( .A1(n9341), .A2(n15104), .ZN(n15103) );
  NAND2_X1 U15033 ( .A1(a_30_), .A2(n8964), .ZN(n15104) );
  AND2_X1 U15034 ( .A1(n15105), .A2(n7953), .ZN(n14863) );
  NOR2_X1 U15035 ( .A1(n8667), .A2(n8963), .ZN(n15105) );
  XOR2_X1 U15036 ( .A(n15106), .B(n15107), .Z(n14843) );
  XOR2_X1 U15037 ( .A(n15108), .B(n15109), .Z(n15106) );
  XNOR2_X1 U15038 ( .A(n15110), .B(n15111), .ZN(n14868) );
  NAND2_X1 U15039 ( .A1(n15112), .A2(n15113), .ZN(n15110) );
  XNOR2_X1 U15040 ( .A(n15114), .B(n15115), .ZN(n14873) );
  NAND2_X1 U15041 ( .A1(n15116), .A2(n15117), .ZN(n15114) );
  XNOR2_X1 U15042 ( .A(n15118), .B(n15119), .ZN(n14877) );
  XNOR2_X1 U15043 ( .A(n15120), .B(n15121), .ZN(n15118) );
  XNOR2_X1 U15044 ( .A(n15122), .B(n15123), .ZN(n14885) );
  NAND2_X1 U15045 ( .A1(n15124), .A2(n15125), .ZN(n15122) );
  XNOR2_X1 U15046 ( .A(n15126), .B(n15127), .ZN(n14888) );
  XNOR2_X1 U15047 ( .A(n15128), .B(n15129), .ZN(n15127) );
  XOR2_X1 U15048 ( .A(n15130), .B(n15131), .Z(n14892) );
  XOR2_X1 U15049 ( .A(n15132), .B(n15133), .Z(n15130) );
  NOR2_X1 U15050 ( .A1(n8944), .A2(n8963), .ZN(n15133) );
  XNOR2_X1 U15051 ( .A(n15134), .B(n15135), .ZN(n14799) );
  XNOR2_X1 U15052 ( .A(n15136), .B(n15137), .ZN(n15134) );
  XOR2_X1 U15053 ( .A(n15138), .B(n15139), .Z(n14792) );
  XOR2_X1 U15054 ( .A(n15140), .B(n15141), .Z(n15138) );
  XNOR2_X1 U15055 ( .A(n15142), .B(n15143), .ZN(n14897) );
  XNOR2_X1 U15056 ( .A(n15144), .B(n15145), .ZN(n15143) );
  XNOR2_X1 U15057 ( .A(n15146), .B(n15147), .ZN(n14901) );
  XNOR2_X1 U15058 ( .A(n15148), .B(n15149), .ZN(n15147) );
  XNOR2_X1 U15059 ( .A(n15150), .B(n15151), .ZN(n14905) );
  XNOR2_X1 U15060 ( .A(n15152), .B(n15153), .ZN(n15151) );
  XNOR2_X1 U15061 ( .A(n15154), .B(n15155), .ZN(n14909) );
  XNOR2_X1 U15062 ( .A(n15156), .B(n15157), .ZN(n15155) );
  XNOR2_X1 U15063 ( .A(n15158), .B(n15159), .ZN(n14913) );
  XNOR2_X1 U15064 ( .A(n15160), .B(n15161), .ZN(n15159) );
  XNOR2_X1 U15065 ( .A(n15162), .B(n15163), .ZN(n14917) );
  XNOR2_X1 U15066 ( .A(n15164), .B(n15165), .ZN(n15163) );
  XNOR2_X1 U15067 ( .A(n15166), .B(n15167), .ZN(n14921) );
  XNOR2_X1 U15068 ( .A(n15168), .B(n15169), .ZN(n15167) );
  XNOR2_X1 U15069 ( .A(n15170), .B(n15171), .ZN(n14925) );
  XNOR2_X1 U15070 ( .A(n15172), .B(n15173), .ZN(n15171) );
  XNOR2_X1 U15071 ( .A(n15174), .B(n15175), .ZN(n14929) );
  XOR2_X1 U15072 ( .A(n15176), .B(n15177), .Z(n15175) );
  NAND2_X1 U15073 ( .A1(b_6_), .A2(a_9_), .ZN(n15177) );
  INV_X1 U15074 ( .A(n8877), .ZN(n14935) );
  NAND2_X1 U15075 ( .A1(b_7_), .A2(a_7_), .ZN(n8877) );
  XOR2_X1 U15076 ( .A(n15178), .B(n15179), .Z(n14937) );
  XOR2_X1 U15077 ( .A(n15180), .B(n15181), .Z(n15178) );
  NOR2_X1 U15078 ( .A1(n8962), .A2(n8963), .ZN(n15181) );
  XOR2_X1 U15079 ( .A(n15182), .B(n15183), .Z(n14941) );
  XOR2_X1 U15080 ( .A(n15184), .B(n15185), .Z(n15182) );
  XOR2_X1 U15081 ( .A(n15186), .B(n15187), .Z(n14945) );
  XOR2_X1 U15082 ( .A(n15188), .B(n15189), .Z(n15186) );
  NOR2_X1 U15083 ( .A1(n8723), .A2(n8963), .ZN(n15189) );
  XOR2_X1 U15084 ( .A(n15190), .B(n15191), .Z(n14949) );
  XOR2_X1 U15085 ( .A(n15192), .B(n15193), .Z(n15190) );
  NOR2_X1 U15086 ( .A1(n8966), .A2(n8963), .ZN(n15193) );
  XOR2_X1 U15087 ( .A(n15194), .B(n15195), .Z(n14953) );
  XOR2_X1 U15088 ( .A(n15196), .B(n15197), .Z(n15194) );
  NOR2_X1 U15089 ( .A1(n8778), .A2(n8963), .ZN(n15197) );
  XNOR2_X1 U15090 ( .A(n15198), .B(n15199), .ZN(n14956) );
  XOR2_X1 U15091 ( .A(n15200), .B(n15201), .Z(n15199) );
  NAND2_X1 U15092 ( .A1(b_6_), .A2(a_2_), .ZN(n15201) );
  XOR2_X1 U15093 ( .A(n15202), .B(n15203), .Z(n14960) );
  XOR2_X1 U15094 ( .A(n15204), .B(n15205), .Z(n15202) );
  NOR2_X1 U15095 ( .A1(n8969), .A2(n8963), .ZN(n15205) );
  XNOR2_X1 U15096 ( .A(n14729), .B(n14728), .ZN(n14967) );
  XNOR2_X1 U15097 ( .A(n15206), .B(n15207), .ZN(n14729) );
  NOR2_X1 U15098 ( .A1(n8974), .A2(n8963), .ZN(n15207) );
  NAND2_X1 U15099 ( .A1(n15208), .A2(n15209), .ZN(n8081) );
  OR2_X1 U15100 ( .A1(n15209), .A2(n15208), .ZN(n8080) );
  NAND2_X1 U15101 ( .A1(n15210), .A2(n15211), .ZN(n15208) );
  NAND2_X1 U15102 ( .A1(n15212), .A2(n15213), .ZN(n15211) );
  XOR2_X1 U15103 ( .A(n15214), .B(n15215), .Z(n15213) );
  INV_X1 U15104 ( .A(n15216), .ZN(n15212) );
  NAND2_X1 U15105 ( .A1(n14966), .A2(n14965), .ZN(n15209) );
  NAND2_X1 U15106 ( .A1(n15217), .A2(n15218), .ZN(n14965) );
  NAND2_X1 U15107 ( .A1(n15219), .A2(b_6_), .ZN(n15218) );
  NOR2_X1 U15108 ( .A1(n15220), .A2(n8974), .ZN(n15219) );
  NOR2_X1 U15109 ( .A1(n15206), .A2(n14728), .ZN(n15220) );
  NAND2_X1 U15110 ( .A1(n14728), .A2(n15206), .ZN(n15217) );
  NAND2_X1 U15111 ( .A1(n15221), .A2(n15222), .ZN(n15206) );
  NAND2_X1 U15112 ( .A1(n15223), .A2(b_6_), .ZN(n15222) );
  NOR2_X1 U15113 ( .A1(n15224), .A2(n8969), .ZN(n15223) );
  NOR2_X1 U15114 ( .A1(n15203), .A2(n15204), .ZN(n15224) );
  NAND2_X1 U15115 ( .A1(n15203), .A2(n15204), .ZN(n15221) );
  NAND2_X1 U15116 ( .A1(n15225), .A2(n15226), .ZN(n15204) );
  NAND2_X1 U15117 ( .A1(n15227), .A2(b_6_), .ZN(n15226) );
  NOR2_X1 U15118 ( .A1(n15228), .A2(n8792), .ZN(n15227) );
  NOR2_X1 U15119 ( .A1(n15198), .A2(n15200), .ZN(n15228) );
  NAND2_X1 U15120 ( .A1(n15198), .A2(n15200), .ZN(n15225) );
  NAND2_X1 U15121 ( .A1(n15229), .A2(n15230), .ZN(n15200) );
  NAND2_X1 U15122 ( .A1(n15231), .A2(b_6_), .ZN(n15230) );
  NOR2_X1 U15123 ( .A1(n15232), .A2(n8778), .ZN(n15231) );
  NOR2_X1 U15124 ( .A1(n15195), .A2(n15196), .ZN(n15232) );
  NAND2_X1 U15125 ( .A1(n15195), .A2(n15196), .ZN(n15229) );
  NAND2_X1 U15126 ( .A1(n15233), .A2(n15234), .ZN(n15196) );
  NAND2_X1 U15127 ( .A1(n15235), .A2(b_6_), .ZN(n15234) );
  NOR2_X1 U15128 ( .A1(n15236), .A2(n8966), .ZN(n15235) );
  NOR2_X1 U15129 ( .A1(n15191), .A2(n15192), .ZN(n15236) );
  NAND2_X1 U15130 ( .A1(n15191), .A2(n15192), .ZN(n15233) );
  NAND2_X1 U15131 ( .A1(n15237), .A2(n15238), .ZN(n15192) );
  NAND2_X1 U15132 ( .A1(n15239), .A2(b_6_), .ZN(n15238) );
  NOR2_X1 U15133 ( .A1(n15240), .A2(n8723), .ZN(n15239) );
  NOR2_X1 U15134 ( .A1(n15187), .A2(n15188), .ZN(n15240) );
  NAND2_X1 U15135 ( .A1(n15187), .A2(n15188), .ZN(n15237) );
  NAND2_X1 U15136 ( .A1(n15241), .A2(n15242), .ZN(n15188) );
  NAND2_X1 U15137 ( .A1(n15183), .A2(n15243), .ZN(n15242) );
  OR2_X1 U15138 ( .A1(n15184), .A2(n15185), .ZN(n15243) );
  XOR2_X1 U15139 ( .A(n15244), .B(n15245), .Z(n15183) );
  XOR2_X1 U15140 ( .A(n15246), .B(n15247), .Z(n15244) );
  NOR2_X1 U15141 ( .A1(n8962), .A2(n8964), .ZN(n15247) );
  NAND2_X1 U15142 ( .A1(n15185), .A2(n15184), .ZN(n15241) );
  NAND2_X1 U15143 ( .A1(n15248), .A2(n15249), .ZN(n15184) );
  NAND2_X1 U15144 ( .A1(n15250), .A2(b_6_), .ZN(n15249) );
  NOR2_X1 U15145 ( .A1(n15251), .A2(n8962), .ZN(n15250) );
  NOR2_X1 U15146 ( .A1(n15179), .A2(n15180), .ZN(n15251) );
  NAND2_X1 U15147 ( .A1(n15179), .A2(n15180), .ZN(n15248) );
  NAND2_X1 U15148 ( .A1(n15252), .A2(n15253), .ZN(n15180) );
  NAND2_X1 U15149 ( .A1(n15254), .A2(b_6_), .ZN(n15253) );
  NOR2_X1 U15150 ( .A1(n15255), .A2(n8619), .ZN(n15254) );
  NOR2_X1 U15151 ( .A1(n14999), .A2(n15000), .ZN(n15255) );
  NAND2_X1 U15152 ( .A1(n14999), .A2(n15000), .ZN(n15252) );
  NAND2_X1 U15153 ( .A1(n15256), .A2(n15257), .ZN(n15000) );
  NAND2_X1 U15154 ( .A1(n15258), .A2(b_6_), .ZN(n15257) );
  NOR2_X1 U15155 ( .A1(n15259), .A2(n8605), .ZN(n15258) );
  NOR2_X1 U15156 ( .A1(n15174), .A2(n15176), .ZN(n15259) );
  NAND2_X1 U15157 ( .A1(n15174), .A2(n15176), .ZN(n15256) );
  NAND2_X1 U15158 ( .A1(n15260), .A2(n15261), .ZN(n15176) );
  NAND2_X1 U15159 ( .A1(n15173), .A2(n15262), .ZN(n15261) );
  OR2_X1 U15160 ( .A1(n15172), .A2(n15170), .ZN(n15262) );
  NOR2_X1 U15161 ( .A1(n8963), .A2(n8959), .ZN(n15173) );
  NAND2_X1 U15162 ( .A1(n15170), .A2(n15172), .ZN(n15260) );
  NAND2_X1 U15163 ( .A1(n15263), .A2(n15264), .ZN(n15172) );
  NAND2_X1 U15164 ( .A1(n15169), .A2(n15265), .ZN(n15264) );
  OR2_X1 U15165 ( .A1(n15168), .A2(n15166), .ZN(n15265) );
  NOR2_X1 U15166 ( .A1(n8963), .A2(n8550), .ZN(n15169) );
  NAND2_X1 U15167 ( .A1(n15166), .A2(n15168), .ZN(n15263) );
  NAND2_X1 U15168 ( .A1(n15266), .A2(n15267), .ZN(n15168) );
  NAND2_X1 U15169 ( .A1(n15165), .A2(n15268), .ZN(n15267) );
  OR2_X1 U15170 ( .A1(n15164), .A2(n15162), .ZN(n15268) );
  NOR2_X1 U15171 ( .A1(n8963), .A2(n8956), .ZN(n15165) );
  NAND2_X1 U15172 ( .A1(n15162), .A2(n15164), .ZN(n15266) );
  NAND2_X1 U15173 ( .A1(n15269), .A2(n15270), .ZN(n15164) );
  NAND2_X1 U15174 ( .A1(n15161), .A2(n15271), .ZN(n15270) );
  OR2_X1 U15175 ( .A1(n15160), .A2(n15158), .ZN(n15271) );
  NOR2_X1 U15176 ( .A1(n8963), .A2(n8495), .ZN(n15161) );
  NAND2_X1 U15177 ( .A1(n15158), .A2(n15160), .ZN(n15269) );
  NAND2_X1 U15178 ( .A1(n15272), .A2(n15273), .ZN(n15160) );
  NAND2_X1 U15179 ( .A1(n15157), .A2(n15274), .ZN(n15273) );
  OR2_X1 U15180 ( .A1(n15154), .A2(n15156), .ZN(n15274) );
  NOR2_X1 U15181 ( .A1(n8963), .A2(n8953), .ZN(n15157) );
  NAND2_X1 U15182 ( .A1(n15154), .A2(n15156), .ZN(n15272) );
  NAND2_X1 U15183 ( .A1(n15275), .A2(n15276), .ZN(n15156) );
  NAND2_X1 U15184 ( .A1(n15153), .A2(n15277), .ZN(n15276) );
  OR2_X1 U15185 ( .A1(n15152), .A2(n15150), .ZN(n15277) );
  NOR2_X1 U15186 ( .A1(n8963), .A2(n8440), .ZN(n15153) );
  NAND2_X1 U15187 ( .A1(n15150), .A2(n15152), .ZN(n15275) );
  NAND2_X1 U15188 ( .A1(n15278), .A2(n15279), .ZN(n15152) );
  NAND2_X1 U15189 ( .A1(n15149), .A2(n15280), .ZN(n15279) );
  OR2_X1 U15190 ( .A1(n15146), .A2(n15148), .ZN(n15280) );
  NOR2_X1 U15191 ( .A1(n8963), .A2(n8950), .ZN(n15149) );
  NAND2_X1 U15192 ( .A1(n15146), .A2(n15148), .ZN(n15278) );
  NAND2_X1 U15193 ( .A1(n15281), .A2(n15282), .ZN(n15148) );
  NAND2_X1 U15194 ( .A1(n15145), .A2(n15283), .ZN(n15282) );
  OR2_X1 U15195 ( .A1(n15144), .A2(n15142), .ZN(n15283) );
  NOR2_X1 U15196 ( .A1(n8963), .A2(n8385), .ZN(n15145) );
  NAND2_X1 U15197 ( .A1(n15142), .A2(n15144), .ZN(n15281) );
  NAND2_X1 U15198 ( .A1(n15284), .A2(n15285), .ZN(n15144) );
  NAND2_X1 U15199 ( .A1(n15141), .A2(n15286), .ZN(n15285) );
  OR2_X1 U15200 ( .A1(n15139), .A2(n15140), .ZN(n15286) );
  NOR2_X1 U15201 ( .A1(n8963), .A2(n8947), .ZN(n15141) );
  NAND2_X1 U15202 ( .A1(n15139), .A2(n15140), .ZN(n15284) );
  NAND2_X1 U15203 ( .A1(n15287), .A2(n15288), .ZN(n15140) );
  NAND2_X1 U15204 ( .A1(n15137), .A2(n15289), .ZN(n15288) );
  NAND2_X1 U15205 ( .A1(n15136), .A2(n15135), .ZN(n15289) );
  NOR2_X1 U15206 ( .A1(n8963), .A2(n8324), .ZN(n15137) );
  OR2_X1 U15207 ( .A1(n15135), .A2(n15136), .ZN(n15287) );
  AND2_X1 U15208 ( .A1(n15290), .A2(n15291), .ZN(n15136) );
  NAND2_X1 U15209 ( .A1(n15292), .A2(b_6_), .ZN(n15291) );
  NOR2_X1 U15210 ( .A1(n15293), .A2(n8944), .ZN(n15292) );
  NOR2_X1 U15211 ( .A1(n15132), .A2(n15131), .ZN(n15293) );
  NAND2_X1 U15212 ( .A1(n15131), .A2(n15132), .ZN(n15290) );
  NAND2_X1 U15213 ( .A1(n15294), .A2(n15295), .ZN(n15132) );
  NAND2_X1 U15214 ( .A1(n15129), .A2(n15296), .ZN(n15295) );
  OR2_X1 U15215 ( .A1(n15126), .A2(n15128), .ZN(n15296) );
  NOR2_X1 U15216 ( .A1(n8963), .A2(n8268), .ZN(n15129) );
  NAND2_X1 U15217 ( .A1(n15126), .A2(n15128), .ZN(n15294) );
  NAND2_X1 U15218 ( .A1(n15124), .A2(n15297), .ZN(n15128) );
  NAND2_X1 U15219 ( .A1(n15123), .A2(n15125), .ZN(n15297) );
  NAND2_X1 U15220 ( .A1(n15298), .A2(n15299), .ZN(n15125) );
  NAND2_X1 U15221 ( .A1(b_6_), .A2(a_22_), .ZN(n15299) );
  INV_X1 U15222 ( .A(n15300), .ZN(n15298) );
  XNOR2_X1 U15223 ( .A(n15301), .B(n15302), .ZN(n15123) );
  XOR2_X1 U15224 ( .A(n15303), .B(n15304), .Z(n15302) );
  NAND2_X1 U15225 ( .A1(b_5_), .A2(a_23_), .ZN(n15304) );
  NAND2_X1 U15226 ( .A1(a_22_), .A2(n15300), .ZN(n15124) );
  NAND2_X1 U15227 ( .A1(n15305), .A2(n15306), .ZN(n15300) );
  NAND2_X1 U15228 ( .A1(n15307), .A2(b_6_), .ZN(n15306) );
  NOR2_X1 U15229 ( .A1(n15308), .A2(n8213), .ZN(n15307) );
  NOR2_X1 U15230 ( .A1(n15065), .A2(n15063), .ZN(n15308) );
  NAND2_X1 U15231 ( .A1(n15063), .A2(n15065), .ZN(n15305) );
  NAND2_X1 U15232 ( .A1(n15309), .A2(n15310), .ZN(n15065) );
  NAND2_X1 U15233 ( .A1(n15121), .A2(n15311), .ZN(n15310) );
  NAND2_X1 U15234 ( .A1(n15120), .A2(n15119), .ZN(n15311) );
  NOR2_X1 U15235 ( .A1(n8963), .A2(n8939), .ZN(n15121) );
  OR2_X1 U15236 ( .A1(n15119), .A2(n15120), .ZN(n15309) );
  AND2_X1 U15237 ( .A1(n15116), .A2(n15312), .ZN(n15120) );
  NAND2_X1 U15238 ( .A1(n15115), .A2(n15117), .ZN(n15312) );
  NAND2_X1 U15239 ( .A1(n15313), .A2(n15314), .ZN(n15117) );
  NAND2_X1 U15240 ( .A1(b_6_), .A2(a_25_), .ZN(n15314) );
  INV_X1 U15241 ( .A(n15315), .ZN(n15313) );
  XNOR2_X1 U15242 ( .A(n15316), .B(n15317), .ZN(n15115) );
  NAND2_X1 U15243 ( .A1(n15318), .A2(n15319), .ZN(n15316) );
  NAND2_X1 U15244 ( .A1(a_25_), .A2(n15315), .ZN(n15116) );
  NAND2_X1 U15245 ( .A1(n15112), .A2(n15320), .ZN(n15315) );
  NAND2_X1 U15246 ( .A1(n15111), .A2(n15113), .ZN(n15320) );
  NAND2_X1 U15247 ( .A1(n15321), .A2(n15322), .ZN(n15113) );
  NAND2_X1 U15248 ( .A1(b_6_), .A2(a_26_), .ZN(n15322) );
  INV_X1 U15249 ( .A(n15323), .ZN(n15321) );
  XNOR2_X1 U15250 ( .A(n15324), .B(n15325), .ZN(n15111) );
  NAND2_X1 U15251 ( .A1(n15326), .A2(n15327), .ZN(n15324) );
  NAND2_X1 U15252 ( .A1(a_26_), .A2(n15323), .ZN(n15112) );
  NAND2_X1 U15253 ( .A1(n15082), .A2(n15328), .ZN(n15323) );
  NAND2_X1 U15254 ( .A1(n15081), .A2(n15083), .ZN(n15328) );
  NAND2_X1 U15255 ( .A1(n15329), .A2(n15330), .ZN(n15083) );
  NAND2_X1 U15256 ( .A1(b_6_), .A2(a_27_), .ZN(n15330) );
  INV_X1 U15257 ( .A(n15331), .ZN(n15329) );
  XOR2_X1 U15258 ( .A(n15332), .B(n15333), .Z(n15081) );
  XNOR2_X1 U15259 ( .A(n15334), .B(n15335), .ZN(n15332) );
  NAND2_X1 U15260 ( .A1(b_5_), .A2(a_28_), .ZN(n15334) );
  NAND2_X1 U15261 ( .A1(a_27_), .A2(n15331), .ZN(n15082) );
  NAND2_X1 U15262 ( .A1(n15336), .A2(n15337), .ZN(n15331) );
  NAND2_X1 U15263 ( .A1(n15338), .A2(b_6_), .ZN(n15337) );
  NOR2_X1 U15264 ( .A1(n15339), .A2(n8055), .ZN(n15338) );
  NOR2_X1 U15265 ( .A1(n15089), .A2(n15091), .ZN(n15339) );
  NAND2_X1 U15266 ( .A1(n15089), .A2(n15091), .ZN(n15336) );
  NAND2_X1 U15267 ( .A1(n15340), .A2(n15341), .ZN(n15091) );
  NAND2_X1 U15268 ( .A1(n15107), .A2(n15342), .ZN(n15341) );
  OR2_X1 U15269 ( .A1(n15108), .A2(n15109), .ZN(n15342) );
  NOR2_X1 U15270 ( .A1(n8963), .A2(n8041), .ZN(n15107) );
  NAND2_X1 U15271 ( .A1(n15109), .A2(n15108), .ZN(n15340) );
  NAND2_X1 U15272 ( .A1(n15343), .A2(n15344), .ZN(n15108) );
  NAND2_X1 U15273 ( .A1(b_4_), .A2(n15345), .ZN(n15344) );
  NAND2_X1 U15274 ( .A1(n8003), .A2(n15346), .ZN(n15345) );
  NAND2_X1 U15275 ( .A1(a_31_), .A2(n8964), .ZN(n15346) );
  NAND2_X1 U15276 ( .A1(b_5_), .A2(n15347), .ZN(n15343) );
  NAND2_X1 U15277 ( .A1(n9341), .A2(n15348), .ZN(n15347) );
  NAND2_X1 U15278 ( .A1(a_30_), .A2(n8965), .ZN(n15348) );
  AND2_X1 U15279 ( .A1(n15349), .A2(n7953), .ZN(n15109) );
  NOR2_X1 U15280 ( .A1(n8963), .A2(n8964), .ZN(n15349) );
  XOR2_X1 U15281 ( .A(n15350), .B(n15351), .Z(n15089) );
  XOR2_X1 U15282 ( .A(n15352), .B(n15353), .Z(n15350) );
  XOR2_X1 U15283 ( .A(n15354), .B(n15355), .Z(n15119) );
  NAND2_X1 U15284 ( .A1(n15356), .A2(n15357), .ZN(n15354) );
  XOR2_X1 U15285 ( .A(n15358), .B(n15359), .Z(n15063) );
  XOR2_X1 U15286 ( .A(n15360), .B(n15361), .Z(n15358) );
  NOR2_X1 U15287 ( .A1(n8939), .A2(n8964), .ZN(n15361) );
  XNOR2_X1 U15288 ( .A(n15362), .B(n15363), .ZN(n15126) );
  XOR2_X1 U15289 ( .A(n15364), .B(n15365), .Z(n15363) );
  NAND2_X1 U15290 ( .A1(b_5_), .A2(a_22_), .ZN(n15365) );
  XOR2_X1 U15291 ( .A(n15366), .B(n15367), .Z(n15131) );
  XOR2_X1 U15292 ( .A(n15368), .B(n15369), .Z(n15366) );
  NOR2_X1 U15293 ( .A1(n8268), .A2(n8964), .ZN(n15369) );
  XNOR2_X1 U15294 ( .A(n15370), .B(n15371), .ZN(n15135) );
  XOR2_X1 U15295 ( .A(n15372), .B(n15373), .Z(n15370) );
  NOR2_X1 U15296 ( .A1(n8944), .A2(n8964), .ZN(n15373) );
  XOR2_X1 U15297 ( .A(n15374), .B(n15375), .Z(n15139) );
  XOR2_X1 U15298 ( .A(n15376), .B(n15377), .Z(n15374) );
  NOR2_X1 U15299 ( .A1(n8324), .A2(n8964), .ZN(n15377) );
  XOR2_X1 U15300 ( .A(n15378), .B(n15379), .Z(n15142) );
  XOR2_X1 U15301 ( .A(n15380), .B(n15381), .Z(n15378) );
  NOR2_X1 U15302 ( .A1(n8947), .A2(n8964), .ZN(n15381) );
  XOR2_X1 U15303 ( .A(n15382), .B(n15383), .Z(n15146) );
  XOR2_X1 U15304 ( .A(n15384), .B(n15385), .Z(n15382) );
  NOR2_X1 U15305 ( .A1(n8385), .A2(n8964), .ZN(n15385) );
  XOR2_X1 U15306 ( .A(n15386), .B(n15387), .Z(n15150) );
  XOR2_X1 U15307 ( .A(n15388), .B(n15389), .Z(n15386) );
  NOR2_X1 U15308 ( .A1(n8950), .A2(n8964), .ZN(n15389) );
  XOR2_X1 U15309 ( .A(n15390), .B(n15391), .Z(n15154) );
  XOR2_X1 U15310 ( .A(n15392), .B(n15393), .Z(n15390) );
  NOR2_X1 U15311 ( .A1(n8440), .A2(n8964), .ZN(n15393) );
  XOR2_X1 U15312 ( .A(n15394), .B(n15395), .Z(n15158) );
  XOR2_X1 U15313 ( .A(n15396), .B(n15397), .Z(n15394) );
  NOR2_X1 U15314 ( .A1(n8953), .A2(n8964), .ZN(n15397) );
  XOR2_X1 U15315 ( .A(n15398), .B(n15399), .Z(n15162) );
  XOR2_X1 U15316 ( .A(n15400), .B(n15401), .Z(n15398) );
  NOR2_X1 U15317 ( .A1(n8495), .A2(n8964), .ZN(n15401) );
  XOR2_X1 U15318 ( .A(n15402), .B(n15403), .Z(n15166) );
  XOR2_X1 U15319 ( .A(n15404), .B(n15405), .Z(n15402) );
  NOR2_X1 U15320 ( .A1(n8956), .A2(n8964), .ZN(n15405) );
  XOR2_X1 U15321 ( .A(n15406), .B(n15407), .Z(n15170) );
  XOR2_X1 U15322 ( .A(n15408), .B(n15409), .Z(n15406) );
  NOR2_X1 U15323 ( .A1(n8550), .A2(n8964), .ZN(n15409) );
  XOR2_X1 U15324 ( .A(n15410), .B(n15411), .Z(n15174) );
  XOR2_X1 U15325 ( .A(n15412), .B(n15413), .Z(n15410) );
  NOR2_X1 U15326 ( .A1(n8959), .A2(n8964), .ZN(n15413) );
  XOR2_X1 U15327 ( .A(n15414), .B(n15415), .Z(n14999) );
  XOR2_X1 U15328 ( .A(n15416), .B(n15417), .Z(n15414) );
  NOR2_X1 U15329 ( .A1(n8605), .A2(n8964), .ZN(n15417) );
  XOR2_X1 U15330 ( .A(n15418), .B(n15419), .Z(n15179) );
  XOR2_X1 U15331 ( .A(n15420), .B(n15421), .Z(n15418) );
  NOR2_X1 U15332 ( .A1(n8619), .A2(n8964), .ZN(n15421) );
  INV_X1 U15333 ( .A(n8701), .ZN(n15185) );
  NAND2_X1 U15334 ( .A1(b_6_), .A2(a_6_), .ZN(n8701) );
  XOR2_X1 U15335 ( .A(n15422), .B(n15423), .Z(n15187) );
  XOR2_X1 U15336 ( .A(n15424), .B(n15425), .Z(n15422) );
  NOR2_X1 U15337 ( .A1(n8681), .A2(n8964), .ZN(n15425) );
  XOR2_X1 U15338 ( .A(n15426), .B(n15427), .Z(n15191) );
  XOR2_X1 U15339 ( .A(n15428), .B(n15429), .Z(n15426) );
  XOR2_X1 U15340 ( .A(n15430), .B(n15431), .Z(n15195) );
  XNOR2_X1 U15341 ( .A(n15432), .B(n15433), .ZN(n15430) );
  NAND2_X1 U15342 ( .A1(b_5_), .A2(a_4_), .ZN(n15432) );
  XOR2_X1 U15343 ( .A(n15434), .B(n15435), .Z(n15198) );
  XOR2_X1 U15344 ( .A(n15436), .B(n15437), .Z(n15434) );
  NOR2_X1 U15345 ( .A1(n8778), .A2(n8964), .ZN(n15437) );
  XOR2_X1 U15346 ( .A(n15438), .B(n15439), .Z(n15203) );
  XOR2_X1 U15347 ( .A(n15440), .B(n15441), .Z(n15438) );
  NOR2_X1 U15348 ( .A1(n8792), .A2(n8964), .ZN(n15441) );
  XOR2_X1 U15349 ( .A(n15442), .B(n15443), .Z(n14728) );
  XOR2_X1 U15350 ( .A(n15444), .B(n15445), .Z(n15442) );
  NOR2_X1 U15351 ( .A1(n8969), .A2(n8964), .ZN(n15445) );
  XOR2_X1 U15352 ( .A(n15446), .B(n15447), .Z(n14966) );
  XOR2_X1 U15353 ( .A(n15448), .B(n15449), .Z(n15446) );
  NAND2_X1 U15354 ( .A1(n15450), .A2(n15210), .ZN(n8363) );
  OR2_X1 U15355 ( .A1(n15210), .A2(n15450), .ZN(n8364) );
  XNOR2_X1 U15356 ( .A(n15451), .B(n15452), .ZN(n15450) );
  NAND2_X1 U15357 ( .A1(n15453), .A2(n15216), .ZN(n15210) );
  NAND2_X1 U15358 ( .A1(n15454), .A2(n15455), .ZN(n15216) );
  NAND2_X1 U15359 ( .A1(n15449), .A2(n15456), .ZN(n15455) );
  OR2_X1 U15360 ( .A1(n15447), .A2(n15448), .ZN(n15456) );
  NOR2_X1 U15361 ( .A1(n8964), .A2(n8974), .ZN(n15449) );
  NAND2_X1 U15362 ( .A1(n15447), .A2(n15448), .ZN(n15454) );
  NAND2_X1 U15363 ( .A1(n15457), .A2(n15458), .ZN(n15448) );
  NAND2_X1 U15364 ( .A1(n15459), .A2(b_5_), .ZN(n15458) );
  NOR2_X1 U15365 ( .A1(n15460), .A2(n8969), .ZN(n15459) );
  NOR2_X1 U15366 ( .A1(n15443), .A2(n15444), .ZN(n15460) );
  NAND2_X1 U15367 ( .A1(n15443), .A2(n15444), .ZN(n15457) );
  NAND2_X1 U15368 ( .A1(n15461), .A2(n15462), .ZN(n15444) );
  NAND2_X1 U15369 ( .A1(n15463), .A2(b_5_), .ZN(n15462) );
  NOR2_X1 U15370 ( .A1(n15464), .A2(n8792), .ZN(n15463) );
  NOR2_X1 U15371 ( .A1(n15440), .A2(n15439), .ZN(n15464) );
  NAND2_X1 U15372 ( .A1(n15439), .A2(n15440), .ZN(n15461) );
  NAND2_X1 U15373 ( .A1(n15465), .A2(n15466), .ZN(n15440) );
  NAND2_X1 U15374 ( .A1(n15467), .A2(b_5_), .ZN(n15466) );
  NOR2_X1 U15375 ( .A1(n15468), .A2(n8778), .ZN(n15467) );
  NOR2_X1 U15376 ( .A1(n15436), .A2(n15435), .ZN(n15468) );
  NAND2_X1 U15377 ( .A1(n15435), .A2(n15436), .ZN(n15465) );
  NAND2_X1 U15378 ( .A1(n15469), .A2(n15470), .ZN(n15436) );
  NAND2_X1 U15379 ( .A1(n15471), .A2(b_5_), .ZN(n15470) );
  NOR2_X1 U15380 ( .A1(n15472), .A2(n8966), .ZN(n15471) );
  NOR2_X1 U15381 ( .A1(n15433), .A2(n15431), .ZN(n15472) );
  NAND2_X1 U15382 ( .A1(n15431), .A2(n15433), .ZN(n15469) );
  NAND2_X1 U15383 ( .A1(n15473), .A2(n15474), .ZN(n15433) );
  NAND2_X1 U15384 ( .A1(n15427), .A2(n15475), .ZN(n15474) );
  OR2_X1 U15385 ( .A1(n15428), .A2(n15429), .ZN(n15475) );
  XOR2_X1 U15386 ( .A(n15476), .B(n15477), .Z(n15427) );
  XOR2_X1 U15387 ( .A(n15478), .B(n15479), .Z(n15476) );
  NOR2_X1 U15388 ( .A1(n8681), .A2(n8965), .ZN(n15479) );
  NAND2_X1 U15389 ( .A1(n15429), .A2(n15428), .ZN(n15473) );
  NAND2_X1 U15390 ( .A1(n15480), .A2(n15481), .ZN(n15428) );
  NAND2_X1 U15391 ( .A1(n15482), .A2(b_5_), .ZN(n15481) );
  NOR2_X1 U15392 ( .A1(n15483), .A2(n8681), .ZN(n15482) );
  NOR2_X1 U15393 ( .A1(n15424), .A2(n15423), .ZN(n15483) );
  NAND2_X1 U15394 ( .A1(n15423), .A2(n15424), .ZN(n15480) );
  NAND2_X1 U15395 ( .A1(n15484), .A2(n15485), .ZN(n15424) );
  NAND2_X1 U15396 ( .A1(n15486), .A2(b_5_), .ZN(n15485) );
  NOR2_X1 U15397 ( .A1(n15487), .A2(n8962), .ZN(n15486) );
  NOR2_X1 U15398 ( .A1(n15246), .A2(n15245), .ZN(n15487) );
  NAND2_X1 U15399 ( .A1(n15245), .A2(n15246), .ZN(n15484) );
  NAND2_X1 U15400 ( .A1(n15488), .A2(n15489), .ZN(n15246) );
  NAND2_X1 U15401 ( .A1(n15490), .A2(b_5_), .ZN(n15489) );
  NOR2_X1 U15402 ( .A1(n15491), .A2(n8619), .ZN(n15490) );
  NOR2_X1 U15403 ( .A1(n15420), .A2(n15419), .ZN(n15491) );
  NAND2_X1 U15404 ( .A1(n15419), .A2(n15420), .ZN(n15488) );
  NAND2_X1 U15405 ( .A1(n15492), .A2(n15493), .ZN(n15420) );
  NAND2_X1 U15406 ( .A1(n15494), .A2(b_5_), .ZN(n15493) );
  NOR2_X1 U15407 ( .A1(n15495), .A2(n8605), .ZN(n15494) );
  NOR2_X1 U15408 ( .A1(n15416), .A2(n15415), .ZN(n15495) );
  NAND2_X1 U15409 ( .A1(n15415), .A2(n15416), .ZN(n15492) );
  NAND2_X1 U15410 ( .A1(n15496), .A2(n15497), .ZN(n15416) );
  NAND2_X1 U15411 ( .A1(n15498), .A2(b_5_), .ZN(n15497) );
  NOR2_X1 U15412 ( .A1(n15499), .A2(n8959), .ZN(n15498) );
  NOR2_X1 U15413 ( .A1(n15412), .A2(n15411), .ZN(n15499) );
  NAND2_X1 U15414 ( .A1(n15411), .A2(n15412), .ZN(n15496) );
  NAND2_X1 U15415 ( .A1(n15500), .A2(n15501), .ZN(n15412) );
  NAND2_X1 U15416 ( .A1(n15502), .A2(b_5_), .ZN(n15501) );
  NOR2_X1 U15417 ( .A1(n15503), .A2(n8550), .ZN(n15502) );
  NOR2_X1 U15418 ( .A1(n15408), .A2(n15407), .ZN(n15503) );
  NAND2_X1 U15419 ( .A1(n15407), .A2(n15408), .ZN(n15500) );
  NAND2_X1 U15420 ( .A1(n15504), .A2(n15505), .ZN(n15408) );
  NAND2_X1 U15421 ( .A1(n15506), .A2(b_5_), .ZN(n15505) );
  NOR2_X1 U15422 ( .A1(n15507), .A2(n8956), .ZN(n15506) );
  NOR2_X1 U15423 ( .A1(n15404), .A2(n15403), .ZN(n15507) );
  NAND2_X1 U15424 ( .A1(n15403), .A2(n15404), .ZN(n15504) );
  NAND2_X1 U15425 ( .A1(n15508), .A2(n15509), .ZN(n15404) );
  NAND2_X1 U15426 ( .A1(n15510), .A2(b_5_), .ZN(n15509) );
  NOR2_X1 U15427 ( .A1(n15511), .A2(n8495), .ZN(n15510) );
  NOR2_X1 U15428 ( .A1(n15400), .A2(n15399), .ZN(n15511) );
  NAND2_X1 U15429 ( .A1(n15399), .A2(n15400), .ZN(n15508) );
  NAND2_X1 U15430 ( .A1(n15512), .A2(n15513), .ZN(n15400) );
  NAND2_X1 U15431 ( .A1(n15514), .A2(b_5_), .ZN(n15513) );
  NOR2_X1 U15432 ( .A1(n15515), .A2(n8953), .ZN(n15514) );
  NOR2_X1 U15433 ( .A1(n15396), .A2(n15395), .ZN(n15515) );
  NAND2_X1 U15434 ( .A1(n15395), .A2(n15396), .ZN(n15512) );
  NAND2_X1 U15435 ( .A1(n15516), .A2(n15517), .ZN(n15396) );
  NAND2_X1 U15436 ( .A1(n15518), .A2(b_5_), .ZN(n15517) );
  NOR2_X1 U15437 ( .A1(n15519), .A2(n8440), .ZN(n15518) );
  NOR2_X1 U15438 ( .A1(n15391), .A2(n15392), .ZN(n15519) );
  NAND2_X1 U15439 ( .A1(n15391), .A2(n15392), .ZN(n15516) );
  NAND2_X1 U15440 ( .A1(n15520), .A2(n15521), .ZN(n15392) );
  NAND2_X1 U15441 ( .A1(n15522), .A2(b_5_), .ZN(n15521) );
  NOR2_X1 U15442 ( .A1(n15523), .A2(n8950), .ZN(n15522) );
  NOR2_X1 U15443 ( .A1(n15388), .A2(n15387), .ZN(n15523) );
  NAND2_X1 U15444 ( .A1(n15387), .A2(n15388), .ZN(n15520) );
  NAND2_X1 U15445 ( .A1(n15524), .A2(n15525), .ZN(n15388) );
  NAND2_X1 U15446 ( .A1(n15526), .A2(b_5_), .ZN(n15525) );
  NOR2_X1 U15447 ( .A1(n15527), .A2(n8385), .ZN(n15526) );
  NOR2_X1 U15448 ( .A1(n15383), .A2(n15384), .ZN(n15527) );
  NAND2_X1 U15449 ( .A1(n15383), .A2(n15384), .ZN(n15524) );
  NAND2_X1 U15450 ( .A1(n15528), .A2(n15529), .ZN(n15384) );
  NAND2_X1 U15451 ( .A1(n15530), .A2(b_5_), .ZN(n15529) );
  NOR2_X1 U15452 ( .A1(n15531), .A2(n8947), .ZN(n15530) );
  NOR2_X1 U15453 ( .A1(n15380), .A2(n15379), .ZN(n15531) );
  NAND2_X1 U15454 ( .A1(n15379), .A2(n15380), .ZN(n15528) );
  NAND2_X1 U15455 ( .A1(n15532), .A2(n15533), .ZN(n15380) );
  NAND2_X1 U15456 ( .A1(n15534), .A2(b_5_), .ZN(n15533) );
  NOR2_X1 U15457 ( .A1(n15535), .A2(n8324), .ZN(n15534) );
  NOR2_X1 U15458 ( .A1(n15375), .A2(n15376), .ZN(n15535) );
  NAND2_X1 U15459 ( .A1(n15375), .A2(n15376), .ZN(n15532) );
  NAND2_X1 U15460 ( .A1(n15536), .A2(n15537), .ZN(n15376) );
  NAND2_X1 U15461 ( .A1(n15538), .A2(b_5_), .ZN(n15537) );
  NOR2_X1 U15462 ( .A1(n15539), .A2(n8944), .ZN(n15538) );
  NOR2_X1 U15463 ( .A1(n15372), .A2(n15371), .ZN(n15539) );
  NAND2_X1 U15464 ( .A1(n15371), .A2(n15372), .ZN(n15536) );
  NAND2_X1 U15465 ( .A1(n15540), .A2(n15541), .ZN(n15372) );
  NAND2_X1 U15466 ( .A1(n15542), .A2(b_5_), .ZN(n15541) );
  NOR2_X1 U15467 ( .A1(n15543), .A2(n8268), .ZN(n15542) );
  NOR2_X1 U15468 ( .A1(n15367), .A2(n15368), .ZN(n15543) );
  NAND2_X1 U15469 ( .A1(n15367), .A2(n15368), .ZN(n15540) );
  NAND2_X1 U15470 ( .A1(n15544), .A2(n15545), .ZN(n15368) );
  NAND2_X1 U15471 ( .A1(n15546), .A2(b_5_), .ZN(n15545) );
  NOR2_X1 U15472 ( .A1(n15547), .A2(n8941), .ZN(n15546) );
  NOR2_X1 U15473 ( .A1(n15362), .A2(n15364), .ZN(n15547) );
  NAND2_X1 U15474 ( .A1(n15362), .A2(n15364), .ZN(n15544) );
  NAND2_X1 U15475 ( .A1(n15548), .A2(n15549), .ZN(n15364) );
  NAND2_X1 U15476 ( .A1(n15550), .A2(b_5_), .ZN(n15549) );
  NOR2_X1 U15477 ( .A1(n15551), .A2(n8213), .ZN(n15550) );
  NOR2_X1 U15478 ( .A1(n15301), .A2(n15303), .ZN(n15551) );
  NAND2_X1 U15479 ( .A1(n15301), .A2(n15303), .ZN(n15548) );
  NAND2_X1 U15480 ( .A1(n15552), .A2(n15553), .ZN(n15303) );
  NAND2_X1 U15481 ( .A1(n15554), .A2(b_5_), .ZN(n15553) );
  NOR2_X1 U15482 ( .A1(n15555), .A2(n8939), .ZN(n15554) );
  NOR2_X1 U15483 ( .A1(n15359), .A2(n15360), .ZN(n15555) );
  NAND2_X1 U15484 ( .A1(n15359), .A2(n15360), .ZN(n15552) );
  NAND2_X1 U15485 ( .A1(n15356), .A2(n15556), .ZN(n15360) );
  NAND2_X1 U15486 ( .A1(n15355), .A2(n15357), .ZN(n15556) );
  NAND2_X1 U15487 ( .A1(n15557), .A2(n15558), .ZN(n15357) );
  NAND2_X1 U15488 ( .A1(b_5_), .A2(a_25_), .ZN(n15558) );
  INV_X1 U15489 ( .A(n15559), .ZN(n15557) );
  XNOR2_X1 U15490 ( .A(n15560), .B(n15561), .ZN(n15355) );
  NAND2_X1 U15491 ( .A1(n15562), .A2(n15563), .ZN(n15560) );
  NAND2_X1 U15492 ( .A1(a_25_), .A2(n15559), .ZN(n15356) );
  NAND2_X1 U15493 ( .A1(n15318), .A2(n15564), .ZN(n15559) );
  NAND2_X1 U15494 ( .A1(n15317), .A2(n15319), .ZN(n15564) );
  NAND2_X1 U15495 ( .A1(n15565), .A2(n15566), .ZN(n15319) );
  NAND2_X1 U15496 ( .A1(b_5_), .A2(a_26_), .ZN(n15566) );
  INV_X1 U15497 ( .A(n15567), .ZN(n15565) );
  XNOR2_X1 U15498 ( .A(n15568), .B(n15569), .ZN(n15317) );
  NAND2_X1 U15499 ( .A1(n15570), .A2(n15571), .ZN(n15568) );
  NAND2_X1 U15500 ( .A1(a_26_), .A2(n15567), .ZN(n15318) );
  NAND2_X1 U15501 ( .A1(n15326), .A2(n15572), .ZN(n15567) );
  NAND2_X1 U15502 ( .A1(n15325), .A2(n15327), .ZN(n15572) );
  NAND2_X1 U15503 ( .A1(n15573), .A2(n15574), .ZN(n15327) );
  NAND2_X1 U15504 ( .A1(b_5_), .A2(a_27_), .ZN(n15574) );
  INV_X1 U15505 ( .A(n15575), .ZN(n15573) );
  XOR2_X1 U15506 ( .A(n15576), .B(n15577), .Z(n15325) );
  XNOR2_X1 U15507 ( .A(n15578), .B(n15579), .ZN(n15576) );
  NAND2_X1 U15508 ( .A1(b_4_), .A2(a_28_), .ZN(n15578) );
  NAND2_X1 U15509 ( .A1(a_27_), .A2(n15575), .ZN(n15326) );
  NAND2_X1 U15510 ( .A1(n15580), .A2(n15581), .ZN(n15575) );
  NAND2_X1 U15511 ( .A1(n15582), .A2(b_5_), .ZN(n15581) );
  NOR2_X1 U15512 ( .A1(n15583), .A2(n8055), .ZN(n15582) );
  NOR2_X1 U15513 ( .A1(n15333), .A2(n15335), .ZN(n15583) );
  NAND2_X1 U15514 ( .A1(n15333), .A2(n15335), .ZN(n15580) );
  NAND2_X1 U15515 ( .A1(n15584), .A2(n15585), .ZN(n15335) );
  NAND2_X1 U15516 ( .A1(n15351), .A2(n15586), .ZN(n15585) );
  OR2_X1 U15517 ( .A1(n15352), .A2(n15353), .ZN(n15586) );
  NOR2_X1 U15518 ( .A1(n8964), .A2(n8041), .ZN(n15351) );
  NAND2_X1 U15519 ( .A1(n15353), .A2(n15352), .ZN(n15584) );
  NAND2_X1 U15520 ( .A1(n15587), .A2(n15588), .ZN(n15352) );
  NAND2_X1 U15521 ( .A1(b_3_), .A2(n15589), .ZN(n15588) );
  NAND2_X1 U15522 ( .A1(n8003), .A2(n15590), .ZN(n15589) );
  NAND2_X1 U15523 ( .A1(a_31_), .A2(n8965), .ZN(n15590) );
  NAND2_X1 U15524 ( .A1(b_4_), .A2(n15591), .ZN(n15587) );
  NAND2_X1 U15525 ( .A1(n9341), .A2(n15592), .ZN(n15591) );
  NAND2_X1 U15526 ( .A1(a_30_), .A2(n8967), .ZN(n15592) );
  AND2_X1 U15527 ( .A1(n15593), .A2(n7953), .ZN(n15353) );
  NOR2_X1 U15528 ( .A1(n8964), .A2(n8965), .ZN(n15593) );
  XOR2_X1 U15529 ( .A(n15594), .B(n15595), .Z(n15333) );
  XOR2_X1 U15530 ( .A(n15596), .B(n15597), .Z(n15594) );
  XNOR2_X1 U15531 ( .A(n15598), .B(n15599), .ZN(n15359) );
  XNOR2_X1 U15532 ( .A(n15600), .B(n15601), .ZN(n15599) );
  XOR2_X1 U15533 ( .A(n15602), .B(n15603), .Z(n15301) );
  XOR2_X1 U15534 ( .A(n15604), .B(n15605), .Z(n15602) );
  XOR2_X1 U15535 ( .A(n15606), .B(n15607), .Z(n15362) );
  XOR2_X1 U15536 ( .A(n15608), .B(n15609), .Z(n15606) );
  XOR2_X1 U15537 ( .A(n15610), .B(n15611), .Z(n15367) );
  XOR2_X1 U15538 ( .A(n15612), .B(n15613), .Z(n15610) );
  XNOR2_X1 U15539 ( .A(n15614), .B(n15615), .ZN(n15371) );
  XNOR2_X1 U15540 ( .A(n15616), .B(n15617), .ZN(n15614) );
  XOR2_X1 U15541 ( .A(n15618), .B(n15619), .Z(n15375) );
  XOR2_X1 U15542 ( .A(n15620), .B(n15621), .Z(n15618) );
  XNOR2_X1 U15543 ( .A(n15622), .B(n15623), .ZN(n15379) );
  XNOR2_X1 U15544 ( .A(n15624), .B(n15625), .ZN(n15622) );
  XNOR2_X1 U15545 ( .A(n15626), .B(n15627), .ZN(n15383) );
  XNOR2_X1 U15546 ( .A(n15628), .B(n15629), .ZN(n15627) );
  XNOR2_X1 U15547 ( .A(n15630), .B(n15631), .ZN(n15387) );
  XNOR2_X1 U15548 ( .A(n15632), .B(n15633), .ZN(n15630) );
  XOR2_X1 U15549 ( .A(n15634), .B(n15635), .Z(n15391) );
  XOR2_X1 U15550 ( .A(n15636), .B(n15637), .Z(n15634) );
  XNOR2_X1 U15551 ( .A(n15638), .B(n15639), .ZN(n15395) );
  XNOR2_X1 U15552 ( .A(n15640), .B(n15641), .ZN(n15638) );
  XNOR2_X1 U15553 ( .A(n15642), .B(n15643), .ZN(n15399) );
  XNOR2_X1 U15554 ( .A(n15644), .B(n15645), .ZN(n15643) );
  XOR2_X1 U15555 ( .A(n15646), .B(n15647), .Z(n15403) );
  XNOR2_X1 U15556 ( .A(n15648), .B(n15649), .ZN(n15646) );
  NAND2_X1 U15557 ( .A1(b_4_), .A2(a_13_), .ZN(n15648) );
  XOR2_X1 U15558 ( .A(n15650), .B(n15651), .Z(n15407) );
  XOR2_X1 U15559 ( .A(n15652), .B(n15653), .Z(n15650) );
  NOR2_X1 U15560 ( .A1(n8956), .A2(n8965), .ZN(n15653) );
  XOR2_X1 U15561 ( .A(n15654), .B(n15655), .Z(n15411) );
  XOR2_X1 U15562 ( .A(n15656), .B(n15657), .Z(n15654) );
  NOR2_X1 U15563 ( .A1(n8550), .A2(n8965), .ZN(n15657) );
  XOR2_X1 U15564 ( .A(n15658), .B(n15659), .Z(n15415) );
  XOR2_X1 U15565 ( .A(n15660), .B(n15661), .Z(n15658) );
  NOR2_X1 U15566 ( .A1(n8959), .A2(n8965), .ZN(n15661) );
  XOR2_X1 U15567 ( .A(n15662), .B(n15663), .Z(n15419) );
  XOR2_X1 U15568 ( .A(n15664), .B(n15665), .Z(n15662) );
  NOR2_X1 U15569 ( .A1(n8605), .A2(n8965), .ZN(n15665) );
  XOR2_X1 U15570 ( .A(n15666), .B(n15667), .Z(n15245) );
  XOR2_X1 U15571 ( .A(n15668), .B(n15669), .Z(n15666) );
  NOR2_X1 U15572 ( .A1(n8619), .A2(n8965), .ZN(n15669) );
  XOR2_X1 U15573 ( .A(n15670), .B(n15671), .Z(n15423) );
  XOR2_X1 U15574 ( .A(n15672), .B(n15673), .Z(n15670) );
  NOR2_X1 U15575 ( .A1(n8962), .A2(n8965), .ZN(n15673) );
  INV_X1 U15576 ( .A(n8873), .ZN(n15429) );
  NAND2_X1 U15577 ( .A1(b_5_), .A2(a_5_), .ZN(n8873) );
  XOR2_X1 U15578 ( .A(n15674), .B(n15675), .Z(n15431) );
  XOR2_X1 U15579 ( .A(n15676), .B(n15677), .Z(n15674) );
  NOR2_X1 U15580 ( .A1(n8723), .A2(n8965), .ZN(n15677) );
  XOR2_X1 U15581 ( .A(n15678), .B(n15679), .Z(n15435) );
  XOR2_X1 U15582 ( .A(n15680), .B(n15681), .Z(n15678) );
  XOR2_X1 U15583 ( .A(n15682), .B(n15683), .Z(n15439) );
  XNOR2_X1 U15584 ( .A(n15684), .B(n15685), .ZN(n15682) );
  NAND2_X1 U15585 ( .A1(b_4_), .A2(a_3_), .ZN(n15684) );
  XOR2_X1 U15586 ( .A(n15686), .B(n15687), .Z(n15443) );
  XNOR2_X1 U15587 ( .A(n15688), .B(n15689), .ZN(n15686) );
  NAND2_X1 U15588 ( .A1(b_4_), .A2(a_2_), .ZN(n15688) );
  XOR2_X1 U15589 ( .A(n15690), .B(n15691), .Z(n15447) );
  XOR2_X1 U15590 ( .A(n15692), .B(n15693), .Z(n15690) );
  NOR2_X1 U15591 ( .A1(n8969), .A2(n8965), .ZN(n15693) );
  XNOR2_X1 U15592 ( .A(n15215), .B(n15214), .ZN(n15453) );
  XNOR2_X1 U15593 ( .A(n15694), .B(n15695), .ZN(n15215) );
  NOR2_X1 U15594 ( .A1(n8974), .A2(n8965), .ZN(n15695) );
  NAND2_X1 U15595 ( .A1(n15696), .A2(n15697), .ZN(n8646) );
  OR2_X1 U15596 ( .A1(n15697), .A2(n15696), .ZN(n8645) );
  NAND2_X1 U15597 ( .A1(n15698), .A2(n15699), .ZN(n15696) );
  NAND2_X1 U15598 ( .A1(n15700), .A2(n15701), .ZN(n15699) );
  INV_X1 U15599 ( .A(n15702), .ZN(n15701) );
  XNOR2_X1 U15600 ( .A(n15703), .B(n15704), .ZN(n15700) );
  NAND2_X1 U15601 ( .A1(n15452), .A2(n15451), .ZN(n15697) );
  NAND2_X1 U15602 ( .A1(n15705), .A2(n15706), .ZN(n15451) );
  NAND2_X1 U15603 ( .A1(n15707), .A2(b_4_), .ZN(n15706) );
  NOR2_X1 U15604 ( .A1(n15708), .A2(n8974), .ZN(n15707) );
  NOR2_X1 U15605 ( .A1(n15694), .A2(n15214), .ZN(n15708) );
  NAND2_X1 U15606 ( .A1(n15214), .A2(n15694), .ZN(n15705) );
  NAND2_X1 U15607 ( .A1(n15709), .A2(n15710), .ZN(n15694) );
  NAND2_X1 U15608 ( .A1(n15711), .A2(b_4_), .ZN(n15710) );
  NOR2_X1 U15609 ( .A1(n15712), .A2(n8969), .ZN(n15711) );
  NOR2_X1 U15610 ( .A1(n15691), .A2(n15692), .ZN(n15712) );
  NAND2_X1 U15611 ( .A1(n15691), .A2(n15692), .ZN(n15709) );
  NAND2_X1 U15612 ( .A1(n15713), .A2(n15714), .ZN(n15692) );
  NAND2_X1 U15613 ( .A1(n15715), .A2(b_4_), .ZN(n15714) );
  NOR2_X1 U15614 ( .A1(n15716), .A2(n8792), .ZN(n15715) );
  NOR2_X1 U15615 ( .A1(n15689), .A2(n15687), .ZN(n15716) );
  NAND2_X1 U15616 ( .A1(n15687), .A2(n15689), .ZN(n15713) );
  NAND2_X1 U15617 ( .A1(n15717), .A2(n15718), .ZN(n15689) );
  NAND2_X1 U15618 ( .A1(n15719), .A2(b_4_), .ZN(n15718) );
  NOR2_X1 U15619 ( .A1(n15720), .A2(n8778), .ZN(n15719) );
  NOR2_X1 U15620 ( .A1(n15683), .A2(n15685), .ZN(n15720) );
  NAND2_X1 U15621 ( .A1(n15683), .A2(n15685), .ZN(n15717) );
  NAND2_X1 U15622 ( .A1(n15721), .A2(n15722), .ZN(n15685) );
  NAND2_X1 U15623 ( .A1(n15679), .A2(n15723), .ZN(n15722) );
  OR2_X1 U15624 ( .A1(n15680), .A2(n15681), .ZN(n15723) );
  XNOR2_X1 U15625 ( .A(n15724), .B(n15725), .ZN(n15679) );
  NAND2_X1 U15626 ( .A1(n15726), .A2(n15727), .ZN(n15724) );
  NAND2_X1 U15627 ( .A1(n15681), .A2(n15680), .ZN(n15721) );
  NAND2_X1 U15628 ( .A1(n15728), .A2(n15729), .ZN(n15680) );
  NAND2_X1 U15629 ( .A1(n15730), .A2(b_4_), .ZN(n15729) );
  NOR2_X1 U15630 ( .A1(n15731), .A2(n8723), .ZN(n15730) );
  NOR2_X1 U15631 ( .A1(n15675), .A2(n15676), .ZN(n15731) );
  NAND2_X1 U15632 ( .A1(n15675), .A2(n15676), .ZN(n15728) );
  NAND2_X1 U15633 ( .A1(n15732), .A2(n15733), .ZN(n15676) );
  NAND2_X1 U15634 ( .A1(n15734), .A2(b_4_), .ZN(n15733) );
  NOR2_X1 U15635 ( .A1(n15735), .A2(n8681), .ZN(n15734) );
  NOR2_X1 U15636 ( .A1(n15477), .A2(n15478), .ZN(n15735) );
  NAND2_X1 U15637 ( .A1(n15477), .A2(n15478), .ZN(n15732) );
  NAND2_X1 U15638 ( .A1(n15736), .A2(n15737), .ZN(n15478) );
  NAND2_X1 U15639 ( .A1(n15738), .A2(b_4_), .ZN(n15737) );
  NOR2_X1 U15640 ( .A1(n15739), .A2(n8962), .ZN(n15738) );
  NOR2_X1 U15641 ( .A1(n15671), .A2(n15672), .ZN(n15739) );
  NAND2_X1 U15642 ( .A1(n15671), .A2(n15672), .ZN(n15736) );
  NAND2_X1 U15643 ( .A1(n15740), .A2(n15741), .ZN(n15672) );
  NAND2_X1 U15644 ( .A1(n15742), .A2(b_4_), .ZN(n15741) );
  NOR2_X1 U15645 ( .A1(n15743), .A2(n8619), .ZN(n15742) );
  NOR2_X1 U15646 ( .A1(n15667), .A2(n15668), .ZN(n15743) );
  NAND2_X1 U15647 ( .A1(n15667), .A2(n15668), .ZN(n15740) );
  NAND2_X1 U15648 ( .A1(n15744), .A2(n15745), .ZN(n15668) );
  NAND2_X1 U15649 ( .A1(n15746), .A2(b_4_), .ZN(n15745) );
  NOR2_X1 U15650 ( .A1(n15747), .A2(n8605), .ZN(n15746) );
  NOR2_X1 U15651 ( .A1(n15663), .A2(n15664), .ZN(n15747) );
  NAND2_X1 U15652 ( .A1(n15663), .A2(n15664), .ZN(n15744) );
  NAND2_X1 U15653 ( .A1(n15748), .A2(n15749), .ZN(n15664) );
  NAND2_X1 U15654 ( .A1(n15750), .A2(b_4_), .ZN(n15749) );
  NOR2_X1 U15655 ( .A1(n15751), .A2(n8959), .ZN(n15750) );
  NOR2_X1 U15656 ( .A1(n15659), .A2(n15660), .ZN(n15751) );
  NAND2_X1 U15657 ( .A1(n15659), .A2(n15660), .ZN(n15748) );
  NAND2_X1 U15658 ( .A1(n15752), .A2(n15753), .ZN(n15660) );
  NAND2_X1 U15659 ( .A1(n15754), .A2(b_4_), .ZN(n15753) );
  NOR2_X1 U15660 ( .A1(n15755), .A2(n8550), .ZN(n15754) );
  NOR2_X1 U15661 ( .A1(n15655), .A2(n15656), .ZN(n15755) );
  NAND2_X1 U15662 ( .A1(n15655), .A2(n15656), .ZN(n15752) );
  NAND2_X1 U15663 ( .A1(n15756), .A2(n15757), .ZN(n15656) );
  NAND2_X1 U15664 ( .A1(n15758), .A2(b_4_), .ZN(n15757) );
  NOR2_X1 U15665 ( .A1(n15759), .A2(n8956), .ZN(n15758) );
  NOR2_X1 U15666 ( .A1(n15651), .A2(n15652), .ZN(n15759) );
  NAND2_X1 U15667 ( .A1(n15651), .A2(n15652), .ZN(n15756) );
  NAND2_X1 U15668 ( .A1(n15760), .A2(n15761), .ZN(n15652) );
  NAND2_X1 U15669 ( .A1(n15762), .A2(b_4_), .ZN(n15761) );
  NOR2_X1 U15670 ( .A1(n15763), .A2(n8495), .ZN(n15762) );
  NOR2_X1 U15671 ( .A1(n15647), .A2(n15649), .ZN(n15763) );
  NAND2_X1 U15672 ( .A1(n15647), .A2(n15649), .ZN(n15760) );
  NAND2_X1 U15673 ( .A1(n15764), .A2(n15765), .ZN(n15649) );
  NAND2_X1 U15674 ( .A1(n15645), .A2(n15766), .ZN(n15765) );
  OR2_X1 U15675 ( .A1(n15644), .A2(n15642), .ZN(n15766) );
  NOR2_X1 U15676 ( .A1(n8965), .A2(n8953), .ZN(n15645) );
  NAND2_X1 U15677 ( .A1(n15642), .A2(n15644), .ZN(n15764) );
  NAND2_X1 U15678 ( .A1(n15767), .A2(n15768), .ZN(n15644) );
  NAND2_X1 U15679 ( .A1(n15641), .A2(n15769), .ZN(n15768) );
  NAND2_X1 U15680 ( .A1(n15640), .A2(n15639), .ZN(n15769) );
  NOR2_X1 U15681 ( .A1(n8965), .A2(n8440), .ZN(n15641) );
  OR2_X1 U15682 ( .A1(n15639), .A2(n15640), .ZN(n15767) );
  AND2_X1 U15683 ( .A1(n15770), .A2(n15771), .ZN(n15640) );
  NAND2_X1 U15684 ( .A1(n15637), .A2(n15772), .ZN(n15771) );
  OR2_X1 U15685 ( .A1(n15635), .A2(n15636), .ZN(n15772) );
  NOR2_X1 U15686 ( .A1(n8965), .A2(n8950), .ZN(n15637) );
  NAND2_X1 U15687 ( .A1(n15635), .A2(n15636), .ZN(n15770) );
  NAND2_X1 U15688 ( .A1(n15773), .A2(n15774), .ZN(n15636) );
  NAND2_X1 U15689 ( .A1(n15633), .A2(n15775), .ZN(n15774) );
  NAND2_X1 U15690 ( .A1(n15632), .A2(n15631), .ZN(n15775) );
  NOR2_X1 U15691 ( .A1(n8965), .A2(n8385), .ZN(n15633) );
  OR2_X1 U15692 ( .A1(n15631), .A2(n15632), .ZN(n15773) );
  AND2_X1 U15693 ( .A1(n15776), .A2(n15777), .ZN(n15632) );
  NAND2_X1 U15694 ( .A1(n15629), .A2(n15778), .ZN(n15777) );
  OR2_X1 U15695 ( .A1(n15626), .A2(n15628), .ZN(n15778) );
  NOR2_X1 U15696 ( .A1(n8965), .A2(n8947), .ZN(n15629) );
  NAND2_X1 U15697 ( .A1(n15626), .A2(n15628), .ZN(n15776) );
  NAND2_X1 U15698 ( .A1(n15779), .A2(n15780), .ZN(n15628) );
  NAND2_X1 U15699 ( .A1(n15625), .A2(n15781), .ZN(n15780) );
  NAND2_X1 U15700 ( .A1(n15624), .A2(n15623), .ZN(n15781) );
  NOR2_X1 U15701 ( .A1(n8965), .A2(n8324), .ZN(n15625) );
  OR2_X1 U15702 ( .A1(n15623), .A2(n15624), .ZN(n15779) );
  AND2_X1 U15703 ( .A1(n15782), .A2(n15783), .ZN(n15624) );
  NAND2_X1 U15704 ( .A1(n15621), .A2(n15784), .ZN(n15783) );
  OR2_X1 U15705 ( .A1(n15619), .A2(n15620), .ZN(n15784) );
  NOR2_X1 U15706 ( .A1(n8965), .A2(n8944), .ZN(n15621) );
  NAND2_X1 U15707 ( .A1(n15619), .A2(n15620), .ZN(n15782) );
  NAND2_X1 U15708 ( .A1(n15785), .A2(n15786), .ZN(n15620) );
  NAND2_X1 U15709 ( .A1(n15617), .A2(n15787), .ZN(n15786) );
  NAND2_X1 U15710 ( .A1(n15616), .A2(n15615), .ZN(n15787) );
  NOR2_X1 U15711 ( .A1(n8965), .A2(n8268), .ZN(n15617) );
  OR2_X1 U15712 ( .A1(n15615), .A2(n15616), .ZN(n15785) );
  AND2_X1 U15713 ( .A1(n15788), .A2(n15789), .ZN(n15616) );
  NAND2_X1 U15714 ( .A1(n15613), .A2(n15790), .ZN(n15789) );
  OR2_X1 U15715 ( .A1(n15611), .A2(n15612), .ZN(n15790) );
  NOR2_X1 U15716 ( .A1(n8965), .A2(n8941), .ZN(n15613) );
  NAND2_X1 U15717 ( .A1(n15611), .A2(n15612), .ZN(n15788) );
  NAND2_X1 U15718 ( .A1(n15791), .A2(n15792), .ZN(n15612) );
  NAND2_X1 U15719 ( .A1(n15609), .A2(n15793), .ZN(n15792) );
  OR2_X1 U15720 ( .A1(n15607), .A2(n15608), .ZN(n15793) );
  NOR2_X1 U15721 ( .A1(n8965), .A2(n8213), .ZN(n15609) );
  NAND2_X1 U15722 ( .A1(n15607), .A2(n15608), .ZN(n15791) );
  NAND2_X1 U15723 ( .A1(n15794), .A2(n15795), .ZN(n15608) );
  NAND2_X1 U15724 ( .A1(n15605), .A2(n15796), .ZN(n15795) );
  OR2_X1 U15725 ( .A1(n15603), .A2(n15604), .ZN(n15796) );
  NOR2_X1 U15726 ( .A1(n8965), .A2(n8939), .ZN(n15605) );
  NAND2_X1 U15727 ( .A1(n15603), .A2(n15604), .ZN(n15794) );
  NAND2_X1 U15728 ( .A1(n15797), .A2(n15798), .ZN(n15604) );
  NAND2_X1 U15729 ( .A1(n15601), .A2(n15799), .ZN(n15798) );
  OR2_X1 U15730 ( .A1(n15598), .A2(n15600), .ZN(n15799) );
  NOR2_X1 U15731 ( .A1(n8965), .A2(n8158), .ZN(n15601) );
  NAND2_X1 U15732 ( .A1(n15598), .A2(n15600), .ZN(n15797) );
  NAND2_X1 U15733 ( .A1(n15562), .A2(n15800), .ZN(n15600) );
  NAND2_X1 U15734 ( .A1(n15561), .A2(n15563), .ZN(n15800) );
  NAND2_X1 U15735 ( .A1(n15801), .A2(n15802), .ZN(n15563) );
  NAND2_X1 U15736 ( .A1(b_4_), .A2(a_26_), .ZN(n15802) );
  INV_X1 U15737 ( .A(n15803), .ZN(n15801) );
  XNOR2_X1 U15738 ( .A(n15804), .B(n15805), .ZN(n15561) );
  NAND2_X1 U15739 ( .A1(n15806), .A2(n15807), .ZN(n15804) );
  NAND2_X1 U15740 ( .A1(a_26_), .A2(n15803), .ZN(n15562) );
  NAND2_X1 U15741 ( .A1(n15570), .A2(n15808), .ZN(n15803) );
  NAND2_X1 U15742 ( .A1(n15569), .A2(n15571), .ZN(n15808) );
  NAND2_X1 U15743 ( .A1(n15809), .A2(n15810), .ZN(n15571) );
  NAND2_X1 U15744 ( .A1(b_4_), .A2(a_27_), .ZN(n15810) );
  INV_X1 U15745 ( .A(n15811), .ZN(n15809) );
  XOR2_X1 U15746 ( .A(n15812), .B(n15813), .Z(n15569) );
  XNOR2_X1 U15747 ( .A(n15814), .B(n15815), .ZN(n15812) );
  NAND2_X1 U15748 ( .A1(b_3_), .A2(a_28_), .ZN(n15814) );
  NAND2_X1 U15749 ( .A1(a_27_), .A2(n15811), .ZN(n15570) );
  NAND2_X1 U15750 ( .A1(n15816), .A2(n15817), .ZN(n15811) );
  NAND2_X1 U15751 ( .A1(n15818), .A2(b_4_), .ZN(n15817) );
  NOR2_X1 U15752 ( .A1(n15819), .A2(n8055), .ZN(n15818) );
  NOR2_X1 U15753 ( .A1(n15577), .A2(n15579), .ZN(n15819) );
  NAND2_X1 U15754 ( .A1(n15577), .A2(n15579), .ZN(n15816) );
  NAND2_X1 U15755 ( .A1(n15820), .A2(n15821), .ZN(n15579) );
  NAND2_X1 U15756 ( .A1(n15595), .A2(n15822), .ZN(n15821) );
  OR2_X1 U15757 ( .A1(n15596), .A2(n15597), .ZN(n15822) );
  NOR2_X1 U15758 ( .A1(n8965), .A2(n8041), .ZN(n15595) );
  NAND2_X1 U15759 ( .A1(n15597), .A2(n15596), .ZN(n15820) );
  NAND2_X1 U15760 ( .A1(n15823), .A2(n15824), .ZN(n15596) );
  NAND2_X1 U15761 ( .A1(b_2_), .A2(n15825), .ZN(n15824) );
  NAND2_X1 U15762 ( .A1(n8003), .A2(n15826), .ZN(n15825) );
  NAND2_X1 U15763 ( .A1(a_31_), .A2(n8967), .ZN(n15826) );
  NAND2_X1 U15764 ( .A1(b_3_), .A2(n15827), .ZN(n15823) );
  NAND2_X1 U15765 ( .A1(n9341), .A2(n15828), .ZN(n15827) );
  NAND2_X1 U15766 ( .A1(a_30_), .A2(n8968), .ZN(n15828) );
  AND2_X1 U15767 ( .A1(n15829), .A2(n7953), .ZN(n15597) );
  NOR2_X1 U15768 ( .A1(n8965), .A2(n8967), .ZN(n15829) );
  XOR2_X1 U15769 ( .A(n15830), .B(n15831), .Z(n15577) );
  XOR2_X1 U15770 ( .A(n15832), .B(n15833), .Z(n15830) );
  XNOR2_X1 U15771 ( .A(n15834), .B(n15835), .ZN(n15598) );
  NAND2_X1 U15772 ( .A1(n15836), .A2(n15837), .ZN(n15834) );
  XNOR2_X1 U15773 ( .A(n15838), .B(n15839), .ZN(n15603) );
  NAND2_X1 U15774 ( .A1(n15840), .A2(n15841), .ZN(n15838) );
  XOR2_X1 U15775 ( .A(n15842), .B(n15843), .Z(n15607) );
  XOR2_X1 U15776 ( .A(n15844), .B(n15845), .Z(n15842) );
  NOR2_X1 U15777 ( .A1(n8939), .A2(n8967), .ZN(n15845) );
  XNOR2_X1 U15778 ( .A(n15846), .B(n15847), .ZN(n15611) );
  NAND2_X1 U15779 ( .A1(n15848), .A2(n15849), .ZN(n15846) );
  XOR2_X1 U15780 ( .A(n15850), .B(n15851), .Z(n15615) );
  XOR2_X1 U15781 ( .A(n15852), .B(n15853), .Z(n15851) );
  NAND2_X1 U15782 ( .A1(b_3_), .A2(a_22_), .ZN(n15853) );
  XNOR2_X1 U15783 ( .A(n15854), .B(n15855), .ZN(n15619) );
  NAND2_X1 U15784 ( .A1(n15856), .A2(n15857), .ZN(n15854) );
  XNOR2_X1 U15785 ( .A(n15858), .B(n15859), .ZN(n15623) );
  XOR2_X1 U15786 ( .A(n15860), .B(n15861), .Z(n15858) );
  NOR2_X1 U15787 ( .A1(n8944), .A2(n8967), .ZN(n15861) );
  XNOR2_X1 U15788 ( .A(n15862), .B(n15863), .ZN(n15626) );
  NAND2_X1 U15789 ( .A1(n15864), .A2(n15865), .ZN(n15862) );
  XNOR2_X1 U15790 ( .A(n15866), .B(n15867), .ZN(n15631) );
  XNOR2_X1 U15791 ( .A(n15868), .B(n15869), .ZN(n15866) );
  NAND2_X1 U15792 ( .A1(b_3_), .A2(a_18_), .ZN(n15868) );
  XNOR2_X1 U15793 ( .A(n15870), .B(n15871), .ZN(n15635) );
  NAND2_X1 U15794 ( .A1(n15872), .A2(n15873), .ZN(n15870) );
  XNOR2_X1 U15795 ( .A(n15874), .B(n15875), .ZN(n15639) );
  XOR2_X1 U15796 ( .A(n15876), .B(n15877), .Z(n15874) );
  NOR2_X1 U15797 ( .A1(n8950), .A2(n8967), .ZN(n15877) );
  XNOR2_X1 U15798 ( .A(n15878), .B(n15879), .ZN(n15642) );
  NAND2_X1 U15799 ( .A1(n15880), .A2(n15881), .ZN(n15878) );
  XNOR2_X1 U15800 ( .A(n15882), .B(n15883), .ZN(n15647) );
  XOR2_X1 U15801 ( .A(n15884), .B(n15885), .Z(n15883) );
  NAND2_X1 U15802 ( .A1(b_3_), .A2(a_14_), .ZN(n15885) );
  XNOR2_X1 U15803 ( .A(n15886), .B(n15887), .ZN(n15651) );
  NAND2_X1 U15804 ( .A1(n15888), .A2(n15889), .ZN(n15886) );
  XOR2_X1 U15805 ( .A(n15890), .B(n15891), .Z(n15655) );
  XOR2_X1 U15806 ( .A(n15892), .B(n15893), .Z(n15890) );
  NOR2_X1 U15807 ( .A1(n8956), .A2(n8967), .ZN(n15893) );
  XNOR2_X1 U15808 ( .A(n15894), .B(n15895), .ZN(n15659) );
  NAND2_X1 U15809 ( .A1(n15896), .A2(n15897), .ZN(n15894) );
  XOR2_X1 U15810 ( .A(n15898), .B(n15899), .Z(n15663) );
  XOR2_X1 U15811 ( .A(n15900), .B(n15901), .Z(n15898) );
  NOR2_X1 U15812 ( .A1(n8959), .A2(n8967), .ZN(n15901) );
  XNOR2_X1 U15813 ( .A(n15902), .B(n15903), .ZN(n15667) );
  NAND2_X1 U15814 ( .A1(n15904), .A2(n15905), .ZN(n15902) );
  XOR2_X1 U15815 ( .A(n15906), .B(n15907), .Z(n15671) );
  XOR2_X1 U15816 ( .A(n15908), .B(n15909), .Z(n15906) );
  NOR2_X1 U15817 ( .A1(n8619), .A2(n8967), .ZN(n15909) );
  XNOR2_X1 U15818 ( .A(n15910), .B(n15911), .ZN(n15477) );
  NAND2_X1 U15819 ( .A1(n15912), .A2(n15913), .ZN(n15910) );
  XOR2_X1 U15820 ( .A(n15914), .B(n15915), .Z(n15675) );
  XOR2_X1 U15821 ( .A(n15916), .B(n15917), .Z(n15914) );
  NOR2_X1 U15822 ( .A1(n8681), .A2(n8967), .ZN(n15917) );
  INV_X1 U15823 ( .A(n8756), .ZN(n15681) );
  NAND2_X1 U15824 ( .A1(b_4_), .A2(a_4_), .ZN(n8756) );
  XOR2_X1 U15825 ( .A(n15918), .B(n15919), .Z(n15683) );
  XOR2_X1 U15826 ( .A(n15920), .B(n15921), .Z(n15918) );
  NOR2_X1 U15827 ( .A1(n8966), .A2(n8967), .ZN(n15921) );
  XOR2_X1 U15828 ( .A(n15922), .B(n15923), .Z(n15687) );
  XOR2_X1 U15829 ( .A(n15924), .B(n15925), .Z(n15922) );
  XOR2_X1 U15830 ( .A(n15926), .B(n15927), .Z(n15691) );
  XOR2_X1 U15831 ( .A(n15928), .B(n15929), .Z(n15926) );
  NOR2_X1 U15832 ( .A1(n8792), .A2(n8967), .ZN(n15929) );
  XNOR2_X1 U15833 ( .A(n15930), .B(n15931), .ZN(n15214) );
  NAND2_X1 U15834 ( .A1(n15932), .A2(n15933), .ZN(n15930) );
  XOR2_X1 U15835 ( .A(n15934), .B(n15935), .Z(n15452) );
  XOR2_X1 U15836 ( .A(n15936), .B(n15937), .Z(n15934) );
  NAND2_X1 U15837 ( .A1(n15938), .A2(n15698), .ZN(n8990) );
  XNOR2_X1 U15838 ( .A(n15939), .B(n15940), .ZN(n15938) );
  OR2_X1 U15839 ( .A1(n15941), .A2(n15698), .ZN(n8991) );
  NAND2_X1 U15840 ( .A1(n15942), .A2(n15702), .ZN(n15698) );
  NAND2_X1 U15841 ( .A1(n15943), .A2(n15944), .ZN(n15702) );
  NAND2_X1 U15842 ( .A1(n15937), .A2(n15945), .ZN(n15944) );
  OR2_X1 U15843 ( .A1(n15935), .A2(n15936), .ZN(n15945) );
  NOR2_X1 U15844 ( .A1(n8967), .A2(n8974), .ZN(n15937) );
  NAND2_X1 U15845 ( .A1(n15935), .A2(n15936), .ZN(n15943) );
  NAND2_X1 U15846 ( .A1(n15932), .A2(n15946), .ZN(n15936) );
  NAND2_X1 U15847 ( .A1(n15931), .A2(n15933), .ZN(n15946) );
  NAND2_X1 U15848 ( .A1(n15947), .A2(n15948), .ZN(n15933) );
  NAND2_X1 U15849 ( .A1(b_3_), .A2(a_1_), .ZN(n15948) );
  INV_X1 U15850 ( .A(n15949), .ZN(n15947) );
  XOR2_X1 U15851 ( .A(n15950), .B(n15951), .Z(n15931) );
  XOR2_X1 U15852 ( .A(n8812), .B(n15952), .Z(n15950) );
  NAND2_X1 U15853 ( .A1(a_1_), .A2(n15949), .ZN(n15932) );
  NAND2_X1 U15854 ( .A1(n15953), .A2(n15954), .ZN(n15949) );
  NAND2_X1 U15855 ( .A1(n15955), .A2(b_3_), .ZN(n15954) );
  NOR2_X1 U15856 ( .A1(n15956), .A2(n8792), .ZN(n15955) );
  NOR2_X1 U15857 ( .A1(n15928), .A2(n15927), .ZN(n15956) );
  NAND2_X1 U15858 ( .A1(n15927), .A2(n15928), .ZN(n15953) );
  NAND2_X1 U15859 ( .A1(n15957), .A2(n15958), .ZN(n15928) );
  NAND2_X1 U15860 ( .A1(n15923), .A2(n15959), .ZN(n15958) );
  OR2_X1 U15861 ( .A1(n15924), .A2(n15925), .ZN(n15959) );
  XNOR2_X1 U15862 ( .A(n15960), .B(n15961), .ZN(n15923) );
  NAND2_X1 U15863 ( .A1(n15962), .A2(n15963), .ZN(n15960) );
  NAND2_X1 U15864 ( .A1(n15925), .A2(n15924), .ZN(n15957) );
  NAND2_X1 U15865 ( .A1(n15964), .A2(n15965), .ZN(n15924) );
  NAND2_X1 U15866 ( .A1(n15966), .A2(b_3_), .ZN(n15965) );
  NOR2_X1 U15867 ( .A1(n15967), .A2(n8966), .ZN(n15966) );
  NOR2_X1 U15868 ( .A1(n15920), .A2(n15919), .ZN(n15967) );
  NAND2_X1 U15869 ( .A1(n15919), .A2(n15920), .ZN(n15964) );
  NAND2_X1 U15870 ( .A1(n15726), .A2(n15968), .ZN(n15920) );
  NAND2_X1 U15871 ( .A1(n15725), .A2(n15727), .ZN(n15968) );
  NAND2_X1 U15872 ( .A1(n15969), .A2(n15970), .ZN(n15727) );
  NAND2_X1 U15873 ( .A1(b_3_), .A2(a_5_), .ZN(n15970) );
  INV_X1 U15874 ( .A(n15971), .ZN(n15969) );
  XNOR2_X1 U15875 ( .A(n15972), .B(n15973), .ZN(n15725) );
  NAND2_X1 U15876 ( .A1(n15974), .A2(n15975), .ZN(n15972) );
  NAND2_X1 U15877 ( .A1(a_5_), .A2(n15971), .ZN(n15726) );
  NAND2_X1 U15878 ( .A1(n15976), .A2(n15977), .ZN(n15971) );
  NAND2_X1 U15879 ( .A1(n15978), .A2(b_3_), .ZN(n15977) );
  NOR2_X1 U15880 ( .A1(n15979), .A2(n8681), .ZN(n15978) );
  NOR2_X1 U15881 ( .A1(n15916), .A2(n15915), .ZN(n15979) );
  NAND2_X1 U15882 ( .A1(n15915), .A2(n15916), .ZN(n15976) );
  NAND2_X1 U15883 ( .A1(n15912), .A2(n15980), .ZN(n15916) );
  NAND2_X1 U15884 ( .A1(n15911), .A2(n15913), .ZN(n15980) );
  NAND2_X1 U15885 ( .A1(n15981), .A2(n15982), .ZN(n15913) );
  NAND2_X1 U15886 ( .A1(b_3_), .A2(a_7_), .ZN(n15982) );
  INV_X1 U15887 ( .A(n15983), .ZN(n15981) );
  XNOR2_X1 U15888 ( .A(n15984), .B(n15985), .ZN(n15911) );
  NAND2_X1 U15889 ( .A1(n15986), .A2(n15987), .ZN(n15984) );
  NAND2_X1 U15890 ( .A1(a_7_), .A2(n15983), .ZN(n15912) );
  NAND2_X1 U15891 ( .A1(n15988), .A2(n15989), .ZN(n15983) );
  NAND2_X1 U15892 ( .A1(n15990), .A2(b_3_), .ZN(n15989) );
  NOR2_X1 U15893 ( .A1(n15991), .A2(n8619), .ZN(n15990) );
  NOR2_X1 U15894 ( .A1(n15908), .A2(n15907), .ZN(n15991) );
  NAND2_X1 U15895 ( .A1(n15907), .A2(n15908), .ZN(n15988) );
  NAND2_X1 U15896 ( .A1(n15904), .A2(n15992), .ZN(n15908) );
  NAND2_X1 U15897 ( .A1(n15903), .A2(n15905), .ZN(n15992) );
  NAND2_X1 U15898 ( .A1(n15993), .A2(n15994), .ZN(n15905) );
  NAND2_X1 U15899 ( .A1(b_3_), .A2(a_9_), .ZN(n15994) );
  INV_X1 U15900 ( .A(n15995), .ZN(n15993) );
  XNOR2_X1 U15901 ( .A(n15996), .B(n15997), .ZN(n15903) );
  NAND2_X1 U15902 ( .A1(n15998), .A2(n15999), .ZN(n15996) );
  NAND2_X1 U15903 ( .A1(a_9_), .A2(n15995), .ZN(n15904) );
  NAND2_X1 U15904 ( .A1(n16000), .A2(n16001), .ZN(n15995) );
  NAND2_X1 U15905 ( .A1(n16002), .A2(b_3_), .ZN(n16001) );
  NOR2_X1 U15906 ( .A1(n16003), .A2(n8959), .ZN(n16002) );
  NOR2_X1 U15907 ( .A1(n15900), .A2(n15899), .ZN(n16003) );
  NAND2_X1 U15908 ( .A1(n15899), .A2(n15900), .ZN(n16000) );
  NAND2_X1 U15909 ( .A1(n15896), .A2(n16004), .ZN(n15900) );
  NAND2_X1 U15910 ( .A1(n15895), .A2(n15897), .ZN(n16004) );
  NAND2_X1 U15911 ( .A1(n16005), .A2(n16006), .ZN(n15897) );
  NAND2_X1 U15912 ( .A1(b_3_), .A2(a_11_), .ZN(n16006) );
  INV_X1 U15913 ( .A(n16007), .ZN(n16005) );
  XNOR2_X1 U15914 ( .A(n16008), .B(n16009), .ZN(n15895) );
  NAND2_X1 U15915 ( .A1(n16010), .A2(n16011), .ZN(n16008) );
  NAND2_X1 U15916 ( .A1(a_11_), .A2(n16007), .ZN(n15896) );
  NAND2_X1 U15917 ( .A1(n16012), .A2(n16013), .ZN(n16007) );
  NAND2_X1 U15918 ( .A1(n16014), .A2(b_3_), .ZN(n16013) );
  NOR2_X1 U15919 ( .A1(n16015), .A2(n8956), .ZN(n16014) );
  NOR2_X1 U15920 ( .A1(n15892), .A2(n15891), .ZN(n16015) );
  NAND2_X1 U15921 ( .A1(n15891), .A2(n15892), .ZN(n16012) );
  NAND2_X1 U15922 ( .A1(n15888), .A2(n16016), .ZN(n15892) );
  NAND2_X1 U15923 ( .A1(n15887), .A2(n15889), .ZN(n16016) );
  NAND2_X1 U15924 ( .A1(n16017), .A2(n16018), .ZN(n15889) );
  NAND2_X1 U15925 ( .A1(b_3_), .A2(a_13_), .ZN(n16018) );
  INV_X1 U15926 ( .A(n16019), .ZN(n16017) );
  XNOR2_X1 U15927 ( .A(n16020), .B(n16021), .ZN(n15887) );
  NAND2_X1 U15928 ( .A1(n16022), .A2(n16023), .ZN(n16020) );
  NAND2_X1 U15929 ( .A1(a_13_), .A2(n16019), .ZN(n15888) );
  NAND2_X1 U15930 ( .A1(n16024), .A2(n16025), .ZN(n16019) );
  NAND2_X1 U15931 ( .A1(n16026), .A2(b_3_), .ZN(n16025) );
  NOR2_X1 U15932 ( .A1(n16027), .A2(n8953), .ZN(n16026) );
  NOR2_X1 U15933 ( .A1(n15884), .A2(n15882), .ZN(n16027) );
  NAND2_X1 U15934 ( .A1(n15882), .A2(n15884), .ZN(n16024) );
  NAND2_X1 U15935 ( .A1(n15880), .A2(n16028), .ZN(n15884) );
  NAND2_X1 U15936 ( .A1(n15879), .A2(n15881), .ZN(n16028) );
  NAND2_X1 U15937 ( .A1(n16029), .A2(n16030), .ZN(n15881) );
  NAND2_X1 U15938 ( .A1(b_3_), .A2(a_15_), .ZN(n16030) );
  INV_X1 U15939 ( .A(n16031), .ZN(n16029) );
  XNOR2_X1 U15940 ( .A(n16032), .B(n16033), .ZN(n15879) );
  NAND2_X1 U15941 ( .A1(n16034), .A2(n16035), .ZN(n16032) );
  NAND2_X1 U15942 ( .A1(a_15_), .A2(n16031), .ZN(n15880) );
  NAND2_X1 U15943 ( .A1(n16036), .A2(n16037), .ZN(n16031) );
  NAND2_X1 U15944 ( .A1(n16038), .A2(b_3_), .ZN(n16037) );
  NOR2_X1 U15945 ( .A1(n16039), .A2(n8950), .ZN(n16038) );
  NOR2_X1 U15946 ( .A1(n15876), .A2(n15875), .ZN(n16039) );
  NAND2_X1 U15947 ( .A1(n15875), .A2(n15876), .ZN(n16036) );
  NAND2_X1 U15948 ( .A1(n15872), .A2(n16040), .ZN(n15876) );
  NAND2_X1 U15949 ( .A1(n15871), .A2(n15873), .ZN(n16040) );
  NAND2_X1 U15950 ( .A1(n16041), .A2(n16042), .ZN(n15873) );
  NAND2_X1 U15951 ( .A1(b_3_), .A2(a_17_), .ZN(n16042) );
  INV_X1 U15952 ( .A(n16043), .ZN(n16041) );
  XNOR2_X1 U15953 ( .A(n16044), .B(n16045), .ZN(n15871) );
  XNOR2_X1 U15954 ( .A(n16046), .B(n16047), .ZN(n16044) );
  NAND2_X1 U15955 ( .A1(a_17_), .A2(n16043), .ZN(n15872) );
  NAND2_X1 U15956 ( .A1(n16048), .A2(n16049), .ZN(n16043) );
  NAND2_X1 U15957 ( .A1(n16050), .A2(b_3_), .ZN(n16049) );
  NOR2_X1 U15958 ( .A1(n16051), .A2(n8947), .ZN(n16050) );
  NOR2_X1 U15959 ( .A1(n15869), .A2(n15867), .ZN(n16051) );
  NAND2_X1 U15960 ( .A1(n15867), .A2(n15869), .ZN(n16048) );
  NAND2_X1 U15961 ( .A1(n15864), .A2(n16052), .ZN(n15869) );
  NAND2_X1 U15962 ( .A1(n15863), .A2(n15865), .ZN(n16052) );
  NAND2_X1 U15963 ( .A1(n16053), .A2(n16054), .ZN(n15865) );
  NAND2_X1 U15964 ( .A1(b_3_), .A2(a_19_), .ZN(n16054) );
  INV_X1 U15965 ( .A(n16055), .ZN(n16053) );
  XNOR2_X1 U15966 ( .A(n16056), .B(n16057), .ZN(n15863) );
  XNOR2_X1 U15967 ( .A(n16058), .B(n16059), .ZN(n16056) );
  NAND2_X1 U15968 ( .A1(a_19_), .A2(n16055), .ZN(n15864) );
  NAND2_X1 U15969 ( .A1(n16060), .A2(n16061), .ZN(n16055) );
  NAND2_X1 U15970 ( .A1(n16062), .A2(b_3_), .ZN(n16061) );
  NOR2_X1 U15971 ( .A1(n16063), .A2(n8944), .ZN(n16062) );
  NOR2_X1 U15972 ( .A1(n15860), .A2(n15859), .ZN(n16063) );
  NAND2_X1 U15973 ( .A1(n15859), .A2(n15860), .ZN(n16060) );
  NAND2_X1 U15974 ( .A1(n15856), .A2(n16064), .ZN(n15860) );
  NAND2_X1 U15975 ( .A1(n15855), .A2(n15857), .ZN(n16064) );
  NAND2_X1 U15976 ( .A1(n16065), .A2(n16066), .ZN(n15857) );
  NAND2_X1 U15977 ( .A1(b_3_), .A2(a_21_), .ZN(n16066) );
  INV_X1 U15978 ( .A(n16067), .ZN(n16065) );
  XNOR2_X1 U15979 ( .A(n16068), .B(n16069), .ZN(n15855) );
  XNOR2_X1 U15980 ( .A(n16070), .B(n16071), .ZN(n16069) );
  NAND2_X1 U15981 ( .A1(a_21_), .A2(n16067), .ZN(n15856) );
  NAND2_X1 U15982 ( .A1(n16072), .A2(n16073), .ZN(n16067) );
  NAND2_X1 U15983 ( .A1(n16074), .A2(b_3_), .ZN(n16073) );
  NOR2_X1 U15984 ( .A1(n16075), .A2(n8941), .ZN(n16074) );
  NOR2_X1 U15985 ( .A1(n15852), .A2(n15850), .ZN(n16075) );
  NAND2_X1 U15986 ( .A1(n15850), .A2(n15852), .ZN(n16072) );
  NAND2_X1 U15987 ( .A1(n15848), .A2(n16076), .ZN(n15852) );
  NAND2_X1 U15988 ( .A1(n15847), .A2(n15849), .ZN(n16076) );
  NAND2_X1 U15989 ( .A1(n16077), .A2(n16078), .ZN(n15849) );
  NAND2_X1 U15990 ( .A1(b_3_), .A2(a_23_), .ZN(n16078) );
  INV_X1 U15991 ( .A(n16079), .ZN(n16077) );
  XNOR2_X1 U15992 ( .A(n16080), .B(n16081), .ZN(n15847) );
  XNOR2_X1 U15993 ( .A(n16082), .B(n16083), .ZN(n16081) );
  NAND2_X1 U15994 ( .A1(a_23_), .A2(n16079), .ZN(n15848) );
  NAND2_X1 U15995 ( .A1(n16084), .A2(n16085), .ZN(n16079) );
  NAND2_X1 U15996 ( .A1(n16086), .A2(b_3_), .ZN(n16085) );
  NOR2_X1 U15997 ( .A1(n16087), .A2(n8939), .ZN(n16086) );
  NOR2_X1 U15998 ( .A1(n15843), .A2(n15844), .ZN(n16087) );
  NAND2_X1 U15999 ( .A1(n15843), .A2(n15844), .ZN(n16084) );
  NAND2_X1 U16000 ( .A1(n15840), .A2(n16088), .ZN(n15844) );
  NAND2_X1 U16001 ( .A1(n15839), .A2(n15841), .ZN(n16088) );
  NAND2_X1 U16002 ( .A1(n16089), .A2(n16090), .ZN(n15841) );
  NAND2_X1 U16003 ( .A1(b_3_), .A2(a_25_), .ZN(n16090) );
  INV_X1 U16004 ( .A(n16091), .ZN(n16089) );
  XOR2_X1 U16005 ( .A(n16092), .B(n16093), .Z(n15839) );
  XNOR2_X1 U16006 ( .A(n16094), .B(n16095), .ZN(n16092) );
  NAND2_X1 U16007 ( .A1(b_2_), .A2(a_26_), .ZN(n16094) );
  NAND2_X1 U16008 ( .A1(a_25_), .A2(n16091), .ZN(n15840) );
  NAND2_X1 U16009 ( .A1(n15836), .A2(n16096), .ZN(n16091) );
  NAND2_X1 U16010 ( .A1(n15835), .A2(n15837), .ZN(n16096) );
  NAND2_X1 U16011 ( .A1(n16097), .A2(n16098), .ZN(n15837) );
  NAND2_X1 U16012 ( .A1(b_3_), .A2(a_26_), .ZN(n16098) );
  INV_X1 U16013 ( .A(n16099), .ZN(n16097) );
  XNOR2_X1 U16014 ( .A(n16100), .B(n16101), .ZN(n15835) );
  XNOR2_X1 U16015 ( .A(n16102), .B(n16103), .ZN(n16101) );
  NAND2_X1 U16016 ( .A1(a_26_), .A2(n16099), .ZN(n15836) );
  NAND2_X1 U16017 ( .A1(n15806), .A2(n16104), .ZN(n16099) );
  NAND2_X1 U16018 ( .A1(n15805), .A2(n15807), .ZN(n16104) );
  NAND2_X1 U16019 ( .A1(n16105), .A2(n16106), .ZN(n15807) );
  NAND2_X1 U16020 ( .A1(b_3_), .A2(a_27_), .ZN(n16106) );
  INV_X1 U16021 ( .A(n16107), .ZN(n16105) );
  XNOR2_X1 U16022 ( .A(n16108), .B(n16109), .ZN(n15805) );
  XOR2_X1 U16023 ( .A(n16110), .B(n16111), .Z(n16109) );
  NAND2_X1 U16024 ( .A1(b_2_), .A2(a_28_), .ZN(n16111) );
  NAND2_X1 U16025 ( .A1(a_27_), .A2(n16107), .ZN(n15806) );
  NAND2_X1 U16026 ( .A1(n16112), .A2(n16113), .ZN(n16107) );
  NAND2_X1 U16027 ( .A1(n16114), .A2(b_3_), .ZN(n16113) );
  NOR2_X1 U16028 ( .A1(n16115), .A2(n8055), .ZN(n16114) );
  NOR2_X1 U16029 ( .A1(n15813), .A2(n15815), .ZN(n16115) );
  NAND2_X1 U16030 ( .A1(n15813), .A2(n15815), .ZN(n16112) );
  NAND2_X1 U16031 ( .A1(n16116), .A2(n16117), .ZN(n15815) );
  NAND2_X1 U16032 ( .A1(n15831), .A2(n16118), .ZN(n16117) );
  OR2_X1 U16033 ( .A1(n15832), .A2(n15833), .ZN(n16118) );
  NOR2_X1 U16034 ( .A1(n8967), .A2(n8041), .ZN(n15831) );
  NAND2_X1 U16035 ( .A1(n15833), .A2(n15832), .ZN(n16116) );
  NAND2_X1 U16036 ( .A1(n16119), .A2(n16120), .ZN(n15832) );
  NAND2_X1 U16037 ( .A1(b_1_), .A2(n16121), .ZN(n16120) );
  NAND2_X1 U16038 ( .A1(n8003), .A2(n16122), .ZN(n16121) );
  NAND2_X1 U16039 ( .A1(a_31_), .A2(n8968), .ZN(n16122) );
  NAND2_X1 U16040 ( .A1(b_2_), .A2(n16123), .ZN(n16119) );
  NAND2_X1 U16041 ( .A1(n9341), .A2(n16124), .ZN(n16123) );
  NAND2_X1 U16042 ( .A1(a_30_), .A2(n8834), .ZN(n16124) );
  AND2_X1 U16043 ( .A1(n16125), .A2(n7953), .ZN(n15833) );
  NOR2_X1 U16044 ( .A1(n8967), .A2(n8968), .ZN(n16125) );
  XOR2_X1 U16045 ( .A(n16126), .B(n16127), .Z(n15813) );
  NOR2_X1 U16046 ( .A1(n8041), .A2(n8968), .ZN(n16127) );
  XOR2_X1 U16047 ( .A(n16128), .B(n16129), .Z(n16126) );
  XNOR2_X1 U16048 ( .A(n16130), .B(n16131), .ZN(n15843) );
  NAND2_X1 U16049 ( .A1(n16132), .A2(n16133), .ZN(n16130) );
  XOR2_X1 U16050 ( .A(n16134), .B(n16135), .Z(n15850) );
  XNOR2_X1 U16051 ( .A(n16136), .B(n16137), .ZN(n16134) );
  NAND2_X1 U16052 ( .A1(b_2_), .A2(a_23_), .ZN(n16136) );
  XOR2_X1 U16053 ( .A(n16138), .B(n16139), .Z(n15859) );
  XOR2_X1 U16054 ( .A(n16140), .B(n16141), .Z(n16138) );
  NOR2_X1 U16055 ( .A1(n8268), .A2(n8968), .ZN(n16141) );
  XOR2_X1 U16056 ( .A(n16142), .B(n16143), .Z(n15867) );
  XNOR2_X1 U16057 ( .A(n16144), .B(n16145), .ZN(n16142) );
  NAND2_X1 U16058 ( .A1(b_2_), .A2(a_19_), .ZN(n16144) );
  XNOR2_X1 U16059 ( .A(n16146), .B(n16147), .ZN(n15875) );
  XNOR2_X1 U16060 ( .A(n16148), .B(n16149), .ZN(n16146) );
  XOR2_X1 U16061 ( .A(n16150), .B(n16151), .Z(n15882) );
  XOR2_X1 U16062 ( .A(n16152), .B(n16153), .Z(n16150) );
  XNOR2_X1 U16063 ( .A(n16154), .B(n16155), .ZN(n15891) );
  XNOR2_X1 U16064 ( .A(n16156), .B(n16157), .ZN(n16154) );
  XNOR2_X1 U16065 ( .A(n16158), .B(n16159), .ZN(n15899) );
  XNOR2_X1 U16066 ( .A(n16160), .B(n16161), .ZN(n16158) );
  XNOR2_X1 U16067 ( .A(n16162), .B(n16163), .ZN(n15907) );
  XNOR2_X1 U16068 ( .A(n16164), .B(n16165), .ZN(n16162) );
  XNOR2_X1 U16069 ( .A(n16166), .B(n16167), .ZN(n15915) );
  XNOR2_X1 U16070 ( .A(n16168), .B(n16169), .ZN(n16166) );
  XNOR2_X1 U16071 ( .A(n16170), .B(n16171), .ZN(n15919) );
  XNOR2_X1 U16072 ( .A(n16172), .B(n16173), .ZN(n16170) );
  INV_X1 U16073 ( .A(n8869), .ZN(n15925) );
  NAND2_X1 U16074 ( .A1(b_3_), .A2(a_3_), .ZN(n8869) );
  XNOR2_X1 U16075 ( .A(n16174), .B(n16175), .ZN(n15927) );
  XNOR2_X1 U16076 ( .A(n16176), .B(n16177), .ZN(n16174) );
  XOR2_X1 U16077 ( .A(n16178), .B(n16179), .Z(n15935) );
  XOR2_X1 U16078 ( .A(n16180), .B(n16181), .Z(n16178) );
  XOR2_X1 U16079 ( .A(n15704), .B(n15703), .Z(n15942) );
  XOR2_X1 U16080 ( .A(n16182), .B(n16183), .Z(n15703) );
  OR2_X1 U16081 ( .A1(n16184), .A2(n16185), .ZN(n15941) );
  NOR2_X1 U16082 ( .A1(n15940), .A2(n15939), .ZN(n16185) );
  AND2_X1 U16083 ( .A1(n16186), .A2(n16184), .ZN(n9056) );
  INV_X1 U16084 ( .A(n9124), .ZN(n16184) );
  NAND2_X1 U16085 ( .A1(n15940), .A2(n15939), .ZN(n9124) );
  NAND2_X1 U16086 ( .A1(n16187), .A2(n16188), .ZN(n15939) );
  NAND2_X1 U16087 ( .A1(n16182), .A2(n16189), .ZN(n16188) );
  OR2_X1 U16088 ( .A1(n16183), .A2(n15704), .ZN(n16189) );
  NOR2_X1 U16089 ( .A1(n8968), .A2(n8974), .ZN(n16182) );
  NAND2_X1 U16090 ( .A1(n15704), .A2(n16183), .ZN(n16187) );
  NAND2_X1 U16091 ( .A1(n16190), .A2(n16191), .ZN(n16183) );
  NAND2_X1 U16092 ( .A1(n16181), .A2(n16192), .ZN(n16191) );
  OR2_X1 U16093 ( .A1(n16180), .A2(n16179), .ZN(n16192) );
  NOR2_X1 U16094 ( .A1(n8968), .A2(n8969), .ZN(n16181) );
  NAND2_X1 U16095 ( .A1(n16179), .A2(n16180), .ZN(n16190) );
  NAND2_X1 U16096 ( .A1(n16193), .A2(n16194), .ZN(n16180) );
  NAND2_X1 U16097 ( .A1(n15951), .A2(n16195), .ZN(n16194) );
  NAND2_X1 U16098 ( .A1(n15952), .A2(n8812), .ZN(n16195) );
  XOR2_X1 U16099 ( .A(n16196), .B(n16197), .Z(n15951) );
  XNOR2_X1 U16100 ( .A(n16198), .B(n16199), .ZN(n16197) );
  NAND2_X1 U16101 ( .A1(b_1_), .A2(a_3_), .ZN(n16196) );
  OR2_X1 U16102 ( .A1(n8812), .A2(n15952), .ZN(n16193) );
  AND2_X1 U16103 ( .A1(n16200), .A2(n16201), .ZN(n15952) );
  NAND2_X1 U16104 ( .A1(n16177), .A2(n16202), .ZN(n16201) );
  NAND2_X1 U16105 ( .A1(n16176), .A2(n16175), .ZN(n16202) );
  NOR2_X1 U16106 ( .A1(n8968), .A2(n8778), .ZN(n16177) );
  OR2_X1 U16107 ( .A1(n16175), .A2(n16176), .ZN(n16200) );
  AND2_X1 U16108 ( .A1(n15962), .A2(n16203), .ZN(n16176) );
  NAND2_X1 U16109 ( .A1(n15961), .A2(n15963), .ZN(n16203) );
  NAND2_X1 U16110 ( .A1(n16204), .A2(n16205), .ZN(n15963) );
  NAND2_X1 U16111 ( .A1(b_2_), .A2(a_4_), .ZN(n16205) );
  INV_X1 U16112 ( .A(n16206), .ZN(n16204) );
  XOR2_X1 U16113 ( .A(n16207), .B(n16208), .Z(n15961) );
  XNOR2_X1 U16114 ( .A(n16209), .B(n16210), .ZN(n16208) );
  NAND2_X1 U16115 ( .A1(b_1_), .A2(a_5_), .ZN(n16207) );
  NAND2_X1 U16116 ( .A1(a_4_), .A2(n16206), .ZN(n15962) );
  NAND2_X1 U16117 ( .A1(n16211), .A2(n16212), .ZN(n16206) );
  NAND2_X1 U16118 ( .A1(n16173), .A2(n16213), .ZN(n16212) );
  NAND2_X1 U16119 ( .A1(n16172), .A2(n16171), .ZN(n16213) );
  NOR2_X1 U16120 ( .A1(n8968), .A2(n8723), .ZN(n16173) );
  OR2_X1 U16121 ( .A1(n16171), .A2(n16172), .ZN(n16211) );
  AND2_X1 U16122 ( .A1(n15974), .A2(n16214), .ZN(n16172) );
  NAND2_X1 U16123 ( .A1(n15973), .A2(n15975), .ZN(n16214) );
  NAND2_X1 U16124 ( .A1(n16215), .A2(n16216), .ZN(n15975) );
  NAND2_X1 U16125 ( .A1(b_2_), .A2(a_6_), .ZN(n16216) );
  INV_X1 U16126 ( .A(n16217), .ZN(n16215) );
  XOR2_X1 U16127 ( .A(n16218), .B(n16219), .Z(n15973) );
  XNOR2_X1 U16128 ( .A(n16220), .B(n16221), .ZN(n16219) );
  NAND2_X1 U16129 ( .A1(b_1_), .A2(a_7_), .ZN(n16218) );
  NAND2_X1 U16130 ( .A1(a_6_), .A2(n16217), .ZN(n15974) );
  NAND2_X1 U16131 ( .A1(n16222), .A2(n16223), .ZN(n16217) );
  NAND2_X1 U16132 ( .A1(n16169), .A2(n16224), .ZN(n16223) );
  NAND2_X1 U16133 ( .A1(n16168), .A2(n16167), .ZN(n16224) );
  NOR2_X1 U16134 ( .A1(n8968), .A2(n8962), .ZN(n16169) );
  OR2_X1 U16135 ( .A1(n16167), .A2(n16168), .ZN(n16222) );
  AND2_X1 U16136 ( .A1(n15986), .A2(n16225), .ZN(n16168) );
  NAND2_X1 U16137 ( .A1(n15985), .A2(n15987), .ZN(n16225) );
  NAND2_X1 U16138 ( .A1(n16226), .A2(n16227), .ZN(n15987) );
  NAND2_X1 U16139 ( .A1(b_2_), .A2(a_8_), .ZN(n16227) );
  INV_X1 U16140 ( .A(n16228), .ZN(n16226) );
  XOR2_X1 U16141 ( .A(n16229), .B(n16230), .Z(n15985) );
  XNOR2_X1 U16142 ( .A(n16231), .B(n16232), .ZN(n16230) );
  NAND2_X1 U16143 ( .A1(b_1_), .A2(a_9_), .ZN(n16229) );
  NAND2_X1 U16144 ( .A1(a_8_), .A2(n16228), .ZN(n15986) );
  NAND2_X1 U16145 ( .A1(n16233), .A2(n16234), .ZN(n16228) );
  NAND2_X1 U16146 ( .A1(n16165), .A2(n16235), .ZN(n16234) );
  NAND2_X1 U16147 ( .A1(n16164), .A2(n16163), .ZN(n16235) );
  NOR2_X1 U16148 ( .A1(n8968), .A2(n8605), .ZN(n16165) );
  OR2_X1 U16149 ( .A1(n16163), .A2(n16164), .ZN(n16233) );
  AND2_X1 U16150 ( .A1(n15998), .A2(n16236), .ZN(n16164) );
  NAND2_X1 U16151 ( .A1(n15997), .A2(n15999), .ZN(n16236) );
  NAND2_X1 U16152 ( .A1(n16237), .A2(n16238), .ZN(n15999) );
  NAND2_X1 U16153 ( .A1(b_2_), .A2(a_10_), .ZN(n16238) );
  INV_X1 U16154 ( .A(n16239), .ZN(n16237) );
  XOR2_X1 U16155 ( .A(n16240), .B(n16241), .Z(n15997) );
  XNOR2_X1 U16156 ( .A(n16242), .B(n16243), .ZN(n16241) );
  NAND2_X1 U16157 ( .A1(b_1_), .A2(a_11_), .ZN(n16240) );
  NAND2_X1 U16158 ( .A1(a_10_), .A2(n16239), .ZN(n15998) );
  NAND2_X1 U16159 ( .A1(n16244), .A2(n16245), .ZN(n16239) );
  NAND2_X1 U16160 ( .A1(n16161), .A2(n16246), .ZN(n16245) );
  NAND2_X1 U16161 ( .A1(n16160), .A2(n16159), .ZN(n16246) );
  NOR2_X1 U16162 ( .A1(n8968), .A2(n8550), .ZN(n16161) );
  OR2_X1 U16163 ( .A1(n16159), .A2(n16160), .ZN(n16244) );
  AND2_X1 U16164 ( .A1(n16010), .A2(n16247), .ZN(n16160) );
  NAND2_X1 U16165 ( .A1(n16009), .A2(n16011), .ZN(n16247) );
  NAND2_X1 U16166 ( .A1(n16248), .A2(n16249), .ZN(n16011) );
  NAND2_X1 U16167 ( .A1(b_2_), .A2(a_12_), .ZN(n16249) );
  INV_X1 U16168 ( .A(n16250), .ZN(n16248) );
  XOR2_X1 U16169 ( .A(n16251), .B(n16252), .Z(n16009) );
  XNOR2_X1 U16170 ( .A(n16253), .B(n16254), .ZN(n16252) );
  NAND2_X1 U16171 ( .A1(b_1_), .A2(a_13_), .ZN(n16251) );
  NAND2_X1 U16172 ( .A1(a_12_), .A2(n16250), .ZN(n16010) );
  NAND2_X1 U16173 ( .A1(n16255), .A2(n16256), .ZN(n16250) );
  NAND2_X1 U16174 ( .A1(n16157), .A2(n16257), .ZN(n16256) );
  NAND2_X1 U16175 ( .A1(n16156), .A2(n16155), .ZN(n16257) );
  NOR2_X1 U16176 ( .A1(n8968), .A2(n8495), .ZN(n16157) );
  OR2_X1 U16177 ( .A1(n16155), .A2(n16156), .ZN(n16255) );
  AND2_X1 U16178 ( .A1(n16022), .A2(n16258), .ZN(n16156) );
  NAND2_X1 U16179 ( .A1(n16021), .A2(n16023), .ZN(n16258) );
  NAND2_X1 U16180 ( .A1(n16259), .A2(n16260), .ZN(n16023) );
  NAND2_X1 U16181 ( .A1(b_2_), .A2(a_14_), .ZN(n16260) );
  INV_X1 U16182 ( .A(n16261), .ZN(n16259) );
  XOR2_X1 U16183 ( .A(n16262), .B(n16263), .Z(n16021) );
  XNOR2_X1 U16184 ( .A(n16264), .B(n16265), .ZN(n16263) );
  NAND2_X1 U16185 ( .A1(b_1_), .A2(a_15_), .ZN(n16262) );
  NAND2_X1 U16186 ( .A1(a_14_), .A2(n16261), .ZN(n16022) );
  NAND2_X1 U16187 ( .A1(n16266), .A2(n16267), .ZN(n16261) );
  NAND2_X1 U16188 ( .A1(n16153), .A2(n16268), .ZN(n16267) );
  OR2_X1 U16189 ( .A1(n16152), .A2(n16151), .ZN(n16268) );
  NOR2_X1 U16190 ( .A1(n8968), .A2(n8440), .ZN(n16153) );
  NAND2_X1 U16191 ( .A1(n16151), .A2(n16152), .ZN(n16266) );
  NAND2_X1 U16192 ( .A1(n16034), .A2(n16269), .ZN(n16152) );
  NAND2_X1 U16193 ( .A1(n16033), .A2(n16035), .ZN(n16269) );
  NAND2_X1 U16194 ( .A1(n16270), .A2(n16271), .ZN(n16035) );
  NAND2_X1 U16195 ( .A1(b_2_), .A2(a_16_), .ZN(n16271) );
  INV_X1 U16196 ( .A(n16272), .ZN(n16270) );
  XOR2_X1 U16197 ( .A(n16273), .B(n16274), .Z(n16033) );
  XNOR2_X1 U16198 ( .A(n16275), .B(n16276), .ZN(n16274) );
  NAND2_X1 U16199 ( .A1(b_1_), .A2(a_17_), .ZN(n16273) );
  NAND2_X1 U16200 ( .A1(a_16_), .A2(n16272), .ZN(n16034) );
  NAND2_X1 U16201 ( .A1(n16277), .A2(n16278), .ZN(n16272) );
  NAND2_X1 U16202 ( .A1(n16149), .A2(n16279), .ZN(n16278) );
  NAND2_X1 U16203 ( .A1(n16148), .A2(n16147), .ZN(n16279) );
  NOR2_X1 U16204 ( .A1(n8968), .A2(n8385), .ZN(n16149) );
  OR2_X1 U16205 ( .A1(n16147), .A2(n16148), .ZN(n16277) );
  AND2_X1 U16206 ( .A1(n16280), .A2(n16281), .ZN(n16148) );
  NAND2_X1 U16207 ( .A1(n16047), .A2(n16282), .ZN(n16281) );
  NAND2_X1 U16208 ( .A1(n16046), .A2(n16045), .ZN(n16282) );
  NOR2_X1 U16209 ( .A1(n8968), .A2(n8947), .ZN(n16047) );
  OR2_X1 U16210 ( .A1(n16045), .A2(n16046), .ZN(n16280) );
  AND2_X1 U16211 ( .A1(n16283), .A2(n16284), .ZN(n16046) );
  NAND2_X1 U16212 ( .A1(n16285), .A2(b_2_), .ZN(n16284) );
  NOR2_X1 U16213 ( .A1(n16286), .A2(n8324), .ZN(n16285) );
  NOR2_X1 U16214 ( .A1(n16143), .A2(n16145), .ZN(n16286) );
  NAND2_X1 U16215 ( .A1(n16143), .A2(n16145), .ZN(n16283) );
  NAND2_X1 U16216 ( .A1(n16287), .A2(n16288), .ZN(n16145) );
  NAND2_X1 U16217 ( .A1(n16059), .A2(n16289), .ZN(n16288) );
  NAND2_X1 U16218 ( .A1(n16058), .A2(n16057), .ZN(n16289) );
  NOR2_X1 U16219 ( .A1(n8968), .A2(n8944), .ZN(n16059) );
  OR2_X1 U16220 ( .A1(n16057), .A2(n16058), .ZN(n16287) );
  AND2_X1 U16221 ( .A1(n16290), .A2(n16291), .ZN(n16058) );
  NAND2_X1 U16222 ( .A1(n16292), .A2(b_2_), .ZN(n16291) );
  NOR2_X1 U16223 ( .A1(n16293), .A2(n8268), .ZN(n16292) );
  NOR2_X1 U16224 ( .A1(n16139), .A2(n16140), .ZN(n16293) );
  NAND2_X1 U16225 ( .A1(n16139), .A2(n16140), .ZN(n16290) );
  NAND2_X1 U16226 ( .A1(n16294), .A2(n16295), .ZN(n16140) );
  NAND2_X1 U16227 ( .A1(n16071), .A2(n16296), .ZN(n16295) );
  OR2_X1 U16228 ( .A1(n16070), .A2(n16068), .ZN(n16296) );
  NOR2_X1 U16229 ( .A1(n8968), .A2(n8941), .ZN(n16071) );
  NAND2_X1 U16230 ( .A1(n16068), .A2(n16070), .ZN(n16294) );
  NAND2_X1 U16231 ( .A1(n16297), .A2(n16298), .ZN(n16070) );
  NAND2_X1 U16232 ( .A1(n16299), .A2(b_2_), .ZN(n16298) );
  NOR2_X1 U16233 ( .A1(n16300), .A2(n8213), .ZN(n16299) );
  NOR2_X1 U16234 ( .A1(n16135), .A2(n16137), .ZN(n16300) );
  NAND2_X1 U16235 ( .A1(n16135), .A2(n16137), .ZN(n16297) );
  NAND2_X1 U16236 ( .A1(n16301), .A2(n16302), .ZN(n16137) );
  NAND2_X1 U16237 ( .A1(n16083), .A2(n16303), .ZN(n16302) );
  OR2_X1 U16238 ( .A1(n16082), .A2(n16080), .ZN(n16303) );
  NOR2_X1 U16239 ( .A1(n8968), .A2(n8939), .ZN(n16083) );
  NAND2_X1 U16240 ( .A1(n16080), .A2(n16082), .ZN(n16301) );
  NAND2_X1 U16241 ( .A1(n16132), .A2(n16304), .ZN(n16082) );
  NAND2_X1 U16242 ( .A1(n16131), .A2(n16133), .ZN(n16304) );
  NAND2_X1 U16243 ( .A1(n16305), .A2(n16306), .ZN(n16133) );
  NAND2_X1 U16244 ( .A1(b_2_), .A2(a_25_), .ZN(n16306) );
  INV_X1 U16245 ( .A(n16307), .ZN(n16305) );
  XNOR2_X1 U16246 ( .A(n16308), .B(n16309), .ZN(n16131) );
  NAND2_X1 U16247 ( .A1(n16310), .A2(n16311), .ZN(n16308) );
  NAND2_X1 U16248 ( .A1(n16312), .A2(n16313), .ZN(n16311) );
  NAND2_X1 U16249 ( .A1(b_0_), .A2(a_27_), .ZN(n16312) );
  NAND2_X1 U16250 ( .A1(a_25_), .A2(n16307), .ZN(n16132) );
  NAND2_X1 U16251 ( .A1(n16314), .A2(n16315), .ZN(n16307) );
  NAND2_X1 U16252 ( .A1(n16316), .A2(b_2_), .ZN(n16315) );
  NOR2_X1 U16253 ( .A1(n16317), .A2(n8116), .ZN(n16316) );
  NOR2_X1 U16254 ( .A1(n16093), .A2(n16095), .ZN(n16317) );
  NAND2_X1 U16255 ( .A1(n16093), .A2(n16095), .ZN(n16314) );
  NAND2_X1 U16256 ( .A1(n16318), .A2(n16319), .ZN(n16095) );
  NAND2_X1 U16257 ( .A1(n16103), .A2(n16320), .ZN(n16319) );
  OR2_X1 U16258 ( .A1(n16102), .A2(n16100), .ZN(n16320) );
  NOR2_X1 U16259 ( .A1(n8968), .A2(n8937), .ZN(n16103) );
  NAND2_X1 U16260 ( .A1(n16100), .A2(n16102), .ZN(n16318) );
  NAND2_X1 U16261 ( .A1(n16321), .A2(n16322), .ZN(n16102) );
  NAND2_X1 U16262 ( .A1(n16323), .A2(b_2_), .ZN(n16322) );
  NOR2_X1 U16263 ( .A1(n16324), .A2(n8055), .ZN(n16323) );
  NOR2_X1 U16264 ( .A1(n16110), .A2(n16108), .ZN(n16324) );
  NAND2_X1 U16265 ( .A1(n16108), .A2(n16110), .ZN(n16321) );
  NAND2_X1 U16266 ( .A1(n16325), .A2(n16326), .ZN(n16110) );
  NAND2_X1 U16267 ( .A1(n16327), .A2(b_2_), .ZN(n16326) );
  NOR2_X1 U16268 ( .A1(n16328), .A2(n8041), .ZN(n16327) );
  NOR2_X1 U16269 ( .A1(n16129), .A2(n16128), .ZN(n16328) );
  NAND2_X1 U16270 ( .A1(n16129), .A2(n16128), .ZN(n16325) );
  NAND2_X1 U16271 ( .A1(n16329), .A2(n16330), .ZN(n16128) );
  NAND2_X1 U16272 ( .A1(b_0_), .A2(n16331), .ZN(n16330) );
  NAND2_X1 U16273 ( .A1(n8003), .A2(n16332), .ZN(n16331) );
  NAND2_X1 U16274 ( .A1(a_31_), .A2(n8834), .ZN(n16332) );
  NAND2_X1 U16275 ( .A1(b_1_), .A2(n16333), .ZN(n16329) );
  NAND2_X1 U16276 ( .A1(n9341), .A2(n16334), .ZN(n16333) );
  NAND2_X1 U16277 ( .A1(a_30_), .A2(n8975), .ZN(n16334) );
  AND2_X1 U16278 ( .A1(n16336), .A2(n7953), .ZN(n16129) );
  NOR2_X1 U16279 ( .A1(n8968), .A2(n8834), .ZN(n16336) );
  XNOR2_X1 U16280 ( .A(n16337), .B(n16338), .ZN(n16108) );
  XOR2_X1 U16281 ( .A(n16339), .B(n16340), .Z(n16337) );
  XOR2_X1 U16282 ( .A(n16341), .B(n16342), .Z(n16100) );
  NOR2_X1 U16283 ( .A1(n8041), .A2(n8975), .ZN(n16342) );
  XOR2_X1 U16284 ( .A(n16343), .B(n16344), .Z(n16341) );
  XOR2_X1 U16285 ( .A(n16345), .B(n16346), .Z(n16093) );
  NOR2_X1 U16286 ( .A1(n8055), .A2(n8975), .ZN(n16346) );
  XOR2_X1 U16287 ( .A(n16347), .B(n16348), .Z(n16345) );
  XOR2_X1 U16288 ( .A(n16349), .B(n16350), .Z(n16080) );
  XNOR2_X1 U16289 ( .A(n16351), .B(n16352), .ZN(n16350) );
  NAND2_X1 U16290 ( .A1(b_0_), .A2(a_26_), .ZN(n16349) );
  XNOR2_X1 U16291 ( .A(n16353), .B(n16354), .ZN(n16135) );
  NAND2_X1 U16292 ( .A1(n16355), .A2(n16356), .ZN(n16353) );
  NAND2_X1 U16293 ( .A1(n16357), .A2(n16358), .ZN(n16356) );
  NAND2_X1 U16294 ( .A1(b_0_), .A2(a_25_), .ZN(n16357) );
  XOR2_X1 U16295 ( .A(n16359), .B(n16360), .Z(n16068) );
  XNOR2_X1 U16296 ( .A(n16361), .B(n16362), .ZN(n16360) );
  NAND2_X1 U16297 ( .A1(b_0_), .A2(a_24_), .ZN(n16359) );
  XNOR2_X1 U16298 ( .A(n16363), .B(n16364), .ZN(n16139) );
  NAND2_X1 U16299 ( .A1(n16365), .A2(n16366), .ZN(n16363) );
  NAND2_X1 U16300 ( .A1(n16367), .A2(n16368), .ZN(n16366) );
  NAND2_X1 U16301 ( .A1(b_0_), .A2(a_23_), .ZN(n16367) );
  XNOR2_X1 U16302 ( .A(n16369), .B(n16370), .ZN(n16057) );
  XNOR2_X1 U16303 ( .A(n16371), .B(n16372), .ZN(n16370) );
  NAND2_X1 U16304 ( .A1(b_0_), .A2(a_22_), .ZN(n16369) );
  XNOR2_X1 U16305 ( .A(n16373), .B(n16374), .ZN(n16143) );
  NAND2_X1 U16306 ( .A1(n16375), .A2(n16376), .ZN(n16373) );
  NAND2_X1 U16307 ( .A1(n16377), .A2(n16378), .ZN(n16376) );
  NAND2_X1 U16308 ( .A1(b_0_), .A2(a_21_), .ZN(n16377) );
  XNOR2_X1 U16309 ( .A(n16379), .B(n16380), .ZN(n16045) );
  XNOR2_X1 U16310 ( .A(n16381), .B(n16382), .ZN(n16380) );
  NAND2_X1 U16311 ( .A1(b_0_), .A2(a_20_), .ZN(n16379) );
  XOR2_X1 U16312 ( .A(n16383), .B(n16384), .Z(n16147) );
  NAND2_X1 U16313 ( .A1(n16385), .A2(n16386), .ZN(n16383) );
  NAND2_X1 U16314 ( .A1(n16387), .A2(n16388), .ZN(n16386) );
  NAND2_X1 U16315 ( .A1(b_0_), .A2(a_19_), .ZN(n16387) );
  XNOR2_X1 U16316 ( .A(n16389), .B(n16390), .ZN(n16151) );
  NAND2_X1 U16317 ( .A1(n16391), .A2(n16392), .ZN(n16389) );
  NAND2_X1 U16318 ( .A1(n16393), .A2(n16394), .ZN(n16392) );
  NAND2_X1 U16319 ( .A1(b_1_), .A2(a_16_), .ZN(n16393) );
  XOR2_X1 U16320 ( .A(n16395), .B(n16396), .Z(n16155) );
  NAND2_X1 U16321 ( .A1(n16397), .A2(n16398), .ZN(n16395) );
  NAND2_X1 U16322 ( .A1(n16399), .A2(n16400), .ZN(n16398) );
  NAND2_X1 U16323 ( .A1(b_1_), .A2(a_14_), .ZN(n16399) );
  XNOR2_X1 U16324 ( .A(n16401), .B(n16402), .ZN(n16159) );
  NOR2_X1 U16325 ( .A1(n16403), .A2(n16404), .ZN(n16402) );
  INV_X1 U16326 ( .A(n16405), .ZN(n16404) );
  NOR2_X1 U16327 ( .A1(n16406), .A2(n16407), .ZN(n16403) );
  XNOR2_X1 U16328 ( .A(n16408), .B(n16409), .ZN(n16163) );
  NOR2_X1 U16329 ( .A1(n16410), .A2(n16411), .ZN(n16409) );
  INV_X1 U16330 ( .A(n16412), .ZN(n16411) );
  NOR2_X1 U16331 ( .A1(n16413), .A2(n16414), .ZN(n16410) );
  XNOR2_X1 U16332 ( .A(n16415), .B(n16416), .ZN(n16167) );
  NOR2_X1 U16333 ( .A1(n16417), .A2(n16418), .ZN(n16416) );
  INV_X1 U16334 ( .A(n16419), .ZN(n16418) );
  NOR2_X1 U16335 ( .A1(n16420), .A2(n16421), .ZN(n16417) );
  XNOR2_X1 U16336 ( .A(n16422), .B(n16423), .ZN(n16171) );
  NOR2_X1 U16337 ( .A1(n16424), .A2(n16425), .ZN(n16423) );
  INV_X1 U16338 ( .A(n16426), .ZN(n16425) );
  NOR2_X1 U16339 ( .A1(n16427), .A2(n16428), .ZN(n16424) );
  XNOR2_X1 U16340 ( .A(n16429), .B(n16430), .ZN(n16175) );
  NOR2_X1 U16341 ( .A1(n16431), .A2(n16432), .ZN(n16430) );
  INV_X1 U16342 ( .A(n16433), .ZN(n16432) );
  NOR2_X1 U16343 ( .A1(n16434), .A2(n16435), .ZN(n16431) );
  NAND2_X1 U16344 ( .A1(b_2_), .A2(a_2_), .ZN(n8812) );
  XOR2_X1 U16345 ( .A(n16436), .B(n16437), .Z(n16179) );
  NOR2_X1 U16346 ( .A1(n16438), .A2(n16439), .ZN(n16437) );
  INV_X1 U16347 ( .A(n16440), .ZN(n16439) );
  NOR2_X1 U16348 ( .A1(n16441), .A2(n16442), .ZN(n16438) );
  XOR2_X1 U16349 ( .A(n16443), .B(n16444), .Z(n15704) );
  XNOR2_X1 U16350 ( .A(n8867), .B(n16445), .ZN(n16444) );
  NAND2_X1 U16351 ( .A1(b_0_), .A2(a_2_), .ZN(n16443) );
  XOR2_X1 U16352 ( .A(n16446), .B(n16447), .Z(n15940) );
  NOR2_X1 U16353 ( .A1(n16448), .A2(n16449), .ZN(n16447) );
  INV_X1 U16354 ( .A(n16450), .ZN(n16449) );
  NOR2_X1 U16355 ( .A1(n16451), .A2(n16452), .ZN(n16448) );
  NOR2_X1 U16356 ( .A1(n8972), .A2(n9121), .ZN(n16186) );
  NAND2_X1 U16357 ( .A1(n16450), .A2(n16453), .ZN(n9121) );
  NAND2_X1 U16358 ( .A1(n16454), .A2(n16446), .ZN(n16453) );
  NAND2_X1 U16359 ( .A1(n16455), .A2(n16456), .ZN(n16446) );
  NAND2_X1 U16360 ( .A1(n16457), .A2(b_0_), .ZN(n16456) );
  NOR2_X1 U16361 ( .A1(n16458), .A2(n8792), .ZN(n16457) );
  NOR2_X1 U16362 ( .A1(n8867), .A2(n16445), .ZN(n16458) );
  NAND2_X1 U16363 ( .A1(n8867), .A2(n16445), .ZN(n16455) );
  NAND2_X1 U16364 ( .A1(n16440), .A2(n16459), .ZN(n16445) );
  NAND2_X1 U16365 ( .A1(n16460), .A2(n16436), .ZN(n16459) );
  NAND2_X1 U16366 ( .A1(n16461), .A2(n16462), .ZN(n16436) );
  NAND2_X1 U16367 ( .A1(n16463), .A2(b_1_), .ZN(n16462) );
  NOR2_X1 U16368 ( .A1(n16464), .A2(n8778), .ZN(n16463) );
  NOR2_X1 U16369 ( .A1(n16198), .A2(n16199), .ZN(n16464) );
  NAND2_X1 U16370 ( .A1(n16198), .A2(n16199), .ZN(n16461) );
  NAND2_X1 U16371 ( .A1(n16433), .A2(n16465), .ZN(n16199) );
  NAND2_X1 U16372 ( .A1(n16466), .A2(n16429), .ZN(n16465) );
  NAND2_X1 U16373 ( .A1(n16467), .A2(n16468), .ZN(n16429) );
  NAND2_X1 U16374 ( .A1(n16469), .A2(b_1_), .ZN(n16468) );
  NOR2_X1 U16375 ( .A1(n16470), .A2(n8723), .ZN(n16469) );
  NOR2_X1 U16376 ( .A1(n16209), .A2(n16210), .ZN(n16470) );
  NAND2_X1 U16377 ( .A1(n16209), .A2(n16210), .ZN(n16467) );
  NAND2_X1 U16378 ( .A1(n16426), .A2(n16471), .ZN(n16210) );
  NAND2_X1 U16379 ( .A1(n16472), .A2(n16422), .ZN(n16471) );
  NAND2_X1 U16380 ( .A1(n16473), .A2(n16474), .ZN(n16422) );
  NAND2_X1 U16381 ( .A1(n16475), .A2(b_1_), .ZN(n16474) );
  NOR2_X1 U16382 ( .A1(n16476), .A2(n8962), .ZN(n16475) );
  NOR2_X1 U16383 ( .A1(n16220), .A2(n16221), .ZN(n16476) );
  NAND2_X1 U16384 ( .A1(n16220), .A2(n16221), .ZN(n16473) );
  NAND2_X1 U16385 ( .A1(n16419), .A2(n16477), .ZN(n16221) );
  NAND2_X1 U16386 ( .A1(n16478), .A2(n16415), .ZN(n16477) );
  NAND2_X1 U16387 ( .A1(n16479), .A2(n16480), .ZN(n16415) );
  NAND2_X1 U16388 ( .A1(n16481), .A2(b_1_), .ZN(n16480) );
  NOR2_X1 U16389 ( .A1(n16482), .A2(n8605), .ZN(n16481) );
  NOR2_X1 U16390 ( .A1(n16231), .A2(n16232), .ZN(n16482) );
  NAND2_X1 U16391 ( .A1(n16231), .A2(n16232), .ZN(n16479) );
  NAND2_X1 U16392 ( .A1(n16412), .A2(n16483), .ZN(n16232) );
  NAND2_X1 U16393 ( .A1(n16484), .A2(n16408), .ZN(n16483) );
  NAND2_X1 U16394 ( .A1(n16485), .A2(n16486), .ZN(n16408) );
  NAND2_X1 U16395 ( .A1(n16487), .A2(b_1_), .ZN(n16486) );
  NOR2_X1 U16396 ( .A1(n16488), .A2(n8550), .ZN(n16487) );
  NOR2_X1 U16397 ( .A1(n16242), .A2(n16243), .ZN(n16488) );
  NAND2_X1 U16398 ( .A1(n16242), .A2(n16243), .ZN(n16485) );
  NAND2_X1 U16399 ( .A1(n16405), .A2(n16489), .ZN(n16243) );
  NAND2_X1 U16400 ( .A1(n16490), .A2(n16401), .ZN(n16489) );
  NAND2_X1 U16401 ( .A1(n16491), .A2(n16492), .ZN(n16401) );
  NAND2_X1 U16402 ( .A1(n16493), .A2(b_1_), .ZN(n16492) );
  NOR2_X1 U16403 ( .A1(n16494), .A2(n8495), .ZN(n16493) );
  NOR2_X1 U16404 ( .A1(n16253), .A2(n16254), .ZN(n16494) );
  NAND2_X1 U16405 ( .A1(n16253), .A2(n16254), .ZN(n16491) );
  NAND2_X1 U16406 ( .A1(n16397), .A2(n16495), .ZN(n16254) );
  NAND2_X1 U16407 ( .A1(n16496), .A2(n16396), .ZN(n16495) );
  NAND2_X1 U16408 ( .A1(n16497), .A2(n16498), .ZN(n16396) );
  NAND2_X1 U16409 ( .A1(n16499), .A2(b_1_), .ZN(n16498) );
  NOR2_X1 U16410 ( .A1(n16500), .A2(n8440), .ZN(n16499) );
  NOR2_X1 U16411 ( .A1(n16264), .A2(n16265), .ZN(n16500) );
  NAND2_X1 U16412 ( .A1(n16264), .A2(n16265), .ZN(n16497) );
  NAND2_X1 U16413 ( .A1(n16391), .A2(n16501), .ZN(n16265) );
  NAND2_X1 U16414 ( .A1(n16502), .A2(n16390), .ZN(n16501) );
  NAND2_X1 U16415 ( .A1(n16503), .A2(n16504), .ZN(n16390) );
  NAND2_X1 U16416 ( .A1(n16505), .A2(b_1_), .ZN(n16504) );
  NOR2_X1 U16417 ( .A1(n16506), .A2(n8385), .ZN(n16505) );
  NOR2_X1 U16418 ( .A1(n16275), .A2(n16276), .ZN(n16506) );
  NAND2_X1 U16419 ( .A1(n16275), .A2(n16276), .ZN(n16503) );
  NAND2_X1 U16420 ( .A1(n16385), .A2(n16507), .ZN(n16276) );
  NAND2_X1 U16421 ( .A1(n16508), .A2(n16384), .ZN(n16507) );
  NAND2_X1 U16422 ( .A1(n16509), .A2(n16510), .ZN(n16384) );
  NAND2_X1 U16423 ( .A1(n16511), .A2(b_0_), .ZN(n16510) );
  NOR2_X1 U16424 ( .A1(n16512), .A2(n8944), .ZN(n16511) );
  NOR2_X1 U16425 ( .A1(n16381), .A2(n16382), .ZN(n16512) );
  NAND2_X1 U16426 ( .A1(n16381), .A2(n16382), .ZN(n16509) );
  NAND2_X1 U16427 ( .A1(n16375), .A2(n16513), .ZN(n16382) );
  NAND2_X1 U16428 ( .A1(n16514), .A2(n16374), .ZN(n16513) );
  NAND2_X1 U16429 ( .A1(n16515), .A2(n16516), .ZN(n16374) );
  NAND2_X1 U16430 ( .A1(n16517), .A2(b_0_), .ZN(n16516) );
  NOR2_X1 U16431 ( .A1(n16518), .A2(n8941), .ZN(n16517) );
  NOR2_X1 U16432 ( .A1(n16371), .A2(n16372), .ZN(n16518) );
  NAND2_X1 U16433 ( .A1(n16371), .A2(n16372), .ZN(n16515) );
  NAND2_X1 U16434 ( .A1(n16365), .A2(n16519), .ZN(n16372) );
  NAND2_X1 U16435 ( .A1(n16520), .A2(n16364), .ZN(n16519) );
  NAND2_X1 U16436 ( .A1(n16521), .A2(n16522), .ZN(n16364) );
  NAND2_X1 U16437 ( .A1(n16523), .A2(b_0_), .ZN(n16522) );
  NOR2_X1 U16438 ( .A1(n16524), .A2(n8939), .ZN(n16523) );
  NOR2_X1 U16439 ( .A1(n16361), .A2(n16362), .ZN(n16524) );
  NAND2_X1 U16440 ( .A1(n16361), .A2(n16362), .ZN(n16521) );
  NAND2_X1 U16441 ( .A1(n16355), .A2(n16525), .ZN(n16362) );
  NAND2_X1 U16442 ( .A1(n16526), .A2(n16354), .ZN(n16525) );
  NAND2_X1 U16443 ( .A1(n16527), .A2(n16528), .ZN(n16354) );
  NAND2_X1 U16444 ( .A1(n16529), .A2(b_0_), .ZN(n16528) );
  NOR2_X1 U16445 ( .A1(n16530), .A2(n8116), .ZN(n16529) );
  NOR2_X1 U16446 ( .A1(n16351), .A2(n16352), .ZN(n16530) );
  NAND2_X1 U16447 ( .A1(n16351), .A2(n16352), .ZN(n16527) );
  NAND2_X1 U16448 ( .A1(n16310), .A2(n16531), .ZN(n16352) );
  NAND2_X1 U16449 ( .A1(n16532), .A2(n16309), .ZN(n16531) );
  NAND2_X1 U16450 ( .A1(n16533), .A2(n16534), .ZN(n16309) );
  NAND2_X1 U16451 ( .A1(n16535), .A2(b_0_), .ZN(n16534) );
  NOR2_X1 U16452 ( .A1(n16536), .A2(n8055), .ZN(n16535) );
  NOR2_X1 U16453 ( .A1(n16347), .A2(n16348), .ZN(n16536) );
  NAND2_X1 U16454 ( .A1(n16347), .A2(n16348), .ZN(n16533) );
  NAND2_X1 U16455 ( .A1(n16537), .A2(n16538), .ZN(n16348) );
  NAND2_X1 U16456 ( .A1(n16539), .A2(b_0_), .ZN(n16538) );
  NOR2_X1 U16457 ( .A1(n16540), .A2(n8041), .ZN(n16539) );
  NOR2_X1 U16458 ( .A1(n16343), .A2(n16344), .ZN(n16540) );
  NAND2_X1 U16459 ( .A1(n16343), .A2(n16344), .ZN(n16537) );
  NAND2_X1 U16460 ( .A1(n16340), .A2(n16541), .ZN(n16344) );
  NAND2_X1 U16461 ( .A1(n16338), .A2(n16339), .ZN(n16541) );
  NOR2_X1 U16462 ( .A1(n8834), .A2(n8041), .ZN(n16339) );
  NOR2_X1 U16463 ( .A1(n8935), .A2(n8975), .ZN(n16338) );
  NAND2_X1 U16464 ( .A1(n16542), .A2(n7953), .ZN(n16340) );
  NOR2_X1 U16465 ( .A1(n8834), .A2(n8975), .ZN(n16542) );
  NOR2_X1 U16466 ( .A1(n8834), .A2(n8055), .ZN(n16343) );
  NOR2_X1 U16467 ( .A1(n8834), .A2(n8937), .ZN(n16347) );
  NAND2_X1 U16468 ( .A1(n16313), .A2(n8937), .ZN(n16532) );
  NAND2_X1 U16469 ( .A1(n16543), .A2(n16544), .ZN(n16310) );
  INV_X1 U16470 ( .A(n16313), .ZN(n16544) );
  NAND2_X1 U16471 ( .A1(b_1_), .A2(a_26_), .ZN(n16313) );
  NOR2_X1 U16472 ( .A1(n8937), .A2(n8975), .ZN(n16543) );
  NOR2_X1 U16473 ( .A1(n8834), .A2(n8158), .ZN(n16351) );
  NAND2_X1 U16474 ( .A1(n16358), .A2(n8158), .ZN(n16526) );
  NAND2_X1 U16475 ( .A1(n16545), .A2(n16546), .ZN(n16355) );
  INV_X1 U16476 ( .A(n16358), .ZN(n16546) );
  NAND2_X1 U16477 ( .A1(b_1_), .A2(a_24_), .ZN(n16358) );
  NOR2_X1 U16478 ( .A1(n8158), .A2(n8975), .ZN(n16545) );
  NOR2_X1 U16479 ( .A1(n8834), .A2(n8213), .ZN(n16361) );
  NAND2_X1 U16480 ( .A1(n16368), .A2(n8213), .ZN(n16520) );
  NAND2_X1 U16481 ( .A1(n16547), .A2(n16548), .ZN(n16365) );
  INV_X1 U16482 ( .A(n16368), .ZN(n16548) );
  NAND2_X1 U16483 ( .A1(b_1_), .A2(a_22_), .ZN(n16368) );
  NOR2_X1 U16484 ( .A1(n8213), .A2(n8975), .ZN(n16547) );
  NOR2_X1 U16485 ( .A1(n8834), .A2(n8268), .ZN(n16371) );
  NAND2_X1 U16486 ( .A1(n16378), .A2(n8268), .ZN(n16514) );
  NAND2_X1 U16487 ( .A1(n16549), .A2(n16550), .ZN(n16375) );
  INV_X1 U16488 ( .A(n16378), .ZN(n16550) );
  NAND2_X1 U16489 ( .A1(b_1_), .A2(a_20_), .ZN(n16378) );
  NOR2_X1 U16490 ( .A1(n8268), .A2(n8975), .ZN(n16549) );
  NOR2_X1 U16491 ( .A1(n8834), .A2(n8324), .ZN(n16381) );
  NAND2_X1 U16492 ( .A1(n16388), .A2(n8324), .ZN(n16508) );
  NAND2_X1 U16493 ( .A1(n16551), .A2(n16552), .ZN(n16385) );
  INV_X1 U16494 ( .A(n16388), .ZN(n16552) );
  NAND2_X1 U16495 ( .A1(b_1_), .A2(a_18_), .ZN(n16388) );
  NOR2_X1 U16496 ( .A1(n8324), .A2(n8975), .ZN(n16551) );
  NOR2_X1 U16497 ( .A1(n8975), .A2(n8947), .ZN(n16275) );
  NAND2_X1 U16498 ( .A1(n16394), .A2(n8950), .ZN(n16502) );
  NAND2_X1 U16499 ( .A1(n16553), .A2(n16554), .ZN(n16391) );
  INV_X1 U16500 ( .A(n16394), .ZN(n16554) );
  NAND2_X1 U16501 ( .A1(b_0_), .A2(a_17_), .ZN(n16394) );
  NOR2_X1 U16502 ( .A1(n8950), .A2(n8834), .ZN(n16553) );
  NOR2_X1 U16503 ( .A1(n8975), .A2(n8950), .ZN(n16264) );
  NAND2_X1 U16504 ( .A1(n16400), .A2(n8953), .ZN(n16496) );
  NAND2_X1 U16505 ( .A1(n16555), .A2(n16556), .ZN(n16397) );
  INV_X1 U16506 ( .A(n16400), .ZN(n16556) );
  NAND2_X1 U16507 ( .A1(b_0_), .A2(a_15_), .ZN(n16400) );
  NOR2_X1 U16508 ( .A1(n8953), .A2(n8834), .ZN(n16555) );
  NOR2_X1 U16509 ( .A1(n8975), .A2(n8953), .ZN(n16253) );
  OR2_X1 U16510 ( .A1(n16406), .A2(a_12_), .ZN(n16490) );
  NAND2_X1 U16511 ( .A1(n16407), .A2(n16406), .ZN(n16405) );
  NOR2_X1 U16512 ( .A1(n8975), .A2(n8495), .ZN(n16406) );
  NOR2_X1 U16513 ( .A1(n8956), .A2(n8834), .ZN(n16407) );
  NOR2_X1 U16514 ( .A1(n8975), .A2(n8956), .ZN(n16242) );
  OR2_X1 U16515 ( .A1(n16413), .A2(a_10_), .ZN(n16484) );
  NAND2_X1 U16516 ( .A1(n16414), .A2(n16413), .ZN(n16412) );
  NOR2_X1 U16517 ( .A1(n8975), .A2(n8550), .ZN(n16413) );
  NOR2_X1 U16518 ( .A1(n8959), .A2(n8834), .ZN(n16414) );
  NOR2_X1 U16519 ( .A1(n8975), .A2(n8959), .ZN(n16231) );
  OR2_X1 U16520 ( .A1(n16420), .A2(a_8_), .ZN(n16478) );
  NAND2_X1 U16521 ( .A1(n16421), .A2(n16420), .ZN(n16419) );
  NOR2_X1 U16522 ( .A1(n8975), .A2(n8605), .ZN(n16420) );
  NOR2_X1 U16523 ( .A1(n8619), .A2(n8834), .ZN(n16421) );
  NOR2_X1 U16524 ( .A1(n8975), .A2(n8619), .ZN(n16220) );
  OR2_X1 U16525 ( .A1(n16427), .A2(a_6_), .ZN(n16472) );
  NAND2_X1 U16526 ( .A1(n16428), .A2(n16427), .ZN(n16426) );
  NOR2_X1 U16527 ( .A1(n8975), .A2(n8962), .ZN(n16427) );
  NOR2_X1 U16528 ( .A1(n8681), .A2(n8834), .ZN(n16428) );
  NOR2_X1 U16529 ( .A1(n8975), .A2(n8681), .ZN(n16209) );
  OR2_X1 U16530 ( .A1(n16434), .A2(a_4_), .ZN(n16466) );
  NAND2_X1 U16531 ( .A1(n16435), .A2(n16434), .ZN(n16433) );
  NOR2_X1 U16532 ( .A1(n8975), .A2(n8723), .ZN(n16434) );
  NOR2_X1 U16533 ( .A1(n8966), .A2(n8834), .ZN(n16435) );
  NOR2_X1 U16534 ( .A1(n8975), .A2(n8966), .ZN(n16198) );
  OR2_X1 U16535 ( .A1(n16441), .A2(a_2_), .ZN(n16460) );
  NAND2_X1 U16536 ( .A1(n16442), .A2(n16441), .ZN(n16440) );
  NOR2_X1 U16537 ( .A1(n8975), .A2(n8778), .ZN(n16441) );
  NOR2_X1 U16538 ( .A1(n8792), .A2(n8834), .ZN(n16442) );
  NOR2_X1 U16539 ( .A1(n8834), .A2(n8969), .ZN(n8867) );
  OR2_X1 U16540 ( .A1(n16451), .A2(a_0_), .ZN(n16454) );
  NAND2_X1 U16541 ( .A1(n16452), .A2(n16451), .ZN(n16450) );
  NOR2_X1 U16542 ( .A1(n8975), .A2(n8969), .ZN(n16451) );
  NOR2_X1 U16543 ( .A1(n8974), .A2(n8834), .ZN(n16452) );
  NAND2_X1 U16544 ( .A1(b_0_), .A2(a_0_), .ZN(n8972) );
  NAND2_X1 U16545 ( .A1(n16559), .A2(n7955), .ZN(n16558) );
  NOR2_X1 U16546 ( .A1(n16561), .A2(n16562), .ZN(n16559) );
  NOR2_X1 U16547 ( .A1(n8970), .A2(n8974), .ZN(n16562) );
  INV_X1 U16548 ( .A(n8857), .ZN(n8970) );
  NOR2_X1 U16549 ( .A1(b_0_), .A2(n16563), .ZN(n16561) );
  NOR2_X1 U16550 ( .A1(a_0_), .A2(n8857), .ZN(n16563) );
  NAND2_X1 U16551 ( .A1(n16564), .A2(n16565), .ZN(n8857) );
  NAND2_X1 U16552 ( .A1(n16566), .A2(n8834), .ZN(n16565) );
  INV_X1 U16553 ( .A(b_1_), .ZN(n8834) );
  NAND2_X1 U16554 ( .A1(n8830), .A2(n8969), .ZN(n16566) );
  INV_X1 U16555 ( .A(n8839), .ZN(n8830) );
  NAND2_X1 U16556 ( .A1(a_1_), .A2(n8839), .ZN(n16564) );
  NAND2_X1 U16557 ( .A1(n16567), .A2(n16568), .ZN(n8839) );
  NAND2_X1 U16558 ( .A1(n16569), .A2(n8968), .ZN(n16568) );
  INV_X1 U16559 ( .A(b_2_), .ZN(n8968) );
  NAND2_X1 U16560 ( .A1(n8810), .A2(n8792), .ZN(n16569) );
  INV_X1 U16561 ( .A(n8802), .ZN(n8810) );
  NAND2_X1 U16562 ( .A1(a_2_), .A2(n8802), .ZN(n16567) );
  NAND2_X1 U16563 ( .A1(n16570), .A2(n16571), .ZN(n8802) );
  NAND2_X1 U16564 ( .A1(n16572), .A2(n8967), .ZN(n16571) );
  INV_X1 U16565 ( .A(b_3_), .ZN(n8967) );
  NAND2_X1 U16566 ( .A1(n8774), .A2(n8778), .ZN(n16572) );
  INV_X1 U16567 ( .A(n8783), .ZN(n8774) );
  NAND2_X1 U16568 ( .A1(a_3_), .A2(n8783), .ZN(n16570) );
  NAND2_X1 U16569 ( .A1(n16573), .A2(n16574), .ZN(n8783) );
  NAND2_X1 U16570 ( .A1(n16575), .A2(n8965), .ZN(n16574) );
  NAND2_X1 U16571 ( .A1(n8754), .A2(n8966), .ZN(n16575) );
  INV_X1 U16572 ( .A(n8746), .ZN(n8754) );
  NAND2_X1 U16573 ( .A1(a_4_), .A2(n8746), .ZN(n16573) );
  NAND2_X1 U16574 ( .A1(n16576), .A2(n16577), .ZN(n8746) );
  NAND2_X1 U16575 ( .A1(n16578), .A2(n8964), .ZN(n16577) );
  NAND2_X1 U16576 ( .A1(n8719), .A2(n8723), .ZN(n16578) );
  INV_X1 U16577 ( .A(n8728), .ZN(n8719) );
  NAND2_X1 U16578 ( .A1(a_5_), .A2(n8728), .ZN(n16576) );
  NAND2_X1 U16579 ( .A1(n16579), .A2(n16580), .ZN(n8728) );
  NAND2_X1 U16580 ( .A1(n16581), .A2(n8963), .ZN(n16580) );
  NAND2_X1 U16581 ( .A1(n8699), .A2(n8681), .ZN(n16581) );
  INV_X1 U16582 ( .A(n8691), .ZN(n8699) );
  NAND2_X1 U16583 ( .A1(a_6_), .A2(n8691), .ZN(n16579) );
  NAND2_X1 U16584 ( .A1(n16582), .A2(n16583), .ZN(n8691) );
  NAND2_X1 U16585 ( .A1(n16584), .A2(n8667), .ZN(n16583) );
  NAND2_X1 U16586 ( .A1(n8663), .A2(n8962), .ZN(n16584) );
  INV_X1 U16587 ( .A(n8672), .ZN(n8663) );
  NAND2_X1 U16588 ( .A1(a_7_), .A2(n8672), .ZN(n16582) );
  NAND2_X1 U16589 ( .A1(n16585), .A2(n16586), .ZN(n8672) );
  NAND2_X1 U16590 ( .A1(n16587), .A2(n8961), .ZN(n16586) );
  NAND2_X1 U16591 ( .A1(n8637), .A2(n8619), .ZN(n16587) );
  INV_X1 U16592 ( .A(n8629), .ZN(n8637) );
  NAND2_X1 U16593 ( .A1(a_8_), .A2(n8629), .ZN(n16585) );
  NAND2_X1 U16594 ( .A1(n16588), .A2(n16589), .ZN(n8629) );
  NAND2_X1 U16595 ( .A1(n16590), .A2(n8960), .ZN(n16589) );
  INV_X1 U16596 ( .A(b_9_), .ZN(n8960) );
  NAND2_X1 U16597 ( .A1(n8601), .A2(n8605), .ZN(n16590) );
  INV_X1 U16598 ( .A(n8610), .ZN(n8601) );
  NAND2_X1 U16599 ( .A1(a_9_), .A2(n8610), .ZN(n16588) );
  NAND2_X1 U16600 ( .A1(n16591), .A2(n16592), .ZN(n8610) );
  NAND2_X1 U16601 ( .A1(n16593), .A2(n8958), .ZN(n16592) );
  INV_X1 U16602 ( .A(b_10_), .ZN(n8958) );
  NAND2_X1 U16603 ( .A1(n8581), .A2(n8959), .ZN(n16593) );
  INV_X1 U16604 ( .A(n8573), .ZN(n8581) );
  NAND2_X1 U16605 ( .A1(a_10_), .A2(n8573), .ZN(n16591) );
  NAND2_X1 U16606 ( .A1(n16594), .A2(n16595), .ZN(n8573) );
  NAND2_X1 U16607 ( .A1(n16596), .A2(n8957), .ZN(n16595) );
  INV_X1 U16608 ( .A(b_11_), .ZN(n8957) );
  NAND2_X1 U16609 ( .A1(n8546), .A2(n8550), .ZN(n16596) );
  INV_X1 U16610 ( .A(n8555), .ZN(n8546) );
  NAND2_X1 U16611 ( .A1(a_11_), .A2(n8555), .ZN(n16594) );
  NAND2_X1 U16612 ( .A1(n16597), .A2(n16598), .ZN(n8555) );
  NAND2_X1 U16613 ( .A1(n16599), .A2(n8955), .ZN(n16598) );
  INV_X1 U16614 ( .A(b_12_), .ZN(n8955) );
  NAND2_X1 U16615 ( .A1(n8526), .A2(n8956), .ZN(n16599) );
  INV_X1 U16616 ( .A(n8518), .ZN(n8526) );
  NAND2_X1 U16617 ( .A1(a_12_), .A2(n8518), .ZN(n16597) );
  NAND2_X1 U16618 ( .A1(n16600), .A2(n16601), .ZN(n8518) );
  NAND2_X1 U16619 ( .A1(n16602), .A2(n8954), .ZN(n16601) );
  NAND2_X1 U16620 ( .A1(n8491), .A2(n8495), .ZN(n16602) );
  INV_X1 U16621 ( .A(n8500), .ZN(n8491) );
  NAND2_X1 U16622 ( .A1(a_13_), .A2(n8500), .ZN(n16600) );
  NAND2_X1 U16623 ( .A1(n16603), .A2(n16604), .ZN(n8500) );
  NAND2_X1 U16624 ( .A1(n16605), .A2(n8952), .ZN(n16604) );
  INV_X1 U16625 ( .A(b_14_), .ZN(n8952) );
  NAND2_X1 U16626 ( .A1(n8471), .A2(n8953), .ZN(n16605) );
  INV_X1 U16627 ( .A(n8463), .ZN(n8471) );
  NAND2_X1 U16628 ( .A1(a_14_), .A2(n8463), .ZN(n16603) );
  NAND2_X1 U16629 ( .A1(n16606), .A2(n16607), .ZN(n8463) );
  NAND2_X1 U16630 ( .A1(n16608), .A2(n8951), .ZN(n16607) );
  NAND2_X1 U16631 ( .A1(n8436), .A2(n8440), .ZN(n16608) );
  INV_X1 U16632 ( .A(n8445), .ZN(n8436) );
  NAND2_X1 U16633 ( .A1(a_15_), .A2(n8445), .ZN(n16606) );
  NAND2_X1 U16634 ( .A1(n16609), .A2(n16610), .ZN(n8445) );
  NAND2_X1 U16635 ( .A1(n16611), .A2(n8949), .ZN(n16610) );
  INV_X1 U16636 ( .A(b_16_), .ZN(n8949) );
  NAND2_X1 U16637 ( .A1(n8416), .A2(n8950), .ZN(n16611) );
  INV_X1 U16638 ( .A(n8408), .ZN(n8416) );
  NAND2_X1 U16639 ( .A1(a_16_), .A2(n8408), .ZN(n16609) );
  NAND2_X1 U16640 ( .A1(n16612), .A2(n16613), .ZN(n8408) );
  NAND2_X1 U16641 ( .A1(n16614), .A2(n8948), .ZN(n16613) );
  NAND2_X1 U16642 ( .A1(n8381), .A2(n8385), .ZN(n16614) );
  INV_X1 U16643 ( .A(n8390), .ZN(n8381) );
  NAND2_X1 U16644 ( .A1(a_17_), .A2(n8390), .ZN(n16612) );
  NAND2_X1 U16645 ( .A1(n16615), .A2(n16616), .ZN(n8390) );
  NAND2_X1 U16646 ( .A1(n16617), .A2(n8946), .ZN(n16616) );
  INV_X1 U16647 ( .A(b_18_), .ZN(n8946) );
  NAND2_X1 U16648 ( .A1(n8355), .A2(n8947), .ZN(n16617) );
  INV_X1 U16649 ( .A(n8347), .ZN(n8355) );
  NAND2_X1 U16650 ( .A1(a_18_), .A2(n8347), .ZN(n16615) );
  NAND2_X1 U16651 ( .A1(n16618), .A2(n16619), .ZN(n8347) );
  NAND2_X1 U16652 ( .A1(n16620), .A2(n8945), .ZN(n16619) );
  NAND2_X1 U16653 ( .A1(n8320), .A2(n8324), .ZN(n16620) );
  INV_X1 U16654 ( .A(n8329), .ZN(n8320) );
  NAND2_X1 U16655 ( .A1(a_19_), .A2(n8329), .ZN(n16618) );
  NAND2_X1 U16656 ( .A1(n16621), .A2(n16622), .ZN(n8329) );
  NAND2_X1 U16657 ( .A1(n16623), .A2(n8943), .ZN(n16622) );
  INV_X1 U16658 ( .A(b_20_), .ZN(n8943) );
  NAND2_X1 U16659 ( .A1(n8300), .A2(n8944), .ZN(n16623) );
  INV_X1 U16660 ( .A(n8291), .ZN(n8300) );
  NAND2_X1 U16661 ( .A1(a_20_), .A2(n8291), .ZN(n16621) );
  NAND2_X1 U16662 ( .A1(n16624), .A2(n16625), .ZN(n8291) );
  NAND2_X1 U16663 ( .A1(n16626), .A2(n8942), .ZN(n16625) );
  NAND2_X1 U16664 ( .A1(n8264), .A2(n8268), .ZN(n16626) );
  INV_X1 U16665 ( .A(n8273), .ZN(n8264) );
  NAND2_X1 U16666 ( .A1(a_21_), .A2(n8273), .ZN(n16624) );
  NAND2_X1 U16667 ( .A1(n16627), .A2(n16628), .ZN(n8273) );
  NAND2_X1 U16668 ( .A1(n16629), .A2(n8240), .ZN(n16628) );
  NAND2_X1 U16669 ( .A1(n8236), .A2(n8941), .ZN(n16629) );
  INV_X1 U16670 ( .A(n8246), .ZN(n8236) );
  NAND2_X1 U16671 ( .A1(a_22_), .A2(n8246), .ZN(n16627) );
  NAND2_X1 U16672 ( .A1(n16630), .A2(n16631), .ZN(n8246) );
  NAND2_X1 U16673 ( .A1(n16632), .A2(n8940), .ZN(n16631) );
  NAND2_X1 U16674 ( .A1(n8209), .A2(n8213), .ZN(n16632) );
  INV_X1 U16675 ( .A(n8218), .ZN(n8209) );
  NAND2_X1 U16676 ( .A1(a_23_), .A2(n8218), .ZN(n16630) );
  NAND2_X1 U16677 ( .A1(n16633), .A2(n16634), .ZN(n8218) );
  NAND2_X1 U16678 ( .A1(n16635), .A2(n8185), .ZN(n16634) );
  NAND2_X1 U16679 ( .A1(n8181), .A2(n8939), .ZN(n16635) );
  INV_X1 U16680 ( .A(n8191), .ZN(n8181) );
  NAND2_X1 U16681 ( .A1(a_24_), .A2(n8191), .ZN(n16633) );
  NAND2_X1 U16682 ( .A1(n16636), .A2(n16637), .ZN(n8191) );
  NAND2_X1 U16683 ( .A1(n16638), .A2(n8938), .ZN(n16637) );
  NAND2_X1 U16684 ( .A1(n8154), .A2(n8158), .ZN(n16638) );
  INV_X1 U16685 ( .A(n8163), .ZN(n8154) );
  NAND2_X1 U16686 ( .A1(a_25_), .A2(n8163), .ZN(n16636) );
  NAND2_X1 U16687 ( .A1(n16639), .A2(n16640), .ZN(n8163) );
  NAND2_X1 U16688 ( .A1(n16641), .A2(n8130), .ZN(n16640) );
  NAND2_X1 U16689 ( .A1(n8126), .A2(n8116), .ZN(n16641) );
  INV_X1 U16690 ( .A(n8136), .ZN(n8126) );
  NAND2_X1 U16691 ( .A1(a_26_), .A2(n8136), .ZN(n16639) );
  NAND2_X1 U16692 ( .A1(n16642), .A2(n16643), .ZN(n8136) );
  NAND2_X1 U16693 ( .A1(n16644), .A2(n8102), .ZN(n16643) );
  NAND2_X1 U16694 ( .A1(n8098), .A2(n8937), .ZN(n16644) );
  INV_X1 U16695 ( .A(n8107), .ZN(n8098) );
  NAND2_X1 U16696 ( .A1(a_27_), .A2(n8107), .ZN(n16642) );
  NAND2_X1 U16697 ( .A1(n16645), .A2(n16646), .ZN(n8107) );
  NAND2_X1 U16698 ( .A1(n16647), .A2(n8069), .ZN(n16646) );
  NAND2_X1 U16699 ( .A1(n8065), .A2(n8055), .ZN(n16647) );
  INV_X1 U16700 ( .A(n8074), .ZN(n8065) );
  NAND2_X1 U16701 ( .A1(a_28_), .A2(n8074), .ZN(n16645) );
  NAND2_X1 U16702 ( .A1(n16648), .A2(n16649), .ZN(n8074) );
  NAND2_X1 U16703 ( .A1(n16650), .A2(n8936), .ZN(n16649) );
  NAND2_X1 U16704 ( .A1(n8037), .A2(n8041), .ZN(n16650) );
  INV_X1 U16705 ( .A(n8046), .ZN(n8037) );
  NAND2_X1 U16706 ( .A1(a_29_), .A2(n8046), .ZN(n16648) );
  NAND2_X1 U16707 ( .A1(n8000), .A2(n16651), .ZN(n8046) );
  NAND2_X1 U16708 ( .A1(n8020), .A2(n7990), .ZN(n16651) );
  NAND2_X1 U16709 ( .A1(b_31_), .A2(n16335), .ZN(n7990) );
  INV_X1 U16710 ( .A(a_31_), .ZN(n16335) );
  NAND2_X1 U16711 ( .A1(n16652), .A2(n7988), .ZN(n16557) );
  INV_X1 U16712 ( .A(n8013), .ZN(n7988) );
  INV_X1 U16713 ( .A(operation_1_), .ZN(n16560) );
  NOR2_X1 U16714 ( .A1(n16653), .A2(n16654), .ZN(n16652) );
  NOR2_X1 U16715 ( .A1(a_0_), .A2(n8858), .ZN(n16654) );
  INV_X1 U16716 ( .A(n8971), .ZN(n8858) );
  NOR2_X1 U16717 ( .A1(n16655), .A2(n8975), .ZN(n16653) );
  NOR2_X1 U16718 ( .A1(n8974), .A2(n8971), .ZN(n16655) );
  NAND2_X1 U16719 ( .A1(n16656), .A2(n16657), .ZN(n8971) );
  NAND2_X1 U16720 ( .A1(b_1_), .A2(n16658), .ZN(n16657) );
  NAND2_X1 U16721 ( .A1(n8840), .A2(a_1_), .ZN(n16658) );
  INV_X1 U16722 ( .A(n8831), .ZN(n8840) );
  NAND2_X1 U16723 ( .A1(n8831), .A2(n8969), .ZN(n16656) );
  NAND2_X1 U16724 ( .A1(n16659), .A2(n16660), .ZN(n8831) );
  NAND2_X1 U16725 ( .A1(b_2_), .A2(n16661), .ZN(n16660) );
  NAND2_X1 U16726 ( .A1(n8803), .A2(a_2_), .ZN(n16661) );
  INV_X1 U16727 ( .A(n8811), .ZN(n8803) );
  NAND2_X1 U16728 ( .A1(n8811), .A2(n8792), .ZN(n16659) );
  NAND2_X1 U16729 ( .A1(n16662), .A2(n16663), .ZN(n8811) );
  NAND2_X1 U16730 ( .A1(b_3_), .A2(n16664), .ZN(n16663) );
  NAND2_X1 U16731 ( .A1(n8784), .A2(a_3_), .ZN(n16664) );
  INV_X1 U16732 ( .A(n8775), .ZN(n8784) );
  NAND2_X1 U16733 ( .A1(n8775), .A2(n8778), .ZN(n16662) );
  NAND2_X1 U16734 ( .A1(n16665), .A2(n16666), .ZN(n8775) );
  NAND2_X1 U16735 ( .A1(b_4_), .A2(n16667), .ZN(n16666) );
  NAND2_X1 U16736 ( .A1(n8747), .A2(a_4_), .ZN(n16667) );
  INV_X1 U16737 ( .A(n8755), .ZN(n8747) );
  NAND2_X1 U16738 ( .A1(n8755), .A2(n8966), .ZN(n16665) );
  NAND2_X1 U16739 ( .A1(n16668), .A2(n16669), .ZN(n8755) );
  NAND2_X1 U16740 ( .A1(b_5_), .A2(n16670), .ZN(n16669) );
  NAND2_X1 U16741 ( .A1(n8729), .A2(a_5_), .ZN(n16670) );
  INV_X1 U16742 ( .A(n8720), .ZN(n8729) );
  NAND2_X1 U16743 ( .A1(n8720), .A2(n8723), .ZN(n16668) );
  NAND2_X1 U16744 ( .A1(n16671), .A2(n16672), .ZN(n8720) );
  NAND2_X1 U16745 ( .A1(b_6_), .A2(n16673), .ZN(n16672) );
  NAND2_X1 U16746 ( .A1(n8692), .A2(a_6_), .ZN(n16673) );
  INV_X1 U16747 ( .A(n8700), .ZN(n8692) );
  NAND2_X1 U16748 ( .A1(n8700), .A2(n8681), .ZN(n16671) );
  NAND2_X1 U16749 ( .A1(n16674), .A2(n16675), .ZN(n8700) );
  NAND2_X1 U16750 ( .A1(b_7_), .A2(n16676), .ZN(n16675) );
  NAND2_X1 U16751 ( .A1(n8673), .A2(a_7_), .ZN(n16676) );
  INV_X1 U16752 ( .A(n8664), .ZN(n8673) );
  NAND2_X1 U16753 ( .A1(n8664), .A2(n8962), .ZN(n16674) );
  NAND2_X1 U16754 ( .A1(n16677), .A2(n16678), .ZN(n8664) );
  NAND2_X1 U16755 ( .A1(b_8_), .A2(n16679), .ZN(n16678) );
  NAND2_X1 U16756 ( .A1(n8630), .A2(a_8_), .ZN(n16679) );
  INV_X1 U16757 ( .A(n8638), .ZN(n8630) );
  NAND2_X1 U16758 ( .A1(n8638), .A2(n8619), .ZN(n16677) );
  NAND2_X1 U16759 ( .A1(n16680), .A2(n16681), .ZN(n8638) );
  NAND2_X1 U16760 ( .A1(b_9_), .A2(n16682), .ZN(n16681) );
  NAND2_X1 U16761 ( .A1(n8611), .A2(a_9_), .ZN(n16682) );
  INV_X1 U16762 ( .A(n8602), .ZN(n8611) );
  NAND2_X1 U16763 ( .A1(n8602), .A2(n8605), .ZN(n16680) );
  NAND2_X1 U16764 ( .A1(n16683), .A2(n16684), .ZN(n8602) );
  NAND2_X1 U16765 ( .A1(b_10_), .A2(n16685), .ZN(n16684) );
  NAND2_X1 U16766 ( .A1(n8574), .A2(a_10_), .ZN(n16685) );
  INV_X1 U16767 ( .A(n8582), .ZN(n8574) );
  NAND2_X1 U16768 ( .A1(n8582), .A2(n8959), .ZN(n16683) );
  NAND2_X1 U16769 ( .A1(n16686), .A2(n16687), .ZN(n8582) );
  NAND2_X1 U16770 ( .A1(b_11_), .A2(n16688), .ZN(n16687) );
  NAND2_X1 U16771 ( .A1(n8556), .A2(a_11_), .ZN(n16688) );
  INV_X1 U16772 ( .A(n8547), .ZN(n8556) );
  NAND2_X1 U16773 ( .A1(n8547), .A2(n8550), .ZN(n16686) );
  NAND2_X1 U16774 ( .A1(n16689), .A2(n16690), .ZN(n8547) );
  NAND2_X1 U16775 ( .A1(b_12_), .A2(n16691), .ZN(n16690) );
  NAND2_X1 U16776 ( .A1(n8519), .A2(a_12_), .ZN(n16691) );
  INV_X1 U16777 ( .A(n8527), .ZN(n8519) );
  NAND2_X1 U16778 ( .A1(n8527), .A2(n8956), .ZN(n16689) );
  NAND2_X1 U16779 ( .A1(n16692), .A2(n16693), .ZN(n8527) );
  NAND2_X1 U16780 ( .A1(b_13_), .A2(n16694), .ZN(n16693) );
  NAND2_X1 U16781 ( .A1(n8501), .A2(a_13_), .ZN(n16694) );
  INV_X1 U16782 ( .A(n8492), .ZN(n8501) );
  NAND2_X1 U16783 ( .A1(n8492), .A2(n8495), .ZN(n16692) );
  NAND2_X1 U16784 ( .A1(n16695), .A2(n16696), .ZN(n8492) );
  NAND2_X1 U16785 ( .A1(b_14_), .A2(n16697), .ZN(n16696) );
  NAND2_X1 U16786 ( .A1(n8464), .A2(a_14_), .ZN(n16697) );
  INV_X1 U16787 ( .A(n8472), .ZN(n8464) );
  NAND2_X1 U16788 ( .A1(n8472), .A2(n8953), .ZN(n16695) );
  NAND2_X1 U16789 ( .A1(n16698), .A2(n16699), .ZN(n8472) );
  NAND2_X1 U16790 ( .A1(b_15_), .A2(n16700), .ZN(n16699) );
  NAND2_X1 U16791 ( .A1(n8446), .A2(a_15_), .ZN(n16700) );
  INV_X1 U16792 ( .A(n8437), .ZN(n8446) );
  NAND2_X1 U16793 ( .A1(n8437), .A2(n8440), .ZN(n16698) );
  NAND2_X1 U16794 ( .A1(n16701), .A2(n16702), .ZN(n8437) );
  NAND2_X1 U16795 ( .A1(b_16_), .A2(n16703), .ZN(n16702) );
  NAND2_X1 U16796 ( .A1(n8409), .A2(a_16_), .ZN(n16703) );
  INV_X1 U16797 ( .A(n8417), .ZN(n8409) );
  NAND2_X1 U16798 ( .A1(n8417), .A2(n8950), .ZN(n16701) );
  NAND2_X1 U16799 ( .A1(n16704), .A2(n16705), .ZN(n8417) );
  NAND2_X1 U16800 ( .A1(b_17_), .A2(n16706), .ZN(n16705) );
  NAND2_X1 U16801 ( .A1(n8391), .A2(a_17_), .ZN(n16706) );
  INV_X1 U16802 ( .A(n8382), .ZN(n8391) );
  NAND2_X1 U16803 ( .A1(n8382), .A2(n8385), .ZN(n16704) );
  NAND2_X1 U16804 ( .A1(n16707), .A2(n16708), .ZN(n8382) );
  NAND2_X1 U16805 ( .A1(b_18_), .A2(n16709), .ZN(n16708) );
  NAND2_X1 U16806 ( .A1(n8348), .A2(a_18_), .ZN(n16709) );
  INV_X1 U16807 ( .A(n8356), .ZN(n8348) );
  NAND2_X1 U16808 ( .A1(n8356), .A2(n8947), .ZN(n16707) );
  NAND2_X1 U16809 ( .A1(n16710), .A2(n16711), .ZN(n8356) );
  NAND2_X1 U16810 ( .A1(b_19_), .A2(n16712), .ZN(n16711) );
  NAND2_X1 U16811 ( .A1(n8330), .A2(a_19_), .ZN(n16712) );
  INV_X1 U16812 ( .A(n8321), .ZN(n8330) );
  NAND2_X1 U16813 ( .A1(n8321), .A2(n8324), .ZN(n16710) );
  NAND2_X1 U16814 ( .A1(n16713), .A2(n16714), .ZN(n8321) );
  NAND2_X1 U16815 ( .A1(b_20_), .A2(n16715), .ZN(n16714) );
  NAND2_X1 U16816 ( .A1(n8292), .A2(a_20_), .ZN(n16715) );
  INV_X1 U16817 ( .A(n8301), .ZN(n8292) );
  NAND2_X1 U16818 ( .A1(n8301), .A2(n8944), .ZN(n16713) );
  NAND2_X1 U16819 ( .A1(n16716), .A2(n16717), .ZN(n8301) );
  NAND2_X1 U16820 ( .A1(b_21_), .A2(n16718), .ZN(n16717) );
  NAND2_X1 U16821 ( .A1(n8274), .A2(a_21_), .ZN(n16718) );
  INV_X1 U16822 ( .A(n8265), .ZN(n8274) );
  NAND2_X1 U16823 ( .A1(n8265), .A2(n8268), .ZN(n16716) );
  NAND2_X1 U16824 ( .A1(n16719), .A2(n16720), .ZN(n8265) );
  NAND2_X1 U16825 ( .A1(b_22_), .A2(n16721), .ZN(n16720) );
  NAND2_X1 U16826 ( .A1(n8247), .A2(a_22_), .ZN(n16721) );
  INV_X1 U16827 ( .A(n8237), .ZN(n8247) );
  NAND2_X1 U16828 ( .A1(n8237), .A2(n8941), .ZN(n16719) );
  NAND2_X1 U16829 ( .A1(n16722), .A2(n16723), .ZN(n8237) );
  NAND2_X1 U16830 ( .A1(b_23_), .A2(n16724), .ZN(n16723) );
  NAND2_X1 U16831 ( .A1(n8219), .A2(a_23_), .ZN(n16724) );
  INV_X1 U16832 ( .A(n8210), .ZN(n8219) );
  NAND2_X1 U16833 ( .A1(n8210), .A2(n8213), .ZN(n16722) );
  NAND2_X1 U16834 ( .A1(n16725), .A2(n16726), .ZN(n8210) );
  NAND2_X1 U16835 ( .A1(b_24_), .A2(n16727), .ZN(n16726) );
  NAND2_X1 U16836 ( .A1(n8192), .A2(a_24_), .ZN(n16727) );
  INV_X1 U16837 ( .A(n8182), .ZN(n8192) );
  NAND2_X1 U16838 ( .A1(n8182), .A2(n8939), .ZN(n16725) );
  NAND2_X1 U16839 ( .A1(n16728), .A2(n16729), .ZN(n8182) );
  NAND2_X1 U16840 ( .A1(b_25_), .A2(n16730), .ZN(n16729) );
  NAND2_X1 U16841 ( .A1(n8164), .A2(a_25_), .ZN(n16730) );
  INV_X1 U16842 ( .A(n8155), .ZN(n8164) );
  NAND2_X1 U16843 ( .A1(n8155), .A2(n8158), .ZN(n16728) );
  NAND2_X1 U16844 ( .A1(n16731), .A2(n16732), .ZN(n8155) );
  NAND2_X1 U16845 ( .A1(b_26_), .A2(n16733), .ZN(n16732) );
  NAND2_X1 U16846 ( .A1(n8137), .A2(a_26_), .ZN(n16733) );
  INV_X1 U16847 ( .A(n8127), .ZN(n8137) );
  NAND2_X1 U16848 ( .A1(n8127), .A2(n8116), .ZN(n16731) );
  INV_X1 U16849 ( .A(a_26_), .ZN(n8116) );
  NAND2_X1 U16850 ( .A1(n16734), .A2(n16735), .ZN(n8127) );
  NAND2_X1 U16851 ( .A1(b_27_), .A2(n16736), .ZN(n16735) );
  NAND2_X1 U16852 ( .A1(n8108), .A2(a_27_), .ZN(n16736) );
  INV_X1 U16853 ( .A(n8099), .ZN(n8108) );
  NAND2_X1 U16854 ( .A1(n8099), .A2(n8937), .ZN(n16734) );
  INV_X1 U16855 ( .A(a_27_), .ZN(n8937) );
  NAND2_X1 U16856 ( .A1(n16737), .A2(n16738), .ZN(n8099) );
  NAND2_X1 U16857 ( .A1(b_28_), .A2(n16739), .ZN(n16738) );
  NAND2_X1 U16858 ( .A1(n8075), .A2(a_28_), .ZN(n16739) );
  INV_X1 U16859 ( .A(n8066), .ZN(n8075) );
  NAND2_X1 U16860 ( .A1(n8066), .A2(n8055), .ZN(n16737) );
  NAND2_X1 U16861 ( .A1(n16740), .A2(n16741), .ZN(n8066) );
  NAND2_X1 U16862 ( .A1(b_29_), .A2(n16742), .ZN(n16741) );
  NAND2_X1 U16863 ( .A1(n8047), .A2(a_29_), .ZN(n16742) );
  INV_X1 U16864 ( .A(n8038), .ZN(n8047) );
  NAND2_X1 U16865 ( .A1(n8038), .A2(n8041), .ZN(n16740) );
  NAND2_X1 U16866 ( .A1(n8020), .A2(n16743), .ZN(n8038) );
  NAND2_X1 U16867 ( .A1(n7989), .A2(n8000), .ZN(n16743) );
  NAND2_X1 U16868 ( .A1(a_30_), .A2(n8002), .ZN(n8000) );
  NAND2_X1 U16869 ( .A1(a_31_), .A2(n7999), .ZN(n7989) );
  NAND2_X1 U16870 ( .A1(b_30_), .A2(n8935), .ZN(n8020) );
  INV_X1 U16871 ( .A(a_30_), .ZN(n8935) );
endmodule

